magic
tech sky130A
magscale 1 2
timestamp 1712639104
<< nwell >>
rect -658 -815 658 815
<< mvpmos >>
rect -400 118 400 518
rect -400 -518 400 -118
<< mvpdiff >>
rect -458 506 -400 518
rect -458 130 -446 506
rect -412 130 -400 506
rect -458 118 -400 130
rect 400 506 458 518
rect 400 130 412 506
rect 446 130 458 506
rect 400 118 458 130
rect -458 -130 -400 -118
rect -458 -506 -446 -130
rect -412 -506 -400 -130
rect -458 -518 -400 -506
rect 400 -130 458 -118
rect 400 -506 412 -130
rect 446 -506 458 -130
rect 400 -518 458 -506
<< mvpdiffc >>
rect -446 130 -412 506
rect 412 130 446 506
rect -446 -506 -412 -130
rect 412 -506 446 -130
<< mvnsubdiff >>
rect -592 737 592 749
rect -592 703 -484 737
rect 484 703 592 737
rect -592 691 592 703
rect -592 641 -534 691
rect -592 -641 -580 641
rect -546 -641 -534 641
rect 534 641 592 691
rect -592 -691 -534 -641
rect 534 -641 546 641
rect 580 -641 592 641
rect 534 -691 592 -641
rect -592 -703 592 -691
rect -592 -737 -484 -703
rect 484 -737 592 -703
rect -592 -749 592 -737
<< mvnsubdiffcont >>
rect -484 703 484 737
rect -580 -641 -546 641
rect 546 -641 580 641
rect -484 -737 484 -703
<< poly >>
rect -400 599 400 615
rect -400 565 -384 599
rect 384 565 400 599
rect -400 518 400 565
rect -400 71 400 118
rect -400 37 -384 71
rect 384 37 400 71
rect -400 21 400 37
rect -400 -37 400 -21
rect -400 -71 -384 -37
rect 384 -71 400 -37
rect -400 -118 400 -71
rect -400 -565 400 -518
rect -400 -599 -384 -565
rect 384 -599 400 -565
rect -400 -615 400 -599
<< polycont >>
rect -384 565 384 599
rect -384 37 384 71
rect -384 -71 384 -37
rect -384 -599 384 -565
<< locali >>
rect -580 703 -484 737
rect 484 703 580 737
rect -580 641 -546 703
rect 546 641 580 703
rect -400 565 -384 599
rect 384 565 400 599
rect -446 506 -412 522
rect -446 114 -412 130
rect 412 506 446 522
rect 412 114 446 130
rect -400 37 -384 71
rect 384 37 400 71
rect -400 -71 -384 -37
rect 384 -71 400 -37
rect -446 -130 -412 -114
rect -446 -522 -412 -506
rect 412 -130 446 -114
rect 412 -522 446 -506
rect -400 -599 -384 -565
rect 384 -599 400 -565
rect -580 -703 -546 -641
rect 546 -703 580 -641
rect -580 -737 -484 -703
rect 484 -737 580 -703
<< viali >>
rect -346 565 346 599
rect -580 -562 -546 562
rect -446 130 -412 506
rect 412 130 446 506
rect -346 37 346 71
rect -346 -71 346 -37
rect -446 -506 -412 -130
rect 412 -506 446 -130
rect -346 -599 346 -565
<< metal1 >>
rect -358 599 358 605
rect -586 562 -540 574
rect -586 -562 -580 562
rect -546 -562 -540 562
rect -358 565 -346 599
rect 346 565 358 599
rect -358 559 358 565
rect -452 506 -406 518
rect -452 130 -446 506
rect -412 130 -406 506
rect -452 118 -406 130
rect 406 506 452 518
rect 406 130 412 506
rect 446 130 452 506
rect 406 118 452 130
rect -358 71 358 77
rect -358 37 -346 71
rect 346 37 358 71
rect -358 31 358 37
rect -358 -37 358 -31
rect -358 -71 -346 -37
rect 346 -71 358 -37
rect -358 -77 358 -71
rect -452 -130 -406 -118
rect -452 -506 -446 -130
rect -412 -506 -406 -130
rect -452 -518 -406 -506
rect 406 -130 452 -118
rect 406 -506 412 -130
rect 446 -506 452 -130
rect 406 -518 452 -506
rect -586 -574 -540 -562
rect -358 -565 358 -559
rect -358 -599 -346 -565
rect 346 -599 358 -565
rect -358 -605 358 -599
<< properties >>
string FIXED_BBOX -563 -720 563 720
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 2 l 4 m 2 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 90 viagb 0 viagr 0 viagl 80 viagt 0
<< end >>
