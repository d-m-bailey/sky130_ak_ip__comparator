magic
tech sky130A
magscale 1 2
timestamp 1713575861
<< nwell >>
rect -1087 -497 1087 497
<< mvpmos >>
rect -829 -200 -29 200
rect 29 -200 829 200
<< mvpdiff >>
rect -887 188 -829 200
rect -887 -188 -875 188
rect -841 -188 -829 188
rect -887 -200 -829 -188
rect -29 188 29 200
rect -29 -188 -17 188
rect 17 -188 29 188
rect -29 -200 29 -188
rect 829 188 887 200
rect 829 -188 841 188
rect 875 -188 887 188
rect 829 -200 887 -188
<< mvpdiffc >>
rect -875 -188 -841 188
rect -17 -188 17 188
rect 841 -188 875 188
<< mvnsubdiff >>
rect -1021 419 1021 431
rect -1021 385 -913 419
rect 913 385 1021 419
rect -1021 373 1021 385
rect -1021 323 -963 373
rect -1021 -323 -1009 323
rect -975 -323 -963 323
rect 963 323 1021 373
rect -1021 -373 -963 -323
rect 963 -323 975 323
rect 1009 -323 1021 323
rect 963 -373 1021 -323
rect -1021 -385 1021 -373
rect -1021 -419 -913 -385
rect 913 -419 1021 -385
rect -1021 -431 1021 -419
<< mvnsubdiffcont >>
rect -913 385 913 419
rect -1009 -323 -975 323
rect 975 -323 1009 323
rect -913 -419 913 -385
<< poly >>
rect -829 281 -29 297
rect -829 247 -813 281
rect -45 247 -29 281
rect -829 200 -29 247
rect 29 281 829 297
rect 29 247 45 281
rect 813 247 829 281
rect 29 200 829 247
rect -829 -247 -29 -200
rect -829 -281 -813 -247
rect -45 -281 -29 -247
rect -829 -297 -29 -281
rect 29 -247 829 -200
rect 29 -281 45 -247
rect 813 -281 829 -247
rect 29 -297 829 -281
<< polycont >>
rect -813 247 -45 281
rect 45 247 813 281
rect -813 -281 -45 -247
rect 45 -281 813 -247
<< locali >>
rect -1009 385 -913 419
rect 913 385 1009 419
rect -1009 323 -975 385
rect 975 323 1009 385
rect -829 247 -813 281
rect -45 247 -29 281
rect 29 247 45 281
rect 813 247 829 281
rect -875 188 -841 204
rect -875 -204 -841 -188
rect -17 188 17 204
rect -17 -204 17 -188
rect 841 188 875 204
rect 841 -204 875 -188
rect -829 -281 -813 -247
rect -45 -281 -29 -247
rect 29 -281 45 -247
rect 813 -281 829 -247
rect -1009 -385 -975 -323
rect 975 -385 1009 -323
rect -1009 -419 -913 -385
rect 913 -419 1009 -385
<< viali >>
rect -780 385 780 419
rect -813 247 -45 281
rect 45 247 813 281
rect -1009 -154 -975 154
rect -875 -188 -841 188
rect -17 -188 17 188
rect 841 -188 875 188
rect 975 -154 1009 154
rect -813 -281 -45 -247
rect 45 -281 813 -247
<< metal1 >>
rect -792 419 792 425
rect -792 385 -780 419
rect 780 385 792 419
rect -792 379 792 385
rect -825 281 -33 287
rect -825 247 -813 281
rect -45 247 -33 281
rect -825 241 -33 247
rect 33 281 825 287
rect 33 247 45 281
rect 813 247 825 281
rect 33 241 825 247
rect -881 188 -835 200
rect -1015 154 -969 166
rect -1015 -154 -1009 154
rect -975 -154 -969 154
rect -1015 -166 -969 -154
rect -881 -188 -875 188
rect -841 -188 -835 188
rect -881 -200 -835 -188
rect -23 188 23 200
rect -23 -188 -17 188
rect 17 -188 23 188
rect -23 -200 23 -188
rect 835 188 881 200
rect 835 -188 841 188
rect 875 -188 881 188
rect 969 154 1015 166
rect 969 -154 975 154
rect 1009 -154 1015 154
rect 969 -166 1015 -154
rect 835 -200 881 -188
rect -825 -247 -33 -241
rect -825 -281 -813 -247
rect -45 -281 -33 -247
rect -825 -287 -33 -281
rect 33 -247 825 -241
rect 33 -281 45 -247
rect 813 -281 825 -247
rect 33 -287 825 -281
<< properties >>
string FIXED_BBOX -992 -402 992 402
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 2 l 4 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 40 viagl 40 viagt 80
<< end >>
