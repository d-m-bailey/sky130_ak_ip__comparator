magic
tech sky130A
magscale 1 2
timestamp 1713576162
<< nwell >>
rect -358 -1215 358 1215
<< mvpmos >>
rect -100 118 100 918
rect -100 -918 100 -118
<< mvpdiff >>
rect -158 906 -100 918
rect -158 130 -146 906
rect -112 130 -100 906
rect -158 118 -100 130
rect 100 906 158 918
rect 100 130 112 906
rect 146 130 158 906
rect 100 118 158 130
rect -158 -130 -100 -118
rect -158 -906 -146 -130
rect -112 -906 -100 -130
rect -158 -918 -100 -906
rect 100 -130 158 -118
rect 100 -906 112 -130
rect 146 -906 158 -130
rect 100 -918 158 -906
<< mvpdiffc >>
rect -146 130 -112 906
rect 112 130 146 906
rect -146 -906 -112 -130
rect 112 -906 146 -130
<< mvnsubdiff >>
rect -292 1137 292 1149
rect -292 1103 -184 1137
rect 184 1103 292 1137
rect -292 1091 292 1103
rect -292 -1091 -234 1091
rect 234 -1091 292 1091
rect -292 -1103 292 -1091
rect -292 -1137 -184 -1103
rect 184 -1137 292 -1103
rect -292 -1149 292 -1137
<< mvnsubdiffcont >>
rect -184 1103 184 1137
rect -184 -1137 184 -1103
<< poly >>
rect -100 999 100 1015
rect -100 965 -84 999
rect 84 965 100 999
rect -100 918 100 965
rect -100 71 100 118
rect -100 37 -84 71
rect 84 37 100 71
rect -100 21 100 37
rect -100 -37 100 -21
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -100 -118 100 -71
rect -100 -965 100 -918
rect -100 -999 -84 -965
rect 84 -999 100 -965
rect -100 -1015 100 -999
<< polycont >>
rect -84 965 84 999
rect -84 37 84 71
rect -84 -71 84 -37
rect -84 -999 84 -965
<< locali >>
rect -280 1103 -184 1137
rect 184 1103 280 1137
rect -280 882 -246 1103
rect -100 965 -84 999
rect 84 965 100 999
rect -146 906 -112 922
rect -146 114 -112 130
rect 112 906 146 922
rect 112 114 146 130
rect 246 882 280 1103
rect -100 37 -84 71
rect 84 37 100 71
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -280 -1103 -246 -882
rect -146 -130 -112 -114
rect -146 -922 -112 -906
rect 112 -130 146 -114
rect 112 -922 146 -906
rect -100 -999 -84 -965
rect 84 -999 100 -965
rect 246 -1103 280 -882
rect -280 -1137 -197 -1103
rect 197 -1137 280 -1103
<< viali >>
rect -50 965 50 999
rect -280 -882 -246 882
rect -146 130 -112 906
rect 112 130 146 906
rect -50 37 50 71
rect -50 -71 50 -37
rect -146 -906 -112 -130
rect 112 -906 146 -130
rect 246 -882 280 882
rect -50 -999 50 -965
rect -197 -1137 -184 -1103
rect -184 -1137 184 -1103
rect 184 -1137 197 -1103
<< metal1 >>
rect -62 999 62 1005
rect -62 965 -50 999
rect 50 965 62 999
rect -62 959 62 965
rect -152 906 -106 918
rect -286 882 -240 894
rect -286 -882 -280 882
rect -246 -882 -240 882
rect -152 130 -146 906
rect -112 130 -106 906
rect -152 118 -106 130
rect 106 906 152 918
rect 106 130 112 906
rect 146 130 152 906
rect 106 118 152 130
rect 240 882 286 894
rect -62 71 62 77
rect -62 37 -50 71
rect 50 37 62 71
rect -62 31 62 37
rect -62 -37 62 -31
rect -62 -71 -50 -37
rect 50 -71 62 -37
rect -62 -77 62 -71
rect -286 -894 -240 -882
rect -152 -130 -106 -118
rect -152 -906 -146 -130
rect -112 -906 -106 -130
rect -152 -918 -106 -906
rect 106 -130 152 -118
rect 106 -906 112 -130
rect 146 -906 152 -130
rect 240 -882 246 882
rect 280 -882 286 882
rect 240 -894 286 -882
rect 106 -918 152 -906
rect -62 -965 62 -959
rect -62 -999 -50 -965
rect 50 -999 62 -965
rect -62 -1005 62 -999
rect -209 -1103 209 -1097
rect -209 -1137 -197 -1103
rect 197 -1137 209 -1103
rect -209 -1143 209 -1137
<< properties >>
string FIXED_BBOX -263 -1120 263 1120
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 4 l 1 m 2 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 0 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 60 viagb 80 viagr 80 viagl 80 viagt 0
<< end >>
