magic
tech sky130A
magscale 1 2
timestamp 1712539494
<< pwell >>
rect -515 -10403 515 10403
<< mvnmos >>
rect -287 6945 -187 10145
rect -129 6945 -29 10145
rect 29 6945 129 10145
rect 187 6945 287 10145
rect -287 3527 -187 6727
rect -129 3527 -29 6727
rect 29 3527 129 6727
rect 187 3527 287 6727
rect -287 109 -187 3309
rect -129 109 -29 3309
rect 29 109 129 3309
rect 187 109 287 3309
rect -287 -3309 -187 -109
rect -129 -3309 -29 -109
rect 29 -3309 129 -109
rect 187 -3309 287 -109
rect -287 -6727 -187 -3527
rect -129 -6727 -29 -3527
rect 29 -6727 129 -3527
rect 187 -6727 287 -3527
rect -287 -10145 -187 -6945
rect -129 -10145 -29 -6945
rect 29 -10145 129 -6945
rect 187 -10145 287 -6945
<< mvndiff >>
rect -345 10133 -287 10145
rect -345 6957 -333 10133
rect -299 6957 -287 10133
rect -345 6945 -287 6957
rect -187 10133 -129 10145
rect -187 6957 -175 10133
rect -141 6957 -129 10133
rect -187 6945 -129 6957
rect -29 10133 29 10145
rect -29 6957 -17 10133
rect 17 6957 29 10133
rect -29 6945 29 6957
rect 129 10133 187 10145
rect 129 6957 141 10133
rect 175 6957 187 10133
rect 129 6945 187 6957
rect 287 10133 345 10145
rect 287 6957 299 10133
rect 333 6957 345 10133
rect 287 6945 345 6957
rect -345 6715 -287 6727
rect -345 3539 -333 6715
rect -299 3539 -287 6715
rect -345 3527 -287 3539
rect -187 6715 -129 6727
rect -187 3539 -175 6715
rect -141 3539 -129 6715
rect -187 3527 -129 3539
rect -29 6715 29 6727
rect -29 3539 -17 6715
rect 17 3539 29 6715
rect -29 3527 29 3539
rect 129 6715 187 6727
rect 129 3539 141 6715
rect 175 3539 187 6715
rect 129 3527 187 3539
rect 287 6715 345 6727
rect 287 3539 299 6715
rect 333 3539 345 6715
rect 287 3527 345 3539
rect -345 3297 -287 3309
rect -345 121 -333 3297
rect -299 121 -287 3297
rect -345 109 -287 121
rect -187 3297 -129 3309
rect -187 121 -175 3297
rect -141 121 -129 3297
rect -187 109 -129 121
rect -29 3297 29 3309
rect -29 121 -17 3297
rect 17 121 29 3297
rect -29 109 29 121
rect 129 3297 187 3309
rect 129 121 141 3297
rect 175 121 187 3297
rect 129 109 187 121
rect 287 3297 345 3309
rect 287 121 299 3297
rect 333 121 345 3297
rect 287 109 345 121
rect -345 -121 -287 -109
rect -345 -3297 -333 -121
rect -299 -3297 -287 -121
rect -345 -3309 -287 -3297
rect -187 -121 -129 -109
rect -187 -3297 -175 -121
rect -141 -3297 -129 -121
rect -187 -3309 -129 -3297
rect -29 -121 29 -109
rect -29 -3297 -17 -121
rect 17 -3297 29 -121
rect -29 -3309 29 -3297
rect 129 -121 187 -109
rect 129 -3297 141 -121
rect 175 -3297 187 -121
rect 129 -3309 187 -3297
rect 287 -121 345 -109
rect 287 -3297 299 -121
rect 333 -3297 345 -121
rect 287 -3309 345 -3297
rect -345 -3539 -287 -3527
rect -345 -6715 -333 -3539
rect -299 -6715 -287 -3539
rect -345 -6727 -287 -6715
rect -187 -3539 -129 -3527
rect -187 -6715 -175 -3539
rect -141 -6715 -129 -3539
rect -187 -6727 -129 -6715
rect -29 -3539 29 -3527
rect -29 -6715 -17 -3539
rect 17 -6715 29 -3539
rect -29 -6727 29 -6715
rect 129 -3539 187 -3527
rect 129 -6715 141 -3539
rect 175 -6715 187 -3539
rect 129 -6727 187 -6715
rect 287 -3539 345 -3527
rect 287 -6715 299 -3539
rect 333 -6715 345 -3539
rect 287 -6727 345 -6715
rect -345 -6957 -287 -6945
rect -345 -10133 -333 -6957
rect -299 -10133 -287 -6957
rect -345 -10145 -287 -10133
rect -187 -6957 -129 -6945
rect -187 -10133 -175 -6957
rect -141 -10133 -129 -6957
rect -187 -10145 -129 -10133
rect -29 -6957 29 -6945
rect -29 -10133 -17 -6957
rect 17 -10133 29 -6957
rect -29 -10145 29 -10133
rect 129 -6957 187 -6945
rect 129 -10133 141 -6957
rect 175 -10133 187 -6957
rect 129 -10145 187 -10133
rect 287 -6957 345 -6945
rect 287 -10133 299 -6957
rect 333 -10133 345 -6957
rect 287 -10145 345 -10133
<< mvndiffc >>
rect -333 6957 -299 10133
rect -175 6957 -141 10133
rect -17 6957 17 10133
rect 141 6957 175 10133
rect 299 6957 333 10133
rect -333 3539 -299 6715
rect -175 3539 -141 6715
rect -17 3539 17 6715
rect 141 3539 175 6715
rect 299 3539 333 6715
rect -333 121 -299 3297
rect -175 121 -141 3297
rect -17 121 17 3297
rect 141 121 175 3297
rect 299 121 333 3297
rect -333 -3297 -299 -121
rect -175 -3297 -141 -121
rect -17 -3297 17 -121
rect 141 -3297 175 -121
rect 299 -3297 333 -121
rect -333 -6715 -299 -3539
rect -175 -6715 -141 -3539
rect -17 -6715 17 -3539
rect 141 -6715 175 -3539
rect 299 -6715 333 -3539
rect -333 -10133 -299 -6957
rect -175 -10133 -141 -6957
rect -17 -10133 17 -6957
rect 141 -10133 175 -6957
rect 299 -10133 333 -6957
<< mvpsubdiff >>
rect -479 10355 479 10367
rect -479 10321 -371 10355
rect 371 10321 479 10355
rect -479 10309 479 10321
rect -479 10259 -421 10309
rect -479 -10259 -467 10259
rect -433 -10259 -421 10259
rect 421 10259 479 10309
rect -479 -10309 -421 -10259
rect 421 -10259 433 10259
rect 467 -10259 479 10259
rect 421 -10309 479 -10259
rect -479 -10321 479 -10309
rect -479 -10355 -371 -10321
rect 371 -10355 479 -10321
rect -479 -10367 479 -10355
<< mvpsubdiffcont >>
rect -371 10321 371 10355
rect -467 -10259 -433 10259
rect 433 -10259 467 10259
rect -371 -10355 371 -10321
<< poly >>
rect -287 10217 -187 10233
rect -287 10183 -271 10217
rect -203 10183 -187 10217
rect -287 10145 -187 10183
rect -129 10217 -29 10233
rect -129 10183 -113 10217
rect -45 10183 -29 10217
rect -129 10145 -29 10183
rect 29 10217 129 10233
rect 29 10183 45 10217
rect 113 10183 129 10217
rect 29 10145 129 10183
rect 187 10217 287 10233
rect 187 10183 203 10217
rect 271 10183 287 10217
rect 187 10145 287 10183
rect -287 6907 -187 6945
rect -287 6873 -271 6907
rect -203 6873 -187 6907
rect -287 6857 -187 6873
rect -129 6907 -29 6945
rect -129 6873 -113 6907
rect -45 6873 -29 6907
rect -129 6857 -29 6873
rect 29 6907 129 6945
rect 29 6873 45 6907
rect 113 6873 129 6907
rect 29 6857 129 6873
rect 187 6907 287 6945
rect 187 6873 203 6907
rect 271 6873 287 6907
rect 187 6857 287 6873
rect -287 6799 -187 6815
rect -287 6765 -271 6799
rect -203 6765 -187 6799
rect -287 6727 -187 6765
rect -129 6799 -29 6815
rect -129 6765 -113 6799
rect -45 6765 -29 6799
rect -129 6727 -29 6765
rect 29 6799 129 6815
rect 29 6765 45 6799
rect 113 6765 129 6799
rect 29 6727 129 6765
rect 187 6799 287 6815
rect 187 6765 203 6799
rect 271 6765 287 6799
rect 187 6727 287 6765
rect -287 3489 -187 3527
rect -287 3455 -271 3489
rect -203 3455 -187 3489
rect -287 3439 -187 3455
rect -129 3489 -29 3527
rect -129 3455 -113 3489
rect -45 3455 -29 3489
rect -129 3439 -29 3455
rect 29 3489 129 3527
rect 29 3455 45 3489
rect 113 3455 129 3489
rect 29 3439 129 3455
rect 187 3489 287 3527
rect 187 3455 203 3489
rect 271 3455 287 3489
rect 187 3439 287 3455
rect -287 3381 -187 3397
rect -287 3347 -271 3381
rect -203 3347 -187 3381
rect -287 3309 -187 3347
rect -129 3381 -29 3397
rect -129 3347 -113 3381
rect -45 3347 -29 3381
rect -129 3309 -29 3347
rect 29 3381 129 3397
rect 29 3347 45 3381
rect 113 3347 129 3381
rect 29 3309 129 3347
rect 187 3381 287 3397
rect 187 3347 203 3381
rect 271 3347 287 3381
rect 187 3309 287 3347
rect -287 71 -187 109
rect -287 37 -271 71
rect -203 37 -187 71
rect -287 21 -187 37
rect -129 71 -29 109
rect -129 37 -113 71
rect -45 37 -29 71
rect -129 21 -29 37
rect 29 71 129 109
rect 29 37 45 71
rect 113 37 129 71
rect 29 21 129 37
rect 187 71 287 109
rect 187 37 203 71
rect 271 37 287 71
rect 187 21 287 37
rect -287 -37 -187 -21
rect -287 -71 -271 -37
rect -203 -71 -187 -37
rect -287 -109 -187 -71
rect -129 -37 -29 -21
rect -129 -71 -113 -37
rect -45 -71 -29 -37
rect -129 -109 -29 -71
rect 29 -37 129 -21
rect 29 -71 45 -37
rect 113 -71 129 -37
rect 29 -109 129 -71
rect 187 -37 287 -21
rect 187 -71 203 -37
rect 271 -71 287 -37
rect 187 -109 287 -71
rect -287 -3347 -187 -3309
rect -287 -3381 -271 -3347
rect -203 -3381 -187 -3347
rect -287 -3397 -187 -3381
rect -129 -3347 -29 -3309
rect -129 -3381 -113 -3347
rect -45 -3381 -29 -3347
rect -129 -3397 -29 -3381
rect 29 -3347 129 -3309
rect 29 -3381 45 -3347
rect 113 -3381 129 -3347
rect 29 -3397 129 -3381
rect 187 -3347 287 -3309
rect 187 -3381 203 -3347
rect 271 -3381 287 -3347
rect 187 -3397 287 -3381
rect -287 -3455 -187 -3439
rect -287 -3489 -271 -3455
rect -203 -3489 -187 -3455
rect -287 -3527 -187 -3489
rect -129 -3455 -29 -3439
rect -129 -3489 -113 -3455
rect -45 -3489 -29 -3455
rect -129 -3527 -29 -3489
rect 29 -3455 129 -3439
rect 29 -3489 45 -3455
rect 113 -3489 129 -3455
rect 29 -3527 129 -3489
rect 187 -3455 287 -3439
rect 187 -3489 203 -3455
rect 271 -3489 287 -3455
rect 187 -3527 287 -3489
rect -287 -6765 -187 -6727
rect -287 -6799 -271 -6765
rect -203 -6799 -187 -6765
rect -287 -6815 -187 -6799
rect -129 -6765 -29 -6727
rect -129 -6799 -113 -6765
rect -45 -6799 -29 -6765
rect -129 -6815 -29 -6799
rect 29 -6765 129 -6727
rect 29 -6799 45 -6765
rect 113 -6799 129 -6765
rect 29 -6815 129 -6799
rect 187 -6765 287 -6727
rect 187 -6799 203 -6765
rect 271 -6799 287 -6765
rect 187 -6815 287 -6799
rect -287 -6873 -187 -6857
rect -287 -6907 -271 -6873
rect -203 -6907 -187 -6873
rect -287 -6945 -187 -6907
rect -129 -6873 -29 -6857
rect -129 -6907 -113 -6873
rect -45 -6907 -29 -6873
rect -129 -6945 -29 -6907
rect 29 -6873 129 -6857
rect 29 -6907 45 -6873
rect 113 -6907 129 -6873
rect 29 -6945 129 -6907
rect 187 -6873 287 -6857
rect 187 -6907 203 -6873
rect 271 -6907 287 -6873
rect 187 -6945 287 -6907
rect -287 -10183 -187 -10145
rect -287 -10217 -271 -10183
rect -203 -10217 -187 -10183
rect -287 -10233 -187 -10217
rect -129 -10183 -29 -10145
rect -129 -10217 -113 -10183
rect -45 -10217 -29 -10183
rect -129 -10233 -29 -10217
rect 29 -10183 129 -10145
rect 29 -10217 45 -10183
rect 113 -10217 129 -10183
rect 29 -10233 129 -10217
rect 187 -10183 287 -10145
rect 187 -10217 203 -10183
rect 271 -10217 287 -10183
rect 187 -10233 287 -10217
<< polycont >>
rect -271 10183 -203 10217
rect -113 10183 -45 10217
rect 45 10183 113 10217
rect 203 10183 271 10217
rect -271 6873 -203 6907
rect -113 6873 -45 6907
rect 45 6873 113 6907
rect 203 6873 271 6907
rect -271 6765 -203 6799
rect -113 6765 -45 6799
rect 45 6765 113 6799
rect 203 6765 271 6799
rect -271 3455 -203 3489
rect -113 3455 -45 3489
rect 45 3455 113 3489
rect 203 3455 271 3489
rect -271 3347 -203 3381
rect -113 3347 -45 3381
rect 45 3347 113 3381
rect 203 3347 271 3381
rect -271 37 -203 71
rect -113 37 -45 71
rect 45 37 113 71
rect 203 37 271 71
rect -271 -71 -203 -37
rect -113 -71 -45 -37
rect 45 -71 113 -37
rect 203 -71 271 -37
rect -271 -3381 -203 -3347
rect -113 -3381 -45 -3347
rect 45 -3381 113 -3347
rect 203 -3381 271 -3347
rect -271 -3489 -203 -3455
rect -113 -3489 -45 -3455
rect 45 -3489 113 -3455
rect 203 -3489 271 -3455
rect -271 -6799 -203 -6765
rect -113 -6799 -45 -6765
rect 45 -6799 113 -6765
rect 203 -6799 271 -6765
rect -271 -6907 -203 -6873
rect -113 -6907 -45 -6873
rect 45 -6907 113 -6873
rect 203 -6907 271 -6873
rect -271 -10217 -203 -10183
rect -113 -10217 -45 -10183
rect 45 -10217 113 -10183
rect 203 -10217 271 -10183
<< locali >>
rect -467 10321 -371 10355
rect 371 10321 467 10355
rect -467 10259 -433 10321
rect 433 10259 467 10321
rect -287 10183 -271 10217
rect -203 10183 -187 10217
rect -129 10183 -113 10217
rect -45 10183 -29 10217
rect 29 10183 45 10217
rect 113 10183 129 10217
rect 187 10183 203 10217
rect 271 10183 287 10217
rect -333 10133 -299 10149
rect -333 6941 -299 6957
rect -175 10133 -141 10149
rect -175 6941 -141 6957
rect -17 10133 17 10149
rect -17 6941 17 6957
rect 141 10133 175 10149
rect 141 6941 175 6957
rect 299 10133 333 10149
rect 299 6941 333 6957
rect -287 6873 -271 6907
rect -203 6873 -187 6907
rect -129 6873 -113 6907
rect -45 6873 -29 6907
rect 29 6873 45 6907
rect 113 6873 129 6907
rect 187 6873 203 6907
rect 271 6873 287 6907
rect -287 6765 -271 6799
rect -203 6765 -187 6799
rect -129 6765 -113 6799
rect -45 6765 -29 6799
rect 29 6765 45 6799
rect 113 6765 129 6799
rect 187 6765 203 6799
rect 271 6765 287 6799
rect -333 6715 -299 6731
rect -333 3523 -299 3539
rect -175 6715 -141 6731
rect -175 3523 -141 3539
rect -17 6715 17 6731
rect -17 3523 17 3539
rect 141 6715 175 6731
rect 141 3523 175 3539
rect 299 6715 333 6731
rect 299 3523 333 3539
rect -287 3455 -271 3489
rect -203 3455 -187 3489
rect -129 3455 -113 3489
rect -45 3455 -29 3489
rect 29 3455 45 3489
rect 113 3455 129 3489
rect 187 3455 203 3489
rect 271 3455 287 3489
rect -287 3347 -271 3381
rect -203 3347 -187 3381
rect -129 3347 -113 3381
rect -45 3347 -29 3381
rect 29 3347 45 3381
rect 113 3347 129 3381
rect 187 3347 203 3381
rect 271 3347 287 3381
rect -333 3297 -299 3313
rect -333 105 -299 121
rect -175 3297 -141 3313
rect -175 105 -141 121
rect -17 3297 17 3313
rect -17 105 17 121
rect 141 3297 175 3313
rect 141 105 175 121
rect 299 3297 333 3313
rect 299 105 333 121
rect -287 37 -271 71
rect -203 37 -187 71
rect -129 37 -113 71
rect -45 37 -29 71
rect 29 37 45 71
rect 113 37 129 71
rect 187 37 203 71
rect 271 37 287 71
rect -287 -71 -271 -37
rect -203 -71 -187 -37
rect -129 -71 -113 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 113 -71 129 -37
rect 187 -71 203 -37
rect 271 -71 287 -37
rect -333 -121 -299 -105
rect -333 -3313 -299 -3297
rect -175 -121 -141 -105
rect -175 -3313 -141 -3297
rect -17 -121 17 -105
rect -17 -3313 17 -3297
rect 141 -121 175 -105
rect 141 -3313 175 -3297
rect 299 -121 333 -105
rect 299 -3313 333 -3297
rect -287 -3381 -271 -3347
rect -203 -3381 -187 -3347
rect -129 -3381 -113 -3347
rect -45 -3381 -29 -3347
rect 29 -3381 45 -3347
rect 113 -3381 129 -3347
rect 187 -3381 203 -3347
rect 271 -3381 287 -3347
rect -287 -3489 -271 -3455
rect -203 -3489 -187 -3455
rect -129 -3489 -113 -3455
rect -45 -3489 -29 -3455
rect 29 -3489 45 -3455
rect 113 -3489 129 -3455
rect 187 -3489 203 -3455
rect 271 -3489 287 -3455
rect -333 -3539 -299 -3523
rect -333 -6731 -299 -6715
rect -175 -3539 -141 -3523
rect -175 -6731 -141 -6715
rect -17 -3539 17 -3523
rect -17 -6731 17 -6715
rect 141 -3539 175 -3523
rect 141 -6731 175 -6715
rect 299 -3539 333 -3523
rect 299 -6731 333 -6715
rect -287 -6799 -271 -6765
rect -203 -6799 -187 -6765
rect -129 -6799 -113 -6765
rect -45 -6799 -29 -6765
rect 29 -6799 45 -6765
rect 113 -6799 129 -6765
rect 187 -6799 203 -6765
rect 271 -6799 287 -6765
rect -287 -6907 -271 -6873
rect -203 -6907 -187 -6873
rect -129 -6907 -113 -6873
rect -45 -6907 -29 -6873
rect 29 -6907 45 -6873
rect 113 -6907 129 -6873
rect 187 -6907 203 -6873
rect 271 -6907 287 -6873
rect -333 -6957 -299 -6941
rect -333 -10149 -299 -10133
rect -175 -6957 -141 -6941
rect -175 -10149 -141 -10133
rect -17 -6957 17 -6941
rect -17 -10149 17 -10133
rect 141 -6957 175 -6941
rect 141 -10149 175 -10133
rect 299 -6957 333 -6941
rect 299 -10149 333 -10133
rect -287 -10217 -271 -10183
rect -203 -10217 -187 -10183
rect -129 -10217 -113 -10183
rect -45 -10217 -29 -10183
rect 29 -10217 45 -10183
rect 113 -10217 129 -10183
rect 187 -10217 203 -10183
rect 271 -10217 287 -10183
rect -467 -10321 -433 -10259
rect 433 -10321 467 -10259
rect -467 -10355 -371 -10321
rect 371 -10355 467 -10321
<< viali >>
rect -271 10183 -203 10217
rect -113 10183 -45 10217
rect 45 10183 113 10217
rect 203 10183 271 10217
rect -333 6957 -299 10133
rect -175 6957 -141 10133
rect -17 6957 17 10133
rect 141 6957 175 10133
rect 299 6957 333 10133
rect -271 6873 -203 6907
rect -113 6873 -45 6907
rect 45 6873 113 6907
rect 203 6873 271 6907
rect -271 6765 -203 6799
rect -113 6765 -45 6799
rect 45 6765 113 6799
rect 203 6765 271 6799
rect -333 3539 -299 6715
rect -175 3539 -141 6715
rect -17 3539 17 6715
rect 141 3539 175 6715
rect 299 3539 333 6715
rect -271 3455 -203 3489
rect -113 3455 -45 3489
rect 45 3455 113 3489
rect 203 3455 271 3489
rect -271 3347 -203 3381
rect -113 3347 -45 3381
rect 45 3347 113 3381
rect 203 3347 271 3381
rect -333 121 -299 3297
rect -175 121 -141 3297
rect -17 121 17 3297
rect 141 121 175 3297
rect 299 121 333 3297
rect -271 37 -203 71
rect -113 37 -45 71
rect 45 37 113 71
rect 203 37 271 71
rect -271 -71 -203 -37
rect -113 -71 -45 -37
rect 45 -71 113 -37
rect 203 -71 271 -37
rect -333 -3297 -299 -121
rect -175 -3297 -141 -121
rect -17 -3297 17 -121
rect 141 -3297 175 -121
rect 299 -3297 333 -121
rect -271 -3381 -203 -3347
rect -113 -3381 -45 -3347
rect 45 -3381 113 -3347
rect 203 -3381 271 -3347
rect -271 -3489 -203 -3455
rect -113 -3489 -45 -3455
rect 45 -3489 113 -3455
rect 203 -3489 271 -3455
rect -333 -6715 -299 -3539
rect -175 -6715 -141 -3539
rect -17 -6715 17 -3539
rect 141 -6715 175 -3539
rect 299 -6715 333 -3539
rect -271 -6799 -203 -6765
rect -113 -6799 -45 -6765
rect 45 -6799 113 -6765
rect 203 -6799 271 -6765
rect -271 -6907 -203 -6873
rect -113 -6907 -45 -6873
rect 45 -6907 113 -6873
rect 203 -6907 271 -6873
rect -333 -10133 -299 -6957
rect -175 -10133 -141 -6957
rect -17 -10133 17 -6957
rect 141 -10133 175 -6957
rect 299 -10133 333 -6957
rect -271 -10217 -203 -10183
rect -113 -10217 -45 -10183
rect 45 -10217 113 -10183
rect 203 -10217 271 -10183
<< metal1 >>
rect -283 10217 -191 10223
rect -283 10183 -271 10217
rect -203 10183 -191 10217
rect -283 10177 -191 10183
rect -125 10217 -33 10223
rect -125 10183 -113 10217
rect -45 10183 -33 10217
rect -125 10177 -33 10183
rect 33 10217 125 10223
rect 33 10183 45 10217
rect 113 10183 125 10217
rect 33 10177 125 10183
rect 191 10217 283 10223
rect 191 10183 203 10217
rect 271 10183 283 10217
rect 191 10177 283 10183
rect -339 10133 -293 10145
rect -339 6957 -333 10133
rect -299 6957 -293 10133
rect -339 6945 -293 6957
rect -181 10133 -135 10145
rect -181 6957 -175 10133
rect -141 6957 -135 10133
rect -181 6945 -135 6957
rect -23 10133 23 10145
rect -23 6957 -17 10133
rect 17 6957 23 10133
rect -23 6945 23 6957
rect 135 10133 181 10145
rect 135 6957 141 10133
rect 175 6957 181 10133
rect 135 6945 181 6957
rect 293 10133 339 10145
rect 293 6957 299 10133
rect 333 6957 339 10133
rect 293 6945 339 6957
rect -283 6907 -191 6913
rect -283 6873 -271 6907
rect -203 6873 -191 6907
rect -283 6867 -191 6873
rect -125 6907 -33 6913
rect -125 6873 -113 6907
rect -45 6873 -33 6907
rect -125 6867 -33 6873
rect 33 6907 125 6913
rect 33 6873 45 6907
rect 113 6873 125 6907
rect 33 6867 125 6873
rect 191 6907 283 6913
rect 191 6873 203 6907
rect 271 6873 283 6907
rect 191 6867 283 6873
rect -283 6799 -191 6805
rect -283 6765 -271 6799
rect -203 6765 -191 6799
rect -283 6759 -191 6765
rect -125 6799 -33 6805
rect -125 6765 -113 6799
rect -45 6765 -33 6799
rect -125 6759 -33 6765
rect 33 6799 125 6805
rect 33 6765 45 6799
rect 113 6765 125 6799
rect 33 6759 125 6765
rect 191 6799 283 6805
rect 191 6765 203 6799
rect 271 6765 283 6799
rect 191 6759 283 6765
rect -339 6715 -293 6727
rect -339 3539 -333 6715
rect -299 3539 -293 6715
rect -339 3527 -293 3539
rect -181 6715 -135 6727
rect -181 3539 -175 6715
rect -141 3539 -135 6715
rect -181 3527 -135 3539
rect -23 6715 23 6727
rect -23 3539 -17 6715
rect 17 3539 23 6715
rect -23 3527 23 3539
rect 135 6715 181 6727
rect 135 3539 141 6715
rect 175 3539 181 6715
rect 135 3527 181 3539
rect 293 6715 339 6727
rect 293 3539 299 6715
rect 333 3539 339 6715
rect 293 3527 339 3539
rect -283 3489 -191 3495
rect -283 3455 -271 3489
rect -203 3455 -191 3489
rect -283 3449 -191 3455
rect -125 3489 -33 3495
rect -125 3455 -113 3489
rect -45 3455 -33 3489
rect -125 3449 -33 3455
rect 33 3489 125 3495
rect 33 3455 45 3489
rect 113 3455 125 3489
rect 33 3449 125 3455
rect 191 3489 283 3495
rect 191 3455 203 3489
rect 271 3455 283 3489
rect 191 3449 283 3455
rect -283 3381 -191 3387
rect -283 3347 -271 3381
rect -203 3347 -191 3381
rect -283 3341 -191 3347
rect -125 3381 -33 3387
rect -125 3347 -113 3381
rect -45 3347 -33 3381
rect -125 3341 -33 3347
rect 33 3381 125 3387
rect 33 3347 45 3381
rect 113 3347 125 3381
rect 33 3341 125 3347
rect 191 3381 283 3387
rect 191 3347 203 3381
rect 271 3347 283 3381
rect 191 3341 283 3347
rect -339 3297 -293 3309
rect -339 121 -333 3297
rect -299 121 -293 3297
rect -339 109 -293 121
rect -181 3297 -135 3309
rect -181 121 -175 3297
rect -141 121 -135 3297
rect -181 109 -135 121
rect -23 3297 23 3309
rect -23 121 -17 3297
rect 17 121 23 3297
rect -23 109 23 121
rect 135 3297 181 3309
rect 135 121 141 3297
rect 175 121 181 3297
rect 135 109 181 121
rect 293 3297 339 3309
rect 293 121 299 3297
rect 333 121 339 3297
rect 293 109 339 121
rect -283 71 -191 77
rect -283 37 -271 71
rect -203 37 -191 71
rect -283 31 -191 37
rect -125 71 -33 77
rect -125 37 -113 71
rect -45 37 -33 71
rect -125 31 -33 37
rect 33 71 125 77
rect 33 37 45 71
rect 113 37 125 71
rect 33 31 125 37
rect 191 71 283 77
rect 191 37 203 71
rect 271 37 283 71
rect 191 31 283 37
rect -283 -37 -191 -31
rect -283 -71 -271 -37
rect -203 -71 -191 -37
rect -283 -77 -191 -71
rect -125 -37 -33 -31
rect -125 -71 -113 -37
rect -45 -71 -33 -37
rect -125 -77 -33 -71
rect 33 -37 125 -31
rect 33 -71 45 -37
rect 113 -71 125 -37
rect 33 -77 125 -71
rect 191 -37 283 -31
rect 191 -71 203 -37
rect 271 -71 283 -37
rect 191 -77 283 -71
rect -339 -121 -293 -109
rect -339 -3297 -333 -121
rect -299 -3297 -293 -121
rect -339 -3309 -293 -3297
rect -181 -121 -135 -109
rect -181 -3297 -175 -121
rect -141 -3297 -135 -121
rect -181 -3309 -135 -3297
rect -23 -121 23 -109
rect -23 -3297 -17 -121
rect 17 -3297 23 -121
rect -23 -3309 23 -3297
rect 135 -121 181 -109
rect 135 -3297 141 -121
rect 175 -3297 181 -121
rect 135 -3309 181 -3297
rect 293 -121 339 -109
rect 293 -3297 299 -121
rect 333 -3297 339 -121
rect 293 -3309 339 -3297
rect -283 -3347 -191 -3341
rect -283 -3381 -271 -3347
rect -203 -3381 -191 -3347
rect -283 -3387 -191 -3381
rect -125 -3347 -33 -3341
rect -125 -3381 -113 -3347
rect -45 -3381 -33 -3347
rect -125 -3387 -33 -3381
rect 33 -3347 125 -3341
rect 33 -3381 45 -3347
rect 113 -3381 125 -3347
rect 33 -3387 125 -3381
rect 191 -3347 283 -3341
rect 191 -3381 203 -3347
rect 271 -3381 283 -3347
rect 191 -3387 283 -3381
rect -283 -3455 -191 -3449
rect -283 -3489 -271 -3455
rect -203 -3489 -191 -3455
rect -283 -3495 -191 -3489
rect -125 -3455 -33 -3449
rect -125 -3489 -113 -3455
rect -45 -3489 -33 -3455
rect -125 -3495 -33 -3489
rect 33 -3455 125 -3449
rect 33 -3489 45 -3455
rect 113 -3489 125 -3455
rect 33 -3495 125 -3489
rect 191 -3455 283 -3449
rect 191 -3489 203 -3455
rect 271 -3489 283 -3455
rect 191 -3495 283 -3489
rect -339 -3539 -293 -3527
rect -339 -6715 -333 -3539
rect -299 -6715 -293 -3539
rect -339 -6727 -293 -6715
rect -181 -3539 -135 -3527
rect -181 -6715 -175 -3539
rect -141 -6715 -135 -3539
rect -181 -6727 -135 -6715
rect -23 -3539 23 -3527
rect -23 -6715 -17 -3539
rect 17 -6715 23 -3539
rect -23 -6727 23 -6715
rect 135 -3539 181 -3527
rect 135 -6715 141 -3539
rect 175 -6715 181 -3539
rect 135 -6727 181 -6715
rect 293 -3539 339 -3527
rect 293 -6715 299 -3539
rect 333 -6715 339 -3539
rect 293 -6727 339 -6715
rect -283 -6765 -191 -6759
rect -283 -6799 -271 -6765
rect -203 -6799 -191 -6765
rect -283 -6805 -191 -6799
rect -125 -6765 -33 -6759
rect -125 -6799 -113 -6765
rect -45 -6799 -33 -6765
rect -125 -6805 -33 -6799
rect 33 -6765 125 -6759
rect 33 -6799 45 -6765
rect 113 -6799 125 -6765
rect 33 -6805 125 -6799
rect 191 -6765 283 -6759
rect 191 -6799 203 -6765
rect 271 -6799 283 -6765
rect 191 -6805 283 -6799
rect -283 -6873 -191 -6867
rect -283 -6907 -271 -6873
rect -203 -6907 -191 -6873
rect -283 -6913 -191 -6907
rect -125 -6873 -33 -6867
rect -125 -6907 -113 -6873
rect -45 -6907 -33 -6873
rect -125 -6913 -33 -6907
rect 33 -6873 125 -6867
rect 33 -6907 45 -6873
rect 113 -6907 125 -6873
rect 33 -6913 125 -6907
rect 191 -6873 283 -6867
rect 191 -6907 203 -6873
rect 271 -6907 283 -6873
rect 191 -6913 283 -6907
rect -339 -6957 -293 -6945
rect -339 -10133 -333 -6957
rect -299 -10133 -293 -6957
rect -339 -10145 -293 -10133
rect -181 -6957 -135 -6945
rect -181 -10133 -175 -6957
rect -141 -10133 -135 -6957
rect -181 -10145 -135 -10133
rect -23 -6957 23 -6945
rect -23 -10133 -17 -6957
rect 17 -10133 23 -6957
rect -23 -10145 23 -10133
rect 135 -6957 181 -6945
rect 135 -10133 141 -6957
rect 175 -10133 181 -6957
rect 135 -10145 181 -10133
rect 293 -6957 339 -6945
rect 293 -10133 299 -6957
rect 333 -10133 339 -6957
rect 293 -10145 339 -10133
rect -283 -10183 -191 -10177
rect -283 -10217 -271 -10183
rect -203 -10217 -191 -10183
rect -283 -10223 -191 -10217
rect -125 -10183 -33 -10177
rect -125 -10217 -113 -10183
rect -45 -10217 -33 -10183
rect -125 -10223 -33 -10217
rect 33 -10183 125 -10177
rect 33 -10217 45 -10183
rect 113 -10217 125 -10183
rect 33 -10223 125 -10217
rect 191 -10183 283 -10177
rect 191 -10217 203 -10183
rect 271 -10217 283 -10183
rect 191 -10223 283 -10217
<< properties >>
string FIXED_BBOX -450 -10338 450 10338
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 16 l 0.5 m 6 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
