magic
tech sky130A
magscale 1 2
timestamp 1713232929
<< pwell >>
rect -278 -1385 278 1385
<< mvnmos >>
rect -50 727 50 1127
rect -50 109 50 509
rect -50 -509 50 -109
rect -50 -1127 50 -727
<< mvndiff >>
rect -108 1115 -50 1127
rect -108 739 -96 1115
rect -62 739 -50 1115
rect -108 727 -50 739
rect 50 1115 108 1127
rect 50 739 62 1115
rect 96 739 108 1115
rect 50 727 108 739
rect -108 497 -50 509
rect -108 121 -96 497
rect -62 121 -50 497
rect -108 109 -50 121
rect 50 497 108 509
rect 50 121 62 497
rect 96 121 108 497
rect 50 109 108 121
rect -108 -121 -50 -109
rect -108 -497 -96 -121
rect -62 -497 -50 -121
rect -108 -509 -50 -497
rect 50 -121 108 -109
rect 50 -497 62 -121
rect 96 -497 108 -121
rect 50 -509 108 -497
rect -108 -739 -50 -727
rect -108 -1115 -96 -739
rect -62 -1115 -50 -739
rect -108 -1127 -50 -1115
rect 50 -739 108 -727
rect 50 -1115 62 -739
rect 96 -1115 108 -739
rect 50 -1127 108 -1115
<< mvndiffc >>
rect -96 739 -62 1115
rect 62 739 96 1115
rect -96 121 -62 497
rect 62 121 96 497
rect -96 -497 -62 -121
rect 62 -497 96 -121
rect -96 -1115 -62 -739
rect 62 -1115 96 -739
<< mvpsubdiff >>
rect -242 1337 242 1349
rect -242 1303 -134 1337
rect 134 1303 242 1337
rect -242 1291 242 1303
rect -242 1241 -184 1291
rect -242 -1241 -230 1241
rect -196 -1241 -184 1241
rect 184 1241 242 1291
rect -242 -1291 -184 -1241
rect 184 -1241 196 1241
rect 230 -1241 242 1241
rect 184 -1291 242 -1241
rect -242 -1303 242 -1291
rect -242 -1337 -134 -1303
rect 134 -1337 242 -1303
rect -242 -1349 242 -1337
<< mvpsubdiffcont >>
rect -134 1303 134 1337
rect -230 -1241 -196 1241
rect 196 -1241 230 1241
rect -134 -1337 134 -1303
<< poly >>
rect -50 1199 50 1215
rect -50 1165 -34 1199
rect 34 1165 50 1199
rect -50 1127 50 1165
rect -50 689 50 727
rect -50 655 -34 689
rect 34 655 50 689
rect -50 639 50 655
rect -50 581 50 597
rect -50 547 -34 581
rect 34 547 50 581
rect -50 509 50 547
rect -50 71 50 109
rect -50 37 -34 71
rect 34 37 50 71
rect -50 21 50 37
rect -50 -37 50 -21
rect -50 -71 -34 -37
rect 34 -71 50 -37
rect -50 -109 50 -71
rect -50 -547 50 -509
rect -50 -581 -34 -547
rect 34 -581 50 -547
rect -50 -597 50 -581
rect -50 -655 50 -639
rect -50 -689 -34 -655
rect 34 -689 50 -655
rect -50 -727 50 -689
rect -50 -1165 50 -1127
rect -50 -1199 -34 -1165
rect 34 -1199 50 -1165
rect -50 -1215 50 -1199
<< polycont >>
rect -34 1165 34 1199
rect -34 655 34 689
rect -34 547 34 581
rect -34 37 34 71
rect -34 -71 34 -37
rect -34 -581 34 -547
rect -34 -689 34 -655
rect -34 -1199 34 -1165
<< locali >>
rect -230 1303 -134 1337
rect 134 1303 230 1337
rect -230 1241 -196 1303
rect 196 1241 230 1303
rect -50 1165 -34 1199
rect 34 1165 50 1199
rect -96 1115 -62 1131
rect -96 723 -62 739
rect 62 1115 96 1131
rect 62 723 96 739
rect -50 655 -34 689
rect 34 655 50 689
rect -50 547 -34 581
rect 34 547 50 581
rect -96 497 -62 513
rect -96 105 -62 121
rect 62 497 96 513
rect 62 105 96 121
rect -50 37 -34 71
rect 34 37 50 71
rect -50 -71 -34 -37
rect 34 -71 50 -37
rect -96 -121 -62 -105
rect -96 -513 -62 -497
rect 62 -121 96 -105
rect 62 -513 96 -497
rect -50 -581 -34 -547
rect 34 -581 50 -547
rect -50 -689 -34 -655
rect 34 -689 50 -655
rect -96 -739 -62 -723
rect -96 -1131 -62 -1115
rect 62 -739 96 -723
rect 62 -1131 96 -1115
rect -50 -1199 -34 -1165
rect 34 -1199 50 -1165
rect -230 -1303 -196 -1241
rect 196 -1303 230 -1241
rect -230 -1337 -134 -1303
rect 134 -1337 230 -1303
<< viali >>
rect -34 1165 34 1199
rect -96 739 -62 1115
rect 62 739 96 1115
rect -34 655 34 689
rect -34 547 34 581
rect -96 121 -62 497
rect 62 121 96 497
rect -34 37 34 71
rect -34 -71 34 -37
rect -96 -497 -62 -121
rect 62 -497 96 -121
rect -34 -581 34 -547
rect -34 -689 34 -655
rect -96 -1115 -62 -739
rect 62 -1115 96 -739
rect -34 -1199 34 -1165
<< metal1 >>
rect -46 1199 46 1205
rect -46 1165 -34 1199
rect 34 1165 46 1199
rect -46 1159 46 1165
rect -102 1115 -56 1127
rect -102 739 -96 1115
rect -62 739 -56 1115
rect -102 727 -56 739
rect 56 1115 102 1127
rect 56 739 62 1115
rect 96 739 102 1115
rect 56 727 102 739
rect -46 689 46 695
rect -46 655 -34 689
rect 34 655 46 689
rect -46 649 46 655
rect -46 581 46 587
rect -46 547 -34 581
rect 34 547 46 581
rect -46 541 46 547
rect -102 497 -56 509
rect -102 121 -96 497
rect -62 121 -56 497
rect -102 109 -56 121
rect 56 497 102 509
rect 56 121 62 497
rect 96 121 102 497
rect 56 109 102 121
rect -46 71 46 77
rect -46 37 -34 71
rect 34 37 46 71
rect -46 31 46 37
rect -46 -37 46 -31
rect -46 -71 -34 -37
rect 34 -71 46 -37
rect -46 -77 46 -71
rect -102 -121 -56 -109
rect -102 -497 -96 -121
rect -62 -497 -56 -121
rect -102 -509 -56 -497
rect 56 -121 102 -109
rect 56 -497 62 -121
rect 96 -497 102 -121
rect 56 -509 102 -497
rect -46 -547 46 -541
rect -46 -581 -34 -547
rect 34 -581 46 -547
rect -46 -587 46 -581
rect -46 -655 46 -649
rect -46 -689 -34 -655
rect 34 -689 46 -655
rect -46 -695 46 -689
rect -102 -739 -56 -727
rect -102 -1115 -96 -739
rect -62 -1115 -56 -739
rect -102 -1127 -56 -1115
rect 56 -739 102 -727
rect 56 -1115 62 -739
rect 96 -1115 102 -739
rect 56 -1127 102 -1115
rect -46 -1165 46 -1159
rect -46 -1199 -34 -1165
rect 34 -1199 46 -1165
rect -46 -1205 46 -1199
<< properties >>
string FIXED_BBOX -213 -1320 213 1320
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 2 l 0.50 m 4 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
