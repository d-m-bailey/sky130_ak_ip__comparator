magic
tech sky130A
magscale 1 2
timestamp 1713585847
<< error_p >>
rect -582 272 -524 278
rect -424 272 -366 278
rect -266 272 -208 278
rect -108 272 -50 278
rect 50 272 108 278
rect 208 272 266 278
rect 366 272 424 278
rect 524 272 582 278
rect -582 238 -570 272
rect -424 238 -412 272
rect -266 238 -254 272
rect -108 238 -96 272
rect 50 238 62 272
rect 208 238 220 272
rect 366 238 378 272
rect 524 238 536 272
rect -582 232 -524 238
rect -424 232 -366 238
rect -266 232 -208 238
rect -108 232 -50 238
rect 50 232 108 238
rect 208 232 266 238
rect 366 232 424 238
rect 524 232 582 238
rect -582 -238 -524 -232
rect -424 -238 -366 -232
rect -266 -238 -208 -232
rect -108 -238 -50 -232
rect 50 -238 108 -232
rect 208 -238 266 -232
rect 366 -238 424 -232
rect 524 -238 582 -232
rect -582 -272 -570 -238
rect -424 -272 -412 -238
rect -266 -272 -254 -238
rect -108 -272 -96 -238
rect 50 -272 62 -238
rect 208 -272 220 -238
rect 366 -272 378 -238
rect 524 -272 536 -238
rect -582 -278 -524 -272
rect -424 -278 -366 -272
rect -266 -278 -208 -272
rect -108 -278 -50 -272
rect 50 -278 108 -272
rect 208 -278 266 -272
rect 366 -278 424 -272
rect 524 -278 582 -272
<< pwell >>
rect -831 -458 831 458
<< mvnmos >>
rect -603 -200 -503 200
rect -445 -200 -345 200
rect -287 -200 -187 200
rect -129 -200 -29 200
rect 29 -200 129 200
rect 187 -200 287 200
rect 345 -200 445 200
rect 503 -200 603 200
<< mvndiff >>
rect -661 188 -603 200
rect -661 -188 -649 188
rect -615 -188 -603 188
rect -661 -200 -603 -188
rect -503 188 -445 200
rect -503 -188 -491 188
rect -457 -188 -445 188
rect -503 -200 -445 -188
rect -345 188 -287 200
rect -345 -188 -333 188
rect -299 -188 -287 188
rect -345 -200 -287 -188
rect -187 188 -129 200
rect -187 -188 -175 188
rect -141 -188 -129 188
rect -187 -200 -129 -188
rect -29 188 29 200
rect -29 -188 -17 188
rect 17 -188 29 188
rect -29 -200 29 -188
rect 129 188 187 200
rect 129 -188 141 188
rect 175 -188 187 188
rect 129 -200 187 -188
rect 287 188 345 200
rect 287 -188 299 188
rect 333 -188 345 188
rect 287 -200 345 -188
rect 445 188 503 200
rect 445 -188 457 188
rect 491 -188 503 188
rect 445 -200 503 -188
rect 603 188 661 200
rect 603 -188 615 188
rect 649 -188 661 188
rect 603 -200 661 -188
<< mvndiffc >>
rect -649 -188 -615 188
rect -491 -188 -457 188
rect -333 -188 -299 188
rect -175 -188 -141 188
rect -17 -188 17 188
rect 141 -188 175 188
rect 299 -188 333 188
rect 457 -188 491 188
rect 615 -188 649 188
<< mvpsubdiff >>
rect -795 410 795 422
rect -795 376 -687 410
rect 687 376 795 410
rect -795 364 795 376
rect -795 314 -737 364
rect -795 -314 -783 314
rect -749 -314 -737 314
rect 737 314 795 364
rect -795 -364 -737 -314
rect 737 -314 749 314
rect 783 -314 795 314
rect 737 -364 795 -314
rect -795 -376 795 -364
rect -795 -410 -687 -376
rect 687 -410 795 -376
rect -795 -422 795 -410
<< mvpsubdiffcont >>
rect -687 376 687 410
rect -783 -314 -749 314
rect 749 -314 783 314
rect -687 -410 687 -376
<< poly >>
rect -603 272 -503 288
rect -603 238 -587 272
rect -519 238 -503 272
rect -603 200 -503 238
rect -445 272 -345 288
rect -445 238 -429 272
rect -361 238 -345 272
rect -445 200 -345 238
rect -287 272 -187 288
rect -287 238 -271 272
rect -203 238 -187 272
rect -287 200 -187 238
rect -129 272 -29 288
rect -129 238 -113 272
rect -45 238 -29 272
rect -129 200 -29 238
rect 29 272 129 288
rect 29 238 45 272
rect 113 238 129 272
rect 29 200 129 238
rect 187 272 287 288
rect 187 238 203 272
rect 271 238 287 272
rect 187 200 287 238
rect 345 272 445 288
rect 345 238 361 272
rect 429 238 445 272
rect 345 200 445 238
rect 503 272 603 288
rect 503 238 519 272
rect 587 238 603 272
rect 503 200 603 238
rect -603 -238 -503 -200
rect -603 -272 -587 -238
rect -519 -272 -503 -238
rect -603 -288 -503 -272
rect -445 -238 -345 -200
rect -445 -272 -429 -238
rect -361 -272 -345 -238
rect -445 -288 -345 -272
rect -287 -238 -187 -200
rect -287 -272 -271 -238
rect -203 -272 -187 -238
rect -287 -288 -187 -272
rect -129 -238 -29 -200
rect -129 -272 -113 -238
rect -45 -272 -29 -238
rect -129 -288 -29 -272
rect 29 -238 129 -200
rect 29 -272 45 -238
rect 113 -272 129 -238
rect 29 -288 129 -272
rect 187 -238 287 -200
rect 187 -272 203 -238
rect 271 -272 287 -238
rect 187 -288 287 -272
rect 345 -238 445 -200
rect 345 -272 361 -238
rect 429 -272 445 -238
rect 345 -288 445 -272
rect 503 -238 603 -200
rect 503 -272 519 -238
rect 587 -272 603 -238
rect 503 -288 603 -272
<< polycont >>
rect -587 238 -519 272
rect -429 238 -361 272
rect -271 238 -203 272
rect -113 238 -45 272
rect 45 238 113 272
rect 203 238 271 272
rect 361 238 429 272
rect 519 238 587 272
rect -587 -272 -519 -238
rect -429 -272 -361 -238
rect -271 -272 -203 -238
rect -113 -272 -45 -238
rect 45 -272 113 -238
rect 203 -272 271 -238
rect 361 -272 429 -238
rect 519 -272 587 -238
<< locali >>
rect -783 376 -687 410
rect 687 376 783 410
rect -783 314 -749 376
rect 749 314 783 376
rect -603 238 -587 272
rect -519 238 -503 272
rect -445 238 -429 272
rect -361 238 -345 272
rect -287 238 -271 272
rect -203 238 -187 272
rect -129 238 -113 272
rect -45 238 -29 272
rect 29 238 45 272
rect 113 238 129 272
rect 187 238 203 272
rect 271 238 287 272
rect 345 238 361 272
rect 429 238 445 272
rect 503 238 519 272
rect 587 238 603 272
rect -649 188 -615 204
rect -649 -204 -615 -188
rect -491 188 -457 204
rect -491 -204 -457 -188
rect -333 188 -299 204
rect -333 -204 -299 -188
rect -175 188 -141 204
rect -175 -204 -141 -188
rect -17 188 17 204
rect -17 -204 17 -188
rect 141 188 175 204
rect 141 -204 175 -188
rect 299 188 333 204
rect 299 -204 333 -188
rect 457 188 491 204
rect 457 -204 491 -188
rect 615 188 649 204
rect 615 -204 649 -188
rect -603 -272 -587 -238
rect -519 -272 -503 -238
rect -445 -272 -429 -238
rect -361 -272 -345 -238
rect -287 -272 -271 -238
rect -203 -272 -187 -238
rect -129 -272 -113 -238
rect -45 -272 -29 -238
rect 29 -272 45 -238
rect 113 -272 129 -238
rect 187 -272 203 -238
rect 271 -272 287 -238
rect 345 -272 361 -238
rect 429 -272 445 -238
rect 503 -272 519 -238
rect 587 -272 603 -238
rect -783 -376 -749 -314
rect 749 -376 783 -314
rect -783 -410 -687 -376
rect 687 -410 783 -376
<< viali >>
rect -599 376 599 410
rect -783 -301 -749 301
rect -570 238 -536 272
rect -412 238 -378 272
rect -254 238 -220 272
rect -96 238 -62 272
rect 62 238 96 272
rect 220 238 254 272
rect 378 238 412 272
rect 536 238 570 272
rect -649 -188 -615 188
rect -491 -188 -457 188
rect -333 -188 -299 188
rect -175 -188 -141 188
rect -17 -188 17 188
rect 141 -188 175 188
rect 299 -188 333 188
rect 457 -188 491 188
rect 615 -188 649 188
rect -570 -272 -536 -238
rect -412 -272 -378 -238
rect -254 -272 -220 -238
rect -96 -272 -62 -238
rect 62 -272 96 -238
rect 220 -272 254 -238
rect 378 -272 412 -238
rect 536 -272 570 -238
rect 749 -301 783 301
<< metal1 >>
rect -611 410 611 416
rect -611 376 -599 410
rect 599 376 611 410
rect -611 370 611 376
rect -789 301 -743 313
rect -789 -301 -783 301
rect -749 -301 -743 301
rect 743 301 789 313
rect -582 272 -524 278
rect -582 238 -570 272
rect -536 238 -524 272
rect -582 232 -524 238
rect -424 272 -366 278
rect -424 238 -412 272
rect -378 238 -366 272
rect -424 232 -366 238
rect -266 272 -208 278
rect -266 238 -254 272
rect -220 238 -208 272
rect -266 232 -208 238
rect -108 272 -50 278
rect -108 238 -96 272
rect -62 238 -50 272
rect -108 232 -50 238
rect 50 272 108 278
rect 50 238 62 272
rect 96 238 108 272
rect 50 232 108 238
rect 208 272 266 278
rect 208 238 220 272
rect 254 238 266 272
rect 208 232 266 238
rect 366 272 424 278
rect 366 238 378 272
rect 412 238 424 272
rect 366 232 424 238
rect 524 272 582 278
rect 524 238 536 272
rect 570 238 582 272
rect 524 232 582 238
rect -655 188 -609 200
rect -655 -188 -649 188
rect -615 -188 -609 188
rect -655 -200 -609 -188
rect -497 188 -451 200
rect -497 -188 -491 188
rect -457 -188 -451 188
rect -497 -200 -451 -188
rect -339 188 -293 200
rect -339 -188 -333 188
rect -299 -188 -293 188
rect -339 -200 -293 -188
rect -181 188 -135 200
rect -181 -188 -175 188
rect -141 -188 -135 188
rect -181 -200 -135 -188
rect -23 188 23 200
rect -23 -188 -17 188
rect 17 -188 23 188
rect -23 -200 23 -188
rect 135 188 181 200
rect 135 -188 141 188
rect 175 -188 181 188
rect 135 -200 181 -188
rect 293 188 339 200
rect 293 -188 299 188
rect 333 -188 339 188
rect 293 -200 339 -188
rect 451 188 497 200
rect 451 -188 457 188
rect 491 -188 497 188
rect 451 -200 497 -188
rect 609 188 655 200
rect 609 -188 615 188
rect 649 -188 655 188
rect 609 -200 655 -188
rect -582 -238 -524 -232
rect -582 -272 -570 -238
rect -536 -272 -524 -238
rect -582 -278 -524 -272
rect -424 -238 -366 -232
rect -424 -272 -412 -238
rect -378 -272 -366 -238
rect -424 -278 -366 -272
rect -266 -238 -208 -232
rect -266 -272 -254 -238
rect -220 -272 -208 -238
rect -266 -278 -208 -272
rect -108 -238 -50 -232
rect -108 -272 -96 -238
rect -62 -272 -50 -238
rect -108 -278 -50 -272
rect 50 -238 108 -232
rect 50 -272 62 -238
rect 96 -272 108 -238
rect 50 -278 108 -272
rect 208 -238 266 -232
rect 208 -272 220 -238
rect 254 -272 266 -238
rect 208 -278 266 -272
rect 366 -238 424 -232
rect 366 -272 378 -238
rect 412 -272 424 -238
rect 366 -278 424 -272
rect 524 -238 582 -232
rect 524 -272 536 -238
rect 570 -272 582 -238
rect 524 -278 582 -272
rect -789 -313 -743 -301
rect 743 -301 749 301
rect 783 -301 789 301
rect 743 -313 789 -301
<< properties >>
string FIXED_BBOX -766 -393 766 393
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 2 l 0.50 m 1 nf 8 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 80 viagl 80 viagt 80
<< end >>
