magic
tech sky130A
magscale 1 2
timestamp 1713107406
<< pwell >>
rect -2782 -3258 2782 3258
<< psubdiff >>
rect -2746 3188 -2650 3222
rect 2650 3188 2746 3222
rect -2746 3126 -2712 3188
rect 2712 3126 2746 3188
rect -2746 -3188 -2712 -3126
rect 2712 -3188 2746 -3126
rect -2746 -3222 -2650 -3188
rect 2650 -3222 2746 -3188
<< psubdiffcont >>
rect -2650 3188 2650 3222
rect -2746 -3126 -2712 3126
rect 2712 -3126 2746 3126
rect -2650 -3222 2650 -3188
<< xpolycontact >>
rect -2616 2660 -2046 3092
rect -2616 -3092 -2046 -2660
rect -1950 2660 -1380 3092
rect -1950 -3092 -1380 -2660
rect -1284 2660 -714 3092
rect -1284 -3092 -714 -2660
rect -618 2660 -48 3092
rect -618 -3092 -48 -2660
rect 48 2660 618 3092
rect 48 -3092 618 -2660
rect 714 2660 1284 3092
rect 714 -3092 1284 -2660
rect 1380 2660 1950 3092
rect 1380 -3092 1950 -2660
rect 2046 2660 2616 3092
rect 2046 -3092 2616 -2660
<< ppolyres >>
rect -2616 -2660 -2046 2660
rect -1950 -2660 -1380 2660
rect -1284 -2660 -714 2660
rect -618 -2660 -48 2660
rect 48 -2660 618 2660
rect 714 -2660 1284 2660
rect 1380 -2660 1950 2660
rect 2046 -2660 2616 2660
<< locali >>
rect -2746 3188 -2650 3222
rect 2650 3188 2746 3222
rect -2746 3126 -2712 3188
rect 2712 3126 2746 3188
rect -2746 -3188 -2712 -3126
rect 2712 -3188 2746 -3126
rect -2746 -3222 -2650 -3188
rect 2650 -3222 2746 -3188
<< viali >>
rect -2441 3188 2441 3222
rect -2746 -2869 -2712 2869
rect -2600 2677 -2062 3074
rect -1934 2677 -1396 3074
rect -1268 2677 -730 3074
rect -602 2677 -64 3074
rect 64 2677 602 3074
rect 730 2677 1268 3074
rect 1396 2677 1934 3074
rect 2062 2677 2600 3074
rect -2600 -3074 -2062 -2677
rect -1934 -3074 -1396 -2677
rect -1268 -3074 -730 -2677
rect -602 -3074 -64 -2677
rect 64 -3074 602 -2677
rect 730 -3074 1268 -2677
rect 1396 -3074 1934 -2677
rect 2062 -3074 2600 -2677
rect 2712 -2869 2746 2869
rect -2441 -3222 2441 -3188
<< metal1 >>
rect -2453 3222 2453 3228
rect -2453 3188 -2441 3222
rect 2441 3188 2453 3222
rect -2453 3182 2453 3188
rect -2612 3074 -2050 3080
rect -2752 2869 -2706 2881
rect -2752 -2869 -2746 2869
rect -2712 -2869 -2706 2869
rect -2612 2677 -2600 3074
rect -2062 2677 -2050 3074
rect -2612 2671 -2050 2677
rect -1946 3074 -1384 3080
rect -1946 2677 -1934 3074
rect -1396 2677 -1384 3074
rect -1946 2671 -1384 2677
rect -1280 3074 -718 3080
rect -1280 2677 -1268 3074
rect -730 2677 -718 3074
rect -1280 2671 -718 2677
rect -614 3074 -52 3080
rect -614 2677 -602 3074
rect -64 2677 -52 3074
rect -614 2671 -52 2677
rect 52 3074 614 3080
rect 52 2677 64 3074
rect 602 2677 614 3074
rect 52 2671 614 2677
rect 718 3074 1280 3080
rect 718 2677 730 3074
rect 1268 2677 1280 3074
rect 718 2671 1280 2677
rect 1384 3074 1946 3080
rect 1384 2677 1396 3074
rect 1934 2677 1946 3074
rect 1384 2671 1946 2677
rect 2050 3074 2612 3080
rect 2050 2677 2062 3074
rect 2600 2677 2612 3074
rect 2050 2671 2612 2677
rect 2706 2869 2752 2881
rect -2752 -2881 -2706 -2869
rect -2612 -2677 -2050 -2671
rect -2612 -3074 -2600 -2677
rect -2062 -3074 -2050 -2677
rect -2612 -3080 -2050 -3074
rect -1946 -2677 -1384 -2671
rect -1946 -3074 -1934 -2677
rect -1396 -3074 -1384 -2677
rect -1946 -3080 -1384 -3074
rect -1280 -2677 -718 -2671
rect -1280 -3074 -1268 -2677
rect -730 -3074 -718 -2677
rect -1280 -3080 -718 -3074
rect -614 -2677 -52 -2671
rect -614 -3074 -602 -2677
rect -64 -3074 -52 -2677
rect -614 -3080 -52 -3074
rect 52 -2677 614 -2671
rect 52 -3074 64 -2677
rect 602 -3074 614 -2677
rect 52 -3080 614 -3074
rect 718 -2677 1280 -2671
rect 718 -3074 730 -2677
rect 1268 -3074 1280 -2677
rect 718 -3080 1280 -3074
rect 1384 -2677 1946 -2671
rect 1384 -3074 1396 -2677
rect 1934 -3074 1946 -2677
rect 1384 -3080 1946 -3074
rect 2050 -2677 2612 -2671
rect 2050 -3074 2062 -2677
rect 2600 -3074 2612 -2677
rect 2706 -2869 2712 2869
rect 2746 -2869 2752 2869
rect 2706 -2881 2752 -2869
rect 2050 -3080 2612 -3074
rect -2453 -3188 2453 -3182
rect -2453 -3222 -2441 -3188
rect 2441 -3222 2453 -3188
rect -2453 -3228 2453 -3222
<< res2p85 >>
rect -2618 -2662 -2044 2662
rect -1952 -2662 -1378 2662
rect -1286 -2662 -712 2662
rect -620 -2662 -46 2662
rect 46 -2662 620 2662
rect 712 -2662 1286 2662
rect 1378 -2662 1952 2662
rect 2044 -2662 2618 2662
<< properties >>
string FIXED_BBOX -2729 -3205 2729 3205
string gencell sky130_fd_pr__res_high_po_2p85
string library sky130
string parameters w 2.85 l 26.6 m 1 nx 8 wmin 2.850 lmin 0.50 rho 319.8 val 3.121k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 2.850 n_guard 0 hv_guard 0 vias 1 viagb 90 viagt 90 viagl 90 viagr 90
<< end >>
