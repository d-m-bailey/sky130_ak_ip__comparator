magic
tech sky130A
magscale 1 2
timestamp 1713548572
<< error_p >>
rect -32 281 32 287
rect -32 247 -20 281
rect -32 241 32 247
rect -32 -247 32 -241
rect -32 -281 -20 -247
rect -32 -287 32 -281
<< nwell >>
rect -308 -497 308 497
<< mvpmos >>
rect -50 -200 50 200
<< mvpdiff >>
rect -108 188 -50 200
rect -108 -188 -96 188
rect -62 -188 -50 188
rect -108 -200 -50 -188
rect 50 188 108 200
rect 50 -188 62 188
rect 96 -188 108 188
rect 50 -200 108 -188
<< mvpdiffc >>
rect -96 -188 -62 188
rect 62 -188 96 188
<< mvnsubdiff >>
rect -242 419 242 431
rect -242 385 -134 419
rect 134 385 242 419
rect -242 373 242 385
rect -242 -373 -184 373
rect 184 -373 242 373
rect -242 -385 242 -373
rect -242 -419 -134 -385
rect 134 -419 242 -385
rect -242 -431 242 -419
<< mvnsubdiffcont >>
rect -134 385 134 419
rect -134 -419 134 -385
<< poly >>
rect -50 281 50 297
rect -50 247 -34 281
rect 34 247 50 281
rect -50 200 50 247
rect -50 -247 50 -200
rect -50 -281 -34 -247
rect 34 -281 50 -247
rect -50 -297 50 -281
<< polycont >>
rect -34 247 34 281
rect -34 -281 34 -247
<< locali >>
rect -230 -385 -196 419
rect -50 247 -34 281
rect 34 247 50 281
rect -96 188 -62 204
rect -96 -204 -62 -188
rect 62 188 96 204
rect 62 -204 96 -188
rect -50 -281 -34 -247
rect 34 -281 50 -247
rect 196 -385 230 419
rect -230 -419 -134 -385
rect 134 -419 230 -385
<< viali >>
rect -196 385 -134 419
rect -134 385 134 419
rect 134 385 196 419
rect -20 247 20 281
rect -96 -188 -62 188
rect 62 -188 96 188
rect -20 -281 20 -247
<< metal1 >>
rect -208 419 208 425
rect -208 385 -196 419
rect 196 385 208 419
rect -208 379 208 385
rect -32 281 32 287
rect -32 247 -20 281
rect 20 247 32 281
rect -32 241 32 247
rect -102 188 -56 200
rect -102 -188 -96 188
rect -62 -188 -56 188
rect -102 -200 -56 -188
rect 56 188 102 200
rect 56 -188 62 188
rect 96 -188 102 188
rect 56 -200 102 -188
rect -32 -247 32 -241
rect -32 -281 -20 -247
rect 20 -281 32 -247
rect -32 -287 32 -281
<< properties >>
string FIXED_BBOX -213 -402 213 402
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 2 l 0.50 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 0 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 60 viagb 0 viagr 0 viagl 0 viagt 100
<< end >>
