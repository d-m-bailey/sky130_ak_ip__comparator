magic
tech sky130A
timestamp 1712377380
<< pwell >>
rect -214 -529 214 529
<< mvnmos >>
rect -100 -400 100 400
<< mvndiff >>
rect -129 394 -100 400
rect -129 -394 -123 394
rect -106 -394 -100 394
rect -129 -400 -100 -394
rect 100 394 129 400
rect 100 -394 106 394
rect 123 -394 129 394
rect 100 -400 129 -394
<< mvndiffc >>
rect -123 -394 -106 394
rect 106 -394 123 394
<< mvpsubdiff >>
rect -196 505 196 511
rect -196 488 -142 505
rect 142 488 196 505
rect -196 482 196 488
rect -196 457 -167 482
rect -196 -457 -190 457
rect -173 -457 -167 457
rect 167 457 196 482
rect -196 -482 -167 -457
rect 167 -457 173 457
rect 190 -457 196 457
rect 167 -482 196 -457
rect -196 -488 196 -482
rect -196 -505 -142 -488
rect 142 -505 196 -488
rect -196 -511 196 -505
<< mvpsubdiffcont >>
rect -142 488 142 505
rect -190 -457 -173 457
rect 173 -457 190 457
rect -142 -505 142 -488
<< poly >>
rect -100 436 100 444
rect -100 419 -92 436
rect 92 419 100 436
rect -100 400 100 419
rect -100 -419 100 -400
rect -100 -436 -92 -419
rect 92 -436 100 -419
rect -100 -444 100 -436
<< polycont >>
rect -92 419 92 436
rect -92 -436 92 -419
<< locali >>
rect -190 488 -142 505
rect 142 488 190 505
rect -190 457 -173 488
rect 173 457 190 488
rect -100 419 -92 436
rect 92 419 100 436
rect -123 394 -106 402
rect -123 -402 -106 -394
rect 106 394 123 402
rect 106 -402 123 -394
rect -100 -436 -92 -419
rect 92 -436 100 -419
rect -190 -488 -173 -457
rect 173 -488 190 -457
rect -190 -505 -142 -488
rect 142 -505 190 -488
<< viali >>
rect -92 419 92 436
rect -123 -394 -106 394
rect 106 -394 123 394
rect -92 -436 92 -419
<< metal1 >>
rect -98 436 98 439
rect -98 419 -92 436
rect 92 419 98 436
rect -98 416 98 419
rect -126 394 -103 400
rect -126 -394 -123 394
rect -106 -394 -103 394
rect -126 -400 -103 -394
rect 103 394 126 400
rect 103 -394 106 394
rect 123 -394 126 394
rect 103 -400 126 -394
rect -98 -419 98 -416
rect -98 -436 -92 -419
rect 92 -436 98 -419
rect -98 -439 98 -436
<< properties >>
string FIXED_BBOX -181 -496 181 496
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 8 l 2 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
