magic
tech sky130A
magscale 1 2
timestamp 1714698820
<< dnwell >>
rect 210 236 1028 1868
<< nwell >>
rect 290 -1560 360 -1060
rect 870 -1560 940 -1060
rect 290 -1650 940 -1560
<< locali >>
rect 390 1660 750 1696
rect 390 1550 450 1660
rect 626 1592 750 1660
rect 390 1442 478 1550
rect 760 1440 850 1540
rect 490 1330 590 1398
rect 790 1330 850 1440
rect 490 1300 850 1330
rect 490 1294 848 1300
rect 392 -1512 476 -1268
rect 760 -1512 844 -1268
rect 392 -1552 844 -1512
<< metal1 >>
rect 290 1700 950 1790
rect 290 1320 370 1700
rect 520 1390 550 1620
rect 600 1470 630 1700
rect 680 1390 710 1620
rect 500 1120 570 1390
rect 410 1050 570 1120
rect 660 1120 730 1390
rect 870 1320 950 1700
rect 660 1050 820 1120
rect 290 410 350 890
rect 410 860 490 1050
rect 740 860 820 1050
rect 410 680 470 860
rect 410 550 460 680
rect 520 520 560 830
rect 380 510 570 520
rect 380 450 390 510
rect 560 450 570 510
rect 380 440 570 450
rect 600 410 630 600
rect 680 520 720 830
rect 760 740 820 860
rect 770 550 820 740
rect 660 510 850 520
rect 660 450 670 510
rect 840 450 850 510
rect 660 440 850 450
rect 880 410 940 890
rect 290 308 940 410
rect 290 -480 940 -382
rect 290 -820 350 -480
rect 530 -580 710 -480
rect 750 -520 840 -510
rect 750 -630 760 -520
rect 450 -670 760 -630
rect 530 -730 590 -710
rect 400 -740 710 -730
rect 400 -1010 410 -740
rect 480 -790 720 -740
rect 750 -790 760 -670
rect 830 -790 840 -520
rect 480 -1010 490 -790
rect 750 -800 840 -790
rect 400 -1020 490 -1010
rect 290 -1560 360 -1060
rect 420 -1470 470 -1020
rect 760 -1170 810 -800
rect 880 -820 940 -480
rect 500 -1230 810 -1170
rect 600 -1390 630 -1290
rect 590 -1560 650 -1390
rect 870 -1560 940 -1060
rect 290 -1650 940 -1560
<< via1 >>
rect 390 450 560 510
rect 670 450 840 510
rect 410 -1010 480 -740
rect 760 -790 830 -520
<< metal2 >>
rect 380 510 570 520
rect 380 450 390 510
rect 560 450 570 510
rect 380 440 570 450
rect 660 510 850 520
rect 660 450 670 510
rect 840 450 850 510
rect 660 440 850 450
rect 400 -740 490 440
rect 400 -1010 410 -740
rect 480 -1010 490 -740
rect 750 -520 840 440
rect 750 -790 760 -520
rect 830 -790 840 -520
rect 750 -800 840 -790
rect 400 -1020 490 -1010
use sky130_fd_pr__nfet_g5v0d10v5_C5EREZ  sky130_fd_pr__nfet_g5v0d10v5_C5EREZ_0
timestamp 1713585847
transform 0 1 618 -1 0 -648
box -278 -358 278 358
use sky130_fd_pr__nfet_g5v0d10v5_S48KL6  sky130_fd_pr__nfet_g5v0d10v5_S48KL6_0
timestamp 1713585847
transform 1 0 617 0 1 658
box -357 -358 357 358
use sky130_fd_pr__pfet_g5v0d10v5_4V4BDM  sky130_fd_pr__pfet_g5v0d10v5_4V4BDM_0
timestamp 1713594760
transform 1 0 619 0 1 1495
box -387 -347 387 347
use sky130_fd_pr__pfet_g5v0d10v5_8T5BGA  sky130_fd_pr__pfet_g5v0d10v5_8T5BGA_0
timestamp 1713585847
transform 1 0 617 0 1 -1338
box -387 -362 387 362
<< labels >>
flabel via1 760 -600 830 -530 0 FreeSans 320 0 0 0 x_lv
port 2 nsew
flabel metal1 860 -1640 930 -1570 0 FreeSans 320 0 0 0 VDD_LV
port 5 nsew
flabel metal1 870 1710 940 1780 0 FreeSans 320 0 0 0 VDD_HV
port 0 nsew
flabel metal1 576 -466 646 -396 0 FreeSans 320 0 0 0 GND_LV
port 6 nsew
flabel metal1 740 1050 810 1120 0 FreeSans 320 0 0 0 xb_hv
port 4 nsew
flabel metal1 420 1050 490 1120 0 FreeSans 320 0 0 0 x_hv
port 3 nsew
flabel metal1 580 330 650 400 0 FreeSans 320 0 0 0 GND_HV
port 1 nsew
<< end >>
