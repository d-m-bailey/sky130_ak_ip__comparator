magic
tech sky130A
magscale 1 2
timestamp 1713548572
<< nwell >>
rect -425 -619 425 619
<< pmos >>
rect -229 -400 -29 400
rect 29 -400 229 400
<< pdiff >>
rect -287 388 -229 400
rect -287 -388 -275 388
rect -241 -388 -229 388
rect -287 -400 -229 -388
rect -29 388 29 400
rect -29 -388 -17 388
rect 17 -388 29 388
rect -29 -400 29 -388
rect 229 388 287 400
rect 229 -388 241 388
rect 275 -388 287 388
rect 229 -400 287 -388
<< pdiffc >>
rect -275 -388 -241 388
rect -17 -388 17 388
rect 241 -388 275 388
<< nsubdiff >>
rect -389 549 -293 583
rect 293 549 389 583
rect -389 487 -355 549
rect 355 487 389 549
rect -389 -549 -355 -487
rect 355 -549 389 -487
rect -389 -583 -293 -549
rect 293 -583 389 -549
<< nsubdiffcont >>
rect -293 549 293 583
rect -389 -487 -355 487
rect 355 -487 389 487
rect -293 -583 293 -549
<< poly >>
rect -229 481 -29 497
rect -229 447 -213 481
rect -45 447 -29 481
rect -229 400 -29 447
rect 29 481 229 497
rect 29 447 45 481
rect 213 447 229 481
rect 29 400 229 447
rect -229 -447 -29 -400
rect -229 -481 -213 -447
rect -45 -481 -29 -447
rect -229 -497 -29 -481
rect 29 -447 229 -400
rect 29 -481 45 -447
rect 213 -481 229 -447
rect 29 -497 229 -481
<< polycont >>
rect -213 447 -45 481
rect 45 447 213 481
rect -213 -481 -45 -447
rect 45 -481 213 -447
<< locali >>
rect -389 487 -355 583
rect 355 487 389 583
rect -229 447 -213 481
rect -45 447 -29 481
rect 29 447 45 481
rect 213 447 229 481
rect -275 388 -241 404
rect -275 -404 -241 -388
rect -17 388 17 404
rect -17 -404 17 -388
rect 241 388 275 404
rect 241 -404 275 -388
rect -229 -481 -213 -447
rect -45 -481 -29 -447
rect 29 -481 45 -447
rect 213 -481 229 -447
rect -389 -549 -355 -487
rect 355 -549 389 -487
rect -389 -583 -293 -549
rect 293 -583 389 -549
<< viali >>
rect -355 549 -293 583
rect -293 549 293 583
rect 293 549 355 583
rect -179 447 -79 481
rect 79 447 179 481
rect -275 -388 -241 388
rect -17 -388 17 388
rect 241 -388 275 388
rect -179 -481 -79 -447
rect 79 -481 179 -447
<< metal1 >>
rect -367 583 367 589
rect -367 549 -355 583
rect 355 549 367 583
rect -367 543 367 549
rect -191 481 -67 487
rect -191 447 -179 481
rect -79 447 -67 481
rect -191 441 -67 447
rect 67 481 191 487
rect 67 447 79 481
rect 179 447 191 481
rect 67 441 191 447
rect -281 388 -235 400
rect -281 -388 -275 388
rect -241 -388 -235 388
rect -281 -400 -235 -388
rect -23 388 23 400
rect -23 -388 -17 388
rect 17 -388 23 388
rect -23 -400 23 -388
rect 235 388 281 400
rect 235 -388 241 388
rect 275 -388 281 388
rect 235 -400 281 -388
rect -191 -447 -67 -441
rect -191 -481 -179 -447
rect -79 -481 -67 -447
rect -191 -487 -67 -481
rect 67 -447 191 -441
rect 67 -481 79 -447
rect 179 -481 191 -447
rect 67 -487 191 -481
<< properties >>
string FIXED_BBOX -372 -566 372 566
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 4 l 1 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 60 viagb 0 viagr 0 viagl 0 viagt 100
<< end >>
