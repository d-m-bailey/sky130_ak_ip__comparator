magic
tech sky130A
magscale 1 2
timestamp 1712377380
<< nwell >>
rect -1058 -697 1058 697
<< mvpmos >>
rect -800 -400 800 400
<< mvpdiff >>
rect -858 388 -800 400
rect -858 -388 -846 388
rect -812 -388 -800 388
rect -858 -400 -800 -388
rect 800 388 858 400
rect 800 -388 812 388
rect 846 -388 858 388
rect 800 -400 858 -388
<< mvpdiffc >>
rect -846 -388 -812 388
rect 812 -388 846 388
<< mvnsubdiff >>
rect -992 619 992 631
rect -992 585 -884 619
rect 884 585 992 619
rect -992 573 992 585
rect -992 523 -934 573
rect -992 -523 -980 523
rect -946 -523 -934 523
rect 934 523 992 573
rect -992 -573 -934 -523
rect 934 -523 946 523
rect 980 -523 992 523
rect 934 -573 992 -523
rect -992 -585 992 -573
rect -992 -619 -884 -585
rect 884 -619 992 -585
rect -992 -631 992 -619
<< mvnsubdiffcont >>
rect -884 585 884 619
rect -980 -523 -946 523
rect 946 -523 980 523
rect -884 -619 884 -585
<< poly >>
rect -800 481 800 497
rect -800 447 -784 481
rect 784 447 800 481
rect -800 400 800 447
rect -800 -447 800 -400
rect -800 -481 -784 -447
rect 784 -481 800 -447
rect -800 -497 800 -481
<< polycont >>
rect -784 447 784 481
rect -784 -481 784 -447
<< locali >>
rect -980 585 -884 619
rect 884 585 980 619
rect -980 523 -946 585
rect 946 523 980 585
rect -800 447 -784 481
rect 784 447 800 481
rect -846 388 -812 404
rect -846 -404 -812 -388
rect 812 388 846 404
rect 812 -404 846 -388
rect -800 -481 -784 -447
rect 784 -481 800 -447
rect -980 -585 -946 -523
rect 946 -585 980 -523
rect -980 -619 -884 -585
rect 884 -619 980 -585
<< viali >>
rect -784 447 784 481
rect -846 -388 -812 388
rect 812 -388 846 388
rect -784 -481 784 -447
<< metal1 >>
rect -796 481 796 487
rect -796 447 -784 481
rect 784 447 796 481
rect -796 441 796 447
rect -852 388 -806 400
rect -852 -388 -846 388
rect -812 -388 -806 388
rect -852 -400 -806 -388
rect 806 388 852 400
rect 806 -388 812 388
rect 846 -388 852 388
rect 806 -400 852 -388
rect -796 -447 796 -441
rect -796 -481 -784 -447
rect 784 -481 796 -447
rect -796 -487 796 -481
<< properties >>
string FIXED_BBOX -963 -602 963 602
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 4 l 8 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
