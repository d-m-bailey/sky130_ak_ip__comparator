magic
tech sky130A
magscale 1 2
timestamp 1713548572
<< error_p >>
rect -1214 281 -1156 287
rect -1056 281 -998 287
rect -898 281 -840 287
rect -740 281 -682 287
rect -582 281 -524 287
rect -424 281 -366 287
rect -266 281 -208 287
rect -108 281 -50 287
rect 50 281 108 287
rect 208 281 266 287
rect 366 281 424 287
rect 524 281 582 287
rect 682 281 740 287
rect 840 281 898 287
rect 998 281 1056 287
rect 1156 281 1214 287
rect -1214 247 -1202 281
rect -1056 247 -1044 281
rect -898 247 -886 281
rect -740 247 -728 281
rect -582 247 -570 281
rect -424 247 -412 281
rect -266 247 -254 281
rect -108 247 -96 281
rect 50 247 62 281
rect 208 247 220 281
rect 366 247 378 281
rect 524 247 536 281
rect 682 247 694 281
rect 840 247 852 281
rect 998 247 1010 281
rect 1156 247 1168 281
rect -1214 241 -1156 247
rect -1056 241 -998 247
rect -898 241 -840 247
rect -740 241 -682 247
rect -582 241 -524 247
rect -424 241 -366 247
rect -266 241 -208 247
rect -108 241 -50 247
rect 50 241 108 247
rect 208 241 266 247
rect 366 241 424 247
rect 524 241 582 247
rect 682 241 740 247
rect 840 241 898 247
rect 998 241 1056 247
rect 1156 241 1214 247
rect -1214 -247 -1156 -241
rect -1056 -247 -998 -241
rect -898 -247 -840 -241
rect -740 -247 -682 -241
rect -582 -247 -524 -241
rect -424 -247 -366 -241
rect -266 -247 -208 -241
rect -108 -247 -50 -241
rect 50 -247 108 -241
rect 208 -247 266 -241
rect 366 -247 424 -241
rect 524 -247 582 -241
rect 682 -247 740 -241
rect 840 -247 898 -241
rect 998 -247 1056 -241
rect 1156 -247 1214 -241
rect -1214 -281 -1202 -247
rect -1056 -281 -1044 -247
rect -898 -281 -886 -247
rect -740 -281 -728 -247
rect -582 -281 -570 -247
rect -424 -281 -412 -247
rect -266 -281 -254 -247
rect -108 -281 -96 -247
rect 50 -281 62 -247
rect 208 -281 220 -247
rect 366 -281 378 -247
rect 524 -281 536 -247
rect 682 -281 694 -247
rect 840 -281 852 -247
rect 998 -281 1010 -247
rect 1156 -281 1168 -247
rect -1214 -287 -1156 -281
rect -1056 -287 -998 -281
rect -898 -287 -840 -281
rect -740 -287 -682 -281
rect -582 -287 -524 -281
rect -424 -287 -366 -281
rect -266 -287 -208 -281
rect -108 -287 -50 -281
rect 50 -287 108 -281
rect 208 -287 266 -281
rect 366 -287 424 -281
rect 524 -287 582 -281
rect 682 -287 740 -281
rect 840 -287 898 -281
rect 998 -287 1056 -281
rect 1156 -287 1214 -281
<< nwell >>
rect -1493 -497 1493 497
<< mvpmos >>
rect -1235 -200 -1135 200
rect -1077 -200 -977 200
rect -919 -200 -819 200
rect -761 -200 -661 200
rect -603 -200 -503 200
rect -445 -200 -345 200
rect -287 -200 -187 200
rect -129 -200 -29 200
rect 29 -200 129 200
rect 187 -200 287 200
rect 345 -200 445 200
rect 503 -200 603 200
rect 661 -200 761 200
rect 819 -200 919 200
rect 977 -200 1077 200
rect 1135 -200 1235 200
<< mvpdiff >>
rect -1293 188 -1235 200
rect -1293 -188 -1281 188
rect -1247 -188 -1235 188
rect -1293 -200 -1235 -188
rect -1135 188 -1077 200
rect -1135 -188 -1123 188
rect -1089 -188 -1077 188
rect -1135 -200 -1077 -188
rect -977 188 -919 200
rect -977 -188 -965 188
rect -931 -188 -919 188
rect -977 -200 -919 -188
rect -819 188 -761 200
rect -819 -188 -807 188
rect -773 -188 -761 188
rect -819 -200 -761 -188
rect -661 188 -603 200
rect -661 -188 -649 188
rect -615 -188 -603 188
rect -661 -200 -603 -188
rect -503 188 -445 200
rect -503 -188 -491 188
rect -457 -188 -445 188
rect -503 -200 -445 -188
rect -345 188 -287 200
rect -345 -188 -333 188
rect -299 -188 -287 188
rect -345 -200 -287 -188
rect -187 188 -129 200
rect -187 -188 -175 188
rect -141 -188 -129 188
rect -187 -200 -129 -188
rect -29 188 29 200
rect -29 -188 -17 188
rect 17 -188 29 188
rect -29 -200 29 -188
rect 129 188 187 200
rect 129 -188 141 188
rect 175 -188 187 188
rect 129 -200 187 -188
rect 287 188 345 200
rect 287 -188 299 188
rect 333 -188 345 188
rect 287 -200 345 -188
rect 445 188 503 200
rect 445 -188 457 188
rect 491 -188 503 188
rect 445 -200 503 -188
rect 603 188 661 200
rect 603 -188 615 188
rect 649 -188 661 188
rect 603 -200 661 -188
rect 761 188 819 200
rect 761 -188 773 188
rect 807 -188 819 188
rect 761 -200 819 -188
rect 919 188 977 200
rect 919 -188 931 188
rect 965 -188 977 188
rect 919 -200 977 -188
rect 1077 188 1135 200
rect 1077 -188 1089 188
rect 1123 -188 1135 188
rect 1077 -200 1135 -188
rect 1235 188 1293 200
rect 1235 -188 1247 188
rect 1281 -188 1293 188
rect 1235 -200 1293 -188
<< mvpdiffc >>
rect -1281 -188 -1247 188
rect -1123 -188 -1089 188
rect -965 -188 -931 188
rect -807 -188 -773 188
rect -649 -188 -615 188
rect -491 -188 -457 188
rect -333 -188 -299 188
rect -175 -188 -141 188
rect -17 -188 17 188
rect 141 -188 175 188
rect 299 -188 333 188
rect 457 -188 491 188
rect 615 -188 649 188
rect 773 -188 807 188
rect 931 -188 965 188
rect 1089 -188 1123 188
rect 1247 -188 1281 188
<< mvnsubdiff >>
rect -1427 419 1427 431
rect -1427 385 -1319 419
rect 1319 385 1427 419
rect -1427 373 1427 385
rect -1427 323 -1369 373
rect -1427 -323 -1415 323
rect -1381 -323 -1369 323
rect 1369 323 1427 373
rect -1427 -373 -1369 -323
rect 1369 -323 1381 323
rect 1415 -323 1427 323
rect 1369 -373 1427 -323
rect -1427 -385 1427 -373
rect -1427 -419 -1319 -385
rect 1319 -419 1427 -385
rect -1427 -431 1427 -419
<< mvnsubdiffcont >>
rect -1319 385 1319 419
rect -1415 -323 -1381 323
rect 1381 -323 1415 323
rect -1319 -419 1319 -385
<< poly >>
rect -1235 281 -1135 297
rect -1235 247 -1219 281
rect -1151 247 -1135 281
rect -1235 200 -1135 247
rect -1077 281 -977 297
rect -1077 247 -1061 281
rect -993 247 -977 281
rect -1077 200 -977 247
rect -919 281 -819 297
rect -919 247 -903 281
rect -835 247 -819 281
rect -919 200 -819 247
rect -761 281 -661 297
rect -761 247 -745 281
rect -677 247 -661 281
rect -761 200 -661 247
rect -603 281 -503 297
rect -603 247 -587 281
rect -519 247 -503 281
rect -603 200 -503 247
rect -445 281 -345 297
rect -445 247 -429 281
rect -361 247 -345 281
rect -445 200 -345 247
rect -287 281 -187 297
rect -287 247 -271 281
rect -203 247 -187 281
rect -287 200 -187 247
rect -129 281 -29 297
rect -129 247 -113 281
rect -45 247 -29 281
rect -129 200 -29 247
rect 29 281 129 297
rect 29 247 45 281
rect 113 247 129 281
rect 29 200 129 247
rect 187 281 287 297
rect 187 247 203 281
rect 271 247 287 281
rect 187 200 287 247
rect 345 281 445 297
rect 345 247 361 281
rect 429 247 445 281
rect 345 200 445 247
rect 503 281 603 297
rect 503 247 519 281
rect 587 247 603 281
rect 503 200 603 247
rect 661 281 761 297
rect 661 247 677 281
rect 745 247 761 281
rect 661 200 761 247
rect 819 281 919 297
rect 819 247 835 281
rect 903 247 919 281
rect 819 200 919 247
rect 977 281 1077 297
rect 977 247 993 281
rect 1061 247 1077 281
rect 977 200 1077 247
rect 1135 281 1235 297
rect 1135 247 1151 281
rect 1219 247 1235 281
rect 1135 200 1235 247
rect -1235 -247 -1135 -200
rect -1235 -281 -1219 -247
rect -1151 -281 -1135 -247
rect -1235 -297 -1135 -281
rect -1077 -247 -977 -200
rect -1077 -281 -1061 -247
rect -993 -281 -977 -247
rect -1077 -297 -977 -281
rect -919 -247 -819 -200
rect -919 -281 -903 -247
rect -835 -281 -819 -247
rect -919 -297 -819 -281
rect -761 -247 -661 -200
rect -761 -281 -745 -247
rect -677 -281 -661 -247
rect -761 -297 -661 -281
rect -603 -247 -503 -200
rect -603 -281 -587 -247
rect -519 -281 -503 -247
rect -603 -297 -503 -281
rect -445 -247 -345 -200
rect -445 -281 -429 -247
rect -361 -281 -345 -247
rect -445 -297 -345 -281
rect -287 -247 -187 -200
rect -287 -281 -271 -247
rect -203 -281 -187 -247
rect -287 -297 -187 -281
rect -129 -247 -29 -200
rect -129 -281 -113 -247
rect -45 -281 -29 -247
rect -129 -297 -29 -281
rect 29 -247 129 -200
rect 29 -281 45 -247
rect 113 -281 129 -247
rect 29 -297 129 -281
rect 187 -247 287 -200
rect 187 -281 203 -247
rect 271 -281 287 -247
rect 187 -297 287 -281
rect 345 -247 445 -200
rect 345 -281 361 -247
rect 429 -281 445 -247
rect 345 -297 445 -281
rect 503 -247 603 -200
rect 503 -281 519 -247
rect 587 -281 603 -247
rect 503 -297 603 -281
rect 661 -247 761 -200
rect 661 -281 677 -247
rect 745 -281 761 -247
rect 661 -297 761 -281
rect 819 -247 919 -200
rect 819 -281 835 -247
rect 903 -281 919 -247
rect 819 -297 919 -281
rect 977 -247 1077 -200
rect 977 -281 993 -247
rect 1061 -281 1077 -247
rect 977 -297 1077 -281
rect 1135 -247 1235 -200
rect 1135 -281 1151 -247
rect 1219 -281 1235 -247
rect 1135 -297 1235 -281
<< polycont >>
rect -1219 247 -1151 281
rect -1061 247 -993 281
rect -903 247 -835 281
rect -745 247 -677 281
rect -587 247 -519 281
rect -429 247 -361 281
rect -271 247 -203 281
rect -113 247 -45 281
rect 45 247 113 281
rect 203 247 271 281
rect 361 247 429 281
rect 519 247 587 281
rect 677 247 745 281
rect 835 247 903 281
rect 993 247 1061 281
rect 1151 247 1219 281
rect -1219 -281 -1151 -247
rect -1061 -281 -993 -247
rect -903 -281 -835 -247
rect -745 -281 -677 -247
rect -587 -281 -519 -247
rect -429 -281 -361 -247
rect -271 -281 -203 -247
rect -113 -281 -45 -247
rect 45 -281 113 -247
rect 203 -281 271 -247
rect 361 -281 429 -247
rect 519 -281 587 -247
rect 677 -281 745 -247
rect 835 -281 903 -247
rect 993 -281 1061 -247
rect 1151 -281 1219 -247
<< locali >>
rect -1415 385 -1319 419
rect 1319 385 1415 419
rect -1415 323 -1381 385
rect 1381 323 1415 385
rect -1235 247 -1219 281
rect -1151 247 -1135 281
rect -1077 247 -1061 281
rect -993 247 -977 281
rect -919 247 -903 281
rect -835 247 -819 281
rect -761 247 -745 281
rect -677 247 -661 281
rect -603 247 -587 281
rect -519 247 -503 281
rect -445 247 -429 281
rect -361 247 -345 281
rect -287 247 -271 281
rect -203 247 -187 281
rect -129 247 -113 281
rect -45 247 -29 281
rect 29 247 45 281
rect 113 247 129 281
rect 187 247 203 281
rect 271 247 287 281
rect 345 247 361 281
rect 429 247 445 281
rect 503 247 519 281
rect 587 247 603 281
rect 661 247 677 281
rect 745 247 761 281
rect 819 247 835 281
rect 903 247 919 281
rect 977 247 993 281
rect 1061 247 1077 281
rect 1135 247 1151 281
rect 1219 247 1235 281
rect -1281 188 -1247 204
rect -1281 -204 -1247 -188
rect -1123 188 -1089 204
rect -1123 -204 -1089 -188
rect -965 188 -931 204
rect -965 -204 -931 -188
rect -807 188 -773 204
rect -807 -204 -773 -188
rect -649 188 -615 204
rect -649 -204 -615 -188
rect -491 188 -457 204
rect -491 -204 -457 -188
rect -333 188 -299 204
rect -333 -204 -299 -188
rect -175 188 -141 204
rect -175 -204 -141 -188
rect -17 188 17 204
rect -17 -204 17 -188
rect 141 188 175 204
rect 141 -204 175 -188
rect 299 188 333 204
rect 299 -204 333 -188
rect 457 188 491 204
rect 457 -204 491 -188
rect 615 188 649 204
rect 615 -204 649 -188
rect 773 188 807 204
rect 773 -204 807 -188
rect 931 188 965 204
rect 931 -204 965 -188
rect 1089 188 1123 204
rect 1089 -204 1123 -188
rect 1247 188 1281 204
rect 1247 -204 1281 -188
rect -1235 -281 -1219 -247
rect -1151 -281 -1135 -247
rect -1077 -281 -1061 -247
rect -993 -281 -977 -247
rect -919 -281 -903 -247
rect -835 -281 -819 -247
rect -761 -281 -745 -247
rect -677 -281 -661 -247
rect -603 -281 -587 -247
rect -519 -281 -503 -247
rect -445 -281 -429 -247
rect -361 -281 -345 -247
rect -287 -281 -271 -247
rect -203 -281 -187 -247
rect -129 -281 -113 -247
rect -45 -281 -29 -247
rect 29 -281 45 -247
rect 113 -281 129 -247
rect 187 -281 203 -247
rect 271 -281 287 -247
rect 345 -281 361 -247
rect 429 -281 445 -247
rect 503 -281 519 -247
rect 587 -281 603 -247
rect 661 -281 677 -247
rect 745 -281 761 -247
rect 819 -281 835 -247
rect 903 -281 919 -247
rect 977 -281 993 -247
rect 1061 -281 1077 -247
rect 1135 -281 1151 -247
rect 1219 -281 1235 -247
rect -1415 -385 -1381 -323
rect 1381 -385 1415 -323
rect -1415 -419 -1319 -385
rect 1319 -419 1415 -385
<< viali >>
rect -1415 -308 -1381 308
rect -1202 247 -1168 281
rect -1044 247 -1010 281
rect -886 247 -852 281
rect -728 247 -694 281
rect -570 247 -536 281
rect -412 247 -378 281
rect -254 247 -220 281
rect -96 247 -62 281
rect 62 247 96 281
rect 220 247 254 281
rect 378 247 412 281
rect 536 247 570 281
rect 694 247 728 281
rect 852 247 886 281
rect 1010 247 1044 281
rect 1168 247 1202 281
rect -1281 -188 -1247 188
rect -1123 -188 -1089 188
rect -965 -188 -931 188
rect -807 -188 -773 188
rect -649 -188 -615 188
rect -491 -188 -457 188
rect -333 -188 -299 188
rect -175 -188 -141 188
rect -17 -188 17 188
rect 141 -188 175 188
rect 299 -188 333 188
rect 457 -188 491 188
rect 615 -188 649 188
rect 773 -188 807 188
rect 931 -188 965 188
rect 1089 -188 1123 188
rect 1247 -188 1281 188
rect -1202 -281 -1168 -247
rect -1044 -281 -1010 -247
rect -886 -281 -852 -247
rect -728 -281 -694 -247
rect -570 -281 -536 -247
rect -412 -281 -378 -247
rect -254 -281 -220 -247
rect -96 -281 -62 -247
rect 62 -281 96 -247
rect 220 -281 254 -247
rect 378 -281 412 -247
rect 536 -281 570 -247
rect 694 -281 728 -247
rect 852 -281 886 -247
rect 1010 -281 1044 -247
rect 1168 -281 1202 -247
rect 1381 -308 1415 308
rect -1105 -419 1105 -385
<< metal1 >>
rect -1421 308 -1375 320
rect -1421 -308 -1415 308
rect -1381 -308 -1375 308
rect 1375 308 1421 320
rect -1214 281 -1156 287
rect -1214 247 -1202 281
rect -1168 247 -1156 281
rect -1214 241 -1156 247
rect -1056 281 -998 287
rect -1056 247 -1044 281
rect -1010 247 -998 281
rect -1056 241 -998 247
rect -898 281 -840 287
rect -898 247 -886 281
rect -852 247 -840 281
rect -898 241 -840 247
rect -740 281 -682 287
rect -740 247 -728 281
rect -694 247 -682 281
rect -740 241 -682 247
rect -582 281 -524 287
rect -582 247 -570 281
rect -536 247 -524 281
rect -582 241 -524 247
rect -424 281 -366 287
rect -424 247 -412 281
rect -378 247 -366 281
rect -424 241 -366 247
rect -266 281 -208 287
rect -266 247 -254 281
rect -220 247 -208 281
rect -266 241 -208 247
rect -108 281 -50 287
rect -108 247 -96 281
rect -62 247 -50 281
rect -108 241 -50 247
rect 50 281 108 287
rect 50 247 62 281
rect 96 247 108 281
rect 50 241 108 247
rect 208 281 266 287
rect 208 247 220 281
rect 254 247 266 281
rect 208 241 266 247
rect 366 281 424 287
rect 366 247 378 281
rect 412 247 424 281
rect 366 241 424 247
rect 524 281 582 287
rect 524 247 536 281
rect 570 247 582 281
rect 524 241 582 247
rect 682 281 740 287
rect 682 247 694 281
rect 728 247 740 281
rect 682 241 740 247
rect 840 281 898 287
rect 840 247 852 281
rect 886 247 898 281
rect 840 241 898 247
rect 998 281 1056 287
rect 998 247 1010 281
rect 1044 247 1056 281
rect 998 241 1056 247
rect 1156 281 1214 287
rect 1156 247 1168 281
rect 1202 247 1214 281
rect 1156 241 1214 247
rect -1287 188 -1241 200
rect -1287 -188 -1281 188
rect -1247 -188 -1241 188
rect -1287 -200 -1241 -188
rect -1129 188 -1083 200
rect -1129 -188 -1123 188
rect -1089 -188 -1083 188
rect -1129 -200 -1083 -188
rect -971 188 -925 200
rect -971 -188 -965 188
rect -931 -188 -925 188
rect -971 -200 -925 -188
rect -813 188 -767 200
rect -813 -188 -807 188
rect -773 -188 -767 188
rect -813 -200 -767 -188
rect -655 188 -609 200
rect -655 -188 -649 188
rect -615 -188 -609 188
rect -655 -200 -609 -188
rect -497 188 -451 200
rect -497 -188 -491 188
rect -457 -188 -451 188
rect -497 -200 -451 -188
rect -339 188 -293 200
rect -339 -188 -333 188
rect -299 -188 -293 188
rect -339 -200 -293 -188
rect -181 188 -135 200
rect -181 -188 -175 188
rect -141 -188 -135 188
rect -181 -200 -135 -188
rect -23 188 23 200
rect -23 -188 -17 188
rect 17 -188 23 188
rect -23 -200 23 -188
rect 135 188 181 200
rect 135 -188 141 188
rect 175 -188 181 188
rect 135 -200 181 -188
rect 293 188 339 200
rect 293 -188 299 188
rect 333 -188 339 188
rect 293 -200 339 -188
rect 451 188 497 200
rect 451 -188 457 188
rect 491 -188 497 188
rect 451 -200 497 -188
rect 609 188 655 200
rect 609 -188 615 188
rect 649 -188 655 188
rect 609 -200 655 -188
rect 767 188 813 200
rect 767 -188 773 188
rect 807 -188 813 188
rect 767 -200 813 -188
rect 925 188 971 200
rect 925 -188 931 188
rect 965 -188 971 188
rect 925 -200 971 -188
rect 1083 188 1129 200
rect 1083 -188 1089 188
rect 1123 -188 1129 188
rect 1083 -200 1129 -188
rect 1241 188 1287 200
rect 1241 -188 1247 188
rect 1281 -188 1287 188
rect 1241 -200 1287 -188
rect -1214 -247 -1156 -241
rect -1214 -281 -1202 -247
rect -1168 -281 -1156 -247
rect -1214 -287 -1156 -281
rect -1056 -247 -998 -241
rect -1056 -281 -1044 -247
rect -1010 -281 -998 -247
rect -1056 -287 -998 -281
rect -898 -247 -840 -241
rect -898 -281 -886 -247
rect -852 -281 -840 -247
rect -898 -287 -840 -281
rect -740 -247 -682 -241
rect -740 -281 -728 -247
rect -694 -281 -682 -247
rect -740 -287 -682 -281
rect -582 -247 -524 -241
rect -582 -281 -570 -247
rect -536 -281 -524 -247
rect -582 -287 -524 -281
rect -424 -247 -366 -241
rect -424 -281 -412 -247
rect -378 -281 -366 -247
rect -424 -287 -366 -281
rect -266 -247 -208 -241
rect -266 -281 -254 -247
rect -220 -281 -208 -247
rect -266 -287 -208 -281
rect -108 -247 -50 -241
rect -108 -281 -96 -247
rect -62 -281 -50 -247
rect -108 -287 -50 -281
rect 50 -247 108 -241
rect 50 -281 62 -247
rect 96 -281 108 -247
rect 50 -287 108 -281
rect 208 -247 266 -241
rect 208 -281 220 -247
rect 254 -281 266 -247
rect 208 -287 266 -281
rect 366 -247 424 -241
rect 366 -281 378 -247
rect 412 -281 424 -247
rect 366 -287 424 -281
rect 524 -247 582 -241
rect 524 -281 536 -247
rect 570 -281 582 -247
rect 524 -287 582 -281
rect 682 -247 740 -241
rect 682 -281 694 -247
rect 728 -281 740 -247
rect 682 -287 740 -281
rect 840 -247 898 -241
rect 840 -281 852 -247
rect 886 -281 898 -247
rect 840 -287 898 -281
rect 998 -247 1056 -241
rect 998 -281 1010 -247
rect 1044 -281 1056 -247
rect 998 -287 1056 -281
rect 1156 -247 1214 -241
rect 1156 -281 1168 -247
rect 1202 -281 1214 -247
rect 1156 -287 1214 -281
rect -1421 -320 -1375 -308
rect 1375 -308 1381 308
rect 1415 -308 1421 308
rect 1375 -320 1421 -308
rect -1117 -385 1117 -379
rect -1117 -419 -1105 -385
rect 1105 -419 1117 -385
rect -1117 -425 1117 -419
<< properties >>
string FIXED_BBOX -1398 -402 1398 402
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 2 l 0.5 m 1 nf 16 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 80 viagr 80 viagl 80 viagt 0
<< end >>
