magic
tech sky130A
timestamp 1712472733
<< properties >>
string gencell sky130_fd_pr__res_high_po_2p85
string library sky130
string parameters w 2.850 l 2.85*56 m 1 nx 1 wmin 2.850 lmin 0.50 rho 319.8 val 18.045k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 2.850 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
