magic
tech sky130A
magscale 1 2
timestamp 1713112495
<< error_p >>
rect -467 -516 -433 -512
rect 433 -516 467 -512
rect -467 -550 -399 -516
rect 399 -550 467 -516
rect -433 -584 -395 -550
rect 395 -584 433 -550
<< nwell >>
rect -545 -662 545 662
<< mvpmos >>
rect -287 -364 -187 436
rect -129 -364 -29 436
rect 29 -364 129 436
rect 187 -364 287 436
<< mvpdiff >>
rect -345 424 -287 436
rect -345 -352 -333 424
rect -299 -352 -287 424
rect -345 -364 -287 -352
rect -187 424 -129 436
rect -187 -352 -175 424
rect -141 -352 -129 424
rect -187 -364 -129 -352
rect -29 424 29 436
rect -29 -352 -17 424
rect 17 -352 29 424
rect -29 -364 29 -352
rect 129 424 187 436
rect 129 -352 141 424
rect 175 -352 187 424
rect 129 -364 187 -352
rect 287 424 345 436
rect 287 -352 299 424
rect 333 -352 345 424
rect 287 -364 345 -352
<< mvpdiffc >>
rect -333 -352 -299 424
rect -175 -352 -141 424
rect -17 -352 17 424
rect 141 -352 175 424
rect 299 -352 333 424
<< mvnsubdiff >>
rect -479 584 479 596
rect -479 550 -371 584
rect 371 550 479 584
rect -479 538 479 550
rect -479 488 -421 538
rect -479 -488 -467 488
rect -433 -488 -421 488
rect 421 488 479 538
rect -479 -538 -421 -488
rect 421 -488 433 488
rect 467 -488 479 488
rect 421 -538 479 -488
rect -479 -550 479 -538
rect -479 -584 -371 -550
rect 371 -584 479 -550
rect -479 -596 479 -584
<< mvnsubdiffcont >>
rect -371 550 371 584
rect -467 -488 -433 488
rect 433 -488 467 488
rect -371 -584 371 -550
<< poly >>
rect -287 436 -187 462
rect -129 436 -29 462
rect 29 436 129 462
rect 187 436 287 462
rect -287 -411 -187 -364
rect -287 -445 -271 -411
rect -203 -445 -187 -411
rect -287 -461 -187 -445
rect -129 -411 -29 -364
rect -129 -445 -113 -411
rect -45 -445 -29 -411
rect -129 -461 -29 -445
rect 29 -411 129 -364
rect 29 -445 45 -411
rect 113 -445 129 -411
rect 29 -461 129 -445
rect 187 -411 287 -364
rect 187 -445 203 -411
rect 271 -445 287 -411
rect 187 -461 287 -445
<< polycont >>
rect -271 -445 -203 -411
rect -113 -445 -45 -411
rect 45 -445 113 -411
rect 203 -445 271 -411
<< locali >>
rect -467 550 -371 584
rect 371 550 467 584
rect -333 424 -299 440
rect -333 -368 -299 -352
rect -175 424 -141 440
rect -175 -368 -141 -352
rect -17 424 17 440
rect -17 -368 17 -352
rect 141 424 175 440
rect 141 -368 175 -352
rect 299 424 333 440
rect 299 -368 333 -352
rect -287 -445 -271 -411
rect -203 -445 -187 -411
rect -129 -445 -113 -411
rect -45 -445 -29 -411
rect 29 -445 45 -411
rect 113 -445 129 -411
rect 187 -445 203 -411
rect 271 -445 287 -411
rect -467 -584 -433 -550
rect 433 -584 467 -550
<< viali >>
rect -467 488 -433 550
rect -467 -488 -433 488
rect 433 488 467 550
rect -333 -352 -299 424
rect -175 -352 -141 424
rect -17 -352 17 424
rect 141 -352 175 424
rect 299 -352 333 424
rect -264 -445 -210 -411
rect -106 -445 -52 -411
rect 52 -445 106 -411
rect 210 -445 264 -411
rect -467 -550 -433 -488
rect 433 -488 467 488
rect 433 -550 467 -488
rect -433 -584 -371 -550
rect -371 -584 371 -550
rect 371 -584 433 -550
<< metal1 >>
rect -473 550 -427 562
rect -473 -550 -467 550
rect -433 -544 -427 550
rect 427 550 473 562
rect -339 424 -293 436
rect -339 -352 -333 424
rect -299 -352 -293 424
rect -339 -364 -293 -352
rect -181 424 -135 436
rect -181 -352 -175 424
rect -141 -352 -135 424
rect -181 -364 -135 -352
rect -23 424 23 436
rect -23 -352 -17 424
rect 17 -352 23 424
rect -23 -364 23 -352
rect 135 424 181 436
rect 135 -352 141 424
rect 175 -352 181 424
rect 135 -364 181 -352
rect 293 424 339 436
rect 293 -352 299 424
rect 333 -352 339 424
rect 293 -364 339 -352
rect -276 -411 -198 -405
rect -276 -445 -264 -411
rect -210 -445 -198 -411
rect -276 -451 -198 -445
rect -118 -411 -40 -405
rect -118 -445 -106 -411
rect -52 -445 -40 -411
rect -118 -451 -40 -445
rect 40 -411 118 -405
rect 40 -445 52 -411
rect 106 -445 118 -411
rect 40 -451 118 -445
rect 198 -411 276 -405
rect 198 -445 210 -411
rect 264 -445 276 -411
rect 198 -451 276 -445
rect 427 -544 433 550
rect -433 -550 433 -544
rect 467 -550 473 550
rect -473 -562 -433 -550
rect -445 -584 -433 -562
rect 433 -562 473 -550
rect 433 -584 445 -562
rect -445 -590 445 -584
<< properties >>
string FIXED_BBOX -450 -567 450 567
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 4 l 0.5 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 80 viagb 100 viagr 100 viagl 100 viagt 0
<< end >>
