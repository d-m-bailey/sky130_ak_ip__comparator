magic
tech sky130A
magscale 1 2
timestamp 1713548572
<< nwell >>
rect -358 -697 358 697
<< mvpmos >>
rect -100 -400 100 400
<< mvpdiff >>
rect -158 388 -100 400
rect -158 -388 -146 388
rect -112 -388 -100 388
rect -158 -400 -100 -388
rect 100 388 158 400
rect 100 -388 112 388
rect 146 -388 158 388
rect 100 -400 158 -388
<< mvpdiffc >>
rect -146 -388 -112 388
rect 112 -388 146 388
<< mvnsubdiff >>
rect -292 619 292 631
rect -292 585 -184 619
rect 184 585 292 619
rect -292 573 292 585
rect -292 -573 -234 573
rect 234 -573 292 573
rect -292 -585 292 -573
rect -292 -619 -184 -585
rect 184 -619 292 -585
rect -292 -631 292 -619
<< mvnsubdiffcont >>
rect -184 585 184 619
rect -184 -619 184 -585
<< poly >>
rect -100 481 100 497
rect -100 447 -84 481
rect 84 447 100 481
rect -100 400 100 447
rect -100 -447 100 -400
rect -100 -481 -84 -447
rect 84 -481 100 -447
rect -100 -497 100 -481
<< polycont >>
rect -84 447 84 481
rect -84 -481 84 -447
<< locali >>
rect -280 585 -184 619
rect 184 585 280 619
rect -280 -585 -246 585
rect -100 447 -84 481
rect 84 447 100 481
rect -146 388 -112 404
rect -146 -404 -112 -388
rect 112 388 146 404
rect 112 -404 146 -388
rect -100 -481 -84 -447
rect 84 -481 100 -447
rect 246 -585 280 585
rect -280 -619 -184 -585
rect 184 -619 280 -585
<< viali >>
rect -50 447 50 481
rect -146 -388 -112 388
rect 112 -388 146 388
rect -50 -481 50 -447
<< metal1 >>
rect -62 481 62 487
rect -62 447 -50 481
rect 50 447 62 481
rect -62 441 62 447
rect -152 388 -106 400
rect -152 -388 -146 388
rect -112 -388 -106 388
rect -152 -400 -106 -388
rect 106 388 152 400
rect 106 -388 112 388
rect 146 -388 152 388
rect 106 -400 152 -388
rect -62 -447 62 -441
rect -62 -481 -50 -447
rect 50 -481 62 -447
rect -62 -487 62 -481
<< properties >>
string FIXED_BBOX -263 -602 263 602
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 4 l 1 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 0 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 60 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
