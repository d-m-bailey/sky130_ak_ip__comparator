magic
tech sky130A
magscale 1 2
timestamp 1713077738
<< nwell >>
rect 29000 9700 30100 9900
rect -1070 -23030 24670 -22130
rect -770 -32850 22950 -23030
<< locali >>
rect -140 11900 22060 12060
rect -140 11620 60 11900
rect 300 11760 500 11900
rect 960 11760 1160 11900
rect 1620 11760 1820 11900
rect 2060 11620 2260 11900
rect 2500 11760 2700 11900
rect 3160 11760 3360 11900
rect 3820 11760 4020 11900
rect 4260 11620 4460 11900
rect 4700 11760 4900 11900
rect 5360 11760 5560 11900
rect 6020 11760 6220 11900
rect 6460 11620 6660 11900
rect 6900 11760 7100 11900
rect 7560 11760 7760 11900
rect 8220 11760 8420 11900
rect 8660 11620 8860 11900
rect 9100 11760 9300 11900
rect 9760 11760 9960 11900
rect 10420 11760 10620 11900
rect 10860 11620 11060 11900
rect 11300 11760 11500 11900
rect 11960 11760 12160 11900
rect 12620 11760 12820 11900
rect 13060 11620 13260 11900
rect 13500 11760 13700 11900
rect 14160 11760 14360 11900
rect 14820 11760 15020 11900
rect 15260 11620 15460 11900
rect 15700 11760 15900 11900
rect 16360 11760 16560 11900
rect 17020 11760 17220 11900
rect 17460 11620 17660 11900
rect 17900 11760 18100 11900
rect 18560 11760 18760 11900
rect 19220 11760 19420 11900
rect 19660 11620 19860 11900
rect 20100 11760 20300 11900
rect 20760 11760 20960 11900
rect 21420 11760 21620 11900
rect 21860 11620 22060 11900
rect -140 11520 200 11620
rect 1920 11520 2400 11620
rect 4120 11520 4600 11620
rect 6320 11520 6800 11620
rect 8520 11520 9000 11620
rect 10720 11520 11200 11620
rect 12920 11520 13400 11620
rect 15120 11520 15600 11620
rect 17320 11520 17800 11620
rect 19520 11520 20000 11620
rect 21720 11520 22060 11620
rect -140 11260 60 11520
rect 280 11260 480 11400
rect 960 11260 1160 11400
rect 1620 11260 1820 11400
rect 2060 11260 2260 11520
rect 2480 11260 2680 11400
rect 3160 11260 3360 11400
rect 3820 11260 4020 11400
rect 4260 11260 4460 11520
rect 4680 11260 4880 11400
rect 5360 11260 5560 11400
rect 6020 11260 6220 11400
rect 6460 11260 6660 11520
rect 6880 11260 7080 11400
rect 7560 11260 7760 11400
rect 8220 11260 8420 11400
rect 8660 11260 8860 11520
rect 9080 11260 9280 11400
rect 9760 11260 9960 11400
rect 10420 11260 10620 11400
rect 10860 11260 11060 11520
rect 11280 11260 11480 11400
rect 11960 11260 12160 11400
rect 12620 11260 12820 11400
rect 13060 11260 13260 11520
rect 13480 11260 13680 11400
rect 14160 11260 14360 11400
rect 14820 11260 15020 11400
rect 15260 11260 15460 11520
rect 15680 11260 15880 11400
rect 16360 11260 16560 11400
rect 17020 11260 17220 11400
rect 17460 11260 17660 11520
rect 17880 11260 18080 11400
rect 18560 11260 18760 11400
rect 19220 11260 19420 11400
rect 19660 11260 19860 11520
rect 20080 11260 20280 11400
rect 20760 11260 20960 11400
rect 21420 11260 21620 11400
rect 21860 11260 22060 11520
rect -140 11100 22060 11260
rect -140 10930 60 11100
rect 300 10960 500 11100
rect 960 10960 1160 11100
rect 1620 10960 1820 11100
rect -140 10870 -70 10930
rect -10 10870 60 10930
rect -140 10820 60 10870
rect 2060 10930 2260 11100
rect 2060 10870 2130 10930
rect 2190 10870 2260 10930
rect 2060 10820 2260 10870
rect -140 10720 200 10820
rect 1920 10720 2260 10820
rect -140 10460 60 10720
rect 280 10460 480 10600
rect 960 10460 1160 10600
rect 1620 10460 1820 10600
rect 2060 10460 2260 10720
rect 4260 10930 4460 11100
rect 4260 10870 4330 10930
rect 4390 10870 4460 10930
rect 4260 10460 4460 10870
rect 6460 10930 6660 11100
rect 6460 10870 6530 10930
rect 6590 10870 6660 10930
rect 6460 10460 6660 10870
rect 8660 10930 8860 11100
rect 8660 10870 8730 10930
rect 8790 10870 8860 10930
rect 8660 10460 8860 10870
rect 10860 10930 11060 11100
rect 10860 10870 10930 10930
rect 10990 10870 11060 10930
rect 10860 10460 11060 10870
rect 13060 10930 13260 11100
rect 13060 10870 13130 10930
rect 13190 10870 13260 10930
rect 13060 10460 13260 10870
rect 15260 10930 15460 11100
rect 15260 10870 15330 10930
rect 15390 10870 15460 10930
rect 15260 10460 15460 10870
rect 17460 10930 17660 11100
rect 17460 10870 17530 10930
rect 17590 10870 17660 10930
rect 17460 10460 17660 10870
rect 19660 10930 19860 11100
rect 20100 10960 20300 11100
rect 20760 10960 20960 11100
rect 21420 10960 21620 11100
rect 19660 10870 19730 10930
rect 19790 10870 19860 10930
rect 19660 10820 19860 10870
rect 21860 10930 22060 11100
rect 21860 10870 21930 10930
rect 21990 10870 22060 10930
rect 21860 10820 22060 10870
rect 19660 10720 20000 10820
rect 21720 10720 22060 10820
rect 19660 10460 19860 10720
rect 20080 10460 20280 10600
rect 20760 10460 20960 10600
rect 21420 10460 21620 10600
rect 21860 10460 22060 10720
rect -140 10300 22060 10460
rect -140 10130 60 10300
rect 300 10160 500 10300
rect 960 10160 1160 10300
rect 1620 10160 1820 10300
rect -140 10070 -70 10130
rect -10 10070 60 10130
rect -140 10020 60 10070
rect 2060 10130 2260 10300
rect 2060 10070 2130 10130
rect 2190 10070 2260 10130
rect 2060 10020 2260 10070
rect -140 9920 200 10020
rect 1920 9920 2260 10020
rect -140 9660 60 9920
rect 280 9660 480 9800
rect 960 9660 1160 9800
rect 1620 9660 1820 9800
rect 2060 9660 2260 9920
rect 4260 10130 4460 10300
rect 4260 10070 4330 10130
rect 4390 10070 4460 10130
rect 4260 9660 4460 10070
rect 6460 10130 6660 10300
rect 6460 10070 6530 10130
rect 6590 10070 6660 10130
rect 6460 9660 6660 10070
rect 8660 10130 8860 10300
rect 8660 10070 8730 10130
rect 8790 10070 8860 10130
rect 8660 9660 8860 10070
rect 10860 10130 11060 10300
rect 10860 10070 10930 10130
rect 10990 10070 11060 10130
rect 10860 9660 11060 10070
rect 13060 10130 13260 10300
rect 13060 10070 13130 10130
rect 13190 10070 13260 10130
rect 13060 9660 13260 10070
rect 15260 10130 15460 10300
rect 15260 10070 15330 10130
rect 15390 10070 15460 10130
rect 15260 9660 15460 10070
rect 17460 10130 17660 10300
rect 17460 10070 17530 10130
rect 17590 10070 17660 10130
rect 17460 9660 17660 10070
rect 19660 10130 19860 10300
rect 20100 10160 20300 10300
rect 20760 10160 20960 10300
rect 21420 10160 21620 10300
rect 19660 10070 19730 10130
rect 19790 10070 19860 10130
rect 19660 10020 19860 10070
rect 21860 10130 22060 10300
rect 21860 10070 21930 10130
rect 21990 10070 22060 10130
rect 21860 10020 22060 10070
rect 19660 9920 20000 10020
rect 21720 9920 22060 10020
rect 19660 9660 19860 9920
rect 20080 9660 20280 9800
rect 20760 9660 20960 9800
rect 21420 9660 21620 9800
rect 21860 9660 22060 9920
rect -140 9500 22060 9660
rect -140 9330 60 9500
rect 300 9360 500 9500
rect 960 9360 1160 9500
rect 1620 9360 1820 9500
rect -140 9270 -70 9330
rect -10 9270 60 9330
rect -140 9220 60 9270
rect 2060 9330 2260 9500
rect 2060 9270 2130 9330
rect 2190 9270 2260 9330
rect 2060 9220 2260 9270
rect -140 9120 200 9220
rect 1920 9120 2260 9220
rect -140 8860 60 9120
rect 280 8860 480 9000
rect 960 8860 1160 9000
rect 1620 8860 1820 9000
rect 2060 8860 2260 9120
rect 4260 9330 4460 9500
rect 4260 9270 4330 9330
rect 4390 9270 4460 9330
rect 4260 8860 4460 9270
rect 6460 9330 6660 9500
rect 6460 9270 6530 9330
rect 6590 9270 6660 9330
rect 6460 8860 6660 9270
rect 8660 9330 8860 9500
rect 8660 9270 8730 9330
rect 8790 9270 8860 9330
rect 8660 8860 8860 9270
rect 10860 9330 11060 9500
rect 10860 9270 10930 9330
rect 10990 9270 11060 9330
rect 10860 8860 11060 9270
rect 13060 9330 13260 9500
rect 13060 9270 13130 9330
rect 13190 9270 13260 9330
rect 13060 8860 13260 9270
rect 15260 9330 15460 9500
rect 15260 9270 15330 9330
rect 15390 9270 15460 9330
rect 15260 8860 15460 9270
rect 17460 9330 17660 9500
rect 17460 9270 17530 9330
rect 17590 9270 17660 9330
rect 17460 8860 17660 9270
rect 19660 9330 19860 9500
rect 20100 9360 20300 9500
rect 20760 9360 20960 9500
rect 21420 9360 21620 9500
rect 19660 9270 19730 9330
rect 19790 9270 19860 9330
rect 19660 9220 19860 9270
rect 21860 9330 22060 9500
rect 21860 9270 21930 9330
rect 21990 9270 22060 9330
rect 21860 9220 22060 9270
rect 19660 9120 20000 9220
rect 21720 9120 22060 9220
rect 19660 8860 19860 9120
rect 20080 8860 20280 9000
rect 20760 8860 20960 9000
rect 21420 8860 21620 9000
rect 21860 8860 22060 9120
rect -140 8700 22060 8860
rect -140 8530 60 8700
rect 300 8560 500 8700
rect 960 8560 1160 8700
rect 1620 8560 1820 8700
rect -140 8470 -70 8530
rect -10 8470 60 8530
rect -140 8420 60 8470
rect 2060 8530 2260 8700
rect 2060 8470 2130 8530
rect 2190 8470 2260 8530
rect 2060 8420 2260 8470
rect -140 8320 200 8420
rect 1920 8320 2260 8420
rect -140 8060 60 8320
rect 280 8060 480 8200
rect 960 8060 1160 8200
rect 1620 8060 1820 8200
rect 2060 8060 2260 8320
rect 4260 8530 4460 8700
rect 4260 8470 4330 8530
rect 4390 8470 4460 8530
rect 4260 8060 4460 8470
rect 6460 8530 6660 8700
rect 6460 8470 6530 8530
rect 6590 8470 6660 8530
rect 6460 8060 6660 8470
rect 8660 8530 8860 8700
rect 8660 8470 8730 8530
rect 8790 8470 8860 8530
rect 8660 8060 8860 8470
rect 10860 8530 11060 8700
rect 10860 8470 10930 8530
rect 10990 8470 11060 8530
rect 10860 8060 11060 8470
rect 13060 8530 13260 8700
rect 13060 8470 13130 8530
rect 13190 8470 13260 8530
rect 13060 8060 13260 8470
rect 15260 8530 15460 8700
rect 15260 8470 15330 8530
rect 15390 8470 15460 8530
rect 15260 8060 15460 8470
rect 17460 8530 17660 8700
rect 17460 8470 17530 8530
rect 17590 8470 17660 8530
rect 17460 8060 17660 8470
rect 19660 8530 19860 8700
rect 20100 8560 20300 8700
rect 20760 8560 20960 8700
rect 21420 8560 21620 8700
rect 19660 8470 19730 8530
rect 19790 8470 19860 8530
rect 19660 8420 19860 8470
rect 21860 8530 22060 8700
rect 21860 8470 21930 8530
rect 21990 8470 22060 8530
rect 21860 8420 22060 8470
rect 19660 8320 20000 8420
rect 21720 8320 22060 8420
rect 19660 8060 19860 8320
rect 20080 8060 20280 8200
rect 20760 8060 20960 8200
rect 21420 8060 21620 8200
rect 21860 8060 22060 8320
rect -140 7900 22060 8060
rect -140 7730 60 7900
rect 300 7760 500 7900
rect 960 7760 1160 7900
rect 1620 7760 1820 7900
rect -140 7670 -70 7730
rect -10 7670 60 7730
rect -140 7620 60 7670
rect 2060 7730 2260 7900
rect 2060 7670 2130 7730
rect 2190 7670 2260 7730
rect 2060 7620 2260 7670
rect -140 7520 200 7620
rect 1920 7520 2260 7620
rect -140 7260 60 7520
rect 280 7260 480 7400
rect 960 7260 1160 7400
rect 1620 7260 1820 7400
rect 2060 7260 2260 7520
rect 4260 7730 4460 7900
rect 4260 7670 4330 7730
rect 4390 7670 4460 7730
rect 4260 7260 4460 7670
rect 6460 7730 6660 7900
rect 6460 7670 6530 7730
rect 6590 7670 6660 7730
rect 6460 7260 6660 7670
rect 8660 7730 8860 7900
rect 8660 7670 8730 7730
rect 8790 7670 8860 7730
rect 8660 7260 8860 7670
rect 10860 7730 11060 7900
rect 10860 7670 10930 7730
rect 10990 7670 11060 7730
rect 10860 7260 11060 7670
rect 13060 7730 13260 7900
rect 13060 7670 13130 7730
rect 13190 7670 13260 7730
rect 13060 7260 13260 7670
rect 15260 7730 15460 7900
rect 15260 7670 15330 7730
rect 15390 7670 15460 7730
rect 15260 7260 15460 7670
rect 17460 7730 17660 7900
rect 17460 7670 17530 7730
rect 17590 7670 17660 7730
rect 17460 7260 17660 7670
rect 19660 7730 19860 7900
rect 20100 7760 20300 7900
rect 20760 7760 20960 7900
rect 21420 7760 21620 7900
rect 19660 7670 19730 7730
rect 19790 7670 19860 7730
rect 19660 7620 19860 7670
rect 21860 7730 22060 7900
rect 21860 7670 21930 7730
rect 21990 7670 22060 7730
rect 21860 7620 22060 7670
rect 19660 7520 20000 7620
rect 21720 7520 22060 7620
rect 19660 7260 19860 7520
rect 20080 7260 20280 7400
rect 20760 7260 20960 7400
rect 21420 7260 21620 7400
rect 21860 7260 22060 7520
rect -140 7100 22060 7260
rect -140 6930 60 7100
rect 300 6960 500 7100
rect 960 6960 1160 7100
rect 1620 6960 1820 7100
rect -140 6870 -70 6930
rect -10 6870 60 6930
rect -140 6820 60 6870
rect 2060 6930 2260 7100
rect 2060 6870 2130 6930
rect 2190 6870 2260 6930
rect 2060 6820 2260 6870
rect -140 6720 200 6820
rect 1920 6720 2260 6820
rect -140 6460 60 6720
rect 280 6460 480 6600
rect 960 6460 1160 6600
rect 1620 6460 1820 6600
rect 2060 6460 2260 6720
rect 4260 6930 4460 7100
rect 4260 6870 4330 6930
rect 4390 6870 4460 6930
rect 4260 6460 4460 6870
rect 6460 6930 6660 7100
rect 6460 6870 6530 6930
rect 6590 6870 6660 6930
rect 6460 6460 6660 6870
rect 8660 6930 8860 7100
rect 8660 6870 8730 6930
rect 8790 6870 8860 6930
rect 8660 6460 8860 6870
rect 10860 6930 11060 7100
rect 10860 6870 10930 6930
rect 10990 6870 11060 6930
rect 10860 6460 11060 6870
rect 13060 6930 13260 7100
rect 13060 6870 13130 6930
rect 13190 6870 13260 6930
rect 13060 6460 13260 6870
rect 15260 6930 15460 7100
rect 15260 6870 15330 6930
rect 15390 6870 15460 6930
rect 15260 6460 15460 6870
rect 17460 6930 17660 7100
rect 17460 6870 17530 6930
rect 17590 6870 17660 6930
rect 17460 6460 17660 6870
rect 19660 6930 19860 7100
rect 20100 6960 20300 7100
rect 20760 6960 20960 7100
rect 21420 6960 21620 7100
rect 19660 6870 19730 6930
rect 19790 6870 19860 6930
rect 19660 6820 19860 6870
rect 21860 6930 22060 7100
rect 21860 6870 21930 6930
rect 21990 6870 22060 6930
rect 21860 6820 22060 6870
rect 19660 6720 20000 6820
rect 21720 6720 22060 6820
rect 19660 6460 19860 6720
rect 20080 6460 20280 6600
rect 20760 6460 20960 6600
rect 21420 6460 21620 6600
rect 21860 6460 22060 6720
rect -140 6300 22060 6460
rect -140 6130 60 6300
rect 300 6160 500 6300
rect 960 6160 1160 6300
rect 1620 6160 1820 6300
rect -140 6070 -70 6130
rect -10 6070 60 6130
rect -140 6020 60 6070
rect 2060 6130 2260 6300
rect 2060 6070 2130 6130
rect 2190 6070 2260 6130
rect 2060 6020 2260 6070
rect -140 5920 200 6020
rect 1920 5920 2260 6020
rect -140 5660 60 5920
rect 280 5660 480 5800
rect 960 5660 1160 5800
rect 1620 5660 1820 5800
rect 2060 5660 2260 5920
rect 4260 6130 4460 6300
rect 4260 6070 4330 6130
rect 4390 6070 4460 6130
rect 4260 5660 4460 6070
rect 6460 6130 6660 6300
rect 6460 6070 6530 6130
rect 6590 6070 6660 6130
rect 6460 5660 6660 6070
rect 8660 6130 8860 6300
rect 8660 6070 8730 6130
rect 8790 6070 8860 6130
rect 8660 5660 8860 6070
rect 10860 6130 11060 6300
rect 10860 6070 10930 6130
rect 10990 6070 11060 6130
rect 10860 5660 11060 6070
rect 13060 6130 13260 6300
rect 13060 6070 13130 6130
rect 13190 6070 13260 6130
rect 13060 5660 13260 6070
rect 15260 6130 15460 6300
rect 15260 6070 15330 6130
rect 15390 6070 15460 6130
rect 15260 5660 15460 6070
rect 17460 6130 17660 6300
rect 17460 6070 17530 6130
rect 17590 6070 17660 6130
rect 17460 5660 17660 6070
rect 19660 6130 19860 6300
rect 20100 6160 20300 6300
rect 20760 6160 20960 6300
rect 21420 6160 21620 6300
rect 19660 6070 19730 6130
rect 19790 6070 19860 6130
rect 19660 6020 19860 6070
rect 21860 6130 22060 6300
rect 21860 6070 21930 6130
rect 21990 6070 22060 6130
rect 21860 6020 22060 6070
rect 19660 5920 20000 6020
rect 21720 5920 22060 6020
rect 19660 5660 19860 5920
rect 20080 5660 20280 5800
rect 20760 5660 20960 5800
rect 21420 5660 21620 5800
rect 21860 5660 22060 5920
rect -140 5500 22060 5660
rect -140 5330 60 5500
rect 300 5360 500 5500
rect 960 5360 1160 5500
rect 1620 5360 1820 5500
rect -140 5270 -70 5330
rect -10 5270 60 5330
rect -140 5220 60 5270
rect 2060 5330 2260 5500
rect 2060 5270 2130 5330
rect 2190 5270 2260 5330
rect 2060 5220 2260 5270
rect -140 5120 200 5220
rect 1920 5120 2260 5220
rect -140 4860 60 5120
rect 280 4860 480 5000
rect 960 4860 1160 5000
rect 1620 4860 1820 5000
rect 2060 4860 2260 5120
rect 4260 5330 4460 5500
rect 4260 5270 4330 5330
rect 4390 5270 4460 5330
rect 4260 4860 4460 5270
rect 6460 5330 6660 5500
rect 6460 5270 6530 5330
rect 6590 5270 6660 5330
rect 6460 4860 6660 5270
rect 8660 5330 8860 5500
rect 8660 5270 8730 5330
rect 8790 5270 8860 5330
rect 8660 4860 8860 5270
rect 10860 5330 11060 5500
rect 10860 5270 10930 5330
rect 10990 5270 11060 5330
rect 10860 4860 11060 5270
rect 13060 5330 13260 5500
rect 13060 5270 13130 5330
rect 13190 5270 13260 5330
rect 13060 4860 13260 5270
rect 15260 5330 15460 5500
rect 15260 5270 15330 5330
rect 15390 5270 15460 5330
rect 15260 4860 15460 5270
rect 17460 5330 17660 5500
rect 17460 5270 17530 5330
rect 17590 5270 17660 5330
rect 17460 4860 17660 5270
rect 19660 5330 19860 5500
rect 20100 5360 20300 5500
rect 20760 5360 20960 5500
rect 21420 5360 21620 5500
rect 19660 5270 19730 5330
rect 19790 5270 19860 5330
rect 19660 5220 19860 5270
rect 21860 5330 22060 5500
rect 21860 5270 21930 5330
rect 21990 5270 22060 5330
rect 21860 5220 22060 5270
rect 19660 5120 20000 5220
rect 21720 5120 22060 5220
rect 19660 4860 19860 5120
rect 20080 4860 20280 5000
rect 20760 4860 20960 5000
rect 21420 4860 21620 5000
rect 21860 4860 22060 5120
rect -140 4700 22060 4860
rect -140 4420 60 4700
rect 300 4560 500 4700
rect 960 4560 1160 4700
rect 1620 4560 1820 4700
rect 2060 4420 2260 4700
rect 2500 4560 2700 4700
rect 3160 4560 3360 4700
rect 3820 4560 4020 4700
rect 4260 4420 4460 4700
rect 4700 4560 4900 4700
rect 5360 4560 5560 4700
rect 6020 4560 6220 4700
rect 6460 4420 6660 4700
rect 6900 4560 7100 4700
rect 7560 4560 7760 4700
rect 8220 4560 8420 4700
rect 8660 4420 8860 4700
rect 9100 4560 9300 4700
rect 9760 4560 9960 4700
rect 10420 4560 10620 4700
rect 10860 4420 11060 4700
rect 11300 4560 11500 4700
rect 11960 4560 12160 4700
rect 12620 4560 12820 4700
rect 13060 4420 13260 4700
rect 13500 4560 13700 4700
rect 14160 4560 14360 4700
rect 14820 4560 15020 4700
rect 15260 4420 15460 4700
rect 15700 4560 15900 4700
rect 16360 4560 16560 4700
rect 17020 4560 17220 4700
rect 17460 4420 17660 4700
rect 17900 4560 18100 4700
rect 18560 4560 18760 4700
rect 19220 4560 19420 4700
rect 19660 4420 19860 4700
rect 20100 4560 20300 4700
rect 20760 4560 20960 4700
rect 21420 4560 21620 4700
rect 21860 4420 22060 4700
rect -140 4320 200 4420
rect 1920 4320 2400 4420
rect 4120 4320 4600 4420
rect 6320 4320 6800 4420
rect 8520 4320 9000 4420
rect 10720 4320 11200 4420
rect 12920 4320 13400 4420
rect 15120 4320 15600 4420
rect 17320 4320 17800 4420
rect 19520 4320 20000 4420
rect 21720 4320 22060 4420
rect -140 4060 60 4320
rect 280 4060 480 4200
rect 960 4060 1160 4200
rect 1620 4060 1820 4200
rect 2060 4060 2260 4320
rect 2480 4060 2680 4200
rect 3160 4060 3360 4200
rect 3820 4060 4020 4200
rect 4260 4060 4460 4320
rect 4680 4060 4880 4200
rect 5360 4060 5560 4200
rect 6020 4060 6220 4200
rect 6460 4060 6660 4320
rect 6880 4060 7080 4200
rect 7560 4060 7760 4200
rect 8220 4060 8420 4200
rect 8660 4060 8860 4320
rect 9080 4060 9280 4200
rect 9760 4060 9960 4200
rect 10420 4060 10620 4200
rect 10860 4060 11060 4320
rect 11280 4060 11480 4200
rect 11960 4060 12160 4200
rect 12620 4060 12820 4200
rect 13060 4060 13260 4320
rect 13480 4060 13680 4200
rect 14160 4060 14360 4200
rect 14820 4060 15020 4200
rect 15260 4060 15460 4320
rect 15680 4060 15880 4200
rect 16360 4060 16560 4200
rect 17020 4060 17220 4200
rect 17460 4060 17660 4320
rect 17880 4060 18080 4200
rect 18560 4060 18760 4200
rect 19220 4060 19420 4200
rect 19660 4060 19860 4320
rect 20080 4060 20280 4200
rect 20760 4060 20960 4200
rect 21420 4060 21620 4200
rect 21860 4060 22060 4320
rect -140 3900 22060 4060
rect -340 2190 38280 2980
rect -340 2113 -117 2190
rect -340 2020 -130 2113
rect 60 2075 450 2190
rect 55 2060 463 2075
rect 55 2041 71 2060
rect 447 2041 463 2060
rect 500 2029 630 2190
rect 680 2075 1070 2190
rect 1253 2113 1470 2190
rect 673 2060 1081 2075
rect 673 2041 689 2060
rect 1065 2041 1081 2060
rect -13 2020 21 2029
rect -340 2013 21 2020
rect 497 2013 639 2029
rect 1115 2020 1149 2029
rect 1260 2020 1470 2113
rect 1115 2013 1470 2020
rect -340 1245 10 2013
rect 500 1245 630 2013
rect 1120 1245 1470 2013
rect -340 1240 21 1245
rect -340 1145 -130 1240
rect -13 1229 21 1240
rect 497 1240 639 1245
rect 497 1229 531 1240
rect 605 1229 639 1240
rect 1115 1240 1470 1245
rect 1115 1229 1149 1240
rect 55 1210 71 1217
rect 55 1183 440 1210
rect 447 1183 463 1217
rect 673 1183 689 1217
rect -340 1110 -117 1145
rect 70 1110 440 1183
rect 690 1110 1060 1210
rect 1065 1183 1081 1217
rect 1260 1145 1470 1240
rect 1253 1110 1470 1145
rect -340 1030 1470 1110
rect -340 987 -117 1030
rect -340 900 -130 987
rect 70 949 440 1030
rect 55 930 440 949
rect 55 915 71 930
rect 447 915 463 949
rect 673 915 689 949
rect 690 930 1060 1030
rect 1253 987 1470 1030
rect 1065 915 1081 949
rect -13 900 21 903
rect -340 887 21 900
rect 497 900 531 903
rect 605 900 639 903
rect 497 887 639 900
rect 1115 887 1149 903
rect -340 719 10 887
rect 500 719 630 887
rect 1260 860 1470 987
rect 1130 750 1470 860
rect -340 710 21 719
rect -340 619 -130 710
rect -13 703 21 710
rect 497 703 639 719
rect 1115 703 1149 719
rect 55 680 71 691
rect 55 657 440 680
rect 447 657 463 691
rect -340 557 -117 619
rect -340 550 -55 557
rect 70 550 440 657
rect 500 550 630 703
rect 673 657 689 691
rect 690 550 1060 680
rect 1065 657 1081 691
rect 1260 619 1470 750
rect 1253 557 1470 619
rect 1191 550 1470 557
rect 2860 550 3070 2190
rect 4460 550 4670 2190
rect 6060 550 6270 2190
rect 7660 550 7870 2190
rect 9260 550 9470 2190
rect 10860 550 11070 2190
rect 12460 550 12670 2190
rect 14060 550 14270 2190
rect 15660 550 15870 2190
rect 17260 550 17470 2190
rect 18860 550 19070 2190
rect 20460 550 20670 2190
rect 22060 550 22270 2190
rect 23660 550 23870 2190
rect 25260 550 25470 2190
rect 26860 550 27070 2190
rect 28460 550 28670 2190
rect 30060 550 30270 2190
rect 31660 550 31870 2190
rect 33260 550 33470 2190
rect 34860 550 35070 2190
rect 36460 2113 36683 2190
rect 36460 2020 36670 2113
rect 36860 2075 37250 2190
rect 36855 2060 37263 2075
rect 36855 2041 36871 2060
rect 37247 2041 37263 2060
rect 37300 2029 37430 2190
rect 37480 2075 37870 2190
rect 38053 2113 38280 2190
rect 37473 2060 37881 2075
rect 37473 2041 37489 2060
rect 37865 2041 37881 2060
rect 36787 2020 36821 2029
rect 36460 2013 36821 2020
rect 37297 2013 37439 2029
rect 37915 2020 37949 2029
rect 38060 2020 38280 2113
rect 37915 2013 38280 2020
rect 36460 1245 36810 2013
rect 37300 1245 37430 2013
rect 37920 1245 38280 2013
rect 36460 1240 36821 1245
rect 36460 1145 36670 1240
rect 36787 1229 36821 1240
rect 37297 1240 37439 1245
rect 37297 1229 37331 1240
rect 37405 1229 37439 1240
rect 37915 1240 38280 1245
rect 37915 1229 37949 1240
rect 36855 1210 36871 1217
rect 36855 1183 37240 1210
rect 37247 1183 37263 1217
rect 37473 1183 37489 1217
rect 36460 1110 36683 1145
rect 36870 1110 37240 1183
rect 37490 1110 37860 1210
rect 37865 1183 37881 1217
rect 38060 1145 38280 1240
rect 38053 1110 38280 1145
rect 36460 1030 38280 1110
rect 36460 987 36683 1030
rect 36460 900 36670 987
rect 36870 949 37240 1030
rect 36855 930 37240 949
rect 36855 915 36871 930
rect 37247 915 37263 949
rect 37473 915 37489 949
rect 37490 930 37860 1030
rect 38053 987 38280 1030
rect 37865 915 37881 949
rect 36787 900 36821 903
rect 36460 887 36821 900
rect 37297 900 37331 903
rect 37405 900 37439 903
rect 37297 887 37439 900
rect 37915 887 37949 903
rect 36460 719 36810 887
rect 37300 719 37430 887
rect 38060 860 38280 987
rect 37930 750 38280 860
rect 36460 710 36821 719
rect 36460 619 36670 710
rect 36787 703 36821 710
rect 37297 703 37439 719
rect 37915 703 37949 719
rect 36855 680 36871 691
rect 36855 657 37240 680
rect 37247 657 37263 691
rect 36460 557 36683 619
rect 36460 550 36745 557
rect 36870 550 37240 657
rect 37300 550 37430 703
rect 37473 657 37489 691
rect 37490 550 37860 680
rect 37865 657 37881 691
rect 38060 619 38280 750
rect 38053 557 38280 619
rect 37991 550 38280 557
rect -340 390 38280 550
rect -340 313 -117 390
rect -340 220 -130 313
rect 60 275 450 390
rect 55 260 463 275
rect 55 241 71 260
rect 447 241 463 260
rect 500 229 630 390
rect 680 275 1070 390
rect 1253 313 1470 390
rect 673 260 1081 275
rect 673 241 689 260
rect 1065 241 1081 260
rect -13 220 21 229
rect -340 213 21 220
rect 497 213 639 229
rect 1115 220 1149 229
rect 1260 220 1470 313
rect 1115 213 1470 220
rect -340 -555 10 213
rect 500 -555 630 213
rect 1120 -555 1470 213
rect -340 -560 21 -555
rect -340 -655 -130 -560
rect -13 -571 21 -560
rect 497 -560 639 -555
rect 497 -571 531 -560
rect 605 -571 639 -560
rect 1115 -560 1470 -555
rect 1115 -571 1149 -560
rect 55 -590 71 -583
rect 55 -617 440 -590
rect 447 -617 463 -583
rect 673 -617 689 -583
rect -340 -690 -117 -655
rect 70 -690 440 -617
rect 690 -690 1060 -590
rect 1065 -617 1081 -583
rect 1260 -655 1470 -560
rect 1253 -690 1470 -655
rect -340 -770 1470 -690
rect -340 -813 -117 -770
rect -340 -900 -130 -813
rect 70 -851 440 -770
rect 55 -870 440 -851
rect 55 -885 71 -870
rect 447 -885 463 -851
rect 673 -885 689 -851
rect 690 -870 1060 -770
rect 1253 -813 1470 -770
rect 1065 -885 1081 -851
rect -13 -900 21 -897
rect -340 -913 21 -900
rect 497 -900 531 -897
rect 605 -900 639 -897
rect 497 -913 639 -900
rect 1115 -913 1149 -897
rect -340 -1081 10 -913
rect 500 -1081 630 -913
rect 1260 -940 1470 -813
rect 1130 -1050 1470 -940
rect -340 -1090 21 -1081
rect -340 -1181 -130 -1090
rect -13 -1097 21 -1090
rect 497 -1097 639 -1081
rect 1115 -1097 1149 -1081
rect 55 -1120 71 -1109
rect 55 -1143 440 -1120
rect 447 -1143 463 -1109
rect -340 -1243 -117 -1181
rect -340 -1250 -55 -1243
rect 70 -1250 440 -1143
rect 500 -1250 630 -1097
rect 673 -1143 689 -1109
rect 690 -1250 1060 -1120
rect 1065 -1143 1081 -1109
rect 1260 -1181 1470 -1050
rect 1253 -1243 1470 -1181
rect 1191 -1250 1470 -1243
rect 2860 -1250 3070 390
rect 4460 -1250 4670 390
rect 6060 -1250 6270 390
rect 7660 -1250 7870 390
rect 9260 -1250 9470 390
rect 10860 -1250 11070 390
rect 12460 -1250 12670 390
rect 14060 -1250 14270 390
rect 15660 -1250 15870 390
rect 17260 -1250 17470 390
rect 18860 -1250 19070 390
rect 20460 -1250 20670 390
rect 22060 -1250 22270 390
rect 23660 -1250 23870 390
rect 25260 -1250 25470 390
rect 26860 -1250 27070 390
rect 28460 -1250 28670 390
rect 30060 -1250 30270 390
rect 31660 -1250 31870 390
rect 33260 -1250 33470 390
rect 34860 -1250 35070 390
rect 36460 313 36683 390
rect 36460 220 36670 313
rect 36860 275 37250 390
rect 36855 260 37263 275
rect 36855 241 36871 260
rect 37247 241 37263 260
rect 37300 229 37430 390
rect 37480 275 37870 390
rect 38053 313 38280 390
rect 37473 260 37881 275
rect 37473 241 37489 260
rect 37865 241 37881 260
rect 36787 220 36821 229
rect 36460 213 36821 220
rect 37297 213 37439 229
rect 37915 220 37949 229
rect 38060 220 38280 313
rect 37915 213 38280 220
rect 36460 -555 36810 213
rect 37300 -555 37430 213
rect 37920 -555 38280 213
rect 36460 -560 36821 -555
rect 36460 -655 36670 -560
rect 36787 -571 36821 -560
rect 37297 -560 37439 -555
rect 37297 -571 37331 -560
rect 37405 -571 37439 -560
rect 37915 -560 38280 -555
rect 37915 -571 37949 -560
rect 36855 -590 36871 -583
rect 36855 -617 37240 -590
rect 37247 -617 37263 -583
rect 37473 -617 37489 -583
rect 36460 -690 36683 -655
rect 36870 -690 37240 -617
rect 37490 -690 37860 -590
rect 37865 -617 37881 -583
rect 38060 -655 38280 -560
rect 38053 -690 38280 -655
rect 36460 -770 38280 -690
rect 36460 -813 36683 -770
rect 36460 -900 36670 -813
rect 36870 -851 37240 -770
rect 36855 -870 37240 -851
rect 36855 -885 36871 -870
rect 37247 -885 37263 -851
rect 37473 -885 37489 -851
rect 37490 -870 37860 -770
rect 38053 -813 38280 -770
rect 37865 -885 37881 -851
rect 36787 -900 36821 -897
rect 36460 -913 36821 -900
rect 37297 -900 37331 -897
rect 37405 -900 37439 -897
rect 37297 -913 37439 -900
rect 37915 -913 37949 -897
rect 36460 -1081 36810 -913
rect 37300 -1081 37430 -913
rect 38060 -940 38280 -813
rect 37930 -1050 38280 -940
rect 36460 -1090 36821 -1081
rect 36460 -1181 36670 -1090
rect 36787 -1097 36821 -1090
rect 37297 -1097 37439 -1081
rect 37915 -1097 37949 -1081
rect 36855 -1120 36871 -1109
rect 36855 -1143 37240 -1120
rect 37247 -1143 37263 -1109
rect 36460 -1243 36683 -1181
rect 36460 -1250 36745 -1243
rect 36870 -1250 37240 -1143
rect 37300 -1250 37430 -1097
rect 37473 -1143 37489 -1109
rect 37490 -1250 37860 -1120
rect 37865 -1143 37881 -1109
rect 38060 -1181 38280 -1050
rect 38053 -1243 38280 -1181
rect 37991 -1250 38280 -1243
rect -340 -1410 38280 -1250
rect -340 -1487 -117 -1410
rect -340 -1580 -130 -1487
rect 60 -1525 450 -1410
rect 55 -1540 463 -1525
rect 55 -1559 71 -1540
rect 447 -1559 463 -1540
rect 500 -1571 630 -1410
rect 680 -1525 1070 -1410
rect 1253 -1487 1470 -1410
rect 673 -1540 1081 -1525
rect 673 -1559 689 -1540
rect 1065 -1559 1081 -1540
rect -13 -1580 21 -1571
rect -340 -1587 21 -1580
rect 497 -1587 639 -1571
rect 1115 -1580 1149 -1571
rect 1260 -1580 1470 -1487
rect 1115 -1587 1470 -1580
rect -340 -2355 10 -1587
rect 500 -2355 630 -1587
rect 1120 -2355 1470 -1587
rect -340 -2360 21 -2355
rect -340 -2455 -130 -2360
rect -13 -2371 21 -2360
rect 497 -2360 639 -2355
rect 497 -2371 531 -2360
rect 605 -2371 639 -2360
rect 1115 -2360 1470 -2355
rect 1115 -2371 1149 -2360
rect 55 -2390 71 -2383
rect 55 -2417 440 -2390
rect 447 -2417 463 -2383
rect 673 -2417 689 -2383
rect -340 -2490 -117 -2455
rect 70 -2490 440 -2417
rect 690 -2490 1060 -2390
rect 1065 -2417 1081 -2383
rect 1260 -2455 1470 -2360
rect 1253 -2490 1470 -2455
rect -340 -2570 1470 -2490
rect -340 -2613 -117 -2570
rect -340 -2700 -130 -2613
rect 70 -2651 440 -2570
rect 55 -2670 440 -2651
rect 55 -2685 71 -2670
rect 447 -2685 463 -2651
rect 673 -2685 689 -2651
rect 690 -2670 1060 -2570
rect 1253 -2613 1470 -2570
rect 1065 -2685 1081 -2651
rect -13 -2700 21 -2697
rect -340 -2713 21 -2700
rect 497 -2700 531 -2697
rect 605 -2700 639 -2697
rect 497 -2713 639 -2700
rect 1115 -2713 1149 -2697
rect -340 -2881 10 -2713
rect 500 -2881 630 -2713
rect 1260 -2740 1470 -2613
rect 1130 -2850 1470 -2740
rect -340 -2890 21 -2881
rect -340 -2981 -130 -2890
rect -13 -2897 21 -2890
rect 497 -2897 639 -2881
rect 1115 -2897 1149 -2881
rect 55 -2920 71 -2909
rect 55 -2943 440 -2920
rect 447 -2943 463 -2909
rect -340 -3043 -117 -2981
rect -340 -3050 -55 -3043
rect 70 -3050 440 -2943
rect 500 -3050 630 -2897
rect 673 -2943 689 -2909
rect 690 -3050 1060 -2920
rect 1065 -2943 1081 -2909
rect 1260 -2981 1470 -2850
rect 1253 -3043 1470 -2981
rect 1191 -3050 1470 -3043
rect 2860 -3050 3070 -1410
rect 4460 -3050 4670 -1410
rect 6060 -3050 6270 -1410
rect 7660 -3050 7870 -1410
rect 9260 -3050 9470 -1410
rect 10860 -3050 11070 -1410
rect 12460 -3050 12670 -1410
rect 14060 -3050 14270 -1410
rect 15660 -3050 15870 -1410
rect 17260 -3050 17470 -1410
rect 18860 -3050 19070 -1410
rect 20460 -3050 20670 -1410
rect 22060 -3050 22270 -1410
rect 23660 -3050 23870 -1410
rect 25260 -3050 25470 -1410
rect 26860 -3050 27070 -1410
rect 28460 -3050 28670 -1410
rect 30060 -3050 30270 -1410
rect 31660 -3050 31870 -1410
rect 33260 -3050 33470 -1410
rect 34860 -3050 35070 -1410
rect 36460 -1487 36683 -1410
rect 36460 -1580 36670 -1487
rect 36860 -1525 37250 -1410
rect 36855 -1540 37263 -1525
rect 36855 -1559 36871 -1540
rect 37247 -1559 37263 -1540
rect 37300 -1571 37430 -1410
rect 37480 -1525 37870 -1410
rect 38053 -1487 38280 -1410
rect 37473 -1540 37881 -1525
rect 37473 -1559 37489 -1540
rect 37865 -1559 37881 -1540
rect 36787 -1580 36821 -1571
rect 36460 -1587 36821 -1580
rect 37297 -1587 37439 -1571
rect 37915 -1580 37949 -1571
rect 38060 -1580 38280 -1487
rect 37915 -1587 38280 -1580
rect 36460 -2355 36810 -1587
rect 37300 -2355 37430 -1587
rect 37920 -2355 38280 -1587
rect 36460 -2360 36821 -2355
rect 36460 -2455 36670 -2360
rect 36787 -2371 36821 -2360
rect 37297 -2360 37439 -2355
rect 37297 -2371 37331 -2360
rect 37405 -2371 37439 -2360
rect 37915 -2360 38280 -2355
rect 37915 -2371 37949 -2360
rect 36855 -2390 36871 -2383
rect 36855 -2417 37240 -2390
rect 37247 -2417 37263 -2383
rect 37473 -2417 37489 -2383
rect 36460 -2490 36683 -2455
rect 36870 -2490 37240 -2417
rect 37490 -2490 37860 -2390
rect 37865 -2417 37881 -2383
rect 38060 -2455 38280 -2360
rect 38053 -2490 38280 -2455
rect 36460 -2570 38280 -2490
rect 36460 -2613 36683 -2570
rect 36460 -2700 36670 -2613
rect 36870 -2651 37240 -2570
rect 36855 -2670 37240 -2651
rect 36855 -2685 36871 -2670
rect 37247 -2685 37263 -2651
rect 37473 -2685 37489 -2651
rect 37490 -2670 37860 -2570
rect 38053 -2613 38280 -2570
rect 37865 -2685 37881 -2651
rect 36787 -2700 36821 -2697
rect 36460 -2713 36821 -2700
rect 37297 -2700 37331 -2697
rect 37405 -2700 37439 -2697
rect 37297 -2713 37439 -2700
rect 37915 -2713 37949 -2697
rect 36460 -2881 36810 -2713
rect 37300 -2881 37430 -2713
rect 38060 -2740 38280 -2613
rect 37930 -2850 38280 -2740
rect 36460 -2890 36821 -2881
rect 36460 -2981 36670 -2890
rect 36787 -2897 36821 -2890
rect 37297 -2897 37439 -2881
rect 37915 -2897 37949 -2881
rect 36855 -2920 36871 -2909
rect 36855 -2943 37240 -2920
rect 37247 -2943 37263 -2909
rect 36460 -3043 36683 -2981
rect 36460 -3050 36745 -3043
rect 36870 -3050 37240 -2943
rect 37300 -3050 37430 -2897
rect 37473 -2943 37489 -2909
rect 37490 -3050 37860 -2920
rect 37865 -2943 37881 -2909
rect 38060 -2981 38280 -2850
rect 38053 -3043 38280 -2981
rect 37991 -3050 38280 -3043
rect -340 -3210 38280 -3050
rect -340 -3380 -130 -3210
rect 60 -3340 450 -3210
rect -340 -4160 10 -3380
rect 500 -4160 630 -3210
rect 680 -3340 1070 -3210
rect 1260 -3380 1470 -3210
rect 1120 -4160 1470 -3380
rect -340 -4290 -130 -4160
rect 70 -4290 440 -4190
rect 690 -4290 1060 -4190
rect 1260 -4290 1470 -4160
rect -340 -4370 1470 -4290
rect -340 -4500 -130 -4370
rect 70 -4470 440 -4370
rect 690 -4470 1060 -4370
rect -340 -4690 10 -4500
rect -340 -4850 -130 -4690
rect 70 -4850 440 -4720
rect 500 -4850 630 -4500
rect 1260 -4540 1470 -4370
rect 1130 -4650 1470 -4540
rect 690 -4850 1060 -4720
rect 1260 -4850 1470 -4650
rect 2860 -4850 3070 -3210
rect 4460 -4850 4670 -3210
rect 6060 -4850 6270 -3210
rect 7660 -4850 7870 -3210
rect 9260 -4850 9470 -3210
rect 10860 -4850 11070 -3210
rect 12460 -4850 12670 -3210
rect 14060 -4850 14270 -3210
rect 15660 -4850 15870 -3210
rect 17260 -4850 17470 -3210
rect 18860 -4850 19070 -3210
rect 20460 -4850 20670 -3210
rect 22060 -4850 22270 -3210
rect 23660 -4850 23870 -3210
rect 25260 -4850 25470 -3210
rect 26860 -4850 27070 -3210
rect 28460 -4850 28670 -3210
rect 30060 -4850 30270 -3210
rect 31660 -4850 31870 -3210
rect 33260 -4850 33470 -3210
rect 34860 -4850 35070 -3210
rect 36460 -3287 36683 -3210
rect 36460 -3380 36670 -3287
rect 36860 -3325 37250 -3210
rect 36855 -3340 37263 -3325
rect 36855 -3359 36871 -3340
rect 37247 -3359 37263 -3340
rect 37300 -3371 37430 -3210
rect 37480 -3325 37870 -3210
rect 38053 -3287 38280 -3210
rect 37473 -3340 37881 -3325
rect 37473 -3359 37489 -3340
rect 37865 -3359 37881 -3340
rect 36787 -3380 36821 -3371
rect 36460 -3387 36821 -3380
rect 37297 -3387 37439 -3371
rect 37915 -3380 37949 -3371
rect 38060 -3380 38280 -3287
rect 37915 -3387 38280 -3380
rect 36460 -4155 36810 -3387
rect 37300 -4155 37430 -3387
rect 37920 -4155 38280 -3387
rect 36460 -4160 36821 -4155
rect 36460 -4255 36670 -4160
rect 36787 -4171 36821 -4160
rect 37297 -4160 37439 -4155
rect 37297 -4171 37331 -4160
rect 37405 -4171 37439 -4160
rect 37915 -4160 38280 -4155
rect 37915 -4171 37949 -4160
rect 36855 -4190 36871 -4183
rect 36855 -4217 37240 -4190
rect 37247 -4217 37263 -4183
rect 37473 -4217 37489 -4183
rect 36460 -4290 36683 -4255
rect 36870 -4290 37240 -4217
rect 37490 -4290 37860 -4190
rect 37865 -4217 37881 -4183
rect 38060 -4255 38280 -4160
rect 38053 -4290 38280 -4255
rect 36460 -4370 38280 -4290
rect 36460 -4413 36683 -4370
rect 36460 -4500 36670 -4413
rect 36870 -4451 37240 -4370
rect 36855 -4470 37240 -4451
rect 36855 -4485 36871 -4470
rect 37247 -4485 37263 -4451
rect 37473 -4485 37489 -4451
rect 37490 -4470 37860 -4370
rect 38053 -4413 38280 -4370
rect 37865 -4485 37881 -4451
rect 36787 -4500 36821 -4497
rect 36460 -4513 36821 -4500
rect 37297 -4500 37331 -4497
rect 37405 -4500 37439 -4497
rect 37297 -4513 37439 -4500
rect 37915 -4513 37949 -4497
rect 36460 -4681 36810 -4513
rect 37300 -4681 37430 -4513
rect 38060 -4540 38280 -4413
rect 37930 -4650 38280 -4540
rect 36460 -4690 36821 -4681
rect 36460 -4781 36670 -4690
rect 36787 -4697 36821 -4690
rect 37297 -4697 37439 -4681
rect 37915 -4697 37949 -4681
rect 36855 -4720 36871 -4709
rect 36855 -4743 37240 -4720
rect 37247 -4743 37263 -4709
rect 36460 -4843 36683 -4781
rect 36460 -4850 36745 -4843
rect 36870 -4850 37240 -4743
rect 37300 -4850 37430 -4697
rect 37473 -4743 37489 -4709
rect 37490 -4850 37860 -4720
rect 37865 -4743 37881 -4709
rect 38060 -4781 38280 -4650
rect 38053 -4843 38280 -4781
rect 37991 -4850 38280 -4843
rect -340 -5520 38280 -4850
rect 14900 -6620 15040 -5520
rect -140 -24180 22060 -24020
rect -140 -24440 60 -24180
rect 300 -24320 500 -24180
rect 960 -24320 1160 -24180
rect 1640 -24320 1840 -24180
rect 2060 -24440 2260 -24180
rect 2500 -24320 2700 -24180
rect 3160 -24320 3360 -24180
rect 3840 -24320 4040 -24180
rect 4260 -24440 4460 -24180
rect 4700 -24320 4900 -24180
rect 5360 -24320 5560 -24180
rect 6040 -24320 6240 -24180
rect 6460 -24440 6660 -24180
rect 6900 -24320 7100 -24180
rect 7560 -24320 7760 -24180
rect 8240 -24320 8440 -24180
rect 8660 -24440 8860 -24180
rect 9100 -24320 9300 -24180
rect 9760 -24320 9960 -24180
rect 10440 -24320 10640 -24180
rect 10860 -24440 11060 -24180
rect 11300 -24320 11500 -24180
rect 11960 -24320 12160 -24180
rect 12640 -24320 12840 -24180
rect 13060 -24440 13260 -24180
rect 13500 -24320 13700 -24180
rect 14160 -24320 14360 -24180
rect 14840 -24320 15040 -24180
rect 15260 -24440 15460 -24180
rect 15700 -24320 15900 -24180
rect 16360 -24320 16560 -24180
rect 17040 -24320 17240 -24180
rect 17460 -24440 17660 -24180
rect 17900 -24320 18100 -24180
rect 18560 -24320 18760 -24180
rect 19240 -24320 19440 -24180
rect 19660 -24440 19860 -24180
rect 20100 -24320 20300 -24180
rect 20760 -24320 20960 -24180
rect 21440 -24320 21640 -24180
rect 21860 -24440 22060 -24180
rect -140 -24540 200 -24440
rect 1920 -24540 2400 -24440
rect 4120 -24540 4600 -24440
rect 6320 -24540 6800 -24440
rect 8520 -24540 9000 -24440
rect 10720 -24540 11200 -24440
rect 12920 -24540 13400 -24440
rect 15120 -24540 15600 -24440
rect 17320 -24540 17800 -24440
rect 19520 -24540 20000 -24440
rect 21720 -24540 22060 -24440
rect -140 -24820 60 -24540
rect 300 -24820 500 -24680
rect 960 -24820 1160 -24680
rect 1620 -24820 1820 -24680
rect 2060 -24820 2260 -24540
rect 2500 -24820 2700 -24680
rect 3160 -24820 3360 -24680
rect 3820 -24820 4020 -24680
rect 4260 -24820 4460 -24540
rect 4700 -24820 4900 -24680
rect 5360 -24820 5560 -24680
rect 6020 -24820 6220 -24680
rect 6460 -24820 6660 -24540
rect 6900 -24820 7100 -24680
rect 7560 -24820 7760 -24680
rect 8220 -24820 8420 -24680
rect 8660 -24820 8860 -24540
rect 9100 -24820 9300 -24680
rect 9760 -24820 9960 -24680
rect 10420 -24820 10620 -24680
rect 10860 -24820 11060 -24540
rect 11300 -24820 11500 -24680
rect 11960 -24820 12160 -24680
rect 12620 -24820 12820 -24680
rect 13060 -24820 13260 -24540
rect 13500 -24820 13700 -24680
rect 14160 -24820 14360 -24680
rect 14820 -24820 15020 -24680
rect 15260 -24820 15460 -24540
rect 15700 -24820 15900 -24680
rect 16360 -24820 16560 -24680
rect 17020 -24820 17220 -24680
rect 17460 -24820 17660 -24540
rect 17900 -24820 18100 -24680
rect 18560 -24820 18760 -24680
rect 19220 -24820 19420 -24680
rect 19660 -24820 19860 -24540
rect 20100 -24820 20300 -24680
rect 20760 -24820 20960 -24680
rect 21420 -24820 21620 -24680
rect 21860 -24820 22060 -24540
rect -140 -24980 22060 -24820
rect -140 -25240 60 -24980
rect 300 -25120 500 -24980
rect 960 -25120 1160 -24980
rect 1640 -25120 1840 -24980
rect 2060 -25240 2260 -24980
rect -140 -25340 200 -25240
rect 1920 -25340 2260 -25240
rect -140 -25390 60 -25340
rect -140 -25450 -70 -25390
rect -10 -25450 60 -25390
rect -140 -25620 60 -25450
rect 2060 -25390 2260 -25340
rect 2060 -25450 2130 -25390
rect 2190 -25450 2260 -25390
rect 300 -25620 500 -25480
rect 960 -25620 1160 -25480
rect 1620 -25620 1820 -25480
rect 2060 -25620 2260 -25450
rect 4260 -25390 4460 -24980
rect 4260 -25450 4330 -25390
rect 4390 -25450 4460 -25390
rect 4260 -25620 4460 -25450
rect 6460 -25390 6660 -24980
rect 6460 -25450 6530 -25390
rect 6590 -25450 6660 -25390
rect 6460 -25620 6660 -25450
rect 8660 -25390 8860 -24980
rect 8660 -25450 8730 -25390
rect 8790 -25450 8860 -25390
rect 8660 -25620 8860 -25450
rect 10860 -25390 11060 -24980
rect 10860 -25450 10930 -25390
rect 10990 -25450 11060 -25390
rect 10860 -25620 11060 -25450
rect 13060 -25390 13260 -24980
rect 13060 -25450 13130 -25390
rect 13190 -25450 13260 -25390
rect 13060 -25620 13260 -25450
rect 15260 -25390 15460 -24980
rect 15260 -25450 15330 -25390
rect 15390 -25450 15460 -25390
rect 15260 -25620 15460 -25450
rect 17460 -25390 17660 -24980
rect 17460 -25450 17530 -25390
rect 17590 -25450 17660 -25390
rect 17460 -25620 17660 -25450
rect 19660 -25240 19860 -24980
rect 20100 -25120 20300 -24980
rect 20760 -25120 20960 -24980
rect 21440 -25120 21640 -24980
rect 21860 -25240 22060 -24980
rect 19660 -25340 20000 -25240
rect 21720 -25340 22060 -25240
rect 19660 -25390 19860 -25340
rect 19660 -25450 19730 -25390
rect 19790 -25450 19860 -25390
rect 19660 -25620 19860 -25450
rect 21860 -25390 22060 -25340
rect 21860 -25450 21930 -25390
rect 21990 -25450 22060 -25390
rect 20100 -25620 20300 -25480
rect 20760 -25620 20960 -25480
rect 21420 -25620 21620 -25480
rect 21860 -25620 22060 -25450
rect -140 -25780 22060 -25620
rect -140 -26040 60 -25780
rect 300 -25920 500 -25780
rect 960 -25920 1160 -25780
rect 1640 -25920 1840 -25780
rect 2060 -26040 2260 -25780
rect -140 -26140 200 -26040
rect 1920 -26140 2260 -26040
rect -140 -26190 60 -26140
rect -140 -26250 -70 -26190
rect -10 -26250 60 -26190
rect -140 -26420 60 -26250
rect 2060 -26190 2260 -26140
rect 2060 -26250 2130 -26190
rect 2190 -26250 2260 -26190
rect 300 -26420 500 -26280
rect 960 -26420 1160 -26280
rect 1620 -26420 1820 -26280
rect 2060 -26420 2260 -26250
rect 4260 -26190 4460 -25780
rect 4260 -26250 4330 -26190
rect 4390 -26250 4460 -26190
rect 4260 -26420 4460 -26250
rect 6460 -26190 6660 -25780
rect 6460 -26250 6530 -26190
rect 6590 -26250 6660 -26190
rect 6460 -26420 6660 -26250
rect 8660 -26190 8860 -25780
rect 8660 -26250 8730 -26190
rect 8790 -26250 8860 -26190
rect 8660 -26420 8860 -26250
rect 10860 -26190 11060 -25780
rect 10860 -26250 10930 -26190
rect 10990 -26250 11060 -26190
rect 10860 -26420 11060 -26250
rect 13060 -26190 13260 -25780
rect 13060 -26250 13130 -26190
rect 13190 -26250 13260 -26190
rect 13060 -26420 13260 -26250
rect 15260 -26190 15460 -25780
rect 15260 -26250 15330 -26190
rect 15390 -26250 15460 -26190
rect 15260 -26420 15460 -26250
rect 17460 -26190 17660 -25780
rect 17460 -26250 17530 -26190
rect 17590 -26250 17660 -26190
rect 17460 -26420 17660 -26250
rect 19660 -26040 19860 -25780
rect 20100 -25920 20300 -25780
rect 20760 -25920 20960 -25780
rect 21440 -25920 21640 -25780
rect 21860 -26040 22060 -25780
rect 19660 -26140 20000 -26040
rect 21720 -26140 22060 -26040
rect 19660 -26190 19860 -26140
rect 19660 -26250 19730 -26190
rect 19790 -26250 19860 -26190
rect 19660 -26420 19860 -26250
rect 21860 -26190 22060 -26140
rect 21860 -26250 21930 -26190
rect 21990 -26250 22060 -26190
rect 20100 -26420 20300 -26280
rect 20760 -26420 20960 -26280
rect 21420 -26420 21620 -26280
rect 21860 -26420 22060 -26250
rect -140 -26580 22060 -26420
rect -140 -26840 60 -26580
rect 300 -26720 500 -26580
rect 960 -26720 1160 -26580
rect 1640 -26720 1840 -26580
rect 2060 -26840 2260 -26580
rect -140 -26940 200 -26840
rect 1920 -26940 2260 -26840
rect -140 -26990 60 -26940
rect -140 -27050 -70 -26990
rect -10 -27050 60 -26990
rect -140 -27220 60 -27050
rect 2060 -26990 2260 -26940
rect 2060 -27050 2130 -26990
rect 2190 -27050 2260 -26990
rect 300 -27220 500 -27080
rect 960 -27220 1160 -27080
rect 1620 -27220 1820 -27080
rect 2060 -27220 2260 -27050
rect 4260 -26990 4460 -26580
rect 4260 -27050 4330 -26990
rect 4390 -27050 4460 -26990
rect 4260 -27220 4460 -27050
rect 6460 -26990 6660 -26580
rect 6460 -27050 6530 -26990
rect 6590 -27050 6660 -26990
rect 6460 -27220 6660 -27050
rect 8660 -26990 8860 -26580
rect 8660 -27050 8730 -26990
rect 8790 -27050 8860 -26990
rect 8660 -27220 8860 -27050
rect 10860 -26990 11060 -26580
rect 10860 -27050 10930 -26990
rect 10990 -27050 11060 -26990
rect 10860 -27220 11060 -27050
rect 13060 -26990 13260 -26580
rect 13060 -27050 13130 -26990
rect 13190 -27050 13260 -26990
rect 13060 -27220 13260 -27050
rect 15260 -26990 15460 -26580
rect 15260 -27050 15330 -26990
rect 15390 -27050 15460 -26990
rect 15260 -27220 15460 -27050
rect 17460 -26990 17660 -26580
rect 17460 -27050 17530 -26990
rect 17590 -27050 17660 -26990
rect 17460 -27220 17660 -27050
rect 19660 -26840 19860 -26580
rect 20100 -26720 20300 -26580
rect 20760 -26720 20960 -26580
rect 21440 -26720 21640 -26580
rect 21860 -26840 22060 -26580
rect 19660 -26940 20000 -26840
rect 21720 -26940 22060 -26840
rect 19660 -26990 19860 -26940
rect 19660 -27050 19730 -26990
rect 19790 -27050 19860 -26990
rect 19660 -27220 19860 -27050
rect 21860 -26990 22060 -26940
rect 21860 -27050 21930 -26990
rect 21990 -27050 22060 -26990
rect 20100 -27220 20300 -27080
rect 20760 -27220 20960 -27080
rect 21420 -27220 21620 -27080
rect 21860 -27220 22060 -27050
rect -140 -27380 22060 -27220
rect -140 -27640 60 -27380
rect 300 -27520 500 -27380
rect 960 -27520 1160 -27380
rect 1640 -27520 1840 -27380
rect 2060 -27640 2260 -27380
rect -140 -27740 200 -27640
rect 1920 -27740 2260 -27640
rect -140 -27790 60 -27740
rect -140 -27850 -70 -27790
rect -10 -27850 60 -27790
rect -140 -28020 60 -27850
rect 2060 -27790 2260 -27740
rect 2060 -27850 2130 -27790
rect 2190 -27850 2260 -27790
rect 300 -28020 500 -27880
rect 960 -28020 1160 -27880
rect 1620 -28020 1820 -27880
rect 2060 -28020 2260 -27850
rect 4260 -27790 4460 -27380
rect 4260 -27850 4330 -27790
rect 4390 -27850 4460 -27790
rect 4260 -28020 4460 -27850
rect 6460 -27790 6660 -27380
rect 6460 -27850 6530 -27790
rect 6590 -27850 6660 -27790
rect 6460 -28020 6660 -27850
rect 8660 -27790 8860 -27380
rect 8660 -27850 8730 -27790
rect 8790 -27850 8860 -27790
rect 8660 -28020 8860 -27850
rect 10860 -27790 11060 -27380
rect 10860 -27850 10930 -27790
rect 10990 -27850 11060 -27790
rect 10860 -28020 11060 -27850
rect 13060 -27790 13260 -27380
rect 13060 -27850 13130 -27790
rect 13190 -27850 13260 -27790
rect 13060 -28020 13260 -27850
rect 15260 -27790 15460 -27380
rect 15260 -27850 15330 -27790
rect 15390 -27850 15460 -27790
rect 15260 -28020 15460 -27850
rect 17460 -27790 17660 -27380
rect 17460 -27850 17530 -27790
rect 17590 -27850 17660 -27790
rect 17460 -28020 17660 -27850
rect 19660 -27640 19860 -27380
rect 20100 -27520 20300 -27380
rect 20760 -27520 20960 -27380
rect 21440 -27520 21640 -27380
rect 21860 -27640 22060 -27380
rect 19660 -27740 20000 -27640
rect 21720 -27740 22060 -27640
rect 19660 -27790 19860 -27740
rect 19660 -27850 19730 -27790
rect 19790 -27850 19860 -27790
rect 19660 -28020 19860 -27850
rect 21860 -27790 22060 -27740
rect 21860 -27850 21930 -27790
rect 21990 -27850 22060 -27790
rect 20100 -28020 20300 -27880
rect 20760 -28020 20960 -27880
rect 21420 -28020 21620 -27880
rect 21860 -28020 22060 -27850
rect -140 -28180 22060 -28020
rect -140 -28440 60 -28180
rect 300 -28320 500 -28180
rect 960 -28320 1160 -28180
rect 1640 -28320 1840 -28180
rect 2060 -28440 2260 -28180
rect -140 -28540 200 -28440
rect 1920 -28540 2260 -28440
rect -140 -28590 60 -28540
rect -140 -28650 -70 -28590
rect -10 -28650 60 -28590
rect -140 -28820 60 -28650
rect 2060 -28590 2260 -28540
rect 2060 -28650 2130 -28590
rect 2190 -28650 2260 -28590
rect 300 -28820 500 -28680
rect 960 -28820 1160 -28680
rect 1620 -28820 1820 -28680
rect 2060 -28820 2260 -28650
rect 4260 -28590 4460 -28180
rect 4260 -28650 4330 -28590
rect 4390 -28650 4460 -28590
rect 4260 -28820 4460 -28650
rect 6460 -28590 6660 -28180
rect 6460 -28650 6530 -28590
rect 6590 -28650 6660 -28590
rect 6460 -28820 6660 -28650
rect 8660 -28590 8860 -28180
rect 8660 -28650 8730 -28590
rect 8790 -28650 8860 -28590
rect 8660 -28820 8860 -28650
rect 10860 -28590 11060 -28180
rect 10860 -28650 10930 -28590
rect 10990 -28650 11060 -28590
rect 10860 -28820 11060 -28650
rect 13060 -28590 13260 -28180
rect 13060 -28650 13130 -28590
rect 13190 -28650 13260 -28590
rect 13060 -28820 13260 -28650
rect 15260 -28590 15460 -28180
rect 15260 -28650 15330 -28590
rect 15390 -28650 15460 -28590
rect 15260 -28820 15460 -28650
rect 17460 -28590 17660 -28180
rect 17460 -28650 17530 -28590
rect 17590 -28650 17660 -28590
rect 17460 -28820 17660 -28650
rect 19660 -28440 19860 -28180
rect 20100 -28320 20300 -28180
rect 20760 -28320 20960 -28180
rect 21440 -28320 21640 -28180
rect 21860 -28440 22060 -28180
rect 19660 -28540 20000 -28440
rect 21720 -28540 22060 -28440
rect 19660 -28590 19860 -28540
rect 19660 -28650 19730 -28590
rect 19790 -28650 19860 -28590
rect 19660 -28820 19860 -28650
rect 21860 -28590 22060 -28540
rect 21860 -28650 21930 -28590
rect 21990 -28650 22060 -28590
rect 20100 -28820 20300 -28680
rect 20760 -28820 20960 -28680
rect 21420 -28820 21620 -28680
rect 21860 -28820 22060 -28650
rect -140 -28980 22060 -28820
rect -140 -29240 60 -28980
rect 300 -29120 500 -28980
rect 960 -29120 1160 -28980
rect 1640 -29120 1840 -28980
rect 2060 -29240 2260 -28980
rect -140 -29340 200 -29240
rect 1920 -29340 2260 -29240
rect -140 -29390 60 -29340
rect -140 -29450 -70 -29390
rect -10 -29450 60 -29390
rect -140 -29620 60 -29450
rect 2060 -29390 2260 -29340
rect 2060 -29450 2130 -29390
rect 2190 -29450 2260 -29390
rect 300 -29620 500 -29480
rect 960 -29620 1160 -29480
rect 1620 -29620 1820 -29480
rect 2060 -29620 2260 -29450
rect 4260 -29390 4460 -28980
rect 4260 -29450 4330 -29390
rect 4390 -29450 4460 -29390
rect 4260 -29620 4460 -29450
rect 6460 -29390 6660 -28980
rect 6460 -29450 6530 -29390
rect 6590 -29450 6660 -29390
rect 6460 -29620 6660 -29450
rect 8660 -29390 8860 -28980
rect 8660 -29450 8730 -29390
rect 8790 -29450 8860 -29390
rect 8660 -29620 8860 -29450
rect 10860 -29390 11060 -28980
rect 10860 -29450 10930 -29390
rect 10990 -29450 11060 -29390
rect 10860 -29620 11060 -29450
rect 13060 -29390 13260 -28980
rect 13060 -29450 13130 -29390
rect 13190 -29450 13260 -29390
rect 13060 -29620 13260 -29450
rect 15260 -29390 15460 -28980
rect 15260 -29450 15330 -29390
rect 15390 -29450 15460 -29390
rect 15260 -29620 15460 -29450
rect 17460 -29390 17660 -28980
rect 17460 -29450 17530 -29390
rect 17590 -29450 17660 -29390
rect 17460 -29620 17660 -29450
rect 19660 -29240 19860 -28980
rect 20100 -29120 20300 -28980
rect 20760 -29120 20960 -28980
rect 21440 -29120 21640 -28980
rect 21860 -29240 22060 -28980
rect 19660 -29340 20000 -29240
rect 21720 -29340 22060 -29240
rect 19660 -29390 19860 -29340
rect 19660 -29450 19730 -29390
rect 19790 -29450 19860 -29390
rect 19660 -29620 19860 -29450
rect 21860 -29390 22060 -29340
rect 21860 -29450 21930 -29390
rect 21990 -29450 22060 -29390
rect 20100 -29620 20300 -29480
rect 20760 -29620 20960 -29480
rect 21420 -29620 21620 -29480
rect 21860 -29620 22060 -29450
rect -140 -29780 22060 -29620
rect -140 -30040 60 -29780
rect 300 -29920 500 -29780
rect 960 -29920 1160 -29780
rect 1640 -29920 1840 -29780
rect 2060 -30040 2260 -29780
rect -140 -30140 200 -30040
rect 1920 -30140 2260 -30040
rect -140 -30190 60 -30140
rect -140 -30250 -70 -30190
rect -10 -30250 60 -30190
rect -140 -30420 60 -30250
rect 2060 -30190 2260 -30140
rect 2060 -30250 2130 -30190
rect 2190 -30250 2260 -30190
rect 300 -30420 500 -30280
rect 960 -30420 1160 -30280
rect 1620 -30420 1820 -30280
rect 2060 -30420 2260 -30250
rect 4260 -30190 4460 -29780
rect 4260 -30250 4330 -30190
rect 4390 -30250 4460 -30190
rect 4260 -30420 4460 -30250
rect 6460 -30190 6660 -29780
rect 6460 -30250 6530 -30190
rect 6590 -30250 6660 -30190
rect 6460 -30420 6660 -30250
rect 8660 -30190 8860 -29780
rect 8660 -30250 8730 -30190
rect 8790 -30250 8860 -30190
rect 8660 -30420 8860 -30250
rect 10860 -30190 11060 -29780
rect 10860 -30250 10930 -30190
rect 10990 -30250 11060 -30190
rect 10860 -30420 11060 -30250
rect 13060 -30190 13260 -29780
rect 13060 -30250 13130 -30190
rect 13190 -30250 13260 -30190
rect 13060 -30420 13260 -30250
rect 15260 -30190 15460 -29780
rect 15260 -30250 15330 -30190
rect 15390 -30250 15460 -30190
rect 15260 -30420 15460 -30250
rect 17460 -30190 17660 -29780
rect 17460 -30250 17530 -30190
rect 17590 -30250 17660 -30190
rect 17460 -30420 17660 -30250
rect 19660 -30040 19860 -29780
rect 20100 -29920 20300 -29780
rect 20760 -29920 20960 -29780
rect 21440 -29920 21640 -29780
rect 21860 -30040 22060 -29780
rect 19660 -30140 20000 -30040
rect 21720 -30140 22060 -30040
rect 19660 -30190 19860 -30140
rect 19660 -30250 19730 -30190
rect 19790 -30250 19860 -30190
rect 19660 -30420 19860 -30250
rect 21860 -30190 22060 -30140
rect 21860 -30250 21930 -30190
rect 21990 -30250 22060 -30190
rect 20100 -30420 20300 -30280
rect 20760 -30420 20960 -30280
rect 21420 -30420 21620 -30280
rect 21860 -30420 22060 -30250
rect -140 -30580 22060 -30420
rect -140 -30840 60 -30580
rect 300 -30720 500 -30580
rect 960 -30720 1160 -30580
rect 1640 -30720 1840 -30580
rect 2060 -30840 2260 -30580
rect -140 -30940 200 -30840
rect 1920 -30940 2260 -30840
rect -140 -30990 60 -30940
rect -140 -31050 -70 -30990
rect -10 -31050 60 -30990
rect -140 -31220 60 -31050
rect 2060 -30990 2260 -30940
rect 2060 -31050 2130 -30990
rect 2190 -31050 2260 -30990
rect 300 -31220 500 -31080
rect 960 -31220 1160 -31080
rect 1620 -31220 1820 -31080
rect 2060 -31220 2260 -31050
rect 4260 -30990 4460 -30580
rect 4260 -31050 4330 -30990
rect 4390 -31050 4460 -30990
rect 4260 -31220 4460 -31050
rect 6460 -30990 6660 -30580
rect 6460 -31050 6530 -30990
rect 6590 -31050 6660 -30990
rect 6460 -31220 6660 -31050
rect 8660 -30990 8860 -30580
rect 8660 -31050 8730 -30990
rect 8790 -31050 8860 -30990
rect 8660 -31220 8860 -31050
rect 10860 -30990 11060 -30580
rect 10860 -31050 10930 -30990
rect 10990 -31050 11060 -30990
rect 10860 -31220 11060 -31050
rect 13060 -30990 13260 -30580
rect 13060 -31050 13130 -30990
rect 13190 -31050 13260 -30990
rect 13060 -31220 13260 -31050
rect 15260 -30990 15460 -30580
rect 15260 -31050 15330 -30990
rect 15390 -31050 15460 -30990
rect 15260 -31220 15460 -31050
rect 17460 -30990 17660 -30580
rect 17460 -31050 17530 -30990
rect 17590 -31050 17660 -30990
rect 17460 -31220 17660 -31050
rect 19660 -30840 19860 -30580
rect 20100 -30720 20300 -30580
rect 20760 -30720 20960 -30580
rect 21440 -30720 21640 -30580
rect 21860 -30840 22060 -30580
rect 19660 -30940 20000 -30840
rect 21720 -30940 22060 -30840
rect 19660 -30990 19860 -30940
rect 19660 -31050 19730 -30990
rect 19790 -31050 19860 -30990
rect 19660 -31220 19860 -31050
rect 21860 -30990 22060 -30940
rect 21860 -31050 21930 -30990
rect 21990 -31050 22060 -30990
rect 20100 -31220 20300 -31080
rect 20760 -31220 20960 -31080
rect 21420 -31220 21620 -31080
rect 21860 -31220 22060 -31050
rect -140 -31380 22060 -31220
rect -140 -31640 60 -31380
rect 300 -31520 500 -31380
rect 960 -31520 1160 -31380
rect 1640 -31520 1840 -31380
rect 2060 -31640 2260 -31380
rect 2500 -31520 2700 -31380
rect 3160 -31520 3360 -31380
rect 3840 -31520 4040 -31380
rect 4260 -31640 4460 -31380
rect 4700 -31520 4900 -31380
rect 5360 -31520 5560 -31380
rect 6040 -31520 6240 -31380
rect 6460 -31640 6660 -31380
rect 6900 -31520 7100 -31380
rect 7560 -31520 7760 -31380
rect 8240 -31520 8440 -31380
rect 8660 -31640 8860 -31380
rect 9100 -31520 9300 -31380
rect 9760 -31520 9960 -31380
rect 10440 -31520 10640 -31380
rect 10860 -31640 11060 -31380
rect 11300 -31520 11500 -31380
rect 11960 -31520 12160 -31380
rect 12640 -31520 12840 -31380
rect 13060 -31640 13260 -31380
rect 13500 -31520 13700 -31380
rect 14160 -31520 14360 -31380
rect 14840 -31520 15040 -31380
rect 15260 -31640 15460 -31380
rect 15700 -31520 15900 -31380
rect 16360 -31520 16560 -31380
rect 17040 -31520 17240 -31380
rect 17460 -31640 17660 -31380
rect 17900 -31520 18100 -31380
rect 18560 -31520 18760 -31380
rect 19240 -31520 19440 -31380
rect 19660 -31640 19860 -31380
rect 20100 -31520 20300 -31380
rect 20760 -31520 20960 -31380
rect 21440 -31520 21640 -31380
rect 21860 -31640 22060 -31380
rect -140 -31740 200 -31640
rect 1920 -31740 2400 -31640
rect 4120 -31740 4600 -31640
rect 6320 -31740 6800 -31640
rect 8520 -31740 9000 -31640
rect 10720 -31740 11200 -31640
rect 12920 -31740 13400 -31640
rect 15120 -31740 15600 -31640
rect 17320 -31740 17800 -31640
rect 19520 -31740 20000 -31640
rect 21720 -31740 22060 -31640
rect -140 -32020 60 -31740
rect 300 -32020 500 -31880
rect 960 -32020 1160 -31880
rect 1620 -32020 1820 -31880
rect 2060 -32020 2260 -31740
rect 2500 -32020 2700 -31880
rect 3160 -32020 3360 -31880
rect 3820 -32020 4020 -31880
rect 4260 -32020 4460 -31740
rect 4700 -32020 4900 -31880
rect 5360 -32020 5560 -31880
rect 6020 -32020 6220 -31880
rect 6460 -32020 6660 -31740
rect 6900 -32020 7100 -31880
rect 7560 -32020 7760 -31880
rect 8220 -32020 8420 -31880
rect 8660 -32020 8860 -31740
rect 9100 -32020 9300 -31880
rect 9760 -32020 9960 -31880
rect 10420 -32020 10620 -31880
rect 10860 -32020 11060 -31740
rect 11300 -32020 11500 -31880
rect 11960 -32020 12160 -31880
rect 12620 -32020 12820 -31880
rect 13060 -32020 13260 -31740
rect 13500 -32020 13700 -31880
rect 14160 -32020 14360 -31880
rect 14820 -32020 15020 -31880
rect 15260 -32020 15460 -31740
rect 15700 -32020 15900 -31880
rect 16360 -32020 16560 -31880
rect 17020 -32020 17220 -31880
rect 17460 -32020 17660 -31740
rect 17900 -32020 18100 -31880
rect 18560 -32020 18760 -31880
rect 19220 -32020 19420 -31880
rect 19660 -32020 19860 -31740
rect 20100 -32020 20300 -31880
rect 20760 -32020 20960 -31880
rect 21420 -32020 21620 -31880
rect 21860 -32020 22060 -31740
rect -140 -32180 22060 -32020
<< viali >>
rect -70 10870 -10 10930
rect 2130 10870 2190 10930
rect 4330 10870 4390 10930
rect 6530 10870 6590 10930
rect 8730 10870 8790 10930
rect 10930 10870 10990 10930
rect 13130 10870 13190 10930
rect 15330 10870 15390 10930
rect 17530 10870 17590 10930
rect 19730 10870 19790 10930
rect 21930 10870 21990 10930
rect -70 10070 -10 10130
rect 2130 10070 2190 10130
rect 4330 10070 4390 10130
rect 6530 10070 6590 10130
rect 8730 10070 8790 10130
rect 10930 10070 10990 10130
rect 13130 10070 13190 10130
rect 15330 10070 15390 10130
rect 17530 10070 17590 10130
rect 19730 10070 19790 10130
rect 21930 10070 21990 10130
rect -70 9270 -10 9330
rect 2130 9270 2190 9330
rect 4330 9270 4390 9330
rect 6530 9270 6590 9330
rect 8730 9270 8790 9330
rect 10930 9270 10990 9330
rect 13130 9270 13190 9330
rect 15330 9270 15390 9330
rect 17530 9270 17590 9330
rect 19730 9270 19790 9330
rect 21930 9270 21990 9330
rect -70 8470 -10 8530
rect 2130 8470 2190 8530
rect 4330 8470 4390 8530
rect 6530 8470 6590 8530
rect 8730 8470 8790 8530
rect 10930 8470 10990 8530
rect 13130 8470 13190 8530
rect 15330 8470 15390 8530
rect 17530 8470 17590 8530
rect 19730 8470 19790 8530
rect 21930 8470 21990 8530
rect -70 7670 -10 7730
rect 2130 7670 2190 7730
rect 4330 7670 4390 7730
rect 6530 7670 6590 7730
rect 8730 7670 8790 7730
rect 10930 7670 10990 7730
rect 13130 7670 13190 7730
rect 15330 7670 15390 7730
rect 17530 7670 17590 7730
rect 19730 7670 19790 7730
rect 21930 7670 21990 7730
rect -70 6870 -10 6930
rect 2130 6870 2190 6930
rect 4330 6870 4390 6930
rect 6530 6870 6590 6930
rect 8730 6870 8790 6930
rect 10930 6870 10990 6930
rect 13130 6870 13190 6930
rect 15330 6870 15390 6930
rect 17530 6870 17590 6930
rect 19730 6870 19790 6930
rect 21930 6870 21990 6930
rect -70 6070 -10 6130
rect 2130 6070 2190 6130
rect 4330 6070 4390 6130
rect 6530 6070 6590 6130
rect 8730 6070 8790 6130
rect 10930 6070 10990 6130
rect 13130 6070 13190 6130
rect 15330 6070 15390 6130
rect 17530 6070 17590 6130
rect 19730 6070 19790 6130
rect 21930 6070 21990 6130
rect -70 5270 -10 5330
rect 2130 5270 2190 5330
rect 4330 5270 4390 5330
rect 6530 5270 6590 5330
rect 8730 5270 8790 5330
rect 10930 5270 10990 5330
rect 13130 5270 13190 5330
rect 15330 5270 15390 5330
rect 17530 5270 17590 5330
rect 19730 5270 19790 5330
rect 21930 5270 21990 5330
rect -70 -25450 -10 -25390
rect 2130 -25450 2190 -25390
rect 4330 -25450 4390 -25390
rect 6530 -25450 6590 -25390
rect 8730 -25450 8790 -25390
rect 10930 -25450 10990 -25390
rect 13130 -25450 13190 -25390
rect 15330 -25450 15390 -25390
rect 17530 -25450 17590 -25390
rect 19730 -25450 19790 -25390
rect 21930 -25450 21990 -25390
rect -70 -26250 -10 -26190
rect 2130 -26250 2190 -26190
rect 4330 -26250 4390 -26190
rect 6530 -26250 6590 -26190
rect 8730 -26250 8790 -26190
rect 10930 -26250 10990 -26190
rect 13130 -26250 13190 -26190
rect 15330 -26250 15390 -26190
rect 17530 -26250 17590 -26190
rect 19730 -26250 19790 -26190
rect 21930 -26250 21990 -26190
rect -70 -27050 -10 -26990
rect 2130 -27050 2190 -26990
rect 4330 -27050 4390 -26990
rect 6530 -27050 6590 -26990
rect 8730 -27050 8790 -26990
rect 10930 -27050 10990 -26990
rect 13130 -27050 13190 -26990
rect 15330 -27050 15390 -26990
rect 17530 -27050 17590 -26990
rect 19730 -27050 19790 -26990
rect 21930 -27050 21990 -26990
rect -70 -27850 -10 -27790
rect 2130 -27850 2190 -27790
rect 4330 -27850 4390 -27790
rect 6530 -27850 6590 -27790
rect 8730 -27850 8790 -27790
rect 10930 -27850 10990 -27790
rect 13130 -27850 13190 -27790
rect 15330 -27850 15390 -27790
rect 17530 -27850 17590 -27790
rect 19730 -27850 19790 -27790
rect 21930 -27850 21990 -27790
rect -70 -28650 -10 -28590
rect 2130 -28650 2190 -28590
rect 4330 -28650 4390 -28590
rect 6530 -28650 6590 -28590
rect 8730 -28650 8790 -28590
rect 10930 -28650 10990 -28590
rect 13130 -28650 13190 -28590
rect 15330 -28650 15390 -28590
rect 17530 -28650 17590 -28590
rect 19730 -28650 19790 -28590
rect 21930 -28650 21990 -28590
rect -70 -29450 -10 -29390
rect 2130 -29450 2190 -29390
rect 4330 -29450 4390 -29390
rect 6530 -29450 6590 -29390
rect 8730 -29450 8790 -29390
rect 10930 -29450 10990 -29390
rect 13130 -29450 13190 -29390
rect 15330 -29450 15390 -29390
rect 17530 -29450 17590 -29390
rect 19730 -29450 19790 -29390
rect 21930 -29450 21990 -29390
rect -70 -30250 -10 -30190
rect 2130 -30250 2190 -30190
rect 4330 -30250 4390 -30190
rect 6530 -30250 6590 -30190
rect 8730 -30250 8790 -30190
rect 10930 -30250 10990 -30190
rect 13130 -30250 13190 -30190
rect 15330 -30250 15390 -30190
rect 17530 -30250 17590 -30190
rect 19730 -30250 19790 -30190
rect 21930 -30250 21990 -30190
rect -70 -31050 -10 -30990
rect 2130 -31050 2190 -30990
rect 4330 -31050 4390 -30990
rect 6530 -31050 6590 -30990
rect 8730 -31050 8790 -30990
rect 10930 -31050 10990 -30990
rect 13130 -31050 13190 -30990
rect 15330 -31050 15390 -30990
rect 17530 -31050 17590 -30990
rect 19730 -31050 19790 -30990
rect 21930 -31050 21990 -30990
<< metal1 >>
rect 2500 11180 2510 11240
rect 2690 11180 2700 11240
rect 2500 10940 2700 11180
rect 3160 11180 3170 11240
rect 3350 11180 3360 11240
rect 3160 10940 3360 11180
rect 3820 11180 3830 11240
rect 4010 11180 4020 11240
rect 3820 10940 4020 11180
rect 4700 11180 4710 11240
rect 4890 11180 4900 11240
rect 4700 10940 4900 11180
rect 5360 11180 5370 11240
rect 5550 11180 5560 11240
rect 5360 10940 5560 11180
rect 6020 11180 6030 11240
rect 6210 11180 6220 11240
rect 6020 10940 6220 11180
rect 6900 11100 7100 11240
rect 6900 11040 6910 11100
rect 7090 11040 7100 11100
rect 6900 10940 7100 11040
rect 7560 11100 7760 11240
rect 7560 11040 7570 11100
rect 7750 11040 7760 11100
rect 7560 10940 7760 11040
rect 8220 11100 8420 11240
rect 8220 11040 8230 11100
rect 8410 11040 8420 11100
rect 8220 10940 8420 11040
rect 9100 11100 9300 11240
rect 9100 11040 9110 11100
rect 9290 11040 9300 11100
rect 9100 10940 9300 11040
rect 9760 11100 9960 11240
rect 9760 11040 9770 11100
rect 9950 11040 9960 11100
rect 9760 10940 9960 11040
rect 10420 11100 10620 11240
rect 10420 11040 10430 11100
rect 10610 11040 10620 11100
rect 10420 10940 10620 11040
rect 11300 11100 11500 11240
rect 11300 11040 11310 11100
rect 11490 11040 11500 11100
rect 11300 10940 11500 11040
rect 11960 11100 12160 11240
rect 11960 11040 11970 11100
rect 12150 11040 12160 11100
rect 11960 10940 12160 11040
rect 12620 11100 12820 11240
rect 12620 11040 12630 11100
rect 12810 11040 12820 11100
rect 12620 10940 12820 11040
rect 13500 11100 13700 11240
rect 13500 11040 13510 11100
rect 13690 11040 13700 11100
rect 13500 10940 13700 11040
rect 14160 11100 14360 11240
rect 14160 11040 14170 11100
rect 14350 11040 14360 11100
rect 14160 10940 14360 11040
rect 14820 11100 15020 11240
rect 14820 11040 14830 11100
rect 15010 11040 15020 11100
rect 14820 10940 15020 11040
rect 15700 11180 15710 11240
rect 15890 11180 15900 11240
rect 15700 10940 15900 11180
rect 16360 11180 16370 11240
rect 16550 11180 16560 11240
rect 16360 10940 16560 11180
rect 17020 11180 17030 11240
rect 17210 11180 17220 11240
rect 17020 10940 17220 11180
rect 17900 11180 17910 11240
rect 18090 11180 18100 11240
rect 17900 10940 18100 11180
rect 18560 11180 18570 11240
rect 18750 11180 18760 11240
rect 18560 10940 18760 11180
rect 19220 11180 19230 11240
rect 19410 11180 19420 11240
rect 19220 10940 19420 11180
rect -90 10930 10 10940
rect -90 10870 -70 10930
rect -10 10870 10 10930
rect -90 10860 10 10870
rect 2110 10930 2210 10940
rect 2110 10870 2130 10930
rect 2190 10870 2210 10930
rect 2110 10860 2210 10870
rect 4310 10930 4410 10940
rect 4310 10870 4330 10930
rect 4390 10870 4410 10930
rect 4310 10860 4410 10870
rect 6510 10930 6610 10940
rect 6510 10870 6530 10930
rect 6590 10870 6610 10930
rect 6510 10860 6610 10870
rect 8710 10930 8810 10940
rect 8710 10870 8730 10930
rect 8790 10870 8810 10930
rect 8710 10860 8810 10870
rect 10910 10930 11010 10940
rect 10910 10870 10930 10930
rect 10990 10870 11010 10930
rect 10910 10860 11010 10870
rect 13110 10930 13210 10940
rect 13110 10870 13130 10930
rect 13190 10870 13210 10930
rect 13110 10860 13210 10870
rect 15310 10930 15410 10940
rect 15310 10870 15330 10930
rect 15390 10870 15410 10930
rect 15310 10860 15410 10870
rect 17510 10930 17610 10940
rect 17510 10870 17530 10930
rect 17590 10870 17610 10930
rect 17510 10860 17610 10870
rect 19710 10930 19810 10940
rect 19710 10870 19730 10930
rect 19790 10870 19810 10930
rect 19710 10860 19810 10870
rect 21910 10930 22010 10940
rect 21910 10870 21930 10930
rect 21990 10870 22010 10930
rect 21910 10860 22010 10870
rect 1900 10760 2310 10820
rect 4100 10760 4220 10820
rect 4280 10760 4510 10820
rect 6300 10760 6420 10820
rect 6480 10760 6710 10820
rect 8500 10760 8840 10820
rect 8900 10760 8910 10820
rect 10700 10760 11040 10820
rect 11100 10760 11110 10820
rect 12900 10760 13240 10820
rect 13300 10760 13310 10820
rect 15100 10760 15440 10820
rect 15500 10760 15510 10820
rect 17300 10760 17420 10820
rect 17480 10760 17710 10820
rect 22770 10810 23330 11120
rect 19500 10740 19620 10800
rect 19680 10740 19910 10800
rect 2010 10650 2020 10710
rect 2080 10650 2420 10710
rect 4210 10650 4220 10710
rect 4280 10650 4620 10710
rect 6410 10650 6640 10710
rect 6700 10650 6820 10710
rect 8610 10650 8840 10710
rect 8900 10650 9020 10710
rect 10810 10650 11040 10710
rect 11100 10650 11220 10710
rect 13010 10650 13240 10710
rect 13300 10650 13420 10710
rect 15210 10650 15220 10710
rect 15280 10650 15620 10710
rect 17410 10650 17420 10710
rect 17480 10650 17820 10710
rect 19610 10650 20020 10710
rect 2500 10610 4020 10620
rect 2500 10550 2510 10610
rect 4010 10550 4020 10610
rect 2500 10540 4020 10550
rect 4700 10610 6220 10622
rect 4700 10550 4710 10610
rect 6210 10550 6220 10610
rect 4700 10540 6220 10550
rect 6900 10610 8420 10622
rect 6900 10550 6910 10610
rect 8410 10550 8420 10610
rect 6900 10540 8420 10550
rect 9100 10610 10620 10622
rect 9100 10550 9110 10610
rect 10610 10550 10620 10610
rect 9100 10540 10620 10550
rect 11300 10610 12820 10622
rect 11300 10550 11310 10610
rect 12810 10550 12820 10610
rect 11300 10540 12820 10550
rect 13500 10610 15020 10622
rect 13500 10550 13510 10610
rect 15010 10550 15020 10610
rect 13500 10540 15020 10550
rect 15700 10610 17220 10622
rect 15700 10550 15710 10610
rect 17210 10550 17220 10610
rect 15700 10540 17220 10550
rect 17900 10610 19420 10622
rect 17900 10550 17910 10610
rect 19410 10550 19420 10610
rect 22630 10570 23330 10810
rect 23440 10570 24660 10970
rect 24770 10570 25990 10970
rect 26100 10570 27320 10970
rect 28100 10810 28660 11120
rect 30309 10912 30387 10913
rect 30467 10912 30545 10913
rect 30625 10912 30703 10913
rect 30783 10912 30861 10913
rect 29270 10868 29820 10912
rect 30309 10868 30861 10912
rect 30309 10867 30387 10868
rect 30467 10867 30545 10868
rect 30625 10867 30703 10868
rect 30783 10867 30861 10868
rect 31349 10912 31427 10913
rect 31507 10912 31585 10913
rect 31665 10912 31743 10913
rect 31823 10912 31901 10913
rect 31349 10868 31901 10912
rect 31349 10867 31427 10868
rect 31507 10867 31585 10868
rect 31665 10867 31743 10868
rect 31823 10867 31901 10868
rect 28100 10570 28790 10810
rect 17900 10540 19420 10550
rect 2500 10300 2700 10440
rect 2500 10240 2510 10300
rect 2690 10240 2700 10300
rect 2500 10140 2700 10240
rect 3160 10300 3360 10440
rect 3160 10240 3170 10300
rect 3350 10240 3360 10300
rect 3160 10140 3360 10240
rect 3820 10300 4020 10440
rect 3820 10240 3830 10300
rect 4010 10240 4020 10300
rect 3820 10140 4020 10240
rect 4700 10300 4900 10440
rect 4700 10240 4710 10300
rect 4890 10240 4900 10300
rect 4700 10140 4900 10240
rect 5360 10300 5560 10440
rect 5360 10240 5370 10300
rect 5550 10240 5560 10300
rect 5360 10140 5560 10240
rect 6020 10300 6220 10440
rect 6020 10240 6030 10300
rect 6210 10240 6220 10300
rect 6020 10140 6220 10240
rect 6900 10380 6910 10440
rect 7090 10380 7100 10440
rect 6900 10140 7100 10380
rect 7560 10380 7570 10440
rect 7750 10380 7760 10440
rect 7560 10140 7760 10380
rect 8220 10380 8230 10440
rect 8410 10380 8420 10440
rect 8220 10140 8420 10380
rect 9100 10380 9110 10440
rect 9290 10380 9300 10440
rect 9100 10140 9300 10380
rect 9760 10380 9770 10440
rect 9950 10380 9960 10440
rect 9760 10140 9960 10380
rect 10420 10380 10430 10440
rect 10610 10380 10620 10440
rect 10420 10140 10620 10380
rect 11300 10380 11310 10440
rect 11490 10380 11500 10440
rect 11300 10140 11500 10380
rect 11960 10380 11970 10440
rect 12150 10380 12160 10440
rect 11960 10140 12160 10380
rect 12620 10380 12630 10440
rect 12810 10380 12820 10440
rect 12620 10140 12820 10380
rect 13500 10380 13510 10440
rect 13690 10380 13700 10440
rect 13500 10140 13700 10380
rect 14160 10380 14170 10440
rect 14350 10380 14360 10440
rect 14160 10140 14360 10380
rect 14820 10380 14830 10440
rect 15010 10380 15020 10440
rect 14820 10140 15020 10380
rect 15700 10300 15900 10440
rect 15700 10240 15710 10300
rect 15890 10240 15900 10300
rect 15700 10140 15900 10240
rect 16360 10300 16560 10440
rect 16360 10240 16370 10300
rect 16550 10240 16560 10300
rect 16360 10140 16560 10240
rect 17020 10300 17220 10440
rect 17020 10240 17030 10300
rect 17210 10240 17220 10300
rect 17020 10140 17220 10240
rect 17900 10300 18100 10440
rect 17900 10240 17910 10300
rect 18090 10240 18100 10300
rect 17900 10140 18100 10240
rect 18560 10300 18760 10440
rect 18560 10240 18570 10300
rect 18750 10240 18760 10300
rect 18560 10140 18760 10240
rect 19220 10300 19420 10440
rect 19220 10240 19230 10300
rect 19410 10240 19420 10300
rect 19220 10140 19420 10240
rect -90 10130 10 10140
rect -90 10070 -70 10130
rect -10 10070 10 10130
rect -90 10060 10 10070
rect 2110 10130 2210 10140
rect 2110 10070 2130 10130
rect 2190 10070 2210 10130
rect 2110 10060 2210 10070
rect 4310 10130 4410 10140
rect 4310 10070 4330 10130
rect 4390 10070 4410 10130
rect 4310 10060 4410 10070
rect 6510 10130 6610 10140
rect 6510 10070 6530 10130
rect 6590 10070 6610 10130
rect 6510 10060 6610 10070
rect 8710 10130 8810 10140
rect 8710 10070 8730 10130
rect 8790 10070 8810 10130
rect 8710 10060 8810 10070
rect 10910 10130 11010 10140
rect 10910 10070 10930 10130
rect 10990 10070 11010 10130
rect 10910 10060 11010 10070
rect 13110 10130 13210 10140
rect 13110 10070 13130 10130
rect 13190 10070 13210 10130
rect 13110 10060 13210 10070
rect 15310 10130 15410 10140
rect 15310 10070 15330 10130
rect 15390 10070 15410 10130
rect 15310 10060 15410 10070
rect 17510 10130 17610 10140
rect 17510 10070 17530 10130
rect 17590 10070 17610 10130
rect 17510 10060 17610 10070
rect 19710 10130 19810 10140
rect 19710 10070 19730 10130
rect 19790 10070 19810 10130
rect 19710 10060 19810 10070
rect 21910 10130 22010 10140
rect 21910 10070 21930 10130
rect 21990 10070 22010 10130
rect 21910 10060 22010 10070
rect 1900 9960 2310 10020
rect 4100 9960 4440 10020
rect 4500 9960 4510 10020
rect 6300 9960 6640 10020
rect 6700 9960 6710 10020
rect 8500 9960 8620 10020
rect 8680 9960 8910 10020
rect 10700 9960 10820 10020
rect 10880 9960 11110 10020
rect 12900 9960 13020 10020
rect 13080 9960 13310 10020
rect 15100 9960 15220 10020
rect 15280 9960 15510 10020
rect 17300 9960 17640 10020
rect 17700 9960 17710 10020
rect 19500 9940 19840 10000
rect 19900 9940 19910 10000
rect 2010 9850 2240 9910
rect 2300 9850 2420 9910
rect 4210 9850 4440 9910
rect 4500 9850 4620 9910
rect 6410 9850 6420 9910
rect 6480 9850 6820 9910
rect 8610 9850 8620 9910
rect 8680 9850 9020 9910
rect 10810 9850 10820 9910
rect 10880 9850 11220 9910
rect 13010 9850 13020 9910
rect 13080 9850 13420 9910
rect 15210 9850 15440 9910
rect 15500 9850 15620 9910
rect 17410 9850 17640 9910
rect 17700 9850 17820 9910
rect 19610 9850 20020 9910
rect 2500 9810 4020 9822
rect 2500 9750 2510 9810
rect 4010 9750 4020 9810
rect 2500 9740 4020 9750
rect 4700 9810 6220 9822
rect 4700 9750 4710 9810
rect 6210 9750 6220 9810
rect 4700 9740 6220 9750
rect 6900 9810 8420 9822
rect 6900 9750 6910 9810
rect 8410 9750 8420 9810
rect 6900 9740 8420 9750
rect 9100 9810 10620 9822
rect 9100 9750 9110 9810
rect 10610 9750 10620 9810
rect 9100 9740 10620 9750
rect 11300 9810 12820 9822
rect 11300 9750 11310 9810
rect 12810 9750 12820 9810
rect 11300 9740 12820 9750
rect 13500 9810 15020 9822
rect 13500 9750 13510 9810
rect 15010 9750 15020 9810
rect 13500 9740 15020 9750
rect 15700 9810 17220 9822
rect 15700 9750 15710 9810
rect 17210 9750 17220 9810
rect 15700 9740 17220 9750
rect 17900 9810 19420 9822
rect 17900 9750 17910 9810
rect 19410 9750 19420 9810
rect 17900 9740 19420 9750
rect 2500 9580 2510 9640
rect 2690 9580 2700 9640
rect 2500 9340 2700 9580
rect 3160 9580 3170 9640
rect 3350 9580 3360 9640
rect 3160 9340 3360 9580
rect 3820 9580 3830 9640
rect 4010 9580 4020 9640
rect 3820 9340 4020 9580
rect 4700 9580 4710 9640
rect 4890 9580 4900 9640
rect 4700 9340 4900 9580
rect 5360 9580 5370 9640
rect 5550 9580 5560 9640
rect 5360 9340 5560 9580
rect 6020 9580 6030 9640
rect 6210 9580 6220 9640
rect 6020 9340 6220 9580
rect 6900 9500 7100 9640
rect 6900 9440 6910 9500
rect 7090 9440 7100 9500
rect 6900 9340 7100 9440
rect 7560 9500 7760 9640
rect 7560 9440 7570 9500
rect 7750 9440 7760 9500
rect 7560 9340 7760 9440
rect 8220 9500 8420 9640
rect 8220 9440 8230 9500
rect 8410 9440 8420 9500
rect 8220 9340 8420 9440
rect 9100 9500 9300 9640
rect 9100 9440 9110 9500
rect 9290 9440 9300 9500
rect 9100 9340 9300 9440
rect 9760 9500 9960 9640
rect 9760 9440 9770 9500
rect 9950 9440 9960 9500
rect 9760 9340 9960 9440
rect 10420 9500 10620 9640
rect 10420 9440 10430 9500
rect 10610 9440 10620 9500
rect 10420 9340 10620 9440
rect 11300 9500 11500 9640
rect 11300 9440 11310 9500
rect 11490 9440 11500 9500
rect 11300 9340 11500 9440
rect 11960 9500 12160 9640
rect 11960 9440 11970 9500
rect 12150 9440 12160 9500
rect 11960 9340 12160 9440
rect 12620 9500 12820 9640
rect 12620 9440 12630 9500
rect 12810 9440 12820 9500
rect 12620 9340 12820 9440
rect 13500 9500 13700 9640
rect 13500 9440 13510 9500
rect 13690 9440 13700 9500
rect 13500 9340 13700 9440
rect 14160 9500 14360 9640
rect 14160 9440 14170 9500
rect 14350 9440 14360 9500
rect 14160 9340 14360 9440
rect 14820 9500 15020 9640
rect 14820 9440 14830 9500
rect 15010 9440 15020 9500
rect 14820 9340 15020 9440
rect 15700 9580 15710 9640
rect 15890 9580 15900 9640
rect 15700 9340 15900 9580
rect 16360 9580 16370 9640
rect 16550 9580 16560 9640
rect 16360 9340 16560 9580
rect 17020 9580 17030 9640
rect 17210 9580 17220 9640
rect 17020 9340 17220 9580
rect 17900 9580 17910 9640
rect 18090 9580 18100 9640
rect 17900 9340 18100 9580
rect 18560 9580 18570 9640
rect 18750 9580 18760 9640
rect 18560 9340 18760 9580
rect 19220 9580 19230 9640
rect 19410 9580 19420 9640
rect 19220 9340 19420 9580
rect -90 9330 10 9340
rect -90 9270 -70 9330
rect -10 9270 10 9330
rect -90 9260 10 9270
rect 2110 9330 2210 9340
rect 2110 9270 2130 9330
rect 2190 9270 2210 9330
rect 2110 9260 2210 9270
rect 4310 9330 4410 9340
rect 4310 9270 4330 9330
rect 4390 9270 4410 9330
rect 4310 9260 4410 9270
rect 6510 9330 6610 9340
rect 6510 9270 6530 9330
rect 6590 9270 6610 9330
rect 6510 9260 6610 9270
rect 8710 9330 8810 9340
rect 8710 9270 8730 9330
rect 8790 9270 8810 9330
rect 8710 9260 8810 9270
rect 10910 9330 11010 9340
rect 10910 9270 10930 9330
rect 10990 9270 11010 9330
rect 10910 9260 11010 9270
rect 13110 9330 13210 9340
rect 13110 9270 13130 9330
rect 13190 9270 13210 9330
rect 13110 9260 13210 9270
rect 15310 9330 15410 9340
rect 15310 9270 15330 9330
rect 15390 9270 15410 9330
rect 15310 9260 15410 9270
rect 17510 9330 17610 9340
rect 17510 9270 17530 9330
rect 17590 9270 17610 9330
rect 17510 9260 17610 9270
rect 19710 9330 19810 9340
rect 19710 9270 19730 9330
rect 19790 9270 19810 9330
rect 19710 9260 19810 9270
rect 21910 9330 22010 9340
rect 21910 9270 21930 9330
rect 21990 9270 22010 9330
rect 21910 9260 22010 9270
rect 1900 9160 2310 9220
rect 4100 9160 4510 9220
rect 6300 9160 6420 9220
rect 6480 9160 6710 9220
rect 8500 9160 8840 9220
rect 8900 9160 8910 9220
rect 10700 9160 11040 9220
rect 11100 9160 11110 9220
rect 12900 9160 13240 9220
rect 13300 9160 13310 9220
rect 15100 9160 15440 9220
rect 15500 9160 15510 9220
rect 17300 9160 17420 9220
rect 17480 9160 17710 9220
rect 19500 9140 19910 9200
rect 2010 9050 2420 9110
rect 4210 9050 4220 9110
rect 4280 9050 4620 9110
rect 6410 9050 6640 9110
rect 6700 9050 6820 9110
rect 8610 9050 8840 9110
rect 8900 9050 9020 9110
rect 10810 9050 11040 9110
rect 11100 9050 11220 9110
rect 13010 9050 13240 9110
rect 13300 9050 13420 9110
rect 15210 9050 15220 9110
rect 15280 9050 15620 9110
rect 17410 9050 17820 9110
rect 19610 9050 20020 9110
rect 4700 9010 6220 9022
rect 420 8990 620 9000
rect 420 8910 430 8990
rect 610 8980 620 8990
rect 610 8920 4040 8980
rect 4700 8950 4710 9010
rect 6210 8950 6220 9010
rect 4700 8940 6220 8950
rect 6900 9010 8420 9022
rect 6900 8950 6910 9010
rect 8410 8950 8420 9010
rect 6900 8940 8420 8950
rect 9100 9010 10620 9022
rect 9100 8950 9110 9010
rect 10610 8950 10620 9010
rect 9100 8940 10620 8950
rect 11300 9010 12820 9022
rect 11300 8950 11310 9010
rect 12810 8950 12820 9010
rect 11300 8940 12820 8950
rect 13500 9010 15020 9022
rect 13500 8950 13510 9010
rect 15010 8950 15020 9010
rect 13500 8940 15020 8950
rect 15700 9010 17220 9022
rect 15700 8950 15710 9010
rect 17210 8950 17220 9010
rect 21300 8990 21500 9000
rect 21300 8980 21310 8990
rect 15700 8940 17220 8950
rect 17880 8920 21310 8980
rect 610 8910 620 8920
rect 420 8900 620 8910
rect 21300 8910 21310 8920
rect 21490 8910 21500 8990
rect 21300 8900 21500 8910
rect 2500 8700 2700 8840
rect 2500 8640 2510 8700
rect 2690 8640 2700 8700
rect 2500 8540 2700 8640
rect 3160 8700 3360 8840
rect 3160 8640 3170 8700
rect 3350 8640 3360 8700
rect 3160 8540 3360 8640
rect 3820 8700 4020 8840
rect 3820 8640 3830 8700
rect 4010 8640 4020 8700
rect 3820 8540 4020 8640
rect 4700 8700 4900 8840
rect 4700 8640 4710 8700
rect 4890 8640 4900 8700
rect 4700 8540 4900 8640
rect 5360 8700 5560 8840
rect 5360 8640 5370 8700
rect 5550 8640 5560 8700
rect 5360 8540 5560 8640
rect 6020 8700 6220 8840
rect 6020 8640 6030 8700
rect 6210 8640 6220 8700
rect 6020 8540 6220 8640
rect 6900 8780 6910 8840
rect 7090 8780 7100 8840
rect 6900 8540 7100 8780
rect 7560 8780 7570 8840
rect 7750 8780 7760 8840
rect 7560 8540 7760 8780
rect 8220 8780 8230 8840
rect 8410 8780 8420 8840
rect 8220 8540 8420 8780
rect 9100 8780 9110 8840
rect 9290 8780 9300 8840
rect 9100 8540 9300 8780
rect 9760 8780 9770 8840
rect 9950 8780 9960 8840
rect 9760 8540 9960 8780
rect 10420 8780 10430 8840
rect 10610 8780 10620 8840
rect 10420 8540 10620 8780
rect 11300 8780 11310 8840
rect 11490 8780 11500 8840
rect 11300 8540 11500 8780
rect 11960 8780 11970 8840
rect 12150 8780 12160 8840
rect 11960 8540 12160 8780
rect 12620 8780 12630 8840
rect 12810 8780 12820 8840
rect 12620 8540 12820 8780
rect 13500 8780 13510 8840
rect 13690 8780 13700 8840
rect 13500 8540 13700 8780
rect 14160 8780 14170 8840
rect 14350 8780 14360 8840
rect 14160 8540 14360 8780
rect 14820 8780 14830 8840
rect 15010 8780 15020 8840
rect 14820 8540 15020 8780
rect 15700 8700 15900 8840
rect 15700 8640 15710 8700
rect 15890 8640 15900 8700
rect 15700 8540 15900 8640
rect 16360 8700 16560 8840
rect 16360 8640 16370 8700
rect 16550 8640 16560 8700
rect 16360 8540 16560 8640
rect 17020 8700 17220 8840
rect 17020 8640 17030 8700
rect 17210 8640 17220 8700
rect 17020 8540 17220 8640
rect 17900 8700 18100 8840
rect 17900 8640 17910 8700
rect 18090 8640 18100 8700
rect 17900 8540 18100 8640
rect 18560 8700 18760 8840
rect 18560 8640 18570 8700
rect 18750 8640 18760 8700
rect 18560 8540 18760 8640
rect 19220 8700 19420 8840
rect 29206 8798 29252 10826
rect 29364 8798 29410 10826
rect 29522 8798 29568 10826
rect 29680 8798 29726 10826
rect 29838 8798 29884 10826
rect 30246 8798 30292 10826
rect 30404 8798 30450 10826
rect 30562 8798 30608 10826
rect 30720 8798 30766 10826
rect 30878 8798 30924 10826
rect 31286 8798 31332 10826
rect 31444 8798 31490 10826
rect 31602 8798 31648 10826
rect 31760 8798 31806 10826
rect 31918 8798 31964 10826
rect 30309 8756 30387 8757
rect 30467 8756 30545 8757
rect 30625 8756 30703 8757
rect 30783 8756 30861 8757
rect 29270 8712 29820 8756
rect 30309 8712 30861 8756
rect 30309 8711 30387 8712
rect 30467 8711 30545 8712
rect 30625 8711 30703 8712
rect 30783 8711 30861 8712
rect 31349 8756 31427 8757
rect 31507 8756 31585 8757
rect 31665 8756 31743 8757
rect 31823 8756 31901 8757
rect 31349 8712 31901 8756
rect 31349 8711 31427 8712
rect 31507 8711 31585 8712
rect 31665 8711 31743 8712
rect 31823 8711 31901 8712
rect 19220 8640 19230 8700
rect 19410 8640 19420 8700
rect 19220 8540 19420 8640
rect -90 8530 10 8540
rect -90 8470 -70 8530
rect -10 8470 10 8530
rect -90 8460 10 8470
rect 2110 8530 2210 8540
rect 2110 8470 2130 8530
rect 2190 8470 2210 8530
rect 2110 8460 2210 8470
rect 4310 8530 4410 8540
rect 4310 8470 4330 8530
rect 4390 8470 4410 8530
rect 4310 8460 4410 8470
rect 6510 8530 6610 8540
rect 6510 8470 6530 8530
rect 6590 8470 6610 8530
rect 6510 8460 6610 8470
rect 8710 8530 8810 8540
rect 8710 8470 8730 8530
rect 8790 8470 8810 8530
rect 8710 8460 8810 8470
rect 10910 8530 11010 8540
rect 10910 8470 10930 8530
rect 10990 8470 11010 8530
rect 10910 8460 11010 8470
rect 13110 8530 13210 8540
rect 13110 8470 13130 8530
rect 13190 8470 13210 8530
rect 13110 8460 13210 8470
rect 15310 8530 15410 8540
rect 15310 8470 15330 8530
rect 15390 8470 15410 8530
rect 15310 8460 15410 8470
rect 17510 8530 17610 8540
rect 17510 8470 17530 8530
rect 17590 8470 17610 8530
rect 17510 8460 17610 8470
rect 19710 8530 19810 8540
rect 19710 8470 19730 8530
rect 19790 8470 19810 8530
rect 19710 8460 19810 8470
rect 21910 8530 22010 8540
rect 21910 8470 21930 8530
rect 21990 8470 22010 8530
rect 21910 8460 22010 8470
rect 1900 8360 2310 8420
rect 4100 8360 4510 8420
rect 6300 8360 6640 8420
rect 6700 8360 6710 8420
rect 8500 8360 8620 8420
rect 8680 8360 8910 8420
rect 10700 8360 10820 8420
rect 10880 8360 11110 8420
rect 12900 8360 13020 8420
rect 13080 8360 13310 8420
rect 15100 8360 15220 8420
rect 15280 8360 15510 8420
rect 17300 8360 17640 8420
rect 17700 8360 17710 8420
rect 19500 8340 19910 8400
rect 2010 8250 2420 8310
rect 4210 8250 4440 8310
rect 4500 8250 4620 8310
rect 6410 8250 6420 8310
rect 6480 8250 6820 8310
rect 8610 8250 8620 8310
rect 8680 8250 9020 8310
rect 10810 8250 10820 8310
rect 10880 8250 11220 8310
rect 13010 8250 13020 8310
rect 13080 8250 13420 8310
rect 15210 8250 15440 8310
rect 15500 8250 15620 8310
rect 17410 8250 17820 8310
rect 19610 8250 20020 8310
rect 4700 8210 6220 8222
rect 420 8190 620 8200
rect 420 8110 430 8190
rect 610 8180 620 8190
rect 610 8120 4040 8180
rect 4700 8150 4710 8210
rect 6210 8150 6220 8210
rect 4700 8140 6220 8150
rect 6900 8210 8420 8222
rect 6900 8150 6910 8210
rect 8410 8150 8420 8210
rect 6900 8140 8420 8150
rect 9100 8210 10620 8222
rect 9100 8150 9110 8210
rect 10610 8150 10620 8210
rect 9100 8140 10620 8150
rect 11300 8210 12820 8222
rect 11300 8150 11310 8210
rect 12810 8150 12820 8210
rect 11300 8140 12820 8150
rect 13500 8210 15020 8222
rect 13500 8150 13510 8210
rect 15010 8150 15020 8210
rect 13500 8140 15020 8150
rect 15700 8210 17220 8222
rect 15700 8150 15710 8210
rect 17210 8150 17220 8210
rect 21300 8190 21500 8200
rect 21300 8180 21310 8190
rect 15700 8140 17220 8150
rect 17880 8120 21310 8180
rect 610 8110 620 8120
rect 420 8100 620 8110
rect 21300 8110 21310 8120
rect 21490 8110 21500 8190
rect 21300 8100 21500 8110
rect 2500 7900 2700 8040
rect 2500 7840 2510 7900
rect 2690 7840 2700 7900
rect 2500 7740 2700 7840
rect 3160 7900 3360 8040
rect 3160 7840 3170 7900
rect 3350 7840 3360 7900
rect 3160 7740 3360 7840
rect 3820 7900 4020 8040
rect 3820 7840 3830 7900
rect 4010 7840 4020 7900
rect 3820 7740 4020 7840
rect 4700 7900 4900 8040
rect 4700 7840 4710 7900
rect 4890 7840 4900 7900
rect 4700 7740 4900 7840
rect 5360 7900 5560 8040
rect 5360 7840 5370 7900
rect 5550 7840 5560 7900
rect 5360 7740 5560 7840
rect 6020 7900 6220 8040
rect 6020 7840 6030 7900
rect 6210 7840 6220 7900
rect 6020 7740 6220 7840
rect 6900 7980 6910 8040
rect 7090 7980 7100 8040
rect 6900 7740 7100 7980
rect 7560 7980 7570 8040
rect 7750 7980 7760 8040
rect 7560 7740 7760 7980
rect 8220 7980 8230 8040
rect 8410 7980 8420 8040
rect 8220 7740 8420 7980
rect 9100 7980 9110 8040
rect 9290 7980 9300 8040
rect 9100 7740 9300 7980
rect 9760 7980 9770 8040
rect 9950 7980 9960 8040
rect 9760 7740 9960 7980
rect 10420 7980 10430 8040
rect 10610 7980 10620 8040
rect 10420 7740 10620 7980
rect 11300 7980 11310 8040
rect 11490 7980 11500 8040
rect 11300 7740 11500 7980
rect 11960 7980 11970 8040
rect 12150 7980 12160 8040
rect 11960 7740 12160 7980
rect 12620 7980 12630 8040
rect 12810 7980 12820 8040
rect 12620 7740 12820 7980
rect 13500 7980 13510 8040
rect 13690 7980 13700 8040
rect 13500 7740 13700 7980
rect 14160 7980 14170 8040
rect 14350 7980 14360 8040
rect 14160 7740 14360 7980
rect 14820 7980 14830 8040
rect 15010 7980 15020 8040
rect 14820 7740 15020 7980
rect 15700 7900 15900 8040
rect 15700 7840 15710 7900
rect 15890 7840 15900 7900
rect 15700 7740 15900 7840
rect 16360 7900 16560 8040
rect 16360 7840 16370 7900
rect 16550 7840 16560 7900
rect 16360 7740 16560 7840
rect 17020 7900 17220 8040
rect 17020 7840 17030 7900
rect 17210 7840 17220 7900
rect 17020 7740 17220 7840
rect 17900 7900 18100 8040
rect 17900 7840 17910 7900
rect 18090 7840 18100 7900
rect 17900 7740 18100 7840
rect 18560 7900 18760 8040
rect 18560 7840 18570 7900
rect 18750 7840 18760 7900
rect 18560 7740 18760 7840
rect 19220 7900 19420 8040
rect 19220 7840 19230 7900
rect 19410 7840 19420 7900
rect 19220 7740 19420 7840
rect -90 7730 10 7740
rect -90 7670 -70 7730
rect -10 7670 10 7730
rect -90 7660 10 7670
rect 2110 7730 2210 7740
rect 2110 7670 2130 7730
rect 2190 7670 2210 7730
rect 2110 7660 2210 7670
rect 4310 7730 4410 7740
rect 4310 7670 4330 7730
rect 4390 7670 4410 7730
rect 4310 7660 4410 7670
rect 6510 7730 6610 7740
rect 6510 7670 6530 7730
rect 6590 7670 6610 7730
rect 6510 7660 6610 7670
rect 8710 7730 8810 7740
rect 8710 7670 8730 7730
rect 8790 7670 8810 7730
rect 8710 7660 8810 7670
rect 10910 7730 11010 7740
rect 10910 7670 10930 7730
rect 10990 7670 11010 7730
rect 10910 7660 11010 7670
rect 13110 7730 13210 7740
rect 13110 7670 13130 7730
rect 13190 7670 13210 7730
rect 13110 7660 13210 7670
rect 15310 7730 15410 7740
rect 15310 7670 15330 7730
rect 15390 7670 15410 7730
rect 15310 7660 15410 7670
rect 17510 7730 17610 7740
rect 17510 7670 17530 7730
rect 17590 7670 17610 7730
rect 17510 7660 17610 7670
rect 19710 7730 19810 7740
rect 19710 7670 19730 7730
rect 19790 7670 19810 7730
rect 19710 7660 19810 7670
rect 21910 7730 22010 7740
rect 21910 7670 21930 7730
rect 21990 7670 22010 7730
rect 21910 7660 22010 7670
rect 1900 7560 2310 7620
rect 4100 7560 4510 7620
rect 6300 7560 6640 7620
rect 6700 7560 6710 7620
rect 8500 7560 8620 7620
rect 8680 7560 8910 7620
rect 10700 7560 10820 7620
rect 10880 7560 11110 7620
rect 12900 7560 13020 7620
rect 13080 7560 13310 7620
rect 15100 7560 15220 7620
rect 15280 7560 15510 7620
rect 17300 7560 17640 7620
rect 17700 7560 17710 7620
rect 19500 7540 19910 7600
rect 2010 7450 2420 7510
rect 4210 7450 4440 7510
rect 4500 7450 4620 7510
rect 6410 7450 6420 7510
rect 6480 7450 6820 7510
rect 8610 7450 8620 7510
rect 8680 7450 9020 7510
rect 10810 7450 10820 7510
rect 10880 7450 11220 7510
rect 13010 7450 13020 7510
rect 13080 7450 13420 7510
rect 15210 7450 15440 7510
rect 15500 7450 15620 7510
rect 17410 7450 17820 7510
rect 19610 7450 20020 7510
rect 4700 7410 6220 7422
rect 420 7390 620 7400
rect 420 7310 430 7390
rect 610 7380 620 7390
rect 610 7320 4040 7380
rect 4700 7350 4710 7410
rect 6210 7350 6220 7410
rect 4700 7340 6220 7350
rect 6900 7410 8420 7422
rect 6900 7350 6910 7410
rect 8410 7350 8420 7410
rect 6900 7340 8420 7350
rect 9100 7410 10620 7422
rect 9100 7350 9110 7410
rect 10610 7350 10620 7410
rect 9100 7340 10620 7350
rect 11300 7410 12820 7422
rect 11300 7350 11310 7410
rect 12810 7350 12820 7410
rect 11300 7340 12820 7350
rect 13500 7410 15020 7422
rect 13500 7350 13510 7410
rect 15010 7350 15020 7410
rect 13500 7340 15020 7350
rect 15700 7410 17220 7422
rect 15700 7350 15710 7410
rect 17210 7350 17220 7410
rect 21300 7390 21500 7400
rect 21300 7380 21310 7390
rect 15700 7340 17220 7350
rect 17880 7320 21310 7380
rect 610 7310 620 7320
rect 420 7300 620 7310
rect 21300 7310 21310 7320
rect 21490 7310 21500 7390
rect 21300 7300 21500 7310
rect 2500 7180 2510 7240
rect 2690 7180 2700 7240
rect 2500 6940 2700 7180
rect 3160 7180 3170 7240
rect 3350 7180 3360 7240
rect 3160 6940 3360 7180
rect 3820 7180 3830 7240
rect 4010 7180 4020 7240
rect 3820 6940 4020 7180
rect 4700 7180 4710 7240
rect 4890 7180 4900 7240
rect 4700 6940 4900 7180
rect 5360 7180 5370 7240
rect 5550 7180 5560 7240
rect 5360 6940 5560 7180
rect 6020 7180 6030 7240
rect 6210 7180 6220 7240
rect 6020 6940 6220 7180
rect 6900 7100 7100 7240
rect 6900 7040 6910 7100
rect 7090 7040 7100 7100
rect 6900 6940 7100 7040
rect 7560 7100 7760 7240
rect 7560 7040 7570 7100
rect 7750 7040 7760 7100
rect 7560 6940 7760 7040
rect 8220 7100 8420 7240
rect 8220 7040 8230 7100
rect 8410 7040 8420 7100
rect 8220 6940 8420 7040
rect 9100 7100 9300 7240
rect 9100 7040 9110 7100
rect 9290 7040 9300 7100
rect 9100 6940 9300 7040
rect 9760 7100 9960 7240
rect 9760 7040 9770 7100
rect 9950 7040 9960 7100
rect 9760 6940 9960 7040
rect 10420 7100 10620 7240
rect 10420 7040 10430 7100
rect 10610 7040 10620 7100
rect 10420 6940 10620 7040
rect 11300 7100 11500 7240
rect 11300 7040 11310 7100
rect 11490 7040 11500 7100
rect 11300 6940 11500 7040
rect 11960 7100 12160 7240
rect 11960 7040 11970 7100
rect 12150 7040 12160 7100
rect 11960 6940 12160 7040
rect 12620 7100 12820 7240
rect 12620 7040 12630 7100
rect 12810 7040 12820 7100
rect 12620 6940 12820 7040
rect 13500 7100 13700 7240
rect 13500 7040 13510 7100
rect 13690 7040 13700 7100
rect 13500 6940 13700 7040
rect 14160 7100 14360 7240
rect 14160 7040 14170 7100
rect 14350 7040 14360 7100
rect 14160 6940 14360 7040
rect 14820 7100 15020 7240
rect 14820 7040 14830 7100
rect 15010 7040 15020 7100
rect 14820 6940 15020 7040
rect 15700 7180 15710 7240
rect 15890 7180 15900 7240
rect 15700 6940 15900 7180
rect 16360 7180 16370 7240
rect 16550 7180 16560 7240
rect 16360 6940 16560 7180
rect 17020 7180 17030 7240
rect 17210 7180 17220 7240
rect 17020 6940 17220 7180
rect 17900 7180 17910 7240
rect 18090 7180 18100 7240
rect 17900 6940 18100 7180
rect 18560 7180 18570 7240
rect 18750 7180 18760 7240
rect 18560 6940 18760 7180
rect 19220 7180 19230 7240
rect 19410 7180 19420 7240
rect 19220 6940 19420 7180
rect -90 6930 10 6940
rect -90 6870 -70 6930
rect -10 6870 10 6930
rect -90 6860 10 6870
rect 2110 6930 2210 6940
rect 2110 6870 2130 6930
rect 2190 6870 2210 6930
rect 2110 6860 2210 6870
rect 4310 6930 4410 6940
rect 4310 6870 4330 6930
rect 4390 6870 4410 6930
rect 4310 6860 4410 6870
rect 6510 6930 6610 6940
rect 6510 6870 6530 6930
rect 6590 6870 6610 6930
rect 6510 6860 6610 6870
rect 8710 6930 8810 6940
rect 8710 6870 8730 6930
rect 8790 6870 8810 6930
rect 8710 6860 8810 6870
rect 10910 6930 11010 6940
rect 10910 6870 10930 6930
rect 10990 6870 11010 6930
rect 10910 6860 11010 6870
rect 13110 6930 13210 6940
rect 13110 6870 13130 6930
rect 13190 6870 13210 6930
rect 13110 6860 13210 6870
rect 15310 6930 15410 6940
rect 15310 6870 15330 6930
rect 15390 6870 15410 6930
rect 15310 6860 15410 6870
rect 17510 6930 17610 6940
rect 17510 6870 17530 6930
rect 17590 6870 17610 6930
rect 17510 6860 17610 6870
rect 19710 6930 19810 6940
rect 19710 6870 19730 6930
rect 19790 6870 19810 6930
rect 19710 6860 19810 6870
rect 21910 6930 22010 6940
rect 21910 6870 21930 6930
rect 21990 6870 22010 6930
rect 21910 6860 22010 6870
rect 1900 6760 2310 6820
rect 4100 6760 4510 6820
rect 6300 6760 6420 6820
rect 6480 6760 6710 6820
rect 8500 6760 8840 6820
rect 8900 6760 8910 6820
rect 10700 6760 11040 6820
rect 11100 6760 11110 6820
rect 12900 6760 13240 6820
rect 13300 6760 13310 6820
rect 15100 6760 15440 6820
rect 15500 6760 15510 6820
rect 17300 6760 17420 6820
rect 17480 6760 17710 6820
rect 19500 6740 19910 6800
rect 2010 6650 2420 6710
rect 4210 6650 4220 6710
rect 4280 6650 4620 6710
rect 6410 6650 6640 6710
rect 6700 6650 6820 6710
rect 8610 6650 8840 6710
rect 8900 6650 9020 6710
rect 10810 6650 11040 6710
rect 11100 6650 11220 6710
rect 13010 6650 13240 6710
rect 13300 6650 13420 6710
rect 15210 6650 15220 6710
rect 15280 6650 15620 6710
rect 17410 6650 17820 6710
rect 19610 6650 20020 6710
rect 4700 6610 6220 6622
rect 420 6590 620 6600
rect 420 6510 430 6590
rect 610 6580 620 6590
rect 610 6520 4040 6580
rect 4700 6550 4710 6610
rect 6210 6550 6220 6610
rect 4700 6540 6220 6550
rect 6900 6610 8420 6622
rect 6900 6550 6910 6610
rect 8410 6550 8420 6610
rect 6900 6540 8420 6550
rect 9100 6610 10620 6622
rect 9100 6550 9110 6610
rect 10610 6550 10620 6610
rect 9100 6540 10620 6550
rect 11300 6610 12820 6622
rect 11300 6550 11310 6610
rect 12810 6550 12820 6610
rect 11300 6540 12820 6550
rect 13500 6610 15020 6622
rect 13500 6550 13510 6610
rect 15010 6550 15020 6610
rect 13500 6540 15020 6550
rect 15700 6610 17220 6622
rect 15700 6550 15710 6610
rect 17210 6550 17220 6610
rect 21300 6590 21500 6600
rect 21300 6580 21310 6590
rect 15700 6540 17220 6550
rect 17880 6520 21310 6580
rect 610 6510 620 6520
rect 420 6500 620 6510
rect 21300 6510 21310 6520
rect 21490 6510 21500 6590
rect 21300 6500 21500 6510
rect 2500 6300 2700 6440
rect 2500 6240 2510 6300
rect 2690 6240 2700 6300
rect 2500 6140 2700 6240
rect 3160 6300 3360 6440
rect 3160 6240 3170 6300
rect 3350 6240 3360 6300
rect 3160 6140 3360 6240
rect 3820 6300 4020 6440
rect 3820 6240 3830 6300
rect 4010 6240 4020 6300
rect 3820 6140 4020 6240
rect 4700 6300 4900 6440
rect 4700 6240 4710 6300
rect 4890 6240 4900 6300
rect 4700 6140 4900 6240
rect 5360 6300 5560 6440
rect 5360 6240 5370 6300
rect 5550 6240 5560 6300
rect 5360 6140 5560 6240
rect 6020 6300 6220 6440
rect 6020 6240 6030 6300
rect 6210 6240 6220 6300
rect 6020 6140 6220 6240
rect 6900 6380 6910 6440
rect 7090 6380 7100 6440
rect 6900 6140 7100 6380
rect 7560 6380 7570 6440
rect 7750 6380 7760 6440
rect 7560 6140 7760 6380
rect 8220 6380 8230 6440
rect 8410 6380 8420 6440
rect 8220 6140 8420 6380
rect 9100 6380 9110 6440
rect 9290 6380 9300 6440
rect 9100 6140 9300 6380
rect 9760 6380 9770 6440
rect 9950 6380 9960 6440
rect 9760 6140 9960 6380
rect 10420 6380 10430 6440
rect 10610 6380 10620 6440
rect 10420 6140 10620 6380
rect 11300 6380 11310 6440
rect 11490 6380 11500 6440
rect 11300 6140 11500 6380
rect 11960 6380 11970 6440
rect 12150 6380 12160 6440
rect 11960 6140 12160 6380
rect 12620 6380 12630 6440
rect 12810 6380 12820 6440
rect 12620 6140 12820 6380
rect 13500 6380 13510 6440
rect 13690 6380 13700 6440
rect 13500 6140 13700 6380
rect 14160 6380 14170 6440
rect 14350 6380 14360 6440
rect 14160 6140 14360 6380
rect 14820 6380 14830 6440
rect 15010 6380 15020 6440
rect 14820 6140 15020 6380
rect 15700 6300 15900 6440
rect 15700 6240 15710 6300
rect 15890 6240 15900 6300
rect 15700 6140 15900 6240
rect 16360 6300 16560 6440
rect 16360 6240 16370 6300
rect 16550 6240 16560 6300
rect 16360 6140 16560 6240
rect 17020 6300 17220 6440
rect 17020 6240 17030 6300
rect 17210 6240 17220 6300
rect 17020 6140 17220 6240
rect 17900 6300 18100 6440
rect 17900 6240 17910 6300
rect 18090 6240 18100 6300
rect 17900 6140 18100 6240
rect 18560 6300 18760 6440
rect 18560 6240 18570 6300
rect 18750 6240 18760 6300
rect 18560 6140 18760 6240
rect 19220 6300 19420 6440
rect 19220 6240 19230 6300
rect 19410 6240 19420 6300
rect 19220 6140 19420 6240
rect -90 6130 10 6140
rect -90 6070 -70 6130
rect -10 6070 10 6130
rect -90 6060 10 6070
rect 2110 6130 2210 6140
rect 2110 6070 2130 6130
rect 2190 6070 2210 6130
rect 2110 6060 2210 6070
rect 4310 6130 4410 6140
rect 4310 6070 4330 6130
rect 4390 6070 4410 6130
rect 4310 6060 4410 6070
rect 6510 6130 6610 6140
rect 6510 6070 6530 6130
rect 6590 6070 6610 6130
rect 6510 6060 6610 6070
rect 8710 6130 8810 6140
rect 8710 6070 8730 6130
rect 8790 6070 8810 6130
rect 8710 6060 8810 6070
rect 10910 6130 11010 6140
rect 10910 6070 10930 6130
rect 10990 6070 11010 6130
rect 10910 6060 11010 6070
rect 13110 6130 13210 6140
rect 13110 6070 13130 6130
rect 13190 6070 13210 6130
rect 13110 6060 13210 6070
rect 15310 6130 15410 6140
rect 15310 6070 15330 6130
rect 15390 6070 15410 6130
rect 15310 6060 15410 6070
rect 17510 6130 17610 6140
rect 17510 6070 17530 6130
rect 17590 6070 17610 6130
rect 17510 6060 17610 6070
rect 19710 6130 19810 6140
rect 19710 6070 19730 6130
rect 19790 6070 19810 6130
rect 19710 6060 19810 6070
rect 21910 6130 22010 6140
rect 21910 6070 21930 6130
rect 21990 6070 22010 6130
rect 21910 6060 22010 6070
rect 1900 5960 2310 6020
rect 4100 5960 4440 6020
rect 4500 5960 4510 6020
rect 6300 5960 6640 6020
rect 6700 5960 6710 6020
rect 8500 5960 8620 6020
rect 8680 5960 8910 6020
rect 10700 5960 10820 6020
rect 10880 5960 11110 6020
rect 12900 5960 13020 6020
rect 13080 5960 13310 6020
rect 15100 5960 15220 6020
rect 15280 5960 15510 6020
rect 17300 5960 17640 6020
rect 17700 5960 17710 6020
rect 19500 5940 19840 6000
rect 19900 5940 19910 6000
rect 2010 5850 2240 5910
rect 2300 5850 2420 5910
rect 4210 5850 4440 5910
rect 4500 5850 4620 5910
rect 6410 5850 6420 5910
rect 6480 5850 6820 5910
rect 8610 5850 8620 5910
rect 8680 5850 9020 5910
rect 10810 5850 10820 5910
rect 10880 5850 11220 5910
rect 13010 5850 13020 5910
rect 13080 5850 13420 5910
rect 15210 5850 15440 5910
rect 15500 5850 15620 5910
rect 17410 5850 17640 5910
rect 17700 5850 17820 5910
rect 19610 5850 20020 5910
rect 2500 5810 4020 5822
rect 2500 5750 2510 5810
rect 4010 5750 4020 5810
rect 2500 5740 4020 5750
rect 4700 5810 6220 5822
rect 4700 5750 4710 5810
rect 6210 5750 6220 5810
rect 4700 5740 6220 5750
rect 6900 5810 8420 5822
rect 6900 5750 6910 5810
rect 8410 5750 8420 5810
rect 6900 5740 8420 5750
rect 9100 5810 10620 5822
rect 9100 5750 9110 5810
rect 10610 5750 10620 5810
rect 9100 5740 10620 5750
rect 11300 5810 12820 5822
rect 11300 5750 11310 5810
rect 12810 5750 12820 5810
rect 11300 5740 12820 5750
rect 13500 5810 15020 5822
rect 13500 5750 13510 5810
rect 15010 5750 15020 5810
rect 13500 5740 15020 5750
rect 15700 5810 17220 5822
rect 15700 5750 15710 5810
rect 17210 5750 17220 5810
rect 15700 5740 17220 5750
rect 17900 5810 19420 5822
rect 17900 5750 17910 5810
rect 19410 5750 19420 5810
rect 17900 5740 19420 5750
rect 22630 5740 23330 5980
rect 2500 5580 2510 5640
rect 2690 5580 2700 5640
rect 2500 5340 2700 5580
rect 3160 5580 3170 5640
rect 3350 5580 3360 5640
rect 3160 5340 3360 5580
rect 3820 5580 3830 5640
rect 4010 5580 4020 5640
rect 3820 5340 4020 5580
rect 4700 5580 4710 5640
rect 4890 5580 4900 5640
rect 4700 5340 4900 5580
rect 5360 5580 5370 5640
rect 5550 5580 5560 5640
rect 5360 5340 5560 5580
rect 6020 5580 6030 5640
rect 6210 5580 6220 5640
rect 6020 5340 6220 5580
rect 6900 5500 7100 5640
rect 6900 5440 6910 5500
rect 7090 5440 7100 5500
rect 6900 5340 7100 5440
rect 7560 5500 7760 5640
rect 7560 5440 7570 5500
rect 7750 5440 7760 5500
rect 7560 5340 7760 5440
rect 8220 5500 8420 5640
rect 8220 5440 8230 5500
rect 8410 5440 8420 5500
rect 8220 5340 8420 5440
rect 9100 5500 9300 5640
rect 9100 5440 9110 5500
rect 9290 5440 9300 5500
rect 9100 5340 9300 5440
rect 9760 5500 9960 5640
rect 9760 5440 9770 5500
rect 9950 5440 9960 5500
rect 9760 5340 9960 5440
rect 10420 5500 10620 5640
rect 10420 5440 10430 5500
rect 10610 5440 10620 5500
rect 10420 5340 10620 5440
rect 11300 5500 11500 5640
rect 11300 5440 11310 5500
rect 11490 5440 11500 5500
rect 11300 5340 11500 5440
rect 11960 5500 12160 5640
rect 11960 5440 11970 5500
rect 12150 5440 12160 5500
rect 11960 5340 12160 5440
rect 12620 5500 12820 5640
rect 12620 5440 12630 5500
rect 12810 5440 12820 5500
rect 12620 5340 12820 5440
rect 13500 5500 13700 5640
rect 13500 5440 13510 5500
rect 13690 5440 13700 5500
rect 13500 5340 13700 5440
rect 14160 5500 14360 5640
rect 14160 5440 14170 5500
rect 14350 5440 14360 5500
rect 14160 5340 14360 5440
rect 14820 5500 15020 5640
rect 14820 5440 14830 5500
rect 15010 5440 15020 5500
rect 14820 5340 15020 5440
rect 15700 5580 15710 5640
rect 15890 5580 15900 5640
rect 15700 5340 15900 5580
rect 16360 5580 16370 5640
rect 16550 5580 16560 5640
rect 16360 5340 16560 5580
rect 17020 5580 17030 5640
rect 17210 5580 17220 5640
rect 17020 5340 17220 5580
rect 17900 5580 17910 5640
rect 18090 5580 18100 5640
rect 17900 5340 18100 5580
rect 18560 5580 18570 5640
rect 18750 5580 18760 5640
rect 18560 5340 18760 5580
rect 19220 5580 19230 5640
rect 19410 5580 19420 5640
rect 19220 5340 19420 5580
rect 22780 5440 23330 5740
rect 24110 5580 25330 5980
rect 25440 5580 26660 5980
rect 26770 5580 27990 5980
rect 28100 5740 28790 5980
rect 28100 5440 28650 5740
rect -90 5330 10 5340
rect -90 5270 -70 5330
rect -10 5270 10 5330
rect -90 5260 10 5270
rect 2110 5330 2210 5340
rect 2110 5270 2130 5330
rect 2190 5270 2210 5330
rect 2110 5260 2210 5270
rect 4310 5330 4410 5340
rect 4310 5270 4330 5330
rect 4390 5270 4410 5330
rect 4310 5260 4410 5270
rect 6510 5330 6610 5340
rect 6510 5270 6530 5330
rect 6590 5270 6610 5330
rect 6510 5260 6610 5270
rect 8710 5330 8810 5340
rect 8710 5270 8730 5330
rect 8790 5270 8810 5330
rect 8710 5260 8810 5270
rect 10910 5330 11010 5340
rect 10910 5270 10930 5330
rect 10990 5270 11010 5330
rect 10910 5260 11010 5270
rect 13110 5330 13210 5340
rect 13110 5270 13130 5330
rect 13190 5270 13210 5330
rect 13110 5260 13210 5270
rect 15310 5330 15410 5340
rect 15310 5270 15330 5330
rect 15390 5270 15410 5330
rect 15310 5260 15410 5270
rect 17510 5330 17610 5340
rect 17510 5270 17530 5330
rect 17590 5270 17610 5330
rect 17510 5260 17610 5270
rect 19710 5330 19810 5340
rect 19710 5270 19730 5330
rect 19790 5270 19810 5330
rect 19710 5260 19810 5270
rect 21910 5330 22010 5340
rect 21910 5270 21930 5330
rect 21990 5270 22010 5330
rect 21910 5260 22010 5270
rect 1900 5160 2310 5220
rect 4100 5160 4220 5220
rect 4280 5160 4510 5220
rect 6300 5160 6420 5220
rect 6480 5160 6710 5220
rect 8500 5160 8840 5220
rect 8900 5160 8910 5220
rect 10700 5160 11040 5220
rect 11100 5160 11110 5220
rect 12900 5160 13240 5220
rect 13300 5160 13310 5220
rect 15100 5160 15440 5220
rect 15500 5160 15510 5220
rect 17300 5160 17420 5220
rect 17480 5160 17710 5220
rect 19500 5140 19620 5200
rect 19680 5140 19910 5200
rect 2010 5050 2020 5110
rect 2080 5050 2420 5110
rect 4210 5050 4220 5110
rect 4280 5050 4620 5110
rect 6410 5050 6640 5110
rect 6700 5050 6820 5110
rect 8610 5050 8840 5110
rect 8900 5050 9020 5110
rect 10810 5050 11040 5110
rect 11100 5050 11220 5110
rect 13010 5050 13240 5110
rect 13300 5050 13420 5110
rect 15210 5050 15220 5110
rect 15280 5050 15620 5110
rect 17410 5050 17420 5110
rect 17480 5050 17820 5110
rect 19610 5050 20020 5110
rect 2500 5010 4020 5022
rect 2500 4950 2510 5010
rect 4010 4950 4020 5010
rect 2500 4940 4020 4950
rect 4700 5010 6220 5022
rect 4700 4950 4710 5010
rect 6210 4950 6220 5010
rect 4700 4940 6220 4950
rect 6900 5010 8420 5022
rect 6900 4950 6910 5010
rect 8410 4950 8420 5010
rect 6900 4940 8420 4950
rect 9100 5010 10620 5022
rect 9100 4950 9110 5010
rect 10610 4950 10620 5010
rect 9100 4940 10620 4950
rect 11300 5010 12820 5022
rect 11300 4950 11310 5010
rect 12810 4950 12820 5010
rect 11300 4940 12820 4950
rect 13500 5010 15020 5022
rect 13500 4950 13510 5010
rect 15010 4950 15020 5010
rect 13500 4940 15020 4950
rect 15700 5010 17220 5022
rect 15700 4950 15710 5010
rect 17210 4950 17220 5010
rect 15700 4940 17220 4950
rect 17900 5010 19420 5022
rect 17900 4950 17910 5010
rect 19410 4950 19420 5010
rect 17900 4940 19420 4950
rect -820 2160 31780 2240
rect -820 2040 11160 2160
rect 11240 2040 12300 2120
rect 12380 2040 12760 2160
rect 12840 2040 13900 2120
rect 13980 2080 31780 2160
rect 13980 2040 14870 2080
rect 15070 2040 31780 2080
rect 2100 1970 2240 1980
rect 2100 1290 2110 1970
rect 2230 1290 2240 1970
rect 2100 1280 2240 1290
rect 3700 1970 3840 1980
rect 3700 1290 3710 1970
rect 3830 1290 3840 1970
rect 3700 1280 3840 1290
rect 5300 1970 5440 1980
rect 5300 1290 5310 1970
rect 5430 1290 5440 1970
rect 5300 1280 5440 1290
rect 6900 1970 7040 1980
rect 6900 1290 6910 1970
rect 7030 1290 7040 1970
rect 6900 1280 7040 1290
rect 8500 1970 8640 1980
rect 8500 1290 8510 1970
rect 8630 1290 8640 1970
rect 8500 1280 8640 1290
rect 10100 1970 10240 1980
rect 10100 1290 10110 1970
rect 10230 1290 10240 1970
rect 11020 1930 11220 1940
rect 11020 1310 11030 1930
rect 11150 1310 11220 1930
rect 11020 1300 11220 1310
rect 10100 1280 10240 1290
rect 11700 1280 11840 1980
rect 12310 1930 12820 1940
rect 12310 1310 12610 1930
rect 12730 1310 12820 1930
rect 12310 1300 12820 1310
rect 13300 1280 13440 1980
rect 14900 1960 15040 1990
rect 13910 1930 14120 1940
rect 13910 1310 13990 1930
rect 14110 1310 14120 1930
rect 13910 1220 14120 1310
rect 14900 1300 14910 1960
rect 15030 1300 15040 1960
rect 14900 1220 15040 1300
rect 16500 1970 16640 1980
rect 16500 1290 16510 1970
rect 16630 1290 16640 1970
rect 16500 1280 16640 1290
rect 18100 1970 18240 1980
rect 18100 1290 18110 1970
rect 18230 1290 18240 1970
rect 18100 1280 18240 1290
rect 19700 1970 19840 1980
rect 19700 1290 19710 1970
rect 19830 1290 19840 1970
rect 19700 1280 19840 1290
rect 21300 1970 21440 1980
rect 21300 1290 21310 1970
rect 21430 1290 21440 1970
rect 21300 1280 21440 1290
rect 22900 1970 23040 1980
rect 22900 1290 22910 1970
rect 23030 1290 23040 1970
rect 22900 1280 23040 1290
rect 24500 1970 24640 1980
rect 24500 1290 24510 1970
rect 24630 1290 24640 1970
rect 24500 1280 24640 1290
rect 26100 1970 26240 1980
rect 26100 1290 26110 1970
rect 26230 1290 26240 1970
rect 26100 1280 26240 1290
rect 27700 1970 27840 1980
rect 27700 1290 27710 1970
rect 27830 1290 27840 1970
rect 27700 1280 27840 1290
rect 28781 1975 28827 1987
rect 28781 1283 28787 1975
rect 28821 1283 28827 1975
rect 28781 1271 28827 1283
rect 29291 1980 29337 1987
rect 29399 1980 29445 1987
rect 29291 1975 29445 1980
rect 29291 1283 29297 1975
rect 29331 1970 29405 1975
rect 29331 1283 29405 1290
rect 29439 1283 29445 1975
rect 29291 1280 29445 1283
rect 29291 1271 29337 1280
rect 29399 1271 29445 1280
rect 29909 1975 29955 1987
rect 29909 1283 29915 1975
rect 29949 1283 29955 1975
rect 29909 1271 29955 1283
rect 30381 1975 30427 1987
rect 30381 1283 30387 1975
rect 30421 1283 30427 1975
rect 30381 1271 30427 1283
rect 30891 1980 30937 1987
rect 30999 1980 31045 1987
rect 30891 1975 31045 1980
rect 30891 1283 30897 1975
rect 30931 1970 31005 1975
rect 30931 1283 31005 1290
rect 31039 1283 31045 1975
rect 30891 1280 31045 1283
rect 30891 1271 30937 1280
rect 30999 1271 31045 1280
rect 31509 1975 31555 1987
rect 32500 1975 32640 1980
rect 34100 1975 34240 1980
rect 35700 1975 35840 1980
rect 31509 1283 31515 1975
rect 31549 1283 31555 1975
rect 32531 1970 32605 1975
rect 32531 1283 32605 1290
rect 32639 1283 32640 1975
rect 34131 1970 34205 1975
rect 34131 1283 34205 1290
rect 34239 1283 34240 1975
rect 35731 1970 35805 1975
rect 35731 1283 35805 1290
rect 35839 1283 35840 1975
rect 31509 1271 31555 1283
rect 32500 1280 32640 1283
rect 34100 1280 34240 1283
rect 35700 1280 35840 1283
rect 11240 1210 11680 1220
rect 1680 1140 2040 1200
rect 2300 1140 2660 1200
rect 3280 1140 3640 1200
rect 3900 1140 4260 1200
rect 4880 1140 5240 1200
rect 5500 1140 5860 1200
rect 6480 1140 6840 1200
rect 7100 1140 7460 1200
rect 8080 1140 8440 1200
rect 8700 1140 9060 1200
rect 9680 1140 10040 1200
rect 10300 1140 10660 1200
rect 1400 1130 10660 1140
rect 1400 1010 1410 1130
rect 1530 1010 3010 1130
rect 3130 1010 4610 1130
rect 4730 1010 6210 1130
rect 6330 1010 7810 1130
rect 7930 1010 9410 1130
rect 9530 1010 10660 1130
rect 11240 1050 11250 1210
rect 11670 1050 11680 1210
rect 11860 1100 13280 1220
rect 13480 1100 14120 1220
rect 14460 1130 15480 1220
rect 16059 1217 16459 1223
rect 16059 1183 16071 1217
rect 16080 1183 16440 1200
rect 16447 1183 16459 1217
rect 16059 1177 16459 1183
rect 16677 1217 17077 1223
rect 16677 1183 16689 1217
rect 16700 1183 17060 1200
rect 17065 1183 17077 1217
rect 16677 1177 17077 1183
rect 17659 1217 18059 1223
rect 17659 1183 17671 1217
rect 17680 1183 18040 1200
rect 18047 1183 18059 1217
rect 17659 1177 18059 1183
rect 18277 1217 18677 1223
rect 18277 1183 18289 1217
rect 18300 1183 18660 1200
rect 18665 1183 18677 1217
rect 18277 1177 18677 1183
rect 19259 1217 19659 1223
rect 19259 1183 19271 1217
rect 19280 1183 19640 1200
rect 19647 1183 19659 1217
rect 19259 1177 19659 1183
rect 19877 1217 20277 1223
rect 19877 1183 19889 1217
rect 19900 1183 20260 1200
rect 20265 1183 20277 1217
rect 19877 1177 20277 1183
rect 20859 1217 21259 1223
rect 20859 1183 20871 1217
rect 20880 1183 21240 1200
rect 21247 1183 21259 1217
rect 20859 1177 21259 1183
rect 21477 1217 21877 1223
rect 21477 1183 21489 1217
rect 21500 1183 21860 1200
rect 21865 1183 21877 1217
rect 21477 1177 21877 1183
rect 22459 1217 22859 1223
rect 22459 1183 22471 1217
rect 22480 1183 22840 1200
rect 22847 1183 22859 1217
rect 22459 1177 22859 1183
rect 23077 1217 23477 1223
rect 23077 1183 23089 1217
rect 23100 1183 23460 1200
rect 23465 1183 23477 1217
rect 23077 1177 23477 1183
rect 24059 1217 24459 1223
rect 24059 1183 24071 1217
rect 24080 1183 24440 1200
rect 24447 1183 24459 1217
rect 24059 1177 24459 1183
rect 24677 1217 25077 1223
rect 24677 1183 24689 1217
rect 24700 1183 25060 1200
rect 25065 1183 25077 1217
rect 24677 1177 25077 1183
rect 25659 1217 26059 1223
rect 25659 1183 25671 1217
rect 25680 1183 26040 1200
rect 26047 1183 26059 1217
rect 25659 1177 26059 1183
rect 26277 1217 26677 1223
rect 26277 1183 26289 1217
rect 26300 1183 26660 1200
rect 26665 1183 26677 1217
rect 26277 1177 26677 1183
rect 27259 1217 27659 1223
rect 27259 1183 27271 1217
rect 27280 1183 27640 1200
rect 27647 1183 27659 1217
rect 27259 1177 27659 1183
rect 27877 1217 28277 1223
rect 27877 1183 27889 1217
rect 27900 1183 28260 1200
rect 28265 1183 28277 1217
rect 27877 1177 28277 1183
rect 28859 1217 29259 1223
rect 28859 1183 28871 1217
rect 28880 1183 29240 1200
rect 29247 1183 29259 1217
rect 28859 1177 29259 1183
rect 29477 1217 29877 1223
rect 29477 1183 29489 1217
rect 29500 1183 29860 1200
rect 29865 1183 29877 1217
rect 29477 1177 29877 1183
rect 30459 1217 30859 1223
rect 30459 1183 30471 1217
rect 30847 1183 30859 1217
rect 30459 1177 30859 1183
rect 31077 1217 31477 1223
rect 31077 1183 31089 1217
rect 31465 1183 31477 1217
rect 33659 1217 34059 1223
rect 31077 1177 31477 1183
rect 32080 1183 32440 1200
rect 32447 1183 32459 1200
rect 32080 1177 32459 1183
rect 32677 1183 32689 1200
rect 32700 1183 33060 1200
rect 32677 1177 33060 1183
rect 33659 1183 33671 1217
rect 33680 1183 34040 1200
rect 34047 1183 34059 1217
rect 33659 1177 34059 1183
rect 34277 1217 34677 1223
rect 34277 1183 34289 1217
rect 34300 1183 34660 1200
rect 34665 1183 34677 1217
rect 34277 1177 34677 1183
rect 35259 1217 35659 1223
rect 35259 1183 35271 1217
rect 35280 1183 35640 1200
rect 35647 1183 35659 1217
rect 35259 1177 35659 1183
rect 35877 1217 36277 1223
rect 35877 1183 35889 1217
rect 35900 1183 36260 1200
rect 36265 1183 36277 1217
rect 35877 1177 36277 1183
rect 16080 1140 16440 1177
rect 16700 1140 17060 1177
rect 17680 1140 18040 1177
rect 18300 1140 18660 1177
rect 19280 1140 19640 1177
rect 19900 1140 20260 1177
rect 20880 1140 21240 1177
rect 21500 1140 21860 1177
rect 22480 1140 22840 1177
rect 23100 1140 23460 1177
rect 24080 1140 24440 1177
rect 24700 1140 25060 1177
rect 25680 1140 26040 1177
rect 26300 1140 26660 1177
rect 27280 1140 27640 1177
rect 27900 1140 28260 1177
rect 28880 1140 29240 1177
rect 29500 1140 29860 1177
rect 30480 1140 30840 1177
rect 31100 1140 31460 1177
rect 15590 1130 17060 1140
rect 11240 1040 11680 1050
rect 1400 1000 10660 1010
rect 15590 1010 15600 1130
rect 15700 1010 17060 1130
rect 15590 1000 17060 1010
rect 17190 1130 18660 1140
rect 17190 1010 17200 1130
rect 17300 1010 18660 1130
rect 17190 1000 18660 1010
rect 18790 1130 20260 1140
rect 18790 1010 18800 1130
rect 18900 1010 20260 1130
rect 18790 1000 20260 1010
rect 20390 1130 21860 1140
rect 20390 1010 20400 1130
rect 20500 1010 21860 1130
rect 20390 1000 21860 1010
rect 21990 1130 23460 1140
rect 21990 1010 22000 1130
rect 22100 1010 23460 1130
rect 21990 1000 23460 1010
rect 23590 1130 25060 1140
rect 23590 1010 23600 1130
rect 23700 1010 25060 1130
rect 23590 1000 25060 1010
rect 25660 1130 28260 1140
rect 25660 1010 26800 1130
rect 26900 1010 28260 1130
rect 25660 1000 28260 1010
rect 28391 1130 31460 1140
rect 28391 1010 28400 1130
rect 28500 1010 31460 1130
rect 28391 1000 31460 1010
rect 1680 940 2040 1000
rect 2300 940 2660 1000
rect 3280 940 3640 1000
rect 3900 940 4260 1000
rect 4880 940 5240 1000
rect 5500 940 5860 1000
rect 6480 940 6840 1000
rect 7100 940 7460 1000
rect 8080 940 8440 1000
rect 8700 940 9060 1000
rect 9680 940 10040 1000
rect 10300 940 10660 1000
rect 16080 955 16440 1000
rect 16700 955 17060 1000
rect 17680 955 18040 1000
rect 18300 955 18660 1000
rect 19280 955 19640 1000
rect 19900 955 20260 1000
rect 20880 955 21240 1000
rect 21500 955 21860 1000
rect 22480 955 22840 1000
rect 23100 955 23460 1000
rect 24080 955 24440 1000
rect 24700 955 25060 1000
rect 25680 955 26040 1000
rect 26300 955 26660 1000
rect 27280 955 27640 1000
rect 27900 955 28260 1000
rect 28880 955 29240 1000
rect 29500 955 29860 1000
rect 30480 955 30840 1000
rect 31100 955 31460 1000
rect 32080 1140 32440 1177
rect 32700 1140 33060 1177
rect 33680 1140 34040 1177
rect 34300 1140 34660 1177
rect 32080 1000 34660 1140
rect 32080 955 32440 1000
rect 32700 955 33060 1000
rect 33680 955 34040 1000
rect 34300 955 34660 1000
rect 35280 1140 35640 1177
rect 35900 1140 36260 1177
rect 35280 1000 36260 1140
rect 35280 955 35640 1000
rect 35900 955 36260 1000
rect 16059 949 16459 955
rect 1690 930 2030 940
rect 2310 930 2650 940
rect 3290 930 3630 940
rect 3910 930 4250 940
rect 4890 930 5230 940
rect 5510 930 5850 940
rect 6490 930 6830 940
rect 7110 930 7450 940
rect 8090 930 8430 940
rect 8710 930 9050 940
rect 9690 930 10030 940
rect 10310 930 10650 940
rect 16059 915 16071 949
rect 16080 940 16440 949
rect 16090 930 16430 940
rect 16447 915 16459 949
rect 16059 909 16459 915
rect 16677 949 17077 955
rect 16677 915 16689 949
rect 16700 940 17060 949
rect 16710 930 17050 940
rect 17065 915 17077 949
rect 16677 909 17077 915
rect 17659 949 18059 955
rect 17659 915 17671 949
rect 17680 940 18040 949
rect 17690 930 18030 940
rect 18047 915 18059 949
rect 17659 909 18059 915
rect 18277 949 18677 955
rect 18277 915 18289 949
rect 18300 940 18660 949
rect 18310 930 18650 940
rect 18665 915 18677 949
rect 18277 909 18677 915
rect 19259 949 19659 955
rect 19259 915 19271 949
rect 19280 940 19640 949
rect 19290 930 19630 940
rect 19647 915 19659 949
rect 19259 909 19659 915
rect 19877 949 20277 955
rect 19877 915 19889 949
rect 19900 940 20260 949
rect 19910 930 20250 940
rect 20265 915 20277 949
rect 19877 909 20277 915
rect 20859 949 21259 955
rect 20859 915 20871 949
rect 20880 940 21240 949
rect 20890 930 21230 940
rect 21247 915 21259 949
rect 20859 909 21259 915
rect 21477 949 21877 955
rect 21477 915 21489 949
rect 21500 940 21860 949
rect 21510 930 21850 940
rect 21865 915 21877 949
rect 21477 909 21877 915
rect 22459 949 22859 955
rect 22459 915 22471 949
rect 22480 940 22840 949
rect 22490 930 22830 940
rect 22847 915 22859 949
rect 22459 909 22859 915
rect 23077 949 23477 955
rect 23077 915 23089 949
rect 23100 940 23460 949
rect 23110 930 23450 940
rect 23465 915 23477 949
rect 23077 909 23477 915
rect 24059 949 24459 955
rect 24059 915 24071 949
rect 24080 940 24440 949
rect 24090 930 24430 940
rect 24447 915 24459 949
rect 24059 909 24459 915
rect 24677 949 25077 955
rect 24677 915 24689 949
rect 24700 940 25060 949
rect 24710 930 25050 940
rect 25065 915 25077 949
rect 24677 909 25077 915
rect 25659 949 26059 955
rect 25659 915 25671 949
rect 25680 940 26040 949
rect 25690 930 26030 940
rect 26047 915 26059 949
rect 25659 909 26059 915
rect 26277 949 26677 955
rect 26277 915 26289 949
rect 26300 940 26660 949
rect 26310 930 26650 940
rect 26665 915 26677 949
rect 26277 909 26677 915
rect 27259 949 27659 955
rect 27259 915 27271 949
rect 27280 940 27640 949
rect 27290 930 27630 940
rect 27647 915 27659 949
rect 27259 909 27659 915
rect 27877 949 28277 955
rect 27877 915 27889 949
rect 27900 940 28260 949
rect 27910 930 28250 940
rect 28265 915 28277 949
rect 27877 909 28277 915
rect 28859 949 29259 955
rect 28859 915 28871 949
rect 28880 940 29240 949
rect 28890 930 29230 940
rect 29247 915 29259 949
rect 28859 909 29259 915
rect 29477 949 29877 955
rect 29477 915 29489 949
rect 29500 940 29860 949
rect 29510 930 29850 940
rect 29865 915 29877 949
rect 29477 909 29877 915
rect 30459 949 30859 955
rect 30459 915 30471 949
rect 30847 915 30859 949
rect 30459 909 30859 915
rect 31077 949 31477 955
rect 31077 915 31089 949
rect 31465 915 31477 949
rect 32080 949 32459 955
rect 32080 940 32440 949
rect 32447 940 32459 949
rect 32677 949 33060 955
rect 32677 940 32689 949
rect 32700 940 33060 949
rect 33659 949 34059 955
rect 31077 909 31477 915
rect 33659 915 33671 949
rect 33680 940 34040 949
rect 34047 915 34059 949
rect 33659 909 34059 915
rect 34277 949 34677 955
rect 34277 915 34289 949
rect 34300 940 34660 949
rect 34665 915 34677 949
rect 34277 909 34677 915
rect 35259 949 35659 955
rect 35259 915 35271 949
rect 35280 940 35640 949
rect 35647 915 35659 949
rect 35259 909 35659 915
rect 35877 949 36277 955
rect 35877 915 35889 949
rect 35900 940 36260 949
rect 36265 915 36277 949
rect 35877 909 36277 915
rect 12320 870 12520 880
rect 1540 750 12390 870
rect 12510 750 36400 870
rect 1540 740 36400 750
rect 30459 691 30859 697
rect 30459 690 30471 691
rect 30847 690 30859 691
rect 31077 691 31477 697
rect 31077 690 31089 691
rect 31465 690 31477 691
rect 1180 680 1320 690
rect 2780 680 2920 690
rect 4380 680 4520 690
rect 5980 680 6120 690
rect 7580 680 7720 690
rect 9180 680 9320 690
rect 15810 680 15930 690
rect 17410 680 17530 690
rect 19010 680 19130 690
rect 20610 680 20730 690
rect 22210 680 22330 690
rect 23810 680 23930 690
rect 27010 680 27130 690
rect 28610 680 31520 690
rect 1180 560 1190 680
rect 1310 560 2790 680
rect 2910 560 4390 680
rect 4510 560 5990 680
rect 6110 560 7590 680
rect 7710 560 9190 680
rect 9310 560 10720 680
rect 15810 560 15820 680
rect 15920 560 17120 680
rect 17410 560 17420 680
rect 17520 560 18720 680
rect 19010 560 19020 680
rect 19120 560 20320 680
rect 20610 560 20620 680
rect 20720 560 21920 680
rect 22210 560 22220 680
rect 22320 560 23520 680
rect 23810 560 23820 680
rect 23920 560 25120 680
rect 25620 560 27020 680
rect 27120 560 28320 680
rect 28610 560 28620 680
rect 28720 560 31520 680
rect 1180 550 1320 560
rect 2780 550 2920 560
rect 4380 550 4520 560
rect 5980 550 6120 560
rect 7580 550 7720 560
rect 9180 550 9320 560
rect 15810 550 15930 560
rect 17410 550 17530 560
rect 19010 550 19130 560
rect 20610 550 20730 560
rect 22210 550 22330 560
rect 23810 550 23930 560
rect 27010 550 27130 560
rect 28610 550 31520 560
rect 31810 680 31930 690
rect 31810 560 31820 680
rect 31920 560 36270 680
rect 31810 550 31930 560
rect -820 240 38090 440
rect 2100 170 2240 180
rect 2100 -510 2110 170
rect 2230 -510 2240 170
rect 2100 -520 2240 -510
rect 3700 170 3840 180
rect 3700 -510 3710 170
rect 3830 -510 3840 170
rect 3700 -520 3840 -510
rect 5300 170 5440 180
rect 5300 -510 5310 170
rect 5430 -510 5440 170
rect 5300 -520 5440 -510
rect 6900 170 7040 180
rect 6900 -510 6910 170
rect 7030 -510 7040 170
rect 6900 -520 7040 -510
rect 8500 170 8640 180
rect 8500 -510 8510 170
rect 8630 -510 8640 170
rect 8500 -520 8640 -510
rect 10100 170 10240 180
rect 10100 -510 10110 170
rect 10230 -510 10240 170
rect 10100 -520 10240 -510
rect 11700 170 11840 180
rect 11700 -580 11710 170
rect 11260 -590 11710 -580
rect 11830 -580 11840 170
rect 13300 170 13440 180
rect 13300 -510 13310 170
rect 13430 -510 13440 170
rect 14900 170 15040 180
rect 13300 -520 13440 -510
rect 14380 -580 14430 -510
rect 14900 -580 14910 170
rect 11830 -590 12280 -580
rect 1680 -660 2040 -600
rect 2300 -660 2660 -600
rect 3280 -660 3640 -600
rect 3900 -660 4260 -600
rect 4880 -660 5240 -600
rect 5500 -660 5860 -600
rect 6480 -660 6840 -600
rect 7100 -660 7460 -600
rect 8080 -660 8440 -600
rect 8700 -660 9060 -600
rect 9680 -660 10040 -600
rect 10300 -660 10660 -600
rect 1400 -670 10660 -660
rect 1400 -790 1410 -670
rect 1530 -790 3010 -670
rect 3130 -790 4610 -670
rect 4730 -790 6210 -670
rect 6330 -790 7810 -670
rect 7930 -790 9410 -670
rect 9530 -790 10660 -670
rect 11260 -750 11270 -590
rect 12270 -750 12280 -590
rect 14380 -590 14910 -580
rect 15030 -580 15040 170
rect 16500 170 16640 180
rect 16500 -510 16510 170
rect 16630 -510 16640 170
rect 15510 -580 15560 -510
rect 16500 -520 16640 -510
rect 18100 170 18240 180
rect 18100 -510 18110 170
rect 18230 -510 18240 170
rect 18100 -520 18240 -510
rect 19700 170 19840 180
rect 19700 -510 19710 170
rect 19830 -510 19840 170
rect 19700 -520 19840 -510
rect 21300 170 21440 180
rect 21300 -510 21310 170
rect 21430 -510 21440 170
rect 21300 -520 21440 -510
rect 22900 170 23040 180
rect 22900 -510 22910 170
rect 23030 -510 23040 170
rect 22900 -520 23040 -510
rect 24500 170 24640 180
rect 24500 -510 24510 170
rect 24630 -510 24640 170
rect 24500 -520 24640 -510
rect 26100 170 26240 180
rect 26100 -510 26110 170
rect 26230 -510 26240 170
rect 26100 -520 26240 -510
rect 27700 170 27840 180
rect 27700 -510 27710 170
rect 27830 -510 27840 170
rect 27700 -520 27840 -510
rect 28781 175 28827 187
rect 28781 -517 28787 175
rect 28821 -517 28827 175
rect 28781 -529 28827 -517
rect 29291 180 29337 187
rect 29399 180 29445 187
rect 29291 175 29445 180
rect 29291 -517 29297 175
rect 29331 170 29405 175
rect 29331 -517 29405 -510
rect 29439 -517 29445 175
rect 29291 -520 29445 -517
rect 29291 -529 29337 -520
rect 29399 -529 29445 -520
rect 29909 175 29955 187
rect 29909 -517 29915 175
rect 29949 -517 29955 175
rect 29909 -529 29955 -517
rect 30381 175 30427 187
rect 30381 -517 30387 175
rect 30421 -517 30427 175
rect 30381 -529 30427 -517
rect 30891 180 30937 187
rect 30999 180 31045 187
rect 30891 175 31045 180
rect 30891 -517 30897 175
rect 30931 170 31005 175
rect 30931 -517 31005 -510
rect 31039 -517 31045 175
rect 30891 -520 31045 -517
rect 30891 -529 30937 -520
rect 30999 -529 31045 -520
rect 31509 175 31555 187
rect 32500 175 32640 180
rect 31509 -517 31515 175
rect 31549 -517 31555 175
rect 32531 170 32605 175
rect 32531 -517 32605 -510
rect 32639 -517 32640 175
rect 34100 170 34240 180
rect 35700 175 35840 180
rect 35731 170 35805 175
rect 34100 140 34110 170
rect 34230 140 34240 170
rect 34131 -517 34205 -510
rect 34239 -517 34240 140
rect 35731 -517 35805 -510
rect 35839 -517 35840 175
rect 31509 -529 31555 -517
rect 32500 -520 32640 -517
rect 34100 -520 34240 -517
rect 35700 -520 35840 -517
rect 15030 -590 15560 -580
rect 12880 -617 13240 -600
rect 13247 -617 13259 -600
rect 12880 -623 13259 -617
rect 13477 -617 13489 -600
rect 13500 -617 13860 -600
rect 13477 -623 13860 -617
rect 12880 -660 13240 -623
rect 13500 -660 13860 -623
rect 11260 -760 12280 -750
rect 12380 -670 14300 -660
rect 1400 -800 10660 -790
rect 1680 -860 2040 -800
rect 2300 -860 2660 -800
rect 3280 -860 3640 -800
rect 3900 -860 4260 -800
rect 4880 -860 5240 -800
rect 5500 -860 5860 -800
rect 6480 -860 6840 -800
rect 7100 -860 7460 -800
rect 8080 -860 8440 -800
rect 8700 -860 9060 -800
rect 9680 -860 10040 -800
rect 10300 -860 10660 -800
rect 1690 -870 2030 -860
rect 2310 -870 2650 -860
rect 3290 -870 3630 -860
rect 3910 -870 4250 -860
rect 4890 -870 5230 -860
rect 5510 -870 5850 -860
rect 6490 -870 6830 -860
rect 7110 -870 7450 -860
rect 8090 -870 8430 -860
rect 8710 -870 9050 -860
rect 9690 -870 10030 -860
rect 10310 -870 10650 -860
rect 12380 -910 12390 -670
rect 12310 -930 12390 -910
rect 1540 -1050 12390 -930
rect 12510 -800 14300 -670
rect 14380 -750 14470 -590
rect 15470 -750 15560 -590
rect 16059 -583 16459 -577
rect 16059 -617 16071 -583
rect 16080 -617 16440 -600
rect 16447 -617 16459 -583
rect 16059 -623 16459 -617
rect 16677 -583 17077 -577
rect 16677 -617 16689 -583
rect 16700 -617 17060 -600
rect 17065 -617 17077 -583
rect 16677 -623 17077 -617
rect 17659 -583 18059 -577
rect 17659 -617 17671 -583
rect 17680 -617 18040 -600
rect 18047 -617 18059 -583
rect 17659 -623 18059 -617
rect 18277 -583 18677 -577
rect 18277 -617 18289 -583
rect 18300 -617 18660 -600
rect 18665 -617 18677 -583
rect 18277 -623 18677 -617
rect 19259 -583 19659 -577
rect 19259 -617 19271 -583
rect 19280 -617 19640 -600
rect 19647 -617 19659 -583
rect 19259 -623 19659 -617
rect 19877 -583 20277 -577
rect 19877 -617 19889 -583
rect 19900 -617 20260 -600
rect 20265 -617 20277 -583
rect 19877 -623 20277 -617
rect 20859 -583 21259 -577
rect 20859 -617 20871 -583
rect 20880 -617 21240 -600
rect 21247 -617 21259 -583
rect 20859 -623 21259 -617
rect 21477 -583 21877 -577
rect 21477 -617 21489 -583
rect 21500 -617 21860 -600
rect 21865 -617 21877 -583
rect 21477 -623 21877 -617
rect 22459 -583 22859 -577
rect 22459 -617 22471 -583
rect 22480 -617 22840 -600
rect 22847 -617 22859 -583
rect 22459 -623 22859 -617
rect 23077 -583 23477 -577
rect 23077 -617 23089 -583
rect 23100 -617 23460 -600
rect 23465 -617 23477 -583
rect 23077 -623 23477 -617
rect 24059 -583 24459 -577
rect 24059 -617 24071 -583
rect 24080 -617 24440 -600
rect 24447 -617 24459 -583
rect 24059 -623 24459 -617
rect 24677 -583 25077 -577
rect 24677 -617 24689 -583
rect 24700 -617 25060 -600
rect 25065 -617 25077 -583
rect 24677 -623 25077 -617
rect 25659 -583 26059 -577
rect 25659 -617 25671 -583
rect 25680 -617 26040 -600
rect 26047 -617 26059 -583
rect 25659 -623 26059 -617
rect 26277 -583 26677 -577
rect 26277 -617 26289 -583
rect 26300 -617 26660 -600
rect 26665 -617 26677 -583
rect 26277 -623 26677 -617
rect 27259 -583 27659 -577
rect 27259 -617 27271 -583
rect 27280 -617 27640 -600
rect 27647 -617 27659 -583
rect 27259 -623 27659 -617
rect 27877 -583 28277 -577
rect 27877 -617 27889 -583
rect 27900 -617 28260 -600
rect 28265 -617 28277 -583
rect 27877 -623 28277 -617
rect 28859 -583 29259 -577
rect 28859 -617 28871 -583
rect 28880 -617 29240 -600
rect 29247 -617 29259 -583
rect 28859 -623 29259 -617
rect 29477 -583 29877 -577
rect 29477 -617 29489 -583
rect 29500 -617 29860 -600
rect 29865 -617 29877 -583
rect 29477 -623 29877 -617
rect 30459 -583 30859 -577
rect 30459 -617 30471 -583
rect 30847 -617 30859 -583
rect 30459 -623 30859 -617
rect 31077 -583 31477 -577
rect 31077 -617 31089 -583
rect 31465 -617 31477 -583
rect 33659 -583 34059 -577
rect 31077 -623 31477 -617
rect 32080 -617 32440 -600
rect 32447 -617 32459 -600
rect 32080 -623 32459 -617
rect 32677 -617 32689 -600
rect 32700 -617 33060 -600
rect 32677 -623 33060 -617
rect 33659 -617 33671 -583
rect 33680 -617 34040 -600
rect 34047 -617 34059 -583
rect 33659 -623 34059 -617
rect 34277 -583 34677 -577
rect 34277 -617 34289 -583
rect 34300 -617 34660 -600
rect 34665 -617 34677 -583
rect 34277 -623 34677 -617
rect 35259 -583 35659 -577
rect 35259 -617 35271 -583
rect 35280 -617 35640 -600
rect 35647 -617 35659 -583
rect 35259 -623 35659 -617
rect 35877 -583 36277 -577
rect 35877 -617 35889 -583
rect 35900 -617 36260 -600
rect 36265 -617 36277 -583
rect 35877 -623 36277 -617
rect 16080 -660 16440 -623
rect 16700 -660 17060 -623
rect 17680 -660 18040 -623
rect 18300 -660 18660 -623
rect 19280 -660 19640 -623
rect 19900 -660 20260 -623
rect 20880 -660 21240 -623
rect 21500 -660 21860 -623
rect 22480 -660 22840 -623
rect 23100 -660 23460 -623
rect 24080 -660 24440 -623
rect 24700 -660 25060 -623
rect 25680 -660 26040 -623
rect 26300 -660 26660 -623
rect 27280 -660 27640 -623
rect 27900 -660 28260 -623
rect 28880 -660 29240 -623
rect 29500 -660 29860 -623
rect 30480 -660 30840 -623
rect 31100 -660 31460 -623
rect 14380 -760 15560 -750
rect 15590 -670 17060 -660
rect 15590 -790 15600 -670
rect 15700 -790 17060 -670
rect 15590 -800 17060 -790
rect 17190 -670 18660 -660
rect 17190 -790 17200 -670
rect 17300 -790 18660 -670
rect 17190 -800 18660 -790
rect 18790 -670 20260 -660
rect 18790 -790 18800 -670
rect 18900 -790 20260 -670
rect 18790 -800 20260 -790
rect 20390 -670 21860 -660
rect 20390 -790 20400 -670
rect 20500 -790 21860 -670
rect 20390 -800 21860 -790
rect 21990 -670 23460 -660
rect 21990 -790 22000 -670
rect 22100 -790 23460 -670
rect 21990 -800 23460 -790
rect 23590 -670 25060 -660
rect 23590 -790 23600 -670
rect 23700 -790 25060 -670
rect 23590 -800 25060 -790
rect 25660 -670 28260 -660
rect 25660 -790 26800 -670
rect 26900 -790 28260 -670
rect 25660 -800 28260 -790
rect 28390 -670 31460 -660
rect 28390 -790 28400 -670
rect 28500 -790 31460 -670
rect 28390 -800 31460 -790
rect 12510 -1050 12520 -800
rect 12880 -845 13240 -800
rect 13500 -845 13860 -800
rect 12880 -851 13259 -845
rect 12880 -860 13240 -851
rect 13247 -860 13259 -851
rect 13477 -851 13860 -845
rect 13477 -860 13489 -851
rect 13500 -860 13860 -851
rect 1540 -1060 12520 -1050
rect 12620 -930 12820 -920
rect 12620 -1070 12630 -930
rect 12750 -1070 12820 -930
rect 12620 -1080 12820 -1070
rect 13920 -930 14100 -920
rect 13920 -1070 13970 -930
rect 14090 -1070 14100 -930
rect 14160 -930 14300 -800
rect 16080 -845 16440 -800
rect 16700 -845 17060 -800
rect 17680 -845 18040 -800
rect 18300 -845 18660 -800
rect 19280 -845 19640 -800
rect 19900 -845 20260 -800
rect 20880 -845 21240 -800
rect 21500 -845 21860 -800
rect 22480 -845 22840 -800
rect 23100 -845 23460 -800
rect 24080 -845 24440 -800
rect 24700 -845 25060 -800
rect 25680 -845 26040 -800
rect 26300 -845 26660 -800
rect 27280 -845 27640 -800
rect 27900 -845 28260 -800
rect 28880 -845 29240 -800
rect 29500 -845 29860 -800
rect 30480 -845 30840 -800
rect 31100 -845 31460 -800
rect 32080 -660 32440 -623
rect 32700 -660 33060 -623
rect 33680 -660 34040 -623
rect 34300 -660 34660 -623
rect 35280 -660 35640 -623
rect 35900 -660 36260 -623
rect 32080 -800 36260 -660
rect 32080 -845 32440 -800
rect 32700 -845 33060 -800
rect 33680 -845 34040 -800
rect 34300 -845 34660 -800
rect 35280 -845 35640 -800
rect 35900 -845 36260 -800
rect 16059 -851 16459 -845
rect 16059 -885 16071 -851
rect 16080 -860 16440 -851
rect 16090 -870 16430 -860
rect 16447 -885 16459 -851
rect 16059 -891 16459 -885
rect 16677 -851 17077 -845
rect 16677 -885 16689 -851
rect 16700 -860 17060 -851
rect 16710 -870 17050 -860
rect 17065 -885 17077 -851
rect 16677 -891 17077 -885
rect 17659 -851 18059 -845
rect 17659 -885 17671 -851
rect 17680 -860 18040 -851
rect 17690 -870 18030 -860
rect 18047 -885 18059 -851
rect 17659 -891 18059 -885
rect 18277 -851 18677 -845
rect 18277 -885 18289 -851
rect 18300 -860 18660 -851
rect 18310 -870 18650 -860
rect 18665 -885 18677 -851
rect 18277 -891 18677 -885
rect 19259 -851 19659 -845
rect 19259 -885 19271 -851
rect 19280 -860 19640 -851
rect 19290 -870 19630 -860
rect 19647 -885 19659 -851
rect 19259 -891 19659 -885
rect 19877 -851 20277 -845
rect 19877 -885 19889 -851
rect 19900 -860 20260 -851
rect 19910 -870 20250 -860
rect 20265 -885 20277 -851
rect 19877 -891 20277 -885
rect 20859 -851 21259 -845
rect 20859 -885 20871 -851
rect 20880 -860 21240 -851
rect 20890 -870 21230 -860
rect 21247 -885 21259 -851
rect 20859 -891 21259 -885
rect 21477 -851 21877 -845
rect 21477 -885 21489 -851
rect 21500 -860 21860 -851
rect 21510 -870 21850 -860
rect 21865 -885 21877 -851
rect 21477 -891 21877 -885
rect 22459 -851 22859 -845
rect 22459 -885 22471 -851
rect 22480 -860 22840 -851
rect 22490 -870 22830 -860
rect 22847 -885 22859 -851
rect 22459 -891 22859 -885
rect 23077 -851 23477 -845
rect 23077 -885 23089 -851
rect 23100 -860 23460 -851
rect 23110 -870 23450 -860
rect 23465 -885 23477 -851
rect 23077 -891 23477 -885
rect 24059 -851 24459 -845
rect 24059 -885 24071 -851
rect 24080 -860 24440 -851
rect 24090 -870 24430 -860
rect 24447 -885 24459 -851
rect 24059 -891 24459 -885
rect 24677 -851 25077 -845
rect 24677 -885 24689 -851
rect 24700 -860 25060 -851
rect 24710 -870 25050 -860
rect 25065 -885 25077 -851
rect 24677 -891 25077 -885
rect 25659 -851 26059 -845
rect 25659 -885 25671 -851
rect 25680 -860 26040 -851
rect 25690 -870 26030 -860
rect 26047 -885 26059 -851
rect 25659 -891 26059 -885
rect 26277 -851 26677 -845
rect 26277 -885 26289 -851
rect 26300 -860 26660 -851
rect 26310 -870 26650 -860
rect 26665 -885 26677 -851
rect 26277 -891 26677 -885
rect 27259 -851 27659 -845
rect 27259 -885 27271 -851
rect 27280 -860 27640 -851
rect 27290 -870 27630 -860
rect 27647 -885 27659 -851
rect 27259 -891 27659 -885
rect 27877 -851 28277 -845
rect 27877 -885 27889 -851
rect 27900 -860 28260 -851
rect 27910 -870 28250 -860
rect 28265 -885 28277 -851
rect 27877 -891 28277 -885
rect 28859 -851 29259 -845
rect 28859 -885 28871 -851
rect 28880 -860 29240 -851
rect 28890 -870 29230 -860
rect 29247 -885 29259 -851
rect 28859 -891 29259 -885
rect 29477 -851 29877 -845
rect 29477 -885 29489 -851
rect 29500 -860 29860 -851
rect 29510 -870 29850 -860
rect 29865 -885 29877 -851
rect 29477 -891 29877 -885
rect 30459 -851 30859 -845
rect 30459 -885 30471 -851
rect 30847 -885 30859 -851
rect 30459 -891 30859 -885
rect 31077 -851 31477 -845
rect 31077 -885 31089 -851
rect 31465 -885 31477 -851
rect 32080 -851 32459 -845
rect 32080 -860 32440 -851
rect 32447 -860 32459 -851
rect 32677 -851 33060 -845
rect 32677 -860 32689 -851
rect 32700 -860 33060 -851
rect 33659 -851 34059 -845
rect 31077 -891 31477 -885
rect 33659 -885 33671 -851
rect 33680 -860 34040 -851
rect 34047 -885 34059 -851
rect 33659 -891 34059 -885
rect 34277 -851 34677 -845
rect 34277 -885 34289 -851
rect 34300 -860 34660 -851
rect 34665 -885 34677 -851
rect 34277 -891 34677 -885
rect 35259 -851 35659 -845
rect 35259 -885 35271 -851
rect 35280 -860 35640 -851
rect 35647 -885 35659 -851
rect 35259 -891 35659 -885
rect 35877 -851 36277 -845
rect 35877 -885 35889 -851
rect 35900 -860 36260 -851
rect 36265 -885 36277 -851
rect 35877 -891 36277 -885
rect 14160 -1060 36400 -930
rect 13920 -1080 14100 -1070
rect 30459 -1109 30859 -1103
rect 30459 -1110 30471 -1109
rect 30847 -1110 30859 -1109
rect 31077 -1109 31477 -1103
rect 31077 -1110 31089 -1109
rect 31465 -1110 31477 -1109
rect 1180 -1120 1320 -1110
rect 2780 -1120 2920 -1110
rect 4380 -1120 4520 -1110
rect 5980 -1120 6120 -1110
rect 7580 -1120 7720 -1110
rect 9180 -1120 9320 -1110
rect 15810 -1120 15930 -1110
rect 17410 -1120 17530 -1110
rect 19010 -1120 19130 -1110
rect 20610 -1120 20730 -1110
rect 22210 -1120 22330 -1110
rect 23810 -1120 23930 -1110
rect 27010 -1120 28270 -1110
rect 1180 -1240 1190 -1120
rect 1310 -1240 2790 -1120
rect 2910 -1240 4390 -1120
rect 4510 -1240 5990 -1120
rect 6110 -1240 7590 -1120
rect 7710 -1240 9190 -1120
rect 9310 -1240 10720 -1120
rect 12860 -1200 13880 -1120
rect 10800 -1210 13880 -1200
rect 1180 -1250 1320 -1240
rect 2780 -1250 2920 -1240
rect 4380 -1250 4520 -1240
rect 5980 -1250 6120 -1240
rect 7580 -1250 7720 -1240
rect 9180 -1250 9320 -1240
rect 10800 -1270 10810 -1210
rect 10990 -1270 13880 -1210
rect 15810 -1240 15820 -1120
rect 15920 -1240 17120 -1120
rect 17410 -1240 17420 -1120
rect 17520 -1240 18720 -1120
rect 19010 -1240 19020 -1120
rect 19120 -1240 20320 -1120
rect 20610 -1240 20620 -1120
rect 20720 -1240 21920 -1120
rect 22210 -1240 22220 -1120
rect 22320 -1240 23520 -1120
rect 23810 -1240 23820 -1120
rect 23920 -1240 25120 -1120
rect 25620 -1240 27020 -1120
rect 27120 -1240 28270 -1120
rect 15810 -1250 15930 -1240
rect 17410 -1250 17530 -1240
rect 19010 -1250 19130 -1240
rect 20610 -1250 20730 -1240
rect 22210 -1250 22330 -1240
rect 23810 -1250 23930 -1240
rect 27010 -1250 28270 -1240
rect 28610 -1120 31520 -1110
rect 28610 -1240 28620 -1120
rect 28720 -1240 31520 -1120
rect 28610 -1250 31520 -1240
rect 31590 -1120 31710 -1110
rect 31590 -1240 31600 -1120
rect 31700 -1240 36270 -1120
rect 31590 -1250 31710 -1240
rect 10800 -1280 13880 -1270
rect -820 -1560 31780 -1360
rect 33660 -1560 36270 -1500
rect 2100 -1630 2240 -1620
rect 2100 -2310 2110 -1630
rect 2230 -2310 2240 -1630
rect 2100 -2320 2240 -2310
rect 3700 -1630 3840 -1620
rect 3700 -2310 3710 -1630
rect 3830 -2310 3840 -1630
rect 3700 -2320 3840 -2310
rect 5300 -1630 5440 -1620
rect 5300 -2310 5310 -1630
rect 5430 -2310 5440 -1630
rect 5300 -2320 5440 -2310
rect 6900 -1630 7040 -1620
rect 6900 -2310 6910 -1630
rect 7030 -2310 7040 -1630
rect 6900 -2320 7040 -2310
rect 8500 -1630 8640 -1620
rect 8500 -2310 8510 -1630
rect 8630 -2310 8640 -1630
rect 8500 -2320 8640 -2310
rect 10100 -1630 10240 -1620
rect 10100 -2310 10110 -1630
rect 10230 -2310 10240 -1630
rect 10100 -2320 10240 -2310
rect 11700 -1630 11840 -1620
rect 11700 -2310 11710 -1630
rect 11830 -2310 11840 -1630
rect 11700 -2320 11840 -2310
rect 13300 -1630 13440 -1620
rect 13300 -2310 13310 -1630
rect 13430 -2310 13440 -1630
rect 13300 -2320 13440 -2310
rect 14900 -1630 15040 -1620
rect 14900 -2310 14910 -1630
rect 15030 -2310 15040 -1630
rect 14900 -2320 15040 -2310
rect 16500 -1630 16640 -1620
rect 16500 -2310 16510 -1630
rect 16630 -2310 16640 -1630
rect 16500 -2320 16640 -2310
rect 18100 -1630 18240 -1620
rect 18100 -2310 18110 -1630
rect 18230 -2310 18240 -1630
rect 18100 -2320 18240 -2310
rect 19700 -1630 19840 -1620
rect 19700 -2310 19710 -1630
rect 19830 -2310 19840 -1630
rect 19700 -2320 19840 -2310
rect 21300 -1630 21440 -1620
rect 21300 -2310 21310 -1630
rect 21430 -2310 21440 -1630
rect 21300 -2320 21440 -2310
rect 22900 -1630 23040 -1620
rect 22900 -2310 22910 -1630
rect 23030 -2310 23040 -1630
rect 22900 -2320 23040 -2310
rect 24500 -1630 24640 -1620
rect 24500 -2310 24510 -1630
rect 24630 -2310 24640 -1630
rect 24500 -2320 24640 -2310
rect 26100 -1630 26240 -1620
rect 26100 -2310 26110 -1630
rect 26230 -2310 26240 -1630
rect 26100 -2320 26240 -2310
rect 27700 -1630 27840 -1620
rect 27700 -2310 27710 -1630
rect 27830 -2310 27840 -1630
rect 27700 -2320 27840 -2310
rect 28781 -1625 28827 -1613
rect 28781 -2317 28787 -1625
rect 28821 -2317 28827 -1625
rect 28781 -2329 28827 -2317
rect 29291 -1620 29337 -1613
rect 29399 -1620 29445 -1613
rect 29291 -1625 29445 -1620
rect 29291 -2317 29297 -1625
rect 29331 -1630 29405 -1625
rect 29331 -2317 29405 -2310
rect 29439 -2317 29445 -1625
rect 29291 -2320 29445 -2317
rect 29291 -2329 29337 -2320
rect 29399 -2329 29445 -2320
rect 29909 -1625 29955 -1613
rect 29909 -2317 29915 -1625
rect 29949 -2317 29955 -1625
rect 29909 -2329 29955 -2317
rect 30381 -1625 30427 -1613
rect 30381 -2317 30387 -1625
rect 30421 -2317 30427 -1625
rect 30381 -2329 30427 -2317
rect 30891 -1620 30937 -1613
rect 30999 -1620 31045 -1613
rect 30891 -1625 31045 -1620
rect 30891 -2317 30897 -1625
rect 30931 -1630 31005 -1625
rect 30931 -2317 31005 -2310
rect 31039 -2317 31045 -1625
rect 30891 -2320 31045 -2317
rect 30891 -2329 30937 -2320
rect 30999 -2329 31045 -2320
rect 31509 -1625 31555 -1613
rect 32500 -1625 32640 -1620
rect 34100 -1625 34240 -1620
rect 35700 -1625 35840 -1620
rect 31509 -2317 31515 -1625
rect 31549 -2317 31555 -1625
rect 32531 -1630 32605 -1625
rect 32531 -2317 32605 -2310
rect 32639 -2317 32640 -1625
rect 34131 -1630 34205 -1625
rect 34131 -2317 34205 -2310
rect 34239 -2317 34240 -1625
rect 35731 -1630 35805 -1625
rect 35731 -2317 35805 -2310
rect 35839 -2317 35840 -1625
rect 31509 -2329 31555 -2317
rect 32500 -2320 32640 -2317
rect 34100 -2320 34240 -2317
rect 35700 -2320 35840 -2317
rect 11260 -2383 11659 -2380
rect 1680 -2460 2040 -2400
rect 2300 -2460 2660 -2400
rect 3280 -2460 3640 -2400
rect 3900 -2460 4260 -2400
rect 4880 -2460 5240 -2400
rect 5500 -2460 5860 -2400
rect 6480 -2460 6840 -2400
rect 7100 -2460 7460 -2400
rect 8080 -2460 8440 -2400
rect 8700 -2460 9060 -2400
rect 9680 -2460 10040 -2400
rect 10300 -2460 10660 -2400
rect 11260 -2417 11271 -2383
rect 11280 -2417 11640 -2400
rect 11647 -2417 11659 -2383
rect 11260 -2423 11659 -2417
rect 11877 -2383 12277 -2380
rect 11877 -2417 11889 -2383
rect 11900 -2417 12260 -2400
rect 12265 -2417 12277 -2383
rect 11877 -2423 12277 -2417
rect 12860 -2383 13259 -2380
rect 12860 -2417 12871 -2383
rect 12880 -2417 13240 -2400
rect 13247 -2417 13259 -2383
rect 12860 -2423 13259 -2417
rect 13477 -2383 13877 -2380
rect 13477 -2417 13489 -2383
rect 13500 -2417 13860 -2400
rect 13865 -2417 13877 -2383
rect 13477 -2423 13877 -2417
rect 14459 -2383 14859 -2377
rect 14459 -2417 14471 -2383
rect 14480 -2417 14840 -2400
rect 14847 -2417 14859 -2383
rect 14459 -2423 14859 -2417
rect 15077 -2383 15477 -2377
rect 15077 -2417 15089 -2383
rect 15100 -2417 15460 -2400
rect 15465 -2417 15477 -2383
rect 15077 -2423 15477 -2417
rect 16059 -2383 16459 -2377
rect 16059 -2417 16071 -2383
rect 16080 -2417 16440 -2400
rect 16447 -2417 16459 -2383
rect 16059 -2423 16459 -2417
rect 16677 -2383 17077 -2377
rect 16677 -2417 16689 -2383
rect 16700 -2417 17060 -2400
rect 17065 -2417 17077 -2383
rect 16677 -2423 17077 -2417
rect 17659 -2383 18059 -2377
rect 17659 -2417 17671 -2383
rect 17680 -2417 18040 -2400
rect 18047 -2417 18059 -2383
rect 17659 -2423 18059 -2417
rect 18277 -2383 18677 -2377
rect 18277 -2417 18289 -2383
rect 18300 -2417 18660 -2400
rect 18665 -2417 18677 -2383
rect 18277 -2423 18677 -2417
rect 19259 -2383 19659 -2377
rect 19259 -2417 19271 -2383
rect 19280 -2417 19640 -2400
rect 19647 -2417 19659 -2383
rect 19259 -2423 19659 -2417
rect 19877 -2383 20277 -2377
rect 19877 -2417 19889 -2383
rect 19900 -2417 20260 -2400
rect 20265 -2417 20277 -2383
rect 19877 -2423 20277 -2417
rect 20859 -2383 21259 -2377
rect 20859 -2417 20871 -2383
rect 20880 -2417 21240 -2400
rect 21247 -2417 21259 -2383
rect 20859 -2423 21259 -2417
rect 21477 -2383 21877 -2377
rect 21477 -2417 21489 -2383
rect 21500 -2417 21860 -2400
rect 21865 -2417 21877 -2383
rect 21477 -2423 21877 -2417
rect 22459 -2383 22859 -2377
rect 22459 -2417 22471 -2383
rect 22480 -2417 22840 -2400
rect 22847 -2417 22859 -2383
rect 22459 -2423 22859 -2417
rect 23077 -2383 23477 -2377
rect 23077 -2417 23089 -2383
rect 23100 -2417 23460 -2400
rect 23465 -2417 23477 -2383
rect 23077 -2423 23477 -2417
rect 24059 -2383 24459 -2377
rect 24059 -2417 24071 -2383
rect 24080 -2417 24440 -2400
rect 24447 -2417 24459 -2383
rect 24059 -2423 24459 -2417
rect 24677 -2383 25077 -2377
rect 24677 -2417 24689 -2383
rect 24700 -2417 25060 -2400
rect 25065 -2417 25077 -2383
rect 24677 -2423 25077 -2417
rect 25659 -2383 26059 -2377
rect 25659 -2417 25671 -2383
rect 25680 -2417 26040 -2400
rect 26047 -2417 26059 -2383
rect 25659 -2423 26059 -2417
rect 26277 -2383 26677 -2377
rect 26277 -2417 26289 -2383
rect 26300 -2417 26660 -2400
rect 26665 -2417 26677 -2383
rect 26277 -2423 26677 -2417
rect 27259 -2383 27659 -2377
rect 27259 -2417 27271 -2383
rect 27280 -2417 27640 -2400
rect 27647 -2417 27659 -2383
rect 27259 -2423 27659 -2417
rect 27877 -2383 28277 -2377
rect 27877 -2417 27889 -2383
rect 27900 -2417 28260 -2400
rect 28265 -2417 28277 -2383
rect 27877 -2423 28277 -2417
rect 28859 -2383 29259 -2377
rect 28859 -2417 28871 -2383
rect 28880 -2417 29240 -2400
rect 29247 -2417 29259 -2383
rect 28859 -2423 29259 -2417
rect 29477 -2383 29877 -2377
rect 29477 -2417 29489 -2383
rect 29500 -2417 29860 -2400
rect 29865 -2417 29877 -2383
rect 29477 -2423 29877 -2417
rect 30459 -2383 30859 -2377
rect 30459 -2417 30471 -2383
rect 30847 -2417 30859 -2383
rect 30459 -2423 30859 -2417
rect 31077 -2383 31477 -2377
rect 31077 -2417 31089 -2383
rect 31465 -2417 31477 -2383
rect 33659 -2383 34059 -2377
rect 31077 -2423 31477 -2417
rect 32080 -2417 32440 -2400
rect 32447 -2417 32459 -2400
rect 32080 -2423 32459 -2417
rect 32677 -2417 32689 -2400
rect 32700 -2417 33060 -2400
rect 32677 -2423 33060 -2417
rect 33659 -2417 33671 -2383
rect 33680 -2417 34040 -2400
rect 34047 -2417 34059 -2383
rect 33659 -2423 34059 -2417
rect 34277 -2383 34677 -2377
rect 34277 -2417 34289 -2383
rect 34300 -2417 34660 -2400
rect 34665 -2417 34677 -2383
rect 34277 -2423 34677 -2417
rect 35259 -2383 35659 -2377
rect 35259 -2417 35271 -2383
rect 35280 -2417 35640 -2400
rect 35647 -2417 35659 -2383
rect 35259 -2423 35659 -2417
rect 35877 -2383 36277 -2377
rect 35877 -2417 35889 -2383
rect 35900 -2417 36260 -2400
rect 36265 -2417 36277 -2383
rect 35877 -2423 36277 -2417
rect 11280 -2460 11640 -2423
rect 11900 -2460 12260 -2423
rect 12880 -2460 13240 -2423
rect 13500 -2460 13860 -2423
rect 14480 -2460 14840 -2423
rect 15100 -2460 15460 -2423
rect 16080 -2460 16440 -2423
rect 16700 -2460 17060 -2423
rect 17680 -2460 18040 -2423
rect 18300 -2460 18660 -2423
rect 19280 -2460 19640 -2423
rect 19900 -2460 20260 -2423
rect 20880 -2460 21240 -2423
rect 21500 -2460 21860 -2423
rect 22480 -2460 22840 -2423
rect 23100 -2460 23460 -2423
rect 24080 -2460 24440 -2423
rect 24700 -2460 25060 -2423
rect 25680 -2460 26040 -2423
rect 26300 -2460 26660 -2423
rect 27280 -2460 27640 -2423
rect 27900 -2460 28260 -2423
rect 28880 -2460 29240 -2423
rect 29500 -2460 29860 -2423
rect 30480 -2460 30840 -2423
rect 31100 -2460 31460 -2423
rect 1400 -2470 10660 -2460
rect 1400 -2590 1410 -2470
rect 1530 -2590 3010 -2470
rect 3130 -2590 4610 -2470
rect 4730 -2590 6210 -2470
rect 6330 -2590 7810 -2470
rect 7930 -2590 9410 -2470
rect 9530 -2590 10660 -2470
rect 1400 -2600 10660 -2590
rect 11260 -2600 12260 -2460
rect 12860 -2600 13860 -2460
rect 14460 -2600 15460 -2460
rect 15590 -2470 17060 -2460
rect 15590 -2590 15600 -2470
rect 15700 -2590 17060 -2470
rect 15590 -2600 17060 -2590
rect 17190 -2470 18660 -2460
rect 17190 -2590 17200 -2470
rect 17300 -2590 18660 -2470
rect 17190 -2600 18660 -2590
rect 18790 -2470 20260 -2460
rect 18790 -2590 18800 -2470
rect 18900 -2590 20260 -2470
rect 18790 -2600 20260 -2590
rect 20390 -2470 21860 -2460
rect 20390 -2590 20400 -2470
rect 20500 -2590 21860 -2470
rect 20390 -2600 21860 -2590
rect 21990 -2470 23460 -2460
rect 21990 -2590 22000 -2470
rect 22100 -2590 23460 -2470
rect 21990 -2600 23460 -2590
rect 23590 -2470 25060 -2460
rect 23590 -2590 23600 -2470
rect 23700 -2590 25060 -2470
rect 23590 -2600 25060 -2590
rect 25190 -2470 26660 -2460
rect 25190 -2590 25200 -2470
rect 25300 -2590 26660 -2470
rect 25190 -2600 26660 -2590
rect 26791 -2470 28260 -2460
rect 26791 -2590 26800 -2470
rect 26900 -2590 28260 -2470
rect 26791 -2600 28260 -2590
rect 28390 -2470 29860 -2460
rect 28390 -2590 28400 -2470
rect 28500 -2590 29860 -2470
rect 28390 -2600 29860 -2590
rect 29990 -2470 31460 -2460
rect 29990 -2590 30000 -2470
rect 30100 -2590 31460 -2470
rect 29990 -2600 31460 -2590
rect 1680 -2660 2040 -2600
rect 2300 -2660 2660 -2600
rect 3280 -2660 3640 -2600
rect 3900 -2660 4260 -2600
rect 4880 -2660 5240 -2600
rect 5500 -2660 5860 -2600
rect 6480 -2660 6840 -2600
rect 7100 -2660 7460 -2600
rect 8080 -2660 8440 -2600
rect 8700 -2660 9060 -2600
rect 9680 -2660 10040 -2600
rect 10300 -2660 10660 -2600
rect 11280 -2645 11640 -2600
rect 11900 -2645 12260 -2600
rect 12880 -2645 13240 -2600
rect 13500 -2645 13860 -2600
rect 14480 -2645 14840 -2600
rect 15100 -2645 15460 -2600
rect 16080 -2645 16440 -2600
rect 16700 -2645 17060 -2600
rect 17680 -2645 18040 -2600
rect 18300 -2645 18660 -2600
rect 19280 -2645 19640 -2600
rect 19900 -2645 20260 -2600
rect 20880 -2645 21240 -2600
rect 21500 -2645 21860 -2600
rect 22480 -2645 22840 -2600
rect 23100 -2645 23460 -2600
rect 24080 -2645 24440 -2600
rect 24700 -2645 25060 -2600
rect 25680 -2645 26040 -2600
rect 26300 -2645 26660 -2600
rect 27280 -2645 27640 -2600
rect 27900 -2645 28260 -2600
rect 28880 -2645 29240 -2600
rect 29500 -2645 29860 -2600
rect 30480 -2645 30840 -2600
rect 31100 -2645 31460 -2600
rect 32080 -2460 32440 -2423
rect 32700 -2460 33060 -2423
rect 33680 -2460 34040 -2423
rect 34300 -2460 34660 -2423
rect 35280 -2460 35640 -2423
rect 35900 -2460 36260 -2423
rect 32080 -2600 33390 -2460
rect 33680 -2600 36260 -2460
rect 32080 -2645 32440 -2600
rect 32700 -2645 33060 -2600
rect 33680 -2645 34040 -2600
rect 34300 -2645 34660 -2600
rect 35280 -2645 35640 -2600
rect 35900 -2645 36260 -2600
rect 11260 -2651 11659 -2645
rect 1690 -2670 2030 -2660
rect 2310 -2670 2650 -2660
rect 3290 -2670 3630 -2660
rect 3910 -2670 4250 -2660
rect 4890 -2670 5230 -2660
rect 5510 -2670 5850 -2660
rect 6490 -2670 6830 -2660
rect 7110 -2670 7450 -2660
rect 8090 -2670 8430 -2660
rect 8710 -2670 9050 -2660
rect 9690 -2670 10030 -2660
rect 10310 -2670 10650 -2660
rect 11260 -2685 11271 -2651
rect 11280 -2660 11640 -2651
rect 11290 -2670 11630 -2660
rect 11647 -2685 11659 -2651
rect 11260 -2691 11659 -2685
rect 11877 -2651 12277 -2645
rect 11877 -2685 11889 -2651
rect 11900 -2660 12260 -2651
rect 11910 -2670 12250 -2660
rect 12265 -2685 12277 -2651
rect 11877 -2691 12277 -2685
rect 12860 -2651 13259 -2645
rect 12860 -2685 12871 -2651
rect 12880 -2660 13240 -2651
rect 12890 -2670 13230 -2660
rect 13247 -2685 13259 -2651
rect 12860 -2691 13259 -2685
rect 13477 -2651 13877 -2645
rect 13477 -2685 13489 -2651
rect 13500 -2660 13860 -2651
rect 13510 -2670 13850 -2660
rect 13865 -2685 13877 -2651
rect 13477 -2691 13877 -2685
rect 14459 -2651 14859 -2645
rect 14459 -2685 14471 -2651
rect 14480 -2660 14840 -2651
rect 14490 -2670 14830 -2660
rect 14847 -2685 14859 -2651
rect 14459 -2691 14859 -2685
rect 15077 -2651 15477 -2645
rect 15077 -2685 15089 -2651
rect 15100 -2660 15460 -2651
rect 15110 -2670 15450 -2660
rect 15465 -2685 15477 -2651
rect 15077 -2691 15477 -2685
rect 16059 -2651 16459 -2645
rect 16059 -2685 16071 -2651
rect 16080 -2660 16440 -2651
rect 16090 -2670 16430 -2660
rect 16447 -2685 16459 -2651
rect 16059 -2691 16459 -2685
rect 16677 -2651 17077 -2645
rect 16677 -2685 16689 -2651
rect 16700 -2660 17060 -2651
rect 16710 -2670 17050 -2660
rect 17065 -2685 17077 -2651
rect 16677 -2691 17077 -2685
rect 17659 -2651 18059 -2645
rect 17659 -2685 17671 -2651
rect 17680 -2660 18040 -2651
rect 17690 -2670 18030 -2660
rect 18047 -2685 18059 -2651
rect 17659 -2691 18059 -2685
rect 18277 -2651 18677 -2645
rect 18277 -2685 18289 -2651
rect 18300 -2660 18660 -2651
rect 18310 -2670 18650 -2660
rect 18665 -2685 18677 -2651
rect 18277 -2691 18677 -2685
rect 19259 -2651 19659 -2645
rect 19259 -2685 19271 -2651
rect 19280 -2660 19640 -2651
rect 19290 -2670 19630 -2660
rect 19647 -2685 19659 -2651
rect 19259 -2691 19659 -2685
rect 19877 -2651 20277 -2645
rect 19877 -2685 19889 -2651
rect 19900 -2660 20260 -2651
rect 19910 -2670 20250 -2660
rect 20265 -2685 20277 -2651
rect 19877 -2691 20277 -2685
rect 20859 -2651 21259 -2645
rect 20859 -2685 20871 -2651
rect 20880 -2660 21240 -2651
rect 20890 -2670 21230 -2660
rect 21247 -2685 21259 -2651
rect 20859 -2691 21259 -2685
rect 21477 -2651 21877 -2645
rect 21477 -2685 21489 -2651
rect 21500 -2660 21860 -2651
rect 21510 -2670 21850 -2660
rect 21865 -2685 21877 -2651
rect 21477 -2691 21877 -2685
rect 22459 -2651 22859 -2645
rect 22459 -2685 22471 -2651
rect 22480 -2660 22840 -2651
rect 22490 -2670 22830 -2660
rect 22847 -2685 22859 -2651
rect 22459 -2691 22859 -2685
rect 23077 -2651 23477 -2645
rect 23077 -2685 23089 -2651
rect 23100 -2660 23460 -2651
rect 23110 -2670 23450 -2660
rect 23465 -2685 23477 -2651
rect 23077 -2691 23477 -2685
rect 24059 -2651 24459 -2645
rect 24059 -2685 24071 -2651
rect 24080 -2660 24440 -2651
rect 24090 -2670 24430 -2660
rect 24447 -2685 24459 -2651
rect 24059 -2691 24459 -2685
rect 24677 -2651 25077 -2645
rect 24677 -2685 24689 -2651
rect 24700 -2660 25060 -2651
rect 24710 -2670 25050 -2660
rect 25065 -2685 25077 -2651
rect 24677 -2691 25077 -2685
rect 25659 -2651 26059 -2645
rect 25659 -2685 25671 -2651
rect 25680 -2660 26040 -2651
rect 25690 -2670 26030 -2660
rect 26047 -2685 26059 -2651
rect 25659 -2691 26059 -2685
rect 26277 -2651 26677 -2645
rect 26277 -2685 26289 -2651
rect 26300 -2660 26660 -2651
rect 26310 -2670 26650 -2660
rect 26665 -2685 26677 -2651
rect 26277 -2691 26677 -2685
rect 27259 -2651 27659 -2645
rect 27259 -2685 27271 -2651
rect 27280 -2660 27640 -2651
rect 27290 -2670 27630 -2660
rect 27647 -2685 27659 -2651
rect 27259 -2691 27659 -2685
rect 27877 -2651 28277 -2645
rect 27877 -2685 27889 -2651
rect 27900 -2660 28260 -2651
rect 27910 -2670 28250 -2660
rect 28265 -2685 28277 -2651
rect 27877 -2691 28277 -2685
rect 28859 -2651 29259 -2645
rect 28859 -2685 28871 -2651
rect 28880 -2660 29240 -2651
rect 28890 -2670 29230 -2660
rect 29247 -2685 29259 -2651
rect 28859 -2691 29259 -2685
rect 29477 -2651 29877 -2645
rect 29477 -2685 29489 -2651
rect 29500 -2660 29860 -2651
rect 29510 -2670 29850 -2660
rect 29865 -2685 29877 -2651
rect 29477 -2691 29877 -2685
rect 30459 -2651 30859 -2645
rect 30459 -2685 30471 -2651
rect 30847 -2685 30859 -2651
rect 30459 -2691 30859 -2685
rect 31077 -2651 31477 -2645
rect 31077 -2685 31089 -2651
rect 31465 -2685 31477 -2651
rect 32080 -2651 32459 -2645
rect 32080 -2660 32440 -2651
rect 32447 -2660 32459 -2651
rect 32677 -2651 33060 -2645
rect 32677 -2660 32689 -2651
rect 32700 -2660 33060 -2651
rect 33659 -2651 34059 -2645
rect 31077 -2691 31477 -2685
rect 33659 -2685 33671 -2651
rect 33680 -2660 34040 -2651
rect 34047 -2685 34059 -2651
rect 33659 -2691 34059 -2685
rect 34277 -2651 34677 -2645
rect 34277 -2685 34289 -2651
rect 34300 -2660 34660 -2651
rect 34665 -2685 34677 -2651
rect 34277 -2691 34677 -2685
rect 35259 -2651 35659 -2645
rect 35259 -2685 35271 -2651
rect 35280 -2660 35640 -2651
rect 35647 -2685 35659 -2651
rect 35259 -2691 35659 -2685
rect 35877 -2651 36277 -2645
rect 35877 -2685 35889 -2651
rect 35900 -2660 36260 -2651
rect 36265 -2685 36277 -2651
rect 35877 -2691 36277 -2685
rect 12320 -2730 12520 -2720
rect 1540 -2850 12390 -2730
rect 12510 -2850 36400 -2730
rect 1540 -2860 36400 -2850
rect 36390 -2910 36510 -2900
rect 1180 -2920 1320 -2910
rect 2780 -2920 2920 -2910
rect 4380 -2920 4520 -2910
rect 5980 -2920 6120 -2910
rect 7580 -2920 7720 -2910
rect 9180 -2920 9320 -2910
rect 11000 -2920 11140 -2910
rect 14200 -2920 14340 -2910
rect 1180 -3040 1190 -2920
rect 1310 -3040 2790 -2920
rect 2910 -3040 4390 -2920
rect 4510 -3040 5990 -2920
rect 6110 -3040 7590 -2920
rect 7710 -3040 9190 -2920
rect 9310 -3040 10720 -2920
rect 11000 -3040 11010 -2920
rect 11130 -3040 12320 -2920
rect 12820 -3040 14210 -2920
rect 14330 -3040 14340 -2920
rect 1180 -3050 1320 -3040
rect 2780 -3050 2920 -3040
rect 4380 -3050 4520 -3040
rect 5980 -3050 6120 -3040
rect 7580 -3050 7720 -3040
rect 9180 -3050 9320 -3040
rect 11000 -3050 11140 -3040
rect 14200 -3050 14340 -3040
rect 14420 -2920 14560 -2910
rect 15810 -2920 15930 -2910
rect 17410 -2920 17530 -2910
rect 19010 -2920 19130 -2910
rect 20610 -2920 20730 -2910
rect 22210 -2920 22330 -2910
rect 23810 -2920 23930 -2910
rect 25410 -2920 25530 -2910
rect 27011 -2920 27130 -2910
rect 28610 -2920 29880 -2910
rect 14420 -3040 14430 -2920
rect 14550 -3040 15520 -2920
rect 15810 -3040 15820 -2920
rect 15920 -3040 17120 -2920
rect 17410 -3040 17420 -2920
rect 17520 -3040 18720 -2920
rect 19010 -3040 19020 -2920
rect 19120 -3040 20320 -2920
rect 20610 -3040 20620 -2920
rect 20720 -3040 21920 -2920
rect 22210 -3040 22220 -2920
rect 22320 -3040 23520 -2920
rect 23810 -3040 23820 -2920
rect 23920 -3040 25120 -2920
rect 25410 -3040 25420 -2920
rect 25520 -3040 26720 -2920
rect 27011 -3040 27020 -2920
rect 27120 -3040 28320 -2920
rect 28610 -3040 28620 -2920
rect 28720 -3040 29880 -2920
rect 14420 -3050 14560 -3040
rect 15810 -3050 15930 -3040
rect 17410 -3050 17530 -3040
rect 19010 -3050 19130 -3040
rect 20610 -3050 20730 -3040
rect 22210 -3050 22330 -3040
rect 23810 -3050 23930 -3040
rect 25410 -3050 25530 -3040
rect 27011 -3050 27130 -3040
rect 28610 -3050 29880 -3040
rect 30210 -2920 30330 -2910
rect 36390 -2920 36400 -2910
rect 30210 -3040 30220 -2920
rect 30320 -3040 31480 -2920
rect 32060 -3030 36400 -2920
rect 36500 -3030 36510 -2910
rect 32060 -3040 36510 -3030
rect 30210 -3050 30330 -3040
rect -820 -3260 38090 -3160
rect -820 -3360 12520 -3260
rect 12600 -3310 13260 -3300
rect 12600 -3410 12610 -3310
rect 12730 -3360 13260 -3310
rect 13380 -3360 14120 -3260
rect 14200 -3310 14860 -3300
rect 12730 -3410 12740 -3360
rect 12600 -3420 12740 -3410
rect 2100 -3430 2240 -3420
rect 2100 -4110 2110 -3430
rect 2230 -4110 2240 -3430
rect 2100 -4120 2240 -4110
rect 3700 -3430 3840 -3420
rect 3700 -4110 3710 -3430
rect 3830 -4110 3840 -3430
rect 3700 -4120 3840 -4110
rect 5300 -3430 5440 -3420
rect 5300 -4110 5310 -3430
rect 5430 -4110 5440 -3430
rect 5300 -4120 5440 -4110
rect 6900 -3430 7040 -3420
rect 6900 -4110 6910 -3430
rect 7030 -4110 7040 -3430
rect 6900 -4120 7040 -4110
rect 8500 -3430 8640 -3420
rect 8500 -4110 8510 -3430
rect 8630 -4110 8640 -3430
rect 8500 -4120 8640 -4110
rect 10100 -3430 10240 -3420
rect 10100 -4110 10110 -3430
rect 10230 -4110 10240 -3430
rect 10100 -4120 10240 -4110
rect 11700 -3430 11840 -3420
rect 11700 -4110 11710 -3430
rect 11830 -4110 11840 -3430
rect 11700 -4120 11840 -4110
rect 13300 -3430 13440 -3420
rect 13300 -4110 13310 -3430
rect 13430 -4110 13440 -3430
rect 14200 -3430 14210 -3310
rect 14330 -3360 14860 -3310
rect 14980 -3360 38090 -3260
rect 14330 -3430 14340 -3360
rect 14200 -3440 14340 -3430
rect 14900 -3430 15040 -3420
rect 13300 -4120 13440 -4110
rect 14900 -4110 14910 -3430
rect 15030 -4110 15040 -3430
rect 14900 -4120 15040 -4110
rect 16500 -3430 16640 -3420
rect 16500 -4110 16510 -3430
rect 16630 -4110 16640 -3430
rect 16500 -4120 16640 -4110
rect 18100 -3430 18240 -3420
rect 18100 -4110 18110 -3430
rect 18230 -4110 18240 -3430
rect 18100 -4120 18240 -4110
rect 19700 -3430 19840 -3420
rect 19700 -4110 19710 -3430
rect 19830 -4110 19840 -3430
rect 19700 -4120 19840 -4110
rect 21300 -3430 21440 -3420
rect 21300 -4110 21310 -3430
rect 21430 -4110 21440 -3430
rect 21300 -4120 21440 -4110
rect 22900 -3430 23040 -3420
rect 22900 -4110 22910 -3430
rect 23030 -4110 23040 -3430
rect 22900 -4120 23040 -4110
rect 24500 -3430 24640 -3420
rect 24500 -4110 24510 -3430
rect 24630 -4110 24640 -3430
rect 24500 -4120 24640 -4110
rect 26100 -3430 26240 -3420
rect 26100 -4110 26110 -3430
rect 26230 -4110 26240 -3430
rect 26100 -4120 26240 -4110
rect 27700 -3430 27840 -3420
rect 27700 -4110 27710 -3430
rect 27830 -4110 27840 -3430
rect 27700 -4120 27840 -4110
rect 28781 -3425 28827 -3413
rect 28781 -4117 28787 -3425
rect 28821 -4117 28827 -3425
rect 28781 -4129 28827 -4117
rect 29291 -3420 29337 -3413
rect 29399 -3420 29445 -3413
rect 29291 -3425 29445 -3420
rect 29291 -4117 29297 -3425
rect 29331 -3430 29405 -3425
rect 29331 -4117 29405 -4110
rect 29439 -4117 29445 -3425
rect 29291 -4120 29445 -4117
rect 29291 -4129 29337 -4120
rect 29399 -4129 29445 -4120
rect 29909 -3425 29955 -3413
rect 29909 -4117 29915 -3425
rect 29949 -4117 29955 -3425
rect 29909 -4129 29955 -4117
rect 30381 -3425 30427 -3413
rect 30381 -4117 30387 -3425
rect 30421 -4117 30427 -3425
rect 30381 -4129 30427 -4117
rect 30891 -3420 30937 -3413
rect 30999 -3420 31045 -3413
rect 30891 -3425 31045 -3420
rect 30891 -4117 30897 -3425
rect 30931 -3430 31005 -3425
rect 30931 -4117 31005 -4110
rect 31039 -4117 31045 -3425
rect 30891 -4120 31045 -4117
rect 30891 -4129 30937 -4120
rect 30999 -4129 31045 -4120
rect 31509 -3425 31555 -3413
rect 31509 -4117 31515 -3425
rect 31549 -4117 31555 -3425
rect 31509 -4129 31555 -4117
rect 32500 -3430 32640 -3420
rect 34100 -3425 34240 -3420
rect 35700 -3425 35840 -3420
rect 34131 -3430 34205 -3425
rect 32500 -4110 32510 -3430
rect 32630 -4110 32640 -3430
rect 32500 -4120 32640 -4110
rect 34131 -4117 34205 -4110
rect 34239 -4117 34240 -3425
rect 35731 -3430 35805 -3425
rect 35731 -4117 35805 -4110
rect 35839 -4117 35840 -3425
rect 34100 -4120 34240 -4117
rect 35700 -4120 35840 -4117
rect 11260 -4183 11659 -4180
rect 1680 -4260 2040 -4200
rect 2300 -4260 2660 -4200
rect 3280 -4260 3640 -4200
rect 3900 -4260 4260 -4200
rect 4880 -4260 5240 -4200
rect 5500 -4260 5860 -4200
rect 6480 -4260 6840 -4200
rect 7100 -4260 7460 -4200
rect 8080 -4260 8440 -4200
rect 8700 -4260 9060 -4200
rect 9680 -4260 10040 -4200
rect 10300 -4260 10660 -4200
rect 11260 -4217 11271 -4183
rect 11280 -4217 11640 -4200
rect 11647 -4217 11659 -4183
rect 11260 -4223 11659 -4217
rect 11877 -4183 12277 -4180
rect 11877 -4217 11889 -4183
rect 11900 -4217 12260 -4200
rect 12265 -4217 12277 -4183
rect 12860 -4183 13259 -4180
rect 12860 -4200 12871 -4183
rect 13247 -4200 13259 -4183
rect 13477 -4183 13877 -4180
rect 13477 -4200 13489 -4183
rect 13865 -4200 13877 -4183
rect 16059 -4183 16459 -4177
rect 11877 -4223 12277 -4217
rect 11280 -4260 11640 -4223
rect 11900 -4260 12260 -4223
rect 1400 -4270 10660 -4260
rect 1400 -4390 1410 -4270
rect 1530 -4390 3010 -4270
rect 3130 -4390 4610 -4270
rect 4730 -4390 6210 -4270
rect 6330 -4390 7810 -4270
rect 7930 -4390 9410 -4270
rect 9530 -4390 10660 -4270
rect 1400 -4400 10660 -4390
rect 11260 -4400 12260 -4260
rect 12840 -4280 13880 -4200
rect 14440 -4280 15480 -4200
rect 16059 -4217 16071 -4183
rect 16080 -4217 16440 -4200
rect 16447 -4217 16459 -4183
rect 16059 -4223 16459 -4217
rect 16677 -4183 17077 -4177
rect 16677 -4217 16689 -4183
rect 16700 -4217 17060 -4200
rect 17065 -4217 17077 -4183
rect 16677 -4223 17077 -4217
rect 17659 -4183 18059 -4177
rect 17659 -4217 17671 -4183
rect 17680 -4217 18040 -4200
rect 18047 -4217 18059 -4183
rect 17659 -4223 18059 -4217
rect 18277 -4183 18677 -4177
rect 18277 -4217 18289 -4183
rect 18300 -4217 18660 -4200
rect 18665 -4217 18677 -4183
rect 18277 -4223 18677 -4217
rect 19259 -4183 19659 -4177
rect 19259 -4217 19271 -4183
rect 19280 -4217 19640 -4200
rect 19647 -4217 19659 -4183
rect 19259 -4223 19659 -4217
rect 19877 -4183 20277 -4177
rect 19877 -4217 19889 -4183
rect 19900 -4217 20260 -4200
rect 20265 -4217 20277 -4183
rect 19877 -4223 20277 -4217
rect 20859 -4183 21259 -4177
rect 20859 -4217 20871 -4183
rect 20880 -4217 21240 -4200
rect 21247 -4217 21259 -4183
rect 20859 -4223 21259 -4217
rect 21477 -4183 21877 -4177
rect 21477 -4217 21489 -4183
rect 21500 -4217 21860 -4200
rect 21865 -4217 21877 -4183
rect 21477 -4223 21877 -4217
rect 22459 -4183 22859 -4177
rect 22459 -4217 22471 -4183
rect 22480 -4217 22840 -4200
rect 22847 -4217 22859 -4183
rect 22459 -4223 22859 -4217
rect 23077 -4183 23477 -4177
rect 23077 -4217 23089 -4183
rect 23100 -4217 23460 -4200
rect 23465 -4217 23477 -4183
rect 23077 -4223 23477 -4217
rect 24059 -4183 24459 -4177
rect 24059 -4217 24071 -4183
rect 24080 -4217 24440 -4200
rect 24447 -4217 24459 -4183
rect 24059 -4223 24459 -4217
rect 24677 -4183 25077 -4177
rect 24677 -4217 24689 -4183
rect 24700 -4217 25060 -4200
rect 25065 -4217 25077 -4183
rect 24677 -4223 25077 -4217
rect 25659 -4183 26059 -4177
rect 25659 -4217 25671 -4183
rect 25680 -4217 26040 -4200
rect 26047 -4217 26059 -4183
rect 25659 -4223 26059 -4217
rect 26277 -4183 26677 -4177
rect 26277 -4217 26289 -4183
rect 26300 -4217 26660 -4200
rect 26665 -4217 26677 -4183
rect 26277 -4223 26677 -4217
rect 27259 -4183 27659 -4177
rect 27259 -4217 27271 -4183
rect 27280 -4217 27640 -4200
rect 27647 -4217 27659 -4183
rect 27259 -4223 27659 -4217
rect 27877 -4183 28277 -4177
rect 27877 -4217 27889 -4183
rect 27900 -4217 28260 -4200
rect 28265 -4217 28277 -4183
rect 27877 -4223 28277 -4217
rect 28859 -4183 29259 -4177
rect 28859 -4217 28871 -4183
rect 28880 -4217 29240 -4200
rect 29247 -4217 29259 -4183
rect 28859 -4223 29259 -4217
rect 29477 -4183 29877 -4177
rect 29477 -4217 29489 -4183
rect 29500 -4217 29860 -4200
rect 29865 -4217 29877 -4183
rect 29477 -4223 29877 -4217
rect 30459 -4183 30859 -4177
rect 30459 -4217 30471 -4183
rect 30847 -4217 30859 -4183
rect 30459 -4223 30859 -4217
rect 31077 -4183 31477 -4177
rect 31077 -4217 31089 -4183
rect 31465 -4217 31477 -4183
rect 33659 -4183 34059 -4177
rect 31077 -4223 31477 -4217
rect 32080 -4217 32440 -4200
rect 32447 -4217 32459 -4200
rect 32080 -4223 32459 -4217
rect 32677 -4217 32689 -4200
rect 32700 -4217 33060 -4200
rect 32677 -4223 33060 -4217
rect 33659 -4217 33671 -4183
rect 33680 -4217 34040 -4200
rect 34047 -4217 34059 -4183
rect 33659 -4223 34059 -4217
rect 34277 -4183 34677 -4177
rect 34277 -4217 34289 -4183
rect 34300 -4217 34660 -4200
rect 34665 -4217 34677 -4183
rect 34277 -4223 34677 -4217
rect 35259 -4183 35659 -4177
rect 35259 -4217 35271 -4183
rect 35280 -4217 35640 -4200
rect 35647 -4217 35659 -4183
rect 35259 -4223 35659 -4217
rect 35877 -4183 36277 -4177
rect 35877 -4217 35889 -4183
rect 35900 -4217 36260 -4200
rect 36265 -4217 36277 -4183
rect 35877 -4223 36277 -4217
rect 16080 -4260 16440 -4223
rect 16700 -4260 17060 -4223
rect 17680 -4260 18040 -4223
rect 18300 -4260 18660 -4223
rect 19280 -4260 19640 -4223
rect 19900 -4260 20260 -4223
rect 20880 -4260 21240 -4223
rect 21500 -4260 21860 -4223
rect 22480 -4260 22840 -4223
rect 23100 -4260 23460 -4223
rect 24080 -4260 24440 -4223
rect 24700 -4260 25060 -4223
rect 25680 -4260 26040 -4223
rect 26300 -4260 26660 -4223
rect 27280 -4260 27640 -4223
rect 27900 -4260 28260 -4223
rect 28880 -4260 29240 -4223
rect 29500 -4260 29860 -4223
rect 30480 -4260 30840 -4223
rect 31100 -4260 31460 -4223
rect 15590 -4270 17060 -4260
rect 15590 -4390 15600 -4270
rect 15700 -4390 17060 -4270
rect 1680 -4460 2040 -4400
rect 2300 -4460 2660 -4400
rect 3280 -4460 3640 -4400
rect 3900 -4460 4260 -4400
rect 4880 -4460 5240 -4400
rect 5500 -4460 5860 -4400
rect 6480 -4460 6840 -4400
rect 7100 -4460 7460 -4400
rect 8080 -4460 8440 -4400
rect 8700 -4460 9060 -4400
rect 9680 -4460 10040 -4400
rect 10300 -4460 10660 -4400
rect 11280 -4445 11640 -4400
rect 11900 -4445 12260 -4400
rect 11260 -4451 11659 -4445
rect 1690 -4470 2030 -4460
rect 2310 -4470 2650 -4460
rect 3290 -4470 3630 -4460
rect 3910 -4470 4250 -4460
rect 4890 -4470 5230 -4460
rect 5510 -4470 5850 -4460
rect 6490 -4470 6830 -4460
rect 7110 -4470 7450 -4460
rect 8090 -4470 8430 -4460
rect 8710 -4470 9050 -4460
rect 9690 -4470 10030 -4460
rect 10310 -4470 10650 -4460
rect 11260 -4485 11271 -4451
rect 11280 -4460 11640 -4451
rect 11290 -4470 11630 -4460
rect 11647 -4485 11659 -4451
rect 11260 -4491 11659 -4485
rect 11877 -4451 12277 -4445
rect 11877 -4485 11889 -4451
rect 11900 -4460 12260 -4451
rect 11910 -4470 12250 -4460
rect 12265 -4485 12277 -4451
rect 12850 -4480 13880 -4390
rect 14450 -4480 15480 -4390
rect 15590 -4400 17060 -4390
rect 17190 -4270 18660 -4260
rect 17190 -4390 17200 -4270
rect 17300 -4390 18660 -4270
rect 17190 -4400 18660 -4390
rect 18790 -4270 20260 -4260
rect 18790 -4390 18800 -4270
rect 18900 -4390 20260 -4270
rect 18790 -4400 20260 -4390
rect 20390 -4270 21860 -4260
rect 20390 -4390 20400 -4270
rect 20500 -4390 21860 -4270
rect 20390 -4400 21860 -4390
rect 21990 -4270 23460 -4260
rect 21990 -4390 22000 -4270
rect 22100 -4390 23460 -4270
rect 21990 -4400 23460 -4390
rect 23590 -4270 25060 -4260
rect 23590 -4390 23600 -4270
rect 23700 -4390 25060 -4270
rect 23590 -4400 25060 -4390
rect 25190 -4270 26660 -4260
rect 25190 -4390 25200 -4270
rect 25300 -4390 26660 -4270
rect 25190 -4400 26660 -4390
rect 26791 -4270 28260 -4260
rect 26791 -4390 26800 -4270
rect 26900 -4390 28260 -4270
rect 26791 -4400 28260 -4390
rect 28391 -4270 29860 -4260
rect 28391 -4390 28400 -4270
rect 28500 -4390 29860 -4270
rect 28391 -4400 29860 -4390
rect 29990 -4270 31460 -4260
rect 29990 -4390 30000 -4270
rect 30100 -4390 31460 -4270
rect 29990 -4400 31460 -4390
rect 16080 -4445 16440 -4400
rect 16700 -4445 17060 -4400
rect 17680 -4445 18040 -4400
rect 18300 -4445 18660 -4400
rect 19280 -4445 19640 -4400
rect 19900 -4445 20260 -4400
rect 20880 -4445 21240 -4400
rect 21500 -4445 21860 -4400
rect 22480 -4445 22840 -4400
rect 23100 -4445 23460 -4400
rect 24080 -4445 24440 -4400
rect 24700 -4445 25060 -4400
rect 25680 -4445 26040 -4400
rect 26300 -4445 26660 -4400
rect 27280 -4445 27640 -4400
rect 27900 -4445 28260 -4400
rect 28880 -4445 29240 -4400
rect 29500 -4445 29860 -4400
rect 30480 -4445 30840 -4400
rect 31100 -4445 31460 -4400
rect 32080 -4260 32440 -4223
rect 32700 -4260 33060 -4223
rect 33680 -4260 34040 -4223
rect 34300 -4260 34660 -4223
rect 35280 -4260 35640 -4223
rect 35900 -4260 36260 -4223
rect 32080 -4400 36260 -4260
rect 32080 -4445 32440 -4400
rect 32700 -4445 33060 -4400
rect 33680 -4445 34040 -4400
rect 34300 -4445 34660 -4400
rect 35280 -4445 35640 -4400
rect 35900 -4445 36260 -4400
rect 16059 -4451 16459 -4445
rect 11877 -4491 12277 -4485
rect 16059 -4485 16071 -4451
rect 16080 -4460 16440 -4451
rect 16090 -4470 16430 -4460
rect 16447 -4485 16459 -4451
rect 16059 -4491 16459 -4485
rect 16677 -4451 17077 -4445
rect 16677 -4485 16689 -4451
rect 16700 -4460 17060 -4451
rect 16710 -4470 17050 -4460
rect 17065 -4485 17077 -4451
rect 16677 -4491 17077 -4485
rect 17659 -4451 18059 -4445
rect 17659 -4485 17671 -4451
rect 17680 -4460 18040 -4451
rect 17690 -4470 18030 -4460
rect 18047 -4485 18059 -4451
rect 17659 -4491 18059 -4485
rect 18277 -4451 18677 -4445
rect 18277 -4485 18289 -4451
rect 18300 -4460 18660 -4451
rect 18310 -4470 18650 -4460
rect 18665 -4485 18677 -4451
rect 18277 -4491 18677 -4485
rect 19259 -4451 19659 -4445
rect 19259 -4485 19271 -4451
rect 19280 -4460 19640 -4451
rect 19290 -4470 19630 -4460
rect 19647 -4485 19659 -4451
rect 19259 -4491 19659 -4485
rect 19877 -4451 20277 -4445
rect 19877 -4485 19889 -4451
rect 19900 -4460 20260 -4451
rect 19910 -4470 20250 -4460
rect 20265 -4485 20277 -4451
rect 19877 -4491 20277 -4485
rect 20859 -4451 21259 -4445
rect 20859 -4485 20871 -4451
rect 20880 -4460 21240 -4451
rect 20890 -4470 21230 -4460
rect 21247 -4485 21259 -4451
rect 20859 -4491 21259 -4485
rect 21477 -4451 21877 -4445
rect 21477 -4485 21489 -4451
rect 21500 -4460 21860 -4451
rect 21510 -4470 21850 -4460
rect 21865 -4485 21877 -4451
rect 21477 -4491 21877 -4485
rect 22459 -4451 22859 -4445
rect 22459 -4485 22471 -4451
rect 22480 -4460 22840 -4451
rect 22490 -4470 22830 -4460
rect 22847 -4485 22859 -4451
rect 22459 -4491 22859 -4485
rect 23077 -4451 23477 -4445
rect 23077 -4485 23089 -4451
rect 23100 -4460 23460 -4451
rect 23110 -4470 23450 -4460
rect 23465 -4485 23477 -4451
rect 23077 -4491 23477 -4485
rect 24059 -4451 24459 -4445
rect 24059 -4485 24071 -4451
rect 24080 -4460 24440 -4451
rect 24090 -4470 24430 -4460
rect 24447 -4485 24459 -4451
rect 24059 -4491 24459 -4485
rect 24677 -4451 25077 -4445
rect 24677 -4485 24689 -4451
rect 24700 -4460 25060 -4451
rect 24710 -4470 25050 -4460
rect 25065 -4485 25077 -4451
rect 24677 -4491 25077 -4485
rect 25659 -4451 26059 -4445
rect 25659 -4485 25671 -4451
rect 25680 -4460 26040 -4451
rect 25690 -4470 26030 -4460
rect 26047 -4485 26059 -4451
rect 25659 -4491 26059 -4485
rect 26277 -4451 26677 -4445
rect 26277 -4485 26289 -4451
rect 26300 -4460 26660 -4451
rect 26310 -4470 26650 -4460
rect 26665 -4485 26677 -4451
rect 26277 -4491 26677 -4485
rect 27259 -4451 27659 -4445
rect 27259 -4485 27271 -4451
rect 27280 -4460 27640 -4451
rect 27290 -4470 27630 -4460
rect 27647 -4485 27659 -4451
rect 27259 -4491 27659 -4485
rect 27877 -4451 28277 -4445
rect 27877 -4485 27889 -4451
rect 27900 -4460 28260 -4451
rect 27910 -4470 28250 -4460
rect 28265 -4485 28277 -4451
rect 27877 -4491 28277 -4485
rect 28859 -4451 29259 -4445
rect 28859 -4485 28871 -4451
rect 28880 -4460 29240 -4451
rect 28890 -4470 29230 -4460
rect 29247 -4485 29259 -4451
rect 28859 -4491 29259 -4485
rect 29477 -4451 29877 -4445
rect 29477 -4485 29489 -4451
rect 29500 -4460 29860 -4451
rect 29510 -4470 29850 -4460
rect 29865 -4485 29877 -4451
rect 29477 -4491 29877 -4485
rect 30459 -4451 30859 -4445
rect 30459 -4485 30471 -4451
rect 30847 -4485 30859 -4451
rect 30459 -4491 30859 -4485
rect 31077 -4451 31477 -4445
rect 31077 -4485 31089 -4451
rect 31465 -4485 31477 -4451
rect 32080 -4451 32459 -4445
rect 32080 -4460 32440 -4451
rect 32447 -4460 32459 -4451
rect 32677 -4451 33060 -4445
rect 32677 -4460 32689 -4451
rect 32700 -4460 33060 -4451
rect 33659 -4451 34059 -4445
rect 31077 -4491 31477 -4485
rect 33659 -4485 33671 -4451
rect 33680 -4460 34040 -4451
rect 34047 -4485 34059 -4451
rect 33659 -4491 34059 -4485
rect 34277 -4451 34677 -4445
rect 34277 -4485 34289 -4451
rect 34300 -4460 34660 -4451
rect 34665 -4485 34677 -4451
rect 34277 -4491 34677 -4485
rect 35259 -4451 35659 -4445
rect 35259 -4485 35271 -4451
rect 35280 -4460 35640 -4451
rect 35647 -4485 35659 -4451
rect 35259 -4491 35659 -4485
rect 35877 -4451 36277 -4445
rect 35877 -4485 35889 -4451
rect 35900 -4460 36260 -4451
rect 36265 -4485 36277 -4451
rect 35877 -4491 36277 -4485
rect 12320 -4530 12520 -4520
rect 1540 -4650 12390 -4530
rect 12510 -4650 36400 -4530
rect 1540 -4660 36400 -4650
rect 30459 -4709 30859 -4703
rect 1180 -4720 1320 -4710
rect 2780 -4720 2920 -4710
rect 4380 -4720 4520 -4710
rect 5980 -4720 6120 -4710
rect 7580 -4720 7720 -4710
rect 9180 -4720 9320 -4710
rect 15810 -4720 15930 -4710
rect 17410 -4720 17530 -4710
rect 19010 -4720 19130 -4710
rect 20610 -4720 20730 -4710
rect 22210 -4720 22330 -4710
rect 23810 -4720 23930 -4710
rect 25410 -4720 25530 -4710
rect 27011 -4720 27130 -4710
rect 28611 -4720 28730 -4710
rect 30211 -4720 30330 -4710
rect 30459 -4720 30471 -4709
rect 30847 -4720 30859 -4709
rect 31077 -4709 31477 -4703
rect 31077 -4720 31089 -4709
rect 1180 -4840 1190 -4720
rect 1310 -4840 2790 -4720
rect 2910 -4840 4390 -4720
rect 4510 -4840 5990 -4720
rect 6110 -4840 7590 -4720
rect 7710 -4840 9190 -4720
rect 9310 -4840 10720 -4720
rect 11220 -4810 12350 -4720
rect 11220 -4840 11710 -4810
rect 1180 -4850 1320 -4840
rect 2780 -4850 2920 -4840
rect 4380 -4850 4520 -4840
rect 5980 -4850 6120 -4840
rect 7580 -4850 7720 -4840
rect 9180 -4850 9320 -4840
rect 11700 -4930 11710 -4840
rect 11830 -4840 12350 -4810
rect 12600 -4730 12740 -4720
rect 11830 -4930 11840 -4840
rect 12600 -4850 12610 -4730
rect 12730 -4740 12740 -4730
rect 12730 -4840 13260 -4740
rect 13470 -4790 13890 -4720
rect 13470 -4840 13630 -4790
rect 12730 -4850 12740 -4840
rect 12600 -4860 12740 -4850
rect 13620 -4910 13630 -4840
rect 13750 -4840 13890 -4790
rect 14200 -4730 14340 -4720
rect 13750 -4910 13760 -4840
rect 14200 -4850 14210 -4730
rect 14330 -4740 14340 -4730
rect 14330 -4840 14860 -4740
rect 15070 -4790 15490 -4720
rect 15070 -4840 15230 -4790
rect 14330 -4850 14340 -4840
rect 14200 -4860 14340 -4850
rect 13620 -4920 13760 -4910
rect 15220 -4910 15230 -4840
rect 15350 -4840 15490 -4790
rect 15810 -4840 15820 -4720
rect 15920 -4840 17120 -4720
rect 17410 -4840 17420 -4720
rect 17520 -4840 18720 -4720
rect 19010 -4840 19020 -4720
rect 19120 -4840 20320 -4720
rect 20610 -4840 20620 -4720
rect 20720 -4840 21920 -4720
rect 22210 -4840 22220 -4720
rect 22320 -4840 23520 -4720
rect 23810 -4840 23820 -4720
rect 23920 -4840 25120 -4720
rect 25410 -4840 25420 -4720
rect 25520 -4840 26720 -4720
rect 27011 -4840 27020 -4720
rect 27120 -4840 28320 -4720
rect 28611 -4840 28620 -4720
rect 28720 -4840 29920 -4720
rect 30211 -4840 30220 -4720
rect 30320 -4743 31089 -4720
rect 31465 -4720 31477 -4709
rect 36390 -4710 36510 -4700
rect 36390 -4720 36400 -4710
rect 31465 -4743 31520 -4720
rect 30320 -4840 31520 -4743
rect 32060 -4830 36400 -4720
rect 36500 -4830 36510 -4710
rect 32060 -4840 36510 -4830
rect 15350 -4910 15360 -4840
rect 15810 -4850 15930 -4840
rect 17410 -4850 17530 -4840
rect 19010 -4850 19130 -4840
rect 20610 -4850 20730 -4840
rect 22210 -4850 22330 -4840
rect 23810 -4850 23930 -4840
rect 25410 -4850 25530 -4840
rect 27011 -4850 27130 -4840
rect 28611 -4850 28730 -4840
rect 30211 -4850 30330 -4840
rect 15220 -4920 15360 -4910
rect 11700 -4940 11840 -4930
rect 11700 -5830 11840 -5820
rect 11700 -5950 11710 -5830
rect 11830 -5840 11840 -5830
rect 13300 -5830 13440 -5820
rect 13300 -5840 13310 -5830
rect 11830 -5940 13310 -5840
rect 11830 -5950 11840 -5940
rect 11700 -5960 11840 -5950
rect 13300 -5950 13310 -5940
rect 13430 -5950 13440 -5830
rect 13300 -5960 13440 -5950
rect 11700 -6050 11840 -6040
rect 11700 -6170 11710 -6050
rect 11830 -6060 11840 -6050
rect 13620 -6050 13760 -6040
rect 13620 -6060 13630 -6050
rect 11830 -6160 13630 -6060
rect 11830 -6170 11840 -6160
rect 11700 -6180 11840 -6170
rect 13620 -6170 13630 -6160
rect 13750 -6170 13760 -6050
rect 13620 -6180 13760 -6170
rect 14220 -6050 14360 -6040
rect 14220 -6170 14230 -6050
rect 14350 -6060 14360 -6050
rect 15220 -6050 15360 -6040
rect 15220 -6060 15230 -6050
rect 14350 -6160 15230 -6060
rect 14350 -6170 14360 -6160
rect 14220 -6180 14360 -6170
rect 15220 -6170 15230 -6160
rect 15350 -6170 15360 -6050
rect 15220 -6180 15360 -6170
rect 12620 -6270 12760 -6260
rect 12620 -6390 12630 -6270
rect 12750 -6280 12760 -6270
rect 16500 -6270 16640 -6260
rect 16500 -6280 16510 -6270
rect 12750 -6380 16510 -6280
rect 12750 -6390 12760 -6380
rect 12620 -6400 12760 -6390
rect 16500 -6390 16510 -6380
rect 16630 -6390 16640 -6270
rect 16500 -6400 16640 -6390
rect 12400 -6490 12540 -6480
rect 12400 -6610 12410 -6490
rect 12530 -6500 12540 -6490
rect 14900 -6490 15040 -6480
rect 14900 -6500 14910 -6490
rect 12530 -6600 14910 -6500
rect 12530 -6610 12540 -6600
rect 12400 -6620 12540 -6610
rect 14900 -6610 14910 -6600
rect 15030 -6610 15040 -6490
rect 14900 -6620 15040 -6610
rect 1200 -8070 1340 -8060
rect 1200 -8190 1210 -8070
rect 1330 -8080 1340 -8070
rect 2800 -8070 2940 -8060
rect 2800 -8080 2810 -8070
rect 1330 -8180 2810 -8080
rect 1330 -8190 1340 -8180
rect 1200 -8200 1340 -8190
rect 2800 -8190 2810 -8180
rect 2930 -8080 2940 -8070
rect 4400 -8070 4540 -8060
rect 4400 -8080 4410 -8070
rect 2930 -8180 4410 -8080
rect 2930 -8190 2940 -8180
rect 2800 -8200 2940 -8190
rect 4400 -8190 4410 -8180
rect 4530 -8080 4540 -8070
rect 6000 -8070 6140 -8060
rect 6000 -8080 6010 -8070
rect 4530 -8180 6010 -8080
rect 4530 -8190 4540 -8180
rect 4400 -8200 4540 -8190
rect 6000 -8190 6010 -8180
rect 6130 -8080 6140 -8070
rect 7600 -8070 7740 -8060
rect 7600 -8080 7610 -8070
rect 6130 -8180 7610 -8080
rect 6130 -8190 6140 -8180
rect 6000 -8200 6140 -8190
rect 7600 -8190 7610 -8180
rect 7730 -8080 7740 -8070
rect 9200 -8070 9340 -8060
rect 9200 -8080 9210 -8070
rect 7730 -8180 9210 -8080
rect 7730 -8190 7740 -8180
rect 7600 -8200 7740 -8190
rect 9200 -8190 9210 -8180
rect 9330 -8080 9340 -8070
rect 15820 -8070 15960 -8060
rect 9330 -8180 10700 -8080
rect 11270 -8110 15480 -8100
rect 9330 -8190 9340 -8180
rect 9200 -8200 9340 -8190
rect 11270 -8200 11710 -8110
rect 11690 -8230 11710 -8200
rect 11840 -8200 15480 -8110
rect 15820 -8190 15830 -8070
rect 15950 -8100 15960 -8070
rect 17420 -8070 17560 -8060
rect 15950 -8190 17090 -8100
rect 15820 -8200 17090 -8190
rect 17420 -8190 17430 -8070
rect 17550 -8100 17560 -8070
rect 19020 -8070 19160 -8060
rect 17550 -8190 18690 -8100
rect 17420 -8200 18690 -8190
rect 19020 -8190 19030 -8070
rect 19150 -8100 19160 -8070
rect 20620 -8070 20760 -8060
rect 19150 -8190 20290 -8100
rect 19020 -8200 20290 -8190
rect 20620 -8190 20630 -8070
rect 20750 -8100 20760 -8070
rect 22220 -8070 22360 -8060
rect 20750 -8190 21890 -8100
rect 20620 -8200 21890 -8190
rect 22220 -8190 22230 -8070
rect 22350 -8100 22360 -8070
rect 23820 -8070 23960 -8060
rect 22350 -8190 23490 -8100
rect 22220 -8200 23490 -8190
rect 23820 -8190 23830 -8070
rect 23950 -8100 23960 -8070
rect 25420 -8070 25560 -8060
rect 23950 -8190 25090 -8100
rect 23820 -8200 25090 -8190
rect 25420 -8190 25430 -8070
rect 25550 -8100 25560 -8070
rect 27020 -8070 27160 -8060
rect 25550 -8190 26680 -8100
rect 25420 -8200 26680 -8190
rect 27020 -8190 27030 -8070
rect 27150 -8100 27160 -8070
rect 28620 -8070 28760 -8060
rect 27150 -8190 28290 -8100
rect 27020 -8200 28290 -8190
rect 28620 -8190 28630 -8070
rect 28750 -8100 28760 -8070
rect 30220 -8070 30360 -8060
rect 28750 -8190 29890 -8100
rect 28620 -8200 29890 -8190
rect 30220 -8190 30230 -8070
rect 30350 -8100 30360 -8070
rect 30350 -8164 31490 -8100
rect 30350 -8190 31493 -8164
rect 30220 -8200 31493 -8190
rect 11840 -8230 11860 -8200
rect 11690 -8240 11860 -8230
rect 13290 -8240 13460 -8200
rect 14890 -8240 15060 -8200
rect 30457 -8204 30469 -8200
rect 30845 -8204 30857 -8200
rect 30457 -8210 30857 -8204
rect 31093 -8204 31105 -8200
rect 31481 -8204 31493 -8200
rect 31093 -8210 31493 -8204
rect 1560 -8380 10790 -8260
rect 11180 -8390 15570 -8240
rect 30370 -8249 30416 -8237
rect 30370 -8260 30376 -8249
rect 30410 -8260 30416 -8249
rect 30898 -8249 30944 -8237
rect 30898 -8260 30904 -8249
rect 30938 -8260 30944 -8249
rect 31006 -8249 31052 -8237
rect 31006 -8260 31012 -8249
rect 31046 -8260 31052 -8249
rect 31534 -8249 31560 -8237
rect 31534 -8260 31540 -8249
rect 15970 -8380 33200 -8260
rect 30370 -8383 30376 -8380
rect 30410 -8383 30416 -8380
rect 30370 -8395 30416 -8383
rect 30898 -8383 30904 -8380
rect 30938 -8383 30944 -8380
rect 30898 -8395 30944 -8383
rect 31006 -8383 31012 -8380
rect 31046 -8383 31052 -8380
rect 31006 -8395 31052 -8383
rect 31534 -8383 31540 -8380
rect 31534 -8395 31560 -8383
rect 30457 -8428 30857 -8422
rect 30457 -8430 30469 -8428
rect 30845 -8430 30857 -8428
rect 1420 -8510 1560 -8500
rect 1420 -8630 1430 -8510
rect 1550 -8520 1560 -8510
rect 1660 -8520 2060 -8430
rect 2290 -8520 2690 -8430
rect 3020 -8510 3160 -8500
rect 3020 -8520 3030 -8510
rect 1550 -8620 3030 -8520
rect 1550 -8630 1560 -8620
rect 1420 -8640 1560 -8630
rect 1660 -8640 2690 -8620
rect 3020 -8630 3030 -8620
rect 3150 -8520 3160 -8510
rect 3260 -8520 3660 -8430
rect 3890 -8520 4290 -8430
rect 4620 -8510 4760 -8500
rect 4620 -8520 4630 -8510
rect 3150 -8620 4630 -8520
rect 3150 -8630 3160 -8620
rect 3020 -8640 3160 -8630
rect 3260 -8640 4290 -8620
rect 4620 -8630 4630 -8620
rect 4750 -8520 4760 -8510
rect 4860 -8520 5260 -8430
rect 5490 -8520 5890 -8430
rect 6220 -8510 6360 -8500
rect 6220 -8520 6230 -8510
rect 4750 -8620 6230 -8520
rect 4750 -8630 4760 -8620
rect 4620 -8640 4760 -8630
rect 4860 -8640 5890 -8620
rect 6220 -8630 6230 -8620
rect 6350 -8520 6360 -8510
rect 6460 -8520 6860 -8430
rect 7090 -8520 7490 -8430
rect 7820 -8510 7960 -8500
rect 7820 -8520 7830 -8510
rect 6350 -8620 7830 -8520
rect 6350 -8630 6360 -8620
rect 6220 -8640 6360 -8630
rect 6460 -8640 7490 -8620
rect 7820 -8630 7830 -8620
rect 7950 -8520 7960 -8510
rect 8060 -8520 8460 -8430
rect 8690 -8520 9090 -8430
rect 9420 -8510 9560 -8500
rect 9420 -8520 9430 -8510
rect 7950 -8620 9430 -8520
rect 7950 -8630 7960 -8620
rect 7820 -8640 7960 -8630
rect 8060 -8640 9090 -8620
rect 9420 -8630 9430 -8620
rect 9550 -8520 9560 -8510
rect 9660 -8520 10060 -8430
rect 10290 -8520 10690 -8430
rect 11260 -8490 15490 -8430
rect 9550 -8620 10690 -8520
rect 9550 -8630 9560 -8620
rect 9420 -8640 9560 -8630
rect 9660 -8640 10690 -8620
rect 1660 -8730 2060 -8640
rect 2290 -8730 2690 -8640
rect 3260 -8730 3660 -8640
rect 3890 -8730 4290 -8640
rect 4860 -8730 5260 -8640
rect 5490 -8730 5890 -8640
rect 6460 -8730 6860 -8640
rect 7090 -8730 7490 -8640
rect 8060 -8730 8460 -8640
rect 8690 -8730 9090 -8640
rect 9660 -8730 10060 -8640
rect 10290 -8730 10690 -8640
rect 11420 -8650 11480 -8490
rect 12070 -8650 12130 -8490
rect 11260 -8730 12290 -8650
rect 2120 -8810 2240 -8800
rect 2120 -9470 2130 -8810
rect 2230 -9470 2240 -8810
rect 2120 -9480 2240 -9470
rect 3720 -8810 3840 -8800
rect 3720 -9470 3730 -8810
rect 3830 -9470 3840 -8810
rect 3720 -9480 3840 -9470
rect 5320 -8810 5440 -8800
rect 5320 -9470 5330 -8810
rect 5430 -9470 5440 -8810
rect 5320 -9480 5440 -9470
rect 6920 -8810 7040 -8800
rect 6920 -9470 6930 -8810
rect 7030 -9470 7040 -8810
rect 6920 -9480 7040 -9470
rect 8520 -8810 8640 -8800
rect 8520 -9470 8530 -8810
rect 8630 -9470 8640 -8810
rect 8520 -9480 8640 -9470
rect 10120 -8810 10240 -8800
rect 10120 -9470 10130 -8810
rect 10230 -9470 10240 -8810
rect 10120 -9480 10240 -9470
rect 11710 -8810 11840 -8800
rect 11710 -9470 11720 -8810
rect 11830 -9470 11840 -8810
rect 11710 -9480 11840 -9470
rect 12480 -9550 12680 -8490
rect 15600 -8520 15740 -8510
rect 12860 -8730 15490 -8630
rect 15600 -8640 15610 -8520
rect 15730 -8530 15740 -8520
rect 16060 -8530 16450 -8430
rect 16700 -8530 17090 -8430
rect 15730 -8630 17090 -8530
rect 15730 -8640 15740 -8630
rect 15600 -8650 15740 -8640
rect 16060 -8730 16450 -8630
rect 16700 -8730 17090 -8630
rect 17200 -8520 17340 -8510
rect 17200 -8640 17210 -8520
rect 17330 -8530 17340 -8520
rect 17660 -8530 18050 -8430
rect 18300 -8530 18690 -8430
rect 17330 -8630 18690 -8530
rect 17330 -8640 17340 -8630
rect 17200 -8650 17340 -8640
rect 17660 -8730 18050 -8630
rect 18300 -8730 18690 -8630
rect 18800 -8520 18940 -8510
rect 18800 -8640 18810 -8520
rect 18930 -8530 18940 -8520
rect 19260 -8530 19650 -8430
rect 19900 -8530 20290 -8430
rect 18930 -8630 20290 -8530
rect 18930 -8640 18940 -8630
rect 18800 -8650 18940 -8640
rect 19260 -8730 19650 -8630
rect 19900 -8730 20290 -8630
rect 20400 -8520 20540 -8510
rect 20400 -8640 20410 -8520
rect 20530 -8530 20540 -8520
rect 20860 -8530 21250 -8430
rect 21500 -8530 21890 -8430
rect 20530 -8630 21890 -8530
rect 20530 -8640 20540 -8630
rect 20400 -8650 20540 -8640
rect 20860 -8730 21250 -8630
rect 21500 -8730 21890 -8630
rect 22000 -8520 22140 -8510
rect 22000 -8640 22010 -8520
rect 22130 -8530 22140 -8520
rect 22460 -8530 22850 -8430
rect 23100 -8530 23490 -8430
rect 22130 -8630 23490 -8530
rect 22130 -8640 22140 -8630
rect 22000 -8650 22140 -8640
rect 22460 -8730 22850 -8630
rect 23100 -8730 23490 -8630
rect 23600 -8520 23740 -8510
rect 23600 -8640 23610 -8520
rect 23730 -8530 23740 -8520
rect 24060 -8530 24450 -8430
rect 24700 -8530 25090 -8430
rect 23730 -8630 25090 -8530
rect 23730 -8640 23740 -8630
rect 23600 -8650 23740 -8640
rect 24060 -8730 24450 -8630
rect 24700 -8730 25090 -8630
rect 25200 -8520 25340 -8510
rect 25200 -8640 25210 -8520
rect 25330 -8530 25340 -8520
rect 25660 -8530 26050 -8430
rect 26300 -8530 26690 -8430
rect 27260 -8468 27657 -8430
rect 27893 -8468 28290 -8430
rect 25330 -8630 26690 -8530
rect 25330 -8640 25340 -8630
rect 25200 -8650 25340 -8640
rect 25660 -8730 26050 -8630
rect 26300 -8730 26690 -8630
rect 26800 -8520 26940 -8510
rect 26800 -8640 26810 -8520
rect 26930 -8530 26940 -8520
rect 27260 -8530 27650 -8468
rect 27900 -8530 28290 -8468
rect 28860 -8468 29257 -8430
rect 29493 -8468 29890 -8430
rect 30457 -8468 30857 -8430
rect 31093 -8428 31493 -8422
rect 31093 -8430 31105 -8428
rect 31481 -8430 31493 -8428
rect 31093 -8468 31493 -8430
rect 26930 -8630 28290 -8530
rect 26930 -8640 26940 -8630
rect 26800 -8650 26940 -8640
rect 27260 -8690 27650 -8630
rect 27900 -8690 28290 -8630
rect 28400 -8520 28540 -8510
rect 28400 -8640 28410 -8520
rect 28530 -8530 28540 -8520
rect 28860 -8530 29250 -8468
rect 29500 -8530 29890 -8468
rect 28530 -8630 29890 -8530
rect 28530 -8640 28540 -8630
rect 28400 -8650 28540 -8640
rect 27260 -8730 27657 -8690
rect 27893 -8730 28290 -8690
rect 28860 -8690 29250 -8630
rect 29500 -8690 29890 -8630
rect 30000 -8520 30140 -8510
rect 30000 -8640 30010 -8520
rect 30130 -8530 30140 -8520
rect 30460 -8530 30850 -8468
rect 31100 -8530 31490 -8468
rect 30130 -8630 31490 -8530
rect 30130 -8640 30140 -8630
rect 30000 -8650 30140 -8640
rect 28860 -8730 29257 -8690
rect 29493 -8730 29890 -8690
rect 30460 -8690 30850 -8630
rect 31100 -8690 31490 -8630
rect 30460 -8730 30857 -8690
rect 31093 -8730 31490 -8690
rect 13310 -8810 13440 -8730
rect 13310 -9470 13320 -8810
rect 13430 -9470 13440 -8810
rect 13310 -9480 13440 -9470
rect 14910 -8810 15040 -8730
rect 14910 -9470 14920 -8810
rect 15030 -9470 15040 -8810
rect 14910 -9480 15040 -9470
rect 16510 -8800 16640 -8790
rect 16510 -9480 16520 -8800
rect 16630 -9480 16640 -8800
rect 16510 -9490 16640 -9480
rect 18110 -8800 18240 -8790
rect 18110 -9480 18120 -8800
rect 18230 -9480 18240 -8800
rect 18110 -9490 18240 -9480
rect 19710 -8800 19840 -8790
rect 19710 -9480 19720 -8800
rect 19830 -9480 19840 -8800
rect 19710 -9490 19840 -9480
rect 21310 -8800 21440 -8790
rect 21310 -9480 21320 -8800
rect 21430 -9480 21440 -8800
rect 21310 -9490 21440 -9480
rect 22910 -8800 23040 -8790
rect 22910 -9480 22920 -8800
rect 23030 -9480 23040 -8800
rect 22910 -9490 23040 -9480
rect 24510 -8800 24640 -8790
rect 24510 -9480 24520 -8800
rect 24630 -9480 24640 -8800
rect 24510 -9490 24640 -9480
rect 26110 -8800 26240 -8790
rect 26110 -9480 26120 -8800
rect 26230 -9480 26240 -8800
rect 26110 -9490 26240 -9480
rect 27710 -8800 27840 -8790
rect 27710 -9480 27720 -8800
rect 27830 -9480 27840 -8800
rect 27710 -9490 27840 -9480
rect 29310 -8800 29440 -8790
rect 29310 -9480 29320 -8800
rect 29430 -9480 29440 -8800
rect 29310 -9490 29440 -9480
rect 30910 -8800 31040 -8790
rect 30910 -9480 30920 -8800
rect 31030 -9480 31040 -8800
rect 30910 -9490 31040 -9480
rect -960 -9670 12390 -9560
rect 12480 -9620 15490 -9550
rect 15680 -9670 36260 -9560
rect -960 -9760 36260 -9670
rect 1200 -9870 1340 -9860
rect 1200 -9990 1210 -9870
rect 1330 -9880 1340 -9870
rect 2800 -9870 2940 -9860
rect 2800 -9880 2810 -9870
rect 1330 -9980 2810 -9880
rect 1330 -9990 1340 -9980
rect 1200 -10000 1340 -9990
rect 2800 -9990 2810 -9980
rect 2930 -9880 2940 -9870
rect 4400 -9870 4540 -9860
rect 4400 -9880 4410 -9870
rect 2930 -9980 4410 -9880
rect 2930 -9990 2940 -9980
rect 2800 -10000 2940 -9990
rect 4400 -9990 4410 -9980
rect 4530 -9880 4540 -9870
rect 6000 -9870 6140 -9860
rect 6000 -9880 6010 -9870
rect 4530 -9980 6010 -9880
rect 4530 -9990 4540 -9980
rect 4400 -10000 4540 -9990
rect 6000 -9990 6010 -9980
rect 6130 -9880 6140 -9870
rect 7600 -9870 7740 -9860
rect 7600 -9880 7610 -9870
rect 6130 -9980 7610 -9880
rect 6130 -9990 6140 -9980
rect 6000 -10000 6140 -9990
rect 7600 -9990 7610 -9980
rect 7730 -9880 7740 -9870
rect 9200 -9870 9340 -9860
rect 9200 -9880 9210 -9870
rect 7730 -9980 9210 -9880
rect 7730 -9990 7740 -9980
rect 7600 -10000 7740 -9990
rect 9200 -9990 9210 -9980
rect 9330 -9880 9340 -9870
rect 15820 -9870 15960 -9860
rect 9330 -9980 10700 -9880
rect 9330 -9990 9340 -9980
rect 9200 -10000 9340 -9990
rect 15820 -9990 15830 -9870
rect 15950 -9900 15960 -9870
rect 17420 -9870 17560 -9860
rect 15950 -9990 17090 -9900
rect 15820 -10000 17090 -9990
rect 17420 -9990 17430 -9870
rect 17550 -9900 17560 -9870
rect 19020 -9870 19160 -9860
rect 17550 -9990 18690 -9900
rect 17420 -10000 18690 -9990
rect 19020 -9990 19030 -9870
rect 19150 -9900 19160 -9870
rect 20620 -9870 20760 -9860
rect 19150 -9990 20290 -9900
rect 19020 -10000 20290 -9990
rect 20620 -9990 20630 -9870
rect 20750 -9900 20760 -9870
rect 22220 -9870 22360 -9860
rect 20750 -9990 21890 -9900
rect 20620 -10000 21890 -9990
rect 22220 -9990 22230 -9870
rect 22350 -9900 22360 -9870
rect 23820 -9870 23960 -9860
rect 22350 -9990 23490 -9900
rect 22220 -10000 23490 -9990
rect 23820 -9990 23830 -9870
rect 23950 -9900 23960 -9870
rect 25420 -9870 25560 -9860
rect 23950 -9990 25090 -9900
rect 23820 -10000 25090 -9990
rect 25420 -9990 25430 -9870
rect 25550 -9900 25560 -9870
rect 27020 -9870 27160 -9860
rect 25550 -9990 26680 -9900
rect 25420 -10000 26680 -9990
rect 27020 -9990 27030 -9870
rect 27150 -9900 27160 -9870
rect 28620 -9870 28760 -9860
rect 27150 -9990 28290 -9900
rect 27020 -10000 28290 -9990
rect 28620 -9990 28630 -9870
rect 28750 -9900 28760 -9870
rect 30220 -9870 30360 -9860
rect 28750 -9990 29890 -9900
rect 28620 -10000 29890 -9990
rect 30220 -9990 30230 -9870
rect 30350 -9900 30360 -9870
rect 30350 -9964 31490 -9900
rect 30350 -9990 31493 -9964
rect 30220 -10000 31493 -9990
rect 30457 -10004 30469 -10000
rect 30845 -10004 30857 -10000
rect 30457 -10010 30857 -10004
rect 31093 -10004 31105 -10000
rect 31481 -10004 31493 -10000
rect 31093 -10010 31493 -10004
rect 30370 -10049 30416 -10037
rect 30370 -10060 30376 -10049
rect 30410 -10060 30416 -10049
rect 30898 -10049 30944 -10037
rect 30898 -10060 30904 -10049
rect 30938 -10060 30944 -10049
rect 31006 -10049 31052 -10037
rect 31006 -10060 31012 -10049
rect 31046 -10060 31052 -10049
rect 31534 -10049 31560 -10037
rect 31534 -10060 31540 -10049
rect 1560 -10180 33200 -10060
rect 30370 -10183 30376 -10180
rect 30410 -10183 30416 -10180
rect 30370 -10195 30416 -10183
rect 30898 -10183 30904 -10180
rect 30938 -10183 30944 -10180
rect 30898 -10195 30944 -10183
rect 31006 -10183 31012 -10180
rect 31046 -10183 31052 -10180
rect 31006 -10195 31052 -10183
rect 31534 -10183 31540 -10180
rect 31534 -10195 31560 -10183
rect 30457 -10228 30857 -10222
rect 30457 -10230 30469 -10228
rect 30845 -10230 30857 -10228
rect 1420 -10310 1560 -10300
rect 1420 -10430 1430 -10310
rect 1550 -10320 1560 -10310
rect 1660 -10320 2060 -10230
rect 2290 -10320 2690 -10230
rect 3020 -10310 3160 -10300
rect 3020 -10320 3030 -10310
rect 1550 -10420 3030 -10320
rect 1550 -10430 1560 -10420
rect 1420 -10440 1560 -10430
rect 1660 -10440 2690 -10420
rect 3020 -10430 3030 -10420
rect 3150 -10320 3160 -10310
rect 3260 -10320 3660 -10230
rect 3890 -10320 4290 -10230
rect 4620 -10310 4760 -10300
rect 4620 -10320 4630 -10310
rect 3150 -10420 4630 -10320
rect 3150 -10430 3160 -10420
rect 3020 -10440 3160 -10430
rect 3260 -10440 4290 -10420
rect 4620 -10430 4630 -10420
rect 4750 -10320 4760 -10310
rect 4860 -10320 5260 -10230
rect 5490 -10320 5890 -10230
rect 6220 -10310 6360 -10300
rect 6220 -10320 6230 -10310
rect 4750 -10420 6230 -10320
rect 4750 -10430 4760 -10420
rect 4620 -10440 4760 -10430
rect 4860 -10440 5890 -10420
rect 6220 -10430 6230 -10420
rect 6350 -10320 6360 -10310
rect 6460 -10320 6860 -10230
rect 7090 -10320 7490 -10230
rect 7820 -10310 7960 -10300
rect 7820 -10320 7830 -10310
rect 6350 -10420 7830 -10320
rect 6350 -10430 6360 -10420
rect 6220 -10440 6360 -10430
rect 6460 -10440 7490 -10420
rect 7820 -10430 7830 -10420
rect 7950 -10320 7960 -10310
rect 8060 -10320 8460 -10230
rect 8690 -10320 9090 -10230
rect 9420 -10310 9560 -10300
rect 9420 -10320 9430 -10310
rect 7950 -10420 9430 -10320
rect 7950 -10430 7960 -10420
rect 7820 -10440 7960 -10430
rect 8060 -10440 9090 -10420
rect 9420 -10430 9430 -10420
rect 9550 -10320 9560 -10310
rect 9660 -10320 10060 -10230
rect 10290 -10320 10690 -10230
rect 9550 -10420 10690 -10320
rect 15600 -10320 15740 -10310
rect 9550 -10430 9560 -10420
rect 9420 -10440 9560 -10430
rect 9660 -10440 10690 -10420
rect 1660 -10530 2060 -10440
rect 2290 -10530 2690 -10440
rect 3260 -10530 3660 -10440
rect 3890 -10530 4290 -10440
rect 4860 -10530 5260 -10440
rect 5490 -10530 5890 -10440
rect 6460 -10530 6860 -10440
rect 7090 -10530 7490 -10440
rect 8060 -10530 8460 -10440
rect 8690 -10530 9090 -10440
rect 9660 -10530 10060 -10440
rect 10290 -10530 10690 -10440
rect 11020 -10410 11160 -10400
rect 11020 -10530 11030 -10410
rect 11150 -10530 13890 -10410
rect 15600 -10440 15610 -10320
rect 15730 -10330 15740 -10320
rect 16060 -10330 16450 -10230
rect 16700 -10330 17090 -10230
rect 15730 -10430 17090 -10330
rect 15730 -10440 15740 -10430
rect 15600 -10450 15740 -10440
rect 16060 -10530 16450 -10430
rect 16700 -10530 17090 -10430
rect 17200 -10320 17340 -10310
rect 17200 -10440 17210 -10320
rect 17330 -10330 17340 -10320
rect 17660 -10330 18050 -10230
rect 18300 -10330 18690 -10230
rect 17330 -10430 18690 -10330
rect 17330 -10440 17340 -10430
rect 17200 -10450 17340 -10440
rect 17660 -10530 18050 -10430
rect 18300 -10530 18690 -10430
rect 18800 -10320 18940 -10310
rect 18800 -10440 18810 -10320
rect 18930 -10330 18940 -10320
rect 19260 -10330 19650 -10230
rect 19900 -10330 20290 -10230
rect 18930 -10430 20290 -10330
rect 18930 -10440 18940 -10430
rect 18800 -10450 18940 -10440
rect 19260 -10530 19650 -10430
rect 19900 -10530 20290 -10430
rect 20400 -10320 20540 -10310
rect 20400 -10440 20410 -10320
rect 20530 -10330 20540 -10320
rect 20860 -10330 21250 -10230
rect 21500 -10330 21890 -10230
rect 20530 -10430 21890 -10330
rect 20530 -10440 20540 -10430
rect 20400 -10450 20540 -10440
rect 20860 -10530 21250 -10430
rect 21500 -10530 21890 -10430
rect 22000 -10320 22140 -10310
rect 22000 -10440 22010 -10320
rect 22130 -10330 22140 -10320
rect 22460 -10330 22850 -10230
rect 23100 -10330 23490 -10230
rect 22130 -10430 23490 -10330
rect 22130 -10440 22140 -10430
rect 22000 -10450 22140 -10440
rect 22460 -10530 22850 -10430
rect 23100 -10530 23490 -10430
rect 23600 -10320 23740 -10310
rect 23600 -10440 23610 -10320
rect 23730 -10330 23740 -10320
rect 24060 -10330 24450 -10230
rect 24700 -10330 25090 -10230
rect 23730 -10430 25090 -10330
rect 23730 -10440 23740 -10430
rect 23600 -10450 23740 -10440
rect 24060 -10530 24450 -10430
rect 24700 -10530 25090 -10430
rect 25200 -10320 25340 -10310
rect 25200 -10440 25210 -10320
rect 25330 -10330 25340 -10320
rect 25660 -10330 26050 -10230
rect 26300 -10330 26690 -10230
rect 27260 -10268 27657 -10230
rect 27893 -10268 28290 -10230
rect 25330 -10430 26690 -10330
rect 25330 -10440 25340 -10430
rect 25200 -10450 25340 -10440
rect 25660 -10530 26050 -10430
rect 26300 -10530 26690 -10430
rect 26800 -10320 26940 -10310
rect 26800 -10440 26810 -10320
rect 26930 -10330 26940 -10320
rect 27260 -10330 27650 -10268
rect 27900 -10330 28290 -10268
rect 28860 -10268 29257 -10230
rect 29493 -10268 29890 -10230
rect 30457 -10268 30857 -10230
rect 31093 -10228 31493 -10222
rect 31093 -10230 31105 -10228
rect 31481 -10230 31493 -10228
rect 31093 -10268 31493 -10230
rect 26930 -10430 28290 -10330
rect 26930 -10440 26940 -10430
rect 26800 -10450 26940 -10440
rect 27260 -10490 27650 -10430
rect 27900 -10490 28290 -10430
rect 28400 -10320 28540 -10310
rect 28400 -10440 28410 -10320
rect 28530 -10330 28540 -10320
rect 28860 -10330 29250 -10268
rect 29500 -10330 29890 -10268
rect 28530 -10430 29890 -10330
rect 28530 -10440 28540 -10430
rect 28400 -10450 28540 -10440
rect 27260 -10530 27657 -10490
rect 27893 -10530 28290 -10490
rect 28860 -10490 29250 -10430
rect 29500 -10490 29890 -10430
rect 30000 -10320 30140 -10310
rect 30000 -10440 30010 -10320
rect 30130 -10330 30140 -10320
rect 30460 -10330 30850 -10268
rect 31100 -10330 31490 -10268
rect 30130 -10430 31490 -10330
rect 30130 -10440 30140 -10430
rect 30000 -10450 30140 -10440
rect 28860 -10530 29257 -10490
rect 29493 -10530 29890 -10490
rect 30460 -10490 30850 -10430
rect 31100 -10490 31490 -10430
rect 30460 -10530 30857 -10490
rect 31093 -10530 31490 -10490
rect 11020 -10540 11160 -10530
rect 2120 -10610 2240 -10600
rect 2120 -11270 2130 -10610
rect 2230 -11270 2240 -10610
rect 2120 -11280 2240 -11270
rect 3720 -10610 3840 -10600
rect 3720 -11270 3730 -10610
rect 3830 -11270 3840 -10610
rect 3720 -11280 3840 -11270
rect 5320 -10610 5440 -10600
rect 5320 -11270 5330 -10610
rect 5430 -11270 5440 -10610
rect 5320 -11280 5440 -11270
rect 6920 -10610 7040 -10600
rect 6920 -11270 6930 -10610
rect 7030 -11270 7040 -10610
rect 6920 -11280 7040 -11270
rect 8520 -10610 8640 -10600
rect 8520 -11270 8530 -10610
rect 8630 -11270 8640 -10610
rect 8520 -11280 8640 -11270
rect 10120 -10610 10240 -10600
rect 10120 -11270 10130 -10610
rect 10230 -11270 10240 -10610
rect 10120 -11280 10240 -11270
rect 11710 -10610 11840 -10530
rect 11710 -11270 11720 -10610
rect 11830 -11270 11840 -10610
rect 11710 -11280 11840 -11270
rect 13310 -10610 13440 -10530
rect 16510 -10600 16640 -10590
rect 13310 -11270 13320 -10610
rect 13430 -11270 13440 -10610
rect 13310 -11280 13440 -11270
rect 14910 -10610 15040 -10600
rect 14910 -11270 14920 -10610
rect 15030 -11270 15040 -10610
rect 14910 -11280 15040 -11270
rect 16510 -11280 16520 -10600
rect 16630 -11280 16640 -10600
rect 16510 -11290 16640 -11280
rect 18110 -10600 18240 -10590
rect 18110 -11280 18120 -10600
rect 18230 -11280 18240 -10600
rect 18110 -11290 18240 -11280
rect 19710 -10600 19840 -10590
rect 19710 -11280 19720 -10600
rect 19830 -11280 19840 -10600
rect 19710 -11290 19840 -11280
rect 21310 -10600 21440 -10590
rect 21310 -11280 21320 -10600
rect 21430 -11280 21440 -10600
rect 21310 -11290 21440 -11280
rect 22910 -10600 23040 -10590
rect 22910 -11280 22920 -10600
rect 23030 -11280 23040 -10600
rect 22910 -11290 23040 -11280
rect 24510 -10600 24640 -10590
rect 24510 -11280 24520 -10600
rect 24630 -11280 24640 -10600
rect 24510 -11290 24640 -11280
rect 26110 -10600 26240 -10590
rect 26110 -11280 26120 -10600
rect 26230 -11280 26240 -10600
rect 26110 -11290 26240 -11280
rect 27710 -10600 27840 -10590
rect 27710 -11280 27720 -10600
rect 27830 -11280 27840 -10600
rect 27710 -11290 27840 -11280
rect 29310 -10600 29440 -10590
rect 29310 -11280 29320 -10600
rect 29430 -11280 29440 -10600
rect 29310 -11290 29440 -11280
rect 30910 -10600 31040 -10590
rect 30910 -11280 30920 -10600
rect 31030 -11280 31040 -10600
rect 30910 -11290 31040 -11280
rect -960 -11560 36260 -11360
rect 1200 -11670 1340 -11660
rect 1200 -11790 1210 -11670
rect 1330 -11680 1340 -11670
rect 2800 -11670 2940 -11660
rect 2800 -11680 2810 -11670
rect 1330 -11780 2810 -11680
rect 1330 -11790 1340 -11780
rect 1200 -11800 1340 -11790
rect 2800 -11790 2810 -11780
rect 2930 -11680 2940 -11670
rect 4400 -11670 4540 -11660
rect 4400 -11680 4410 -11670
rect 2930 -11780 4410 -11680
rect 2930 -11790 2940 -11780
rect 2800 -11800 2940 -11790
rect 4400 -11790 4410 -11780
rect 4530 -11680 4540 -11670
rect 6000 -11670 6140 -11660
rect 6000 -11680 6010 -11670
rect 4530 -11780 6010 -11680
rect 4530 -11790 4540 -11780
rect 4400 -11800 4540 -11790
rect 6000 -11790 6010 -11780
rect 6130 -11680 6140 -11670
rect 7600 -11670 7740 -11660
rect 7600 -11680 7610 -11670
rect 6130 -11780 7610 -11680
rect 6130 -11790 6140 -11780
rect 6000 -11800 6140 -11790
rect 7600 -11790 7610 -11780
rect 7730 -11680 7740 -11670
rect 9200 -11670 9340 -11660
rect 13300 -11670 13440 -11660
rect 14220 -11670 14360 -11660
rect 14900 -11670 15040 -11660
rect 15820 -11670 15960 -11660
rect 9200 -11680 9210 -11670
rect 7730 -11780 9210 -11680
rect 7730 -11790 7740 -11780
rect 7600 -11800 7740 -11790
rect 9200 -11790 9210 -11780
rect 9330 -11680 9340 -11670
rect 9330 -11780 10700 -11680
rect 9330 -11790 9340 -11780
rect 9200 -11800 9340 -11790
rect 12860 -11790 13310 -11670
rect 13430 -11790 14230 -11670
rect 14350 -11790 14910 -11670
rect 15030 -11790 15490 -11670
rect 12860 -11800 15490 -11790
rect 15820 -11790 15830 -11670
rect 15950 -11700 15960 -11670
rect 17420 -11670 17560 -11660
rect 15950 -11790 17090 -11700
rect 15820 -11800 17090 -11790
rect 17420 -11790 17430 -11670
rect 17550 -11700 17560 -11670
rect 19020 -11670 19160 -11660
rect 17550 -11790 18690 -11700
rect 17420 -11800 18690 -11790
rect 19020 -11790 19030 -11670
rect 19150 -11700 19160 -11670
rect 20620 -11670 20760 -11660
rect 19150 -11790 20290 -11700
rect 19020 -11800 20290 -11790
rect 20620 -11790 20630 -11670
rect 20750 -11700 20760 -11670
rect 22220 -11670 22360 -11660
rect 20750 -11790 21890 -11700
rect 20620 -11800 21890 -11790
rect 22220 -11790 22230 -11670
rect 22350 -11700 22360 -11670
rect 23820 -11670 23960 -11660
rect 22350 -11790 23490 -11700
rect 22220 -11800 23490 -11790
rect 23820 -11790 23830 -11670
rect 23950 -11700 23960 -11670
rect 25420 -11670 25560 -11660
rect 23950 -11790 25090 -11700
rect 23820 -11800 25090 -11790
rect 25420 -11790 25430 -11670
rect 25550 -11700 25560 -11670
rect 27020 -11670 27160 -11660
rect 25550 -11790 26680 -11700
rect 25420 -11800 26680 -11790
rect 27020 -11790 27030 -11670
rect 27150 -11700 27160 -11670
rect 28620 -11670 28760 -11660
rect 27150 -11790 28290 -11700
rect 27020 -11800 28290 -11790
rect 28620 -11790 28630 -11670
rect 28750 -11700 28760 -11670
rect 30220 -11670 30360 -11660
rect 28750 -11790 29890 -11700
rect 28620 -11800 29890 -11790
rect 30220 -11790 30230 -11670
rect 30350 -11700 30360 -11670
rect 30350 -11764 31490 -11700
rect 30350 -11790 31493 -11764
rect 30220 -11800 31493 -11790
rect 30457 -11804 30469 -11800
rect 30845 -11804 30857 -11800
rect 30457 -11810 30857 -11804
rect 31093 -11804 31105 -11800
rect 31481 -11804 31493 -11800
rect 31093 -11810 31493 -11804
rect 30370 -11849 30416 -11837
rect 30370 -11860 30376 -11849
rect 30410 -11860 30416 -11849
rect 30898 -11849 30944 -11837
rect 30898 -11860 30904 -11849
rect 30938 -11860 30944 -11849
rect 31006 -11849 31052 -11837
rect 31006 -11860 31012 -11849
rect 31046 -11860 31052 -11849
rect 31534 -11849 31560 -11837
rect 31534 -11860 31540 -11849
rect 1560 -11980 33200 -11860
rect 30370 -11983 30376 -11980
rect 30410 -11983 30416 -11980
rect 30370 -11995 30416 -11983
rect 30898 -11983 30904 -11980
rect 30938 -11983 30944 -11980
rect 30898 -11995 30944 -11983
rect 31006 -11983 31012 -11980
rect 31046 -11983 31052 -11980
rect 31006 -11995 31052 -11983
rect 31534 -11983 31540 -11980
rect 31534 -11995 31560 -11983
rect 30457 -12028 30857 -12022
rect 30457 -12030 30469 -12028
rect 30845 -12030 30857 -12028
rect 1420 -12110 1560 -12100
rect 1420 -12230 1430 -12110
rect 1550 -12120 1560 -12110
rect 1660 -12120 2060 -12030
rect 2290 -12120 2690 -12030
rect 3020 -12110 3160 -12100
rect 3020 -12120 3030 -12110
rect 1550 -12220 3030 -12120
rect 1550 -12230 1560 -12220
rect 1420 -12240 1560 -12230
rect 1660 -12240 2690 -12220
rect 3020 -12230 3030 -12220
rect 3150 -12120 3160 -12110
rect 3260 -12120 3660 -12030
rect 3890 -12120 4290 -12030
rect 4620 -12110 4760 -12100
rect 4620 -12120 4630 -12110
rect 3150 -12220 4630 -12120
rect 3150 -12230 3160 -12220
rect 3020 -12240 3160 -12230
rect 3260 -12240 4290 -12220
rect 4620 -12230 4630 -12220
rect 4750 -12120 4760 -12110
rect 4860 -12120 5260 -12030
rect 5490 -12120 5890 -12030
rect 6220 -12110 6360 -12100
rect 6220 -12120 6230 -12110
rect 4750 -12220 6230 -12120
rect 4750 -12230 4760 -12220
rect 4620 -12240 4760 -12230
rect 4860 -12240 5890 -12220
rect 6220 -12230 6230 -12220
rect 6350 -12120 6360 -12110
rect 6460 -12120 6860 -12030
rect 7090 -12120 7490 -12030
rect 7820 -12110 7960 -12100
rect 7820 -12120 7830 -12110
rect 6350 -12220 7830 -12120
rect 6350 -12230 6360 -12220
rect 6220 -12240 6360 -12230
rect 6460 -12240 7490 -12220
rect 7820 -12230 7830 -12220
rect 7950 -12120 7960 -12110
rect 8060 -12120 8460 -12030
rect 8690 -12120 9090 -12030
rect 9420 -12110 9560 -12100
rect 9420 -12120 9430 -12110
rect 7950 -12220 9430 -12120
rect 7950 -12230 7960 -12220
rect 7820 -12240 7960 -12230
rect 8060 -12240 9090 -12220
rect 9420 -12230 9430 -12220
rect 9550 -12120 9560 -12110
rect 9660 -12120 10060 -12030
rect 10290 -12120 10690 -12030
rect 12857 -12068 13260 -12030
rect 12860 -12120 13260 -12068
rect 13490 -12068 13893 -12030
rect 14457 -12068 14860 -12030
rect 13490 -12120 13890 -12068
rect 14460 -12120 14860 -12068
rect 15090 -12068 15493 -12030
rect 15090 -12120 15490 -12068
rect 9550 -12220 10690 -12120
rect 9550 -12230 9560 -12220
rect 9420 -12240 9560 -12230
rect 9660 -12240 10690 -12220
rect 1660 -12330 2060 -12240
rect 2290 -12330 2690 -12240
rect 3260 -12330 3660 -12240
rect 3890 -12330 4290 -12240
rect 4860 -12330 5260 -12240
rect 5490 -12330 5890 -12240
rect 6460 -12330 6860 -12240
rect 7090 -12330 7490 -12240
rect 8060 -12330 8460 -12240
rect 8690 -12330 9090 -12240
rect 9660 -12330 10060 -12240
rect 10290 -12330 10690 -12240
rect 10800 -12220 10940 -12210
rect 10800 -12330 10810 -12220
rect 10930 -12230 10940 -12220
rect 11260 -12230 15490 -12120
rect 10930 -12240 15490 -12230
rect 10930 -12320 12290 -12240
rect 12860 -12290 13260 -12240
rect 10930 -12330 10940 -12320
rect 11260 -12330 12290 -12320
rect 12857 -12330 13260 -12290
rect 13490 -12290 13890 -12240
rect 14460 -12290 14860 -12240
rect 13490 -12330 13893 -12290
rect 14457 -12330 14860 -12290
rect 15090 -12290 15490 -12240
rect 15600 -12120 15740 -12110
rect 15600 -12240 15610 -12120
rect 15730 -12130 15740 -12120
rect 16060 -12130 16450 -12030
rect 16700 -12130 17090 -12030
rect 15730 -12230 17090 -12130
rect 15730 -12240 15740 -12230
rect 15600 -12250 15740 -12240
rect 15090 -12330 15493 -12290
rect 16060 -12330 16450 -12230
rect 16700 -12330 17090 -12230
rect 17200 -12120 17340 -12110
rect 17200 -12240 17210 -12120
rect 17330 -12130 17340 -12120
rect 17660 -12130 18050 -12030
rect 18300 -12130 18690 -12030
rect 17330 -12230 18690 -12130
rect 17330 -12240 17340 -12230
rect 17200 -12250 17340 -12240
rect 17660 -12330 18050 -12230
rect 18300 -12330 18690 -12230
rect 18800 -12120 18940 -12110
rect 18800 -12240 18810 -12120
rect 18930 -12130 18940 -12120
rect 19260 -12130 19650 -12030
rect 19900 -12130 20290 -12030
rect 18930 -12230 20290 -12130
rect 18930 -12240 18940 -12230
rect 18800 -12250 18940 -12240
rect 19260 -12330 19650 -12230
rect 19900 -12330 20290 -12230
rect 20400 -12120 20540 -12110
rect 20400 -12240 20410 -12120
rect 20530 -12130 20540 -12120
rect 20860 -12130 21250 -12030
rect 21500 -12130 21890 -12030
rect 20530 -12230 21890 -12130
rect 20530 -12240 20540 -12230
rect 20400 -12250 20540 -12240
rect 20860 -12330 21250 -12230
rect 21500 -12330 21890 -12230
rect 22000 -12120 22140 -12110
rect 22000 -12240 22010 -12120
rect 22130 -12130 22140 -12120
rect 22460 -12130 22850 -12030
rect 23100 -12130 23490 -12030
rect 22130 -12230 23490 -12130
rect 22130 -12240 22140 -12230
rect 22000 -12250 22140 -12240
rect 22460 -12330 22850 -12230
rect 23100 -12330 23490 -12230
rect 23600 -12120 23740 -12110
rect 23600 -12240 23610 -12120
rect 23730 -12130 23740 -12120
rect 24060 -12130 24450 -12030
rect 24700 -12130 25090 -12030
rect 23730 -12230 25090 -12130
rect 23730 -12240 23740 -12230
rect 23600 -12250 23740 -12240
rect 24060 -12330 24450 -12230
rect 24700 -12330 25090 -12230
rect 25200 -12120 25340 -12110
rect 25200 -12240 25210 -12120
rect 25330 -12130 25340 -12120
rect 25660 -12130 26050 -12030
rect 26300 -12130 26690 -12030
rect 27260 -12068 27657 -12030
rect 27893 -12068 28290 -12030
rect 25330 -12230 26690 -12130
rect 25330 -12240 25340 -12230
rect 25200 -12250 25340 -12240
rect 25660 -12330 26050 -12230
rect 26300 -12330 26690 -12230
rect 26800 -12120 26940 -12110
rect 26800 -12240 26810 -12120
rect 26930 -12130 26940 -12120
rect 27260 -12130 27650 -12068
rect 27900 -12130 28290 -12068
rect 28860 -12068 29257 -12030
rect 29493 -12068 29890 -12030
rect 30457 -12068 30857 -12030
rect 31093 -12028 31493 -12022
rect 31093 -12030 31105 -12028
rect 31481 -12030 31493 -12028
rect 31093 -12068 31493 -12030
rect 26930 -12230 28290 -12130
rect 26930 -12240 26940 -12230
rect 26800 -12250 26940 -12240
rect 27260 -12290 27650 -12230
rect 27900 -12290 28290 -12230
rect 28400 -12120 28540 -12110
rect 28400 -12240 28410 -12120
rect 28530 -12130 28540 -12120
rect 28860 -12130 29250 -12068
rect 29500 -12130 29890 -12068
rect 28530 -12230 29890 -12130
rect 28530 -12240 28540 -12230
rect 28400 -12250 28540 -12240
rect 27260 -12330 27657 -12290
rect 27893 -12330 28290 -12290
rect 28860 -12290 29250 -12230
rect 29500 -12290 29890 -12230
rect 30000 -12120 30140 -12110
rect 30000 -12240 30010 -12120
rect 30130 -12130 30140 -12120
rect 30460 -12130 30850 -12068
rect 31100 -12130 31490 -12068
rect 30130 -12230 31490 -12130
rect 30130 -12240 30140 -12230
rect 30000 -12250 30140 -12240
rect 28860 -12330 29257 -12290
rect 29493 -12330 29890 -12290
rect 30460 -12290 30850 -12230
rect 31100 -12290 31490 -12230
rect 30460 -12330 30857 -12290
rect 31093 -12330 31490 -12290
rect 10800 -12340 10940 -12330
rect 16510 -12400 16640 -12390
rect 2120 -12410 2240 -12400
rect 2120 -13070 2130 -12410
rect 2230 -13070 2240 -12410
rect 2120 -13080 2240 -13070
rect 3720 -12410 3840 -12400
rect 3720 -13070 3730 -12410
rect 3830 -13070 3840 -12410
rect 3720 -13080 3840 -13070
rect 5320 -12410 5440 -12400
rect 5320 -13070 5330 -12410
rect 5430 -13070 5440 -12410
rect 5320 -13080 5440 -13070
rect 6920 -12410 7040 -12400
rect 6920 -13070 6930 -12410
rect 7030 -13070 7040 -12410
rect 6920 -13080 7040 -13070
rect 8520 -12410 8640 -12400
rect 8520 -13070 8530 -12410
rect 8630 -13070 8640 -12410
rect 8520 -13080 8640 -13070
rect 10120 -12410 10240 -12400
rect 10120 -13070 10130 -12410
rect 10230 -13070 10240 -12410
rect 10120 -13080 10240 -13070
rect 11710 -12410 11840 -12400
rect 11710 -13070 11720 -12410
rect 11830 -13070 11840 -12410
rect 11710 -13080 11840 -13070
rect 13310 -12410 13440 -12400
rect 13310 -13070 13320 -12410
rect 13430 -13070 13440 -12410
rect 13310 -13080 13440 -13070
rect 14910 -12410 15040 -12400
rect 14910 -13070 14920 -12410
rect 15030 -13070 15040 -12410
rect 14910 -13080 15040 -13070
rect 16510 -13080 16520 -12400
rect 16630 -13080 16640 -12400
rect 16510 -13090 16640 -13080
rect 18110 -12400 18240 -12390
rect 18110 -13080 18120 -12400
rect 18230 -13080 18240 -12400
rect 18110 -13090 18240 -13080
rect 19710 -12400 19840 -12390
rect 19710 -13080 19720 -12400
rect 19830 -13080 19840 -12400
rect 19710 -13090 19840 -13080
rect 21310 -12400 21440 -12390
rect 21310 -13080 21320 -12400
rect 21430 -13080 21440 -12400
rect 21310 -13090 21440 -13080
rect 22910 -12400 23040 -12390
rect 22910 -13080 22920 -12400
rect 23030 -13080 23040 -12400
rect 22910 -13090 23040 -13080
rect 24510 -12400 24640 -12390
rect 24510 -13080 24520 -12400
rect 24630 -13080 24640 -12400
rect 24510 -13090 24640 -13080
rect 26110 -12400 26240 -12390
rect 26110 -13080 26120 -12400
rect 26230 -13080 26240 -12400
rect 26110 -13090 26240 -13080
rect 27710 -12400 27840 -12390
rect 27710 -13080 27720 -12400
rect 27830 -13080 27840 -12400
rect 27710 -13090 27840 -13080
rect 29310 -12400 29440 -12390
rect 29310 -13080 29320 -12400
rect 29430 -13080 29440 -12400
rect 29310 -13090 29440 -13080
rect 30910 -12400 31040 -12390
rect 30910 -13080 30920 -12400
rect 31030 -13080 31040 -12400
rect 30910 -13090 31040 -13080
rect -960 -13260 11190 -13160
rect 11260 -13210 11270 -13150
rect 11650 -13210 12300 -13150
rect 12400 -13260 36260 -13160
rect -960 -13360 36260 -13260
rect 11030 -13440 12530 -13360
rect 1200 -13470 1340 -13460
rect 1200 -13590 1210 -13470
rect 1330 -13480 1340 -13470
rect 2800 -13470 2940 -13460
rect 2800 -13480 2810 -13470
rect 1330 -13580 2810 -13480
rect 1330 -13590 1340 -13580
rect 1200 -13600 1340 -13590
rect 2800 -13590 2810 -13580
rect 2930 -13480 2940 -13470
rect 4400 -13470 4540 -13460
rect 4400 -13480 4410 -13470
rect 2930 -13580 4410 -13480
rect 2930 -13590 2940 -13580
rect 2800 -13600 2940 -13590
rect 4400 -13590 4410 -13580
rect 4530 -13480 4540 -13470
rect 6000 -13470 6140 -13460
rect 6000 -13480 6010 -13470
rect 4530 -13580 6010 -13480
rect 4530 -13590 4540 -13580
rect 4400 -13600 4540 -13590
rect 6000 -13590 6010 -13580
rect 6130 -13480 6140 -13470
rect 7600 -13470 7740 -13460
rect 7600 -13480 7610 -13470
rect 6130 -13580 7610 -13480
rect 6130 -13590 6140 -13580
rect 6000 -13600 6140 -13590
rect 7600 -13590 7610 -13580
rect 7730 -13480 7740 -13470
rect 9200 -13470 9340 -13460
rect 15820 -13470 15960 -13460
rect 9200 -13480 9210 -13470
rect 7730 -13580 9210 -13480
rect 7730 -13590 7740 -13580
rect 7600 -13600 7740 -13590
rect 9200 -13590 9210 -13580
rect 9330 -13480 9340 -13470
rect 14000 -13480 14140 -13470
rect 9330 -13580 10700 -13480
rect 14000 -13520 14010 -13480
rect 9330 -13590 9340 -13580
rect 9200 -13600 9340 -13590
rect 12860 -13600 14010 -13520
rect 14130 -13520 14140 -13480
rect 14130 -13600 15490 -13520
rect 15820 -13590 15830 -13470
rect 15950 -13500 15960 -13470
rect 17420 -13470 17560 -13460
rect 15950 -13590 17090 -13500
rect 15820 -13600 17090 -13590
rect 17420 -13590 17430 -13470
rect 17550 -13500 17560 -13470
rect 19020 -13470 19160 -13460
rect 17550 -13590 18690 -13500
rect 17420 -13600 18690 -13590
rect 19020 -13590 19030 -13470
rect 19150 -13500 19160 -13470
rect 20620 -13470 20760 -13460
rect 19150 -13590 20290 -13500
rect 19020 -13600 20290 -13590
rect 20620 -13590 20630 -13470
rect 20750 -13500 20760 -13470
rect 22220 -13470 22360 -13460
rect 20750 -13590 21890 -13500
rect 20620 -13600 21890 -13590
rect 22220 -13590 22230 -13470
rect 22350 -13500 22360 -13470
rect 23820 -13470 23960 -13460
rect 22350 -13590 23490 -13500
rect 22220 -13600 23490 -13590
rect 23820 -13590 23830 -13470
rect 23950 -13500 23960 -13470
rect 25420 -13470 25560 -13460
rect 23950 -13590 25090 -13500
rect 23820 -13600 25090 -13590
rect 25420 -13590 25430 -13470
rect 25550 -13500 25560 -13470
rect 27020 -13470 27160 -13460
rect 25550 -13590 26680 -13500
rect 25420 -13600 26680 -13590
rect 27020 -13590 27030 -13470
rect 27150 -13500 27160 -13470
rect 28620 -13470 28760 -13460
rect 27150 -13590 28290 -13500
rect 27020 -13600 28290 -13590
rect 28620 -13590 28630 -13470
rect 28750 -13500 28760 -13470
rect 30220 -13470 30360 -13460
rect 28750 -13590 29890 -13500
rect 28620 -13600 29890 -13590
rect 30220 -13590 30230 -13470
rect 30350 -13500 30360 -13470
rect 30350 -13564 31490 -13500
rect 30350 -13590 31493 -13564
rect 30220 -13600 31493 -13590
rect 14000 -13610 14140 -13600
rect 30457 -13604 30469 -13600
rect 30845 -13604 30857 -13600
rect 30457 -13610 30857 -13604
rect 31093 -13604 31105 -13600
rect 31481 -13604 31493 -13600
rect 31093 -13610 31493 -13604
rect 30370 -13649 30416 -13637
rect 30370 -13660 30376 -13649
rect 30410 -13660 30416 -13649
rect 30898 -13649 30944 -13637
rect 30898 -13660 30904 -13649
rect 30938 -13660 30944 -13649
rect 31006 -13649 31052 -13637
rect 31006 -13660 31012 -13649
rect 31046 -13660 31052 -13649
rect 31534 -13649 31560 -13637
rect 31534 -13660 31540 -13649
rect 1560 -13780 33200 -13660
rect 30370 -13783 30376 -13780
rect 30410 -13783 30416 -13780
rect 30370 -13795 30416 -13783
rect 30898 -13783 30904 -13780
rect 30938 -13783 30944 -13780
rect 30898 -13795 30944 -13783
rect 31006 -13783 31012 -13780
rect 31046 -13783 31052 -13780
rect 31006 -13795 31052 -13783
rect 31534 -13783 31540 -13780
rect 31534 -13795 31560 -13783
rect 30457 -13828 30857 -13822
rect 30457 -13830 30469 -13828
rect 30845 -13830 30857 -13828
rect 1420 -13910 1560 -13900
rect 1420 -14030 1430 -13910
rect 1550 -13920 1560 -13910
rect 1660 -13920 2060 -13830
rect 2290 -13920 2690 -13830
rect 3020 -13910 3160 -13900
rect 3020 -13920 3030 -13910
rect 1550 -14020 3030 -13920
rect 1550 -14030 1560 -14020
rect 1420 -14040 1560 -14030
rect 1660 -14040 2690 -14020
rect 3020 -14030 3030 -14020
rect 3150 -13920 3160 -13910
rect 3260 -13920 3660 -13830
rect 3890 -13920 4290 -13830
rect 4620 -13910 4760 -13900
rect 4620 -13920 4630 -13910
rect 3150 -14020 4630 -13920
rect 3150 -14030 3160 -14020
rect 3020 -14040 3160 -14030
rect 3260 -14040 4290 -14020
rect 4620 -14030 4630 -14020
rect 4750 -13920 4760 -13910
rect 4860 -13920 5260 -13830
rect 5490 -13920 5890 -13830
rect 6220 -13910 6360 -13900
rect 6220 -13920 6230 -13910
rect 4750 -14020 6230 -13920
rect 4750 -14030 4760 -14020
rect 4620 -14040 4760 -14030
rect 4860 -14040 5890 -14020
rect 6220 -14030 6230 -14020
rect 6350 -13920 6360 -13910
rect 6460 -13920 6860 -13830
rect 7090 -13920 7490 -13830
rect 7820 -13910 7960 -13900
rect 7820 -13920 7830 -13910
rect 6350 -14020 7830 -13920
rect 6350 -14030 6360 -14020
rect 6220 -14040 6360 -14030
rect 6460 -14040 7490 -14020
rect 7820 -14030 7830 -14020
rect 7950 -13920 7960 -13910
rect 8060 -13920 8460 -13830
rect 8690 -13920 9090 -13830
rect 9420 -13910 9560 -13900
rect 9420 -13920 9430 -13910
rect 7950 -14020 9430 -13920
rect 7950 -14030 7960 -14020
rect 7820 -14040 7960 -14030
rect 8060 -14040 9090 -14020
rect 9420 -14030 9430 -14020
rect 9550 -13920 9560 -13910
rect 9660 -13920 10060 -13830
rect 10290 -13920 10690 -13830
rect 9550 -14020 10690 -13920
rect 9550 -14030 9560 -14020
rect 9420 -14040 9560 -14030
rect 9660 -14040 10690 -14020
rect 1660 -14130 2060 -14040
rect 2290 -14130 2690 -14040
rect 3260 -14130 3660 -14040
rect 3890 -14130 4290 -14040
rect 4860 -14130 5260 -14040
rect 5490 -14130 5890 -14040
rect 6460 -14130 6860 -14040
rect 7090 -14130 7490 -14040
rect 8060 -14130 8460 -14040
rect 8690 -14130 9090 -14040
rect 9660 -14130 10060 -14040
rect 10290 -14130 10690 -14040
rect 12860 -13920 13260 -13830
rect 13490 -13920 13890 -13830
rect 14460 -13920 14860 -13830
rect 15090 -13920 15490 -13830
rect 12860 -14040 15490 -13920
rect 11260 -14060 12290 -14050
rect 11260 -14120 11270 -14060
rect 11650 -14120 12290 -14060
rect 11260 -14130 11660 -14120
rect 12860 -14130 13260 -14040
rect 13490 -14130 13890 -14040
rect 14460 -14130 14860 -14040
rect 15090 -14130 15490 -14040
rect 15600 -13920 15740 -13910
rect 15600 -14040 15610 -13920
rect 15730 -13930 15740 -13920
rect 16060 -13930 16450 -13830
rect 16700 -13930 17090 -13830
rect 15730 -14030 17090 -13930
rect 15730 -14040 15740 -14030
rect 15600 -14050 15740 -14040
rect 16060 -14130 16450 -14030
rect 16700 -14130 17090 -14030
rect 17200 -13920 17340 -13910
rect 17200 -14040 17210 -13920
rect 17330 -13930 17340 -13920
rect 17660 -13930 18050 -13830
rect 18300 -13930 18690 -13830
rect 17330 -14030 18690 -13930
rect 17330 -14040 17340 -14030
rect 17200 -14050 17340 -14040
rect 17660 -14130 18050 -14030
rect 18300 -14130 18690 -14030
rect 18800 -13920 18940 -13910
rect 18800 -14040 18810 -13920
rect 18930 -13930 18940 -13920
rect 19260 -13930 19650 -13830
rect 19900 -13930 20290 -13830
rect 18930 -14030 20290 -13930
rect 18930 -14040 18940 -14030
rect 18800 -14050 18940 -14040
rect 19260 -14130 19650 -14030
rect 19900 -14130 20290 -14030
rect 20400 -13920 20540 -13910
rect 20400 -14040 20410 -13920
rect 20530 -13930 20540 -13920
rect 20860 -13930 21250 -13830
rect 21500 -13930 21890 -13830
rect 20530 -14030 21890 -13930
rect 20530 -14040 20540 -14030
rect 20400 -14050 20540 -14040
rect 20860 -14130 21250 -14030
rect 21500 -14130 21890 -14030
rect 22000 -13920 22140 -13910
rect 22000 -14040 22010 -13920
rect 22130 -13930 22140 -13920
rect 22460 -13930 22850 -13830
rect 23100 -13930 23490 -13830
rect 22130 -14030 23490 -13930
rect 22130 -14040 22140 -14030
rect 22000 -14050 22140 -14040
rect 22460 -14130 22850 -14030
rect 23100 -14130 23490 -14030
rect 23600 -13920 23740 -13910
rect 23600 -14040 23610 -13920
rect 23730 -13930 23740 -13920
rect 24060 -13930 24450 -13830
rect 24700 -13930 25090 -13830
rect 23730 -14030 25090 -13930
rect 23730 -14040 23740 -14030
rect 23600 -14050 23740 -14040
rect 24060 -14130 24450 -14030
rect 24700 -14130 25090 -14030
rect 25200 -13920 25340 -13910
rect 25200 -14040 25210 -13920
rect 25330 -13930 25340 -13920
rect 25660 -13930 26050 -13830
rect 26300 -13930 26690 -13830
rect 27260 -13868 27657 -13830
rect 27893 -13868 28290 -13830
rect 25330 -14030 26690 -13930
rect 25330 -14040 25340 -14030
rect 25200 -14050 25340 -14040
rect 25660 -14130 26050 -14030
rect 26300 -14130 26690 -14030
rect 26800 -13920 26940 -13910
rect 26800 -14040 26810 -13920
rect 26930 -13930 26940 -13920
rect 27260 -13930 27650 -13868
rect 27900 -13930 28290 -13868
rect 28860 -13868 29257 -13830
rect 29493 -13868 29890 -13830
rect 30457 -13868 30857 -13830
rect 31093 -13828 31493 -13822
rect 31093 -13830 31105 -13828
rect 31481 -13830 31493 -13828
rect 31093 -13868 31493 -13830
rect 26930 -14030 28290 -13930
rect 26930 -14040 26940 -14030
rect 26800 -14050 26940 -14040
rect 27260 -14090 27650 -14030
rect 27900 -14090 28290 -14030
rect 28400 -13920 28540 -13910
rect 28400 -14040 28410 -13920
rect 28530 -13930 28540 -13920
rect 28860 -13930 29250 -13868
rect 29500 -13930 29890 -13868
rect 28530 -14030 29890 -13930
rect 28530 -14040 28540 -14030
rect 28400 -14050 28540 -14040
rect 27260 -14130 27657 -14090
rect 27893 -14130 28290 -14090
rect 28860 -14090 29250 -14030
rect 29500 -14090 29890 -14030
rect 30000 -13920 30140 -13910
rect 30000 -14040 30010 -13920
rect 30130 -13930 30140 -13920
rect 30460 -13930 30850 -13868
rect 31100 -13930 31490 -13868
rect 30130 -14030 31490 -13930
rect 30130 -14040 30140 -14030
rect 30000 -14050 30140 -14040
rect 28860 -14130 29257 -14090
rect 29493 -14130 29890 -14090
rect 30460 -14090 30850 -14030
rect 31100 -14090 31490 -14030
rect 30460 -14130 30857 -14090
rect 31093 -14130 31490 -14090
rect 16510 -14200 16640 -14190
rect 2120 -14210 2240 -14200
rect 2120 -14870 2130 -14210
rect 2230 -14870 2240 -14210
rect 2120 -14880 2240 -14870
rect 3720 -14210 3840 -14200
rect 3720 -14870 3730 -14210
rect 3830 -14870 3840 -14210
rect 3720 -14880 3840 -14870
rect 5320 -14210 5440 -14200
rect 5320 -14870 5330 -14210
rect 5430 -14870 5440 -14210
rect 5320 -14880 5440 -14870
rect 6920 -14210 7040 -14200
rect 6920 -14870 6930 -14210
rect 7030 -14870 7040 -14210
rect 6920 -14880 7040 -14870
rect 8520 -14210 8640 -14200
rect 8520 -14870 8530 -14210
rect 8630 -14870 8640 -14210
rect 8520 -14880 8640 -14870
rect 10120 -14210 10240 -14200
rect 10120 -14870 10130 -14210
rect 10230 -14870 10240 -14210
rect 10120 -14880 10240 -14870
rect 11710 -14210 11840 -14200
rect 11710 -14870 11720 -14210
rect 11830 -14870 11840 -14210
rect 11710 -14880 11840 -14870
rect 13310 -14210 13440 -14200
rect 13310 -14870 13320 -14210
rect 13430 -14870 13440 -14210
rect 13310 -14880 13440 -14870
rect 14910 -14210 15040 -14200
rect 14910 -14870 14920 -14210
rect 15030 -14870 15040 -14210
rect 14910 -14880 15040 -14870
rect 16510 -14880 16520 -14200
rect 16630 -14880 16640 -14200
rect 16510 -14890 16640 -14880
rect 18110 -14200 18240 -14190
rect 18110 -14880 18120 -14200
rect 18230 -14880 18240 -14200
rect 18110 -14890 18240 -14880
rect 19710 -14200 19840 -14190
rect 19710 -14880 19720 -14200
rect 19830 -14880 19840 -14200
rect 19710 -14890 19840 -14880
rect 21310 -14200 21440 -14190
rect 21310 -14880 21320 -14200
rect 21430 -14880 21440 -14200
rect 21310 -14890 21440 -14880
rect 22910 -14200 23040 -14190
rect 22910 -14880 22920 -14200
rect 23030 -14880 23040 -14200
rect 22910 -14890 23040 -14880
rect 24510 -14200 24640 -14190
rect 24510 -14880 24520 -14200
rect 24630 -14880 24640 -14200
rect 24510 -14890 24640 -14880
rect 26110 -14200 26240 -14190
rect 26110 -14880 26120 -14200
rect 26230 -14880 26240 -14200
rect 26110 -14890 26240 -14880
rect 27710 -14200 27840 -14190
rect 27710 -14880 27720 -14200
rect 27830 -14880 27840 -14200
rect 27710 -14890 27840 -14880
rect 29310 -14200 29440 -14190
rect 29310 -14880 29320 -14200
rect 29430 -14880 29440 -14200
rect 29310 -14890 29440 -14880
rect 30910 -14200 31040 -14190
rect 30910 -14880 30920 -14200
rect 31030 -14880 31040 -14200
rect 30910 -14890 31040 -14880
rect -960 -15160 36260 -14960
rect 1200 -15270 1340 -15260
rect 1200 -15390 1210 -15270
rect 1330 -15280 1340 -15270
rect 2800 -15270 2940 -15260
rect 2800 -15280 2810 -15270
rect 1330 -15380 2810 -15280
rect 1330 -15390 1340 -15380
rect 1200 -15400 1340 -15390
rect 2800 -15390 2810 -15380
rect 2930 -15280 2940 -15270
rect 4400 -15270 4540 -15260
rect 4400 -15280 4410 -15270
rect 2930 -15380 4410 -15280
rect 2930 -15390 2940 -15380
rect 2800 -15400 2940 -15390
rect 4400 -15390 4410 -15380
rect 4530 -15280 4540 -15270
rect 6000 -15270 6140 -15260
rect 6000 -15280 6010 -15270
rect 4530 -15380 6010 -15280
rect 4530 -15390 4540 -15380
rect 4400 -15400 4540 -15390
rect 6000 -15390 6010 -15380
rect 6130 -15280 6140 -15270
rect 7600 -15270 7740 -15260
rect 7600 -15280 7610 -15270
rect 6130 -15380 7610 -15280
rect 6130 -15390 6140 -15380
rect 6000 -15400 6140 -15390
rect 7600 -15390 7610 -15380
rect 7730 -15280 7740 -15270
rect 9200 -15270 9340 -15260
rect 9200 -15280 9210 -15270
rect 7730 -15380 9210 -15280
rect 7730 -15390 7740 -15380
rect 7600 -15400 7740 -15390
rect 9200 -15390 9210 -15380
rect 9330 -15280 9340 -15270
rect 15820 -15270 15960 -15260
rect 9330 -15380 10700 -15280
rect 13320 -15290 13440 -15280
rect 13320 -15320 13330 -15290
rect 9330 -15390 9340 -15380
rect 9200 -15400 9340 -15390
rect 12860 -15390 13330 -15320
rect 13430 -15320 13440 -15290
rect 14920 -15290 15040 -15280
rect 14010 -15310 14130 -15300
rect 14010 -15320 14020 -15310
rect 13430 -15390 14020 -15320
rect 12860 -15400 14020 -15390
rect 14010 -15410 14020 -15400
rect 14120 -15320 14130 -15310
rect 14920 -15320 14930 -15290
rect 14120 -15390 14930 -15320
rect 15030 -15320 15040 -15290
rect 15030 -15390 15490 -15320
rect 14120 -15400 15490 -15390
rect 15820 -15390 15830 -15270
rect 15950 -15300 15960 -15270
rect 17420 -15270 17560 -15260
rect 15950 -15390 17090 -15300
rect 15820 -15400 17090 -15390
rect 17420 -15390 17430 -15270
rect 17550 -15300 17560 -15270
rect 19020 -15270 19160 -15260
rect 17550 -15390 18690 -15300
rect 17420 -15400 18690 -15390
rect 19020 -15390 19030 -15270
rect 19150 -15300 19160 -15270
rect 20620 -15270 20760 -15260
rect 19150 -15390 20290 -15300
rect 19020 -15400 20290 -15390
rect 20620 -15390 20630 -15270
rect 20750 -15300 20760 -15270
rect 22220 -15270 22360 -15260
rect 20750 -15390 21890 -15300
rect 20620 -15400 21890 -15390
rect 22220 -15390 22230 -15270
rect 22350 -15300 22360 -15270
rect 23820 -15270 23960 -15260
rect 22350 -15390 23490 -15300
rect 22220 -15400 23490 -15390
rect 23820 -15390 23830 -15270
rect 23950 -15300 23960 -15270
rect 27020 -15270 27160 -15260
rect 27020 -15300 27030 -15270
rect 23950 -15390 25090 -15300
rect 23820 -15400 25090 -15390
rect 25660 -15390 27030 -15300
rect 27150 -15300 27160 -15270
rect 28620 -15270 28760 -15260
rect 27150 -15390 28290 -15300
rect 25660 -15400 28290 -15390
rect 28620 -15390 28630 -15270
rect 28750 -15300 28760 -15270
rect 28750 -15390 31490 -15300
rect 28620 -15400 31490 -15390
rect 14120 -15410 14130 -15400
rect 14010 -15420 14130 -15410
rect 1560 -15580 33200 -15460
rect 1420 -15710 1560 -15700
rect 1420 -15830 1430 -15710
rect 1550 -15720 1560 -15710
rect 1660 -15720 2060 -15630
rect 2290 -15720 2690 -15630
rect 3020 -15710 3160 -15700
rect 3020 -15720 3030 -15710
rect 1550 -15820 3030 -15720
rect 1550 -15830 1560 -15820
rect 1420 -15840 1560 -15830
rect 1660 -15840 2690 -15820
rect 3020 -15830 3030 -15820
rect 3150 -15720 3160 -15710
rect 3260 -15720 3660 -15630
rect 3890 -15720 4290 -15630
rect 4620 -15710 4760 -15700
rect 4620 -15720 4630 -15710
rect 3150 -15820 4630 -15720
rect 3150 -15830 3160 -15820
rect 3020 -15840 3160 -15830
rect 3260 -15840 4290 -15820
rect 4620 -15830 4630 -15820
rect 4750 -15720 4760 -15710
rect 4860 -15720 5260 -15630
rect 5490 -15720 5890 -15630
rect 6220 -15710 6360 -15700
rect 6220 -15720 6230 -15710
rect 4750 -15820 6230 -15720
rect 4750 -15830 4760 -15820
rect 4620 -15840 4760 -15830
rect 4860 -15840 5890 -15820
rect 6220 -15830 6230 -15820
rect 6350 -15720 6360 -15710
rect 6460 -15720 6860 -15630
rect 7090 -15720 7490 -15630
rect 7820 -15710 7960 -15700
rect 7820 -15720 7830 -15710
rect 6350 -15820 7830 -15720
rect 6350 -15830 6360 -15820
rect 6220 -15840 6360 -15830
rect 6460 -15840 7490 -15820
rect 7820 -15830 7830 -15820
rect 7950 -15720 7960 -15710
rect 8060 -15720 8460 -15630
rect 8690 -15720 9090 -15630
rect 9420 -15710 9560 -15700
rect 9420 -15720 9430 -15710
rect 7950 -15820 9430 -15720
rect 7950 -15830 7960 -15820
rect 7820 -15840 7960 -15830
rect 8060 -15840 9090 -15820
rect 9420 -15830 9430 -15820
rect 9550 -15720 9560 -15710
rect 9660 -15720 10060 -15630
rect 10290 -15720 10690 -15630
rect 9550 -15820 10690 -15720
rect 9550 -15830 9560 -15820
rect 9420 -15840 9560 -15830
rect 9660 -15840 10690 -15820
rect 1660 -15930 2060 -15840
rect 2290 -15930 2690 -15840
rect 3260 -15930 3660 -15840
rect 3890 -15930 4290 -15840
rect 4860 -15930 5260 -15840
rect 5490 -15930 5890 -15840
rect 6460 -15930 6860 -15840
rect 7090 -15930 7490 -15840
rect 8060 -15930 8460 -15840
rect 8690 -15930 9090 -15840
rect 9660 -15930 10060 -15840
rect 10290 -15930 10690 -15840
rect 12860 -15710 13260 -15630
rect 13490 -15710 13890 -15630
rect 14460 -15710 14860 -15630
rect 12860 -15720 15050 -15710
rect 15090 -15720 15490 -15630
rect 12860 -15830 15490 -15720
rect 12860 -15840 13890 -15830
rect 12860 -15930 13260 -15840
rect 13490 -15930 13890 -15840
rect 14460 -15840 15490 -15830
rect 14460 -15930 14860 -15840
rect 15090 -15930 15490 -15840
rect 15600 -15720 15740 -15710
rect 15600 -15840 15610 -15720
rect 15730 -15730 15740 -15720
rect 16060 -15730 16450 -15630
rect 16700 -15730 17090 -15630
rect 15730 -15830 17090 -15730
rect 15730 -15840 15740 -15830
rect 15600 -15850 15740 -15840
rect 16060 -15930 16450 -15830
rect 16700 -15930 17090 -15830
rect 17200 -15720 17340 -15710
rect 17200 -15840 17210 -15720
rect 17330 -15730 17340 -15720
rect 17660 -15730 18050 -15630
rect 18300 -15730 18690 -15630
rect 17330 -15830 18690 -15730
rect 17330 -15840 17340 -15830
rect 17200 -15850 17340 -15840
rect 17660 -15930 18050 -15830
rect 18300 -15930 18690 -15830
rect 18800 -15720 18940 -15710
rect 18800 -15840 18810 -15720
rect 18930 -15730 18940 -15720
rect 19260 -15730 19650 -15630
rect 19900 -15730 20290 -15630
rect 18930 -15830 20290 -15730
rect 18930 -15840 18940 -15830
rect 18800 -15850 18940 -15840
rect 19260 -15930 19650 -15830
rect 19900 -15930 20290 -15830
rect 20400 -15720 20540 -15710
rect 20400 -15840 20410 -15720
rect 20530 -15730 20540 -15720
rect 20860 -15730 21250 -15630
rect 21500 -15730 21890 -15630
rect 20530 -15830 21890 -15730
rect 20530 -15840 20540 -15830
rect 20400 -15850 20540 -15840
rect 20860 -15930 21250 -15830
rect 21500 -15930 21890 -15830
rect 22000 -15720 22140 -15710
rect 22000 -15840 22010 -15720
rect 22130 -15730 22140 -15720
rect 22460 -15730 22850 -15630
rect 23100 -15730 23490 -15630
rect 22130 -15830 23490 -15730
rect 22130 -15840 22140 -15830
rect 22000 -15850 22140 -15840
rect 22460 -15930 22850 -15830
rect 23100 -15930 23490 -15830
rect 23600 -15720 23740 -15710
rect 23600 -15840 23610 -15720
rect 23730 -15730 23740 -15720
rect 24060 -15730 24450 -15630
rect 24700 -15730 25090 -15630
rect 23730 -15830 25090 -15730
rect 23730 -15840 23740 -15830
rect 23600 -15850 23740 -15840
rect 24060 -15930 24450 -15830
rect 24700 -15930 25090 -15830
rect 25660 -15730 26050 -15630
rect 26300 -15730 26690 -15630
rect 27260 -15668 27657 -15630
rect 27893 -15668 28290 -15630
rect 26800 -15720 26940 -15710
rect 26800 -15730 26810 -15720
rect 25660 -15830 26810 -15730
rect 25660 -15930 26050 -15830
rect 26300 -15930 26690 -15830
rect 26800 -15840 26810 -15830
rect 26930 -15730 26940 -15720
rect 27260 -15730 27650 -15668
rect 27900 -15730 28290 -15668
rect 28860 -15668 29257 -15630
rect 29493 -15668 29890 -15630
rect 26930 -15830 28290 -15730
rect 26930 -15840 26940 -15830
rect 26800 -15850 26940 -15840
rect 27260 -15890 27650 -15830
rect 27900 -15890 28290 -15830
rect 28400 -15720 28540 -15710
rect 28400 -15840 28410 -15720
rect 28530 -15730 28540 -15720
rect 28860 -15730 29250 -15668
rect 29500 -15730 29890 -15668
rect 30460 -15668 30857 -15630
rect 31093 -15668 31490 -15630
rect 30460 -15730 30850 -15668
rect 31100 -15730 31490 -15668
rect 28530 -15830 31490 -15730
rect 28530 -15840 28540 -15830
rect 28400 -15850 28540 -15840
rect 27260 -15930 27657 -15890
rect 27893 -15930 28290 -15890
rect 28860 -15890 29250 -15830
rect 29500 -15890 29890 -15830
rect 28860 -15930 29257 -15890
rect 29493 -15930 29890 -15890
rect 30460 -15890 30850 -15830
rect 31100 -15890 31490 -15830
rect 30460 -15930 30857 -15890
rect 31093 -15930 31490 -15890
rect 16510 -16000 16640 -15990
rect 2120 -16010 2240 -16000
rect 2120 -16430 2130 -16010
rect 2120 -16670 2130 -16630
rect 2230 -16430 2240 -16010
rect 3720 -16010 3840 -16000
rect 3720 -16430 3730 -16010
rect 2230 -16670 2240 -16630
rect 2120 -16680 2240 -16670
rect 3720 -16670 3730 -16630
rect 3830 -16430 3840 -16010
rect 5320 -16010 5440 -16000
rect 5320 -16430 5330 -16010
rect 3830 -16670 3840 -16630
rect 3720 -16680 3840 -16670
rect 5320 -16670 5330 -16630
rect 5430 -16430 5440 -16010
rect 6920 -16010 7040 -16000
rect 6920 -16430 6930 -16010
rect 5430 -16670 5440 -16630
rect 5320 -16680 5440 -16670
rect 6920 -16670 6930 -16630
rect 7030 -16430 7040 -16010
rect 8520 -16010 8640 -16000
rect 7030 -16670 7040 -16630
rect 6920 -16680 7040 -16670
rect 8520 -16670 8530 -16010
rect 8630 -16670 8640 -16010
rect 8520 -16680 8640 -16670
rect 10120 -16010 10240 -16000
rect 10120 -16670 10130 -16010
rect 10230 -16670 10240 -16010
rect 10120 -16680 10240 -16670
rect 11710 -16010 11840 -16000
rect 11710 -16670 11720 -16010
rect 11830 -16670 11840 -16010
rect 11710 -16680 11840 -16670
rect 13310 -16010 13440 -16000
rect 13310 -16670 13320 -16010
rect 13430 -16670 13440 -16010
rect 13310 -16680 13440 -16670
rect 14910 -16010 15040 -16000
rect 14910 -16670 14920 -16010
rect 15030 -16670 15040 -16010
rect 14910 -16680 15040 -16670
rect 16510 -16680 16520 -16000
rect 16630 -16680 16640 -16000
rect 16510 -16690 16640 -16680
rect 18110 -16000 18240 -15990
rect 18110 -16680 18120 -16000
rect 18230 -16680 18240 -16000
rect 18110 -16690 18240 -16680
rect 19710 -16000 19840 -15990
rect 19710 -16680 19720 -16000
rect 19830 -16680 19840 -16000
rect 19710 -16690 19840 -16680
rect 21310 -16000 21440 -15990
rect 21310 -16680 21320 -16000
rect 21430 -16680 21440 -16000
rect 21310 -16690 21440 -16680
rect 22910 -16000 23040 -15990
rect 22910 -16680 22920 -16000
rect 23030 -16680 23040 -16000
rect 22910 -16690 23040 -16680
rect 24510 -16000 24640 -15990
rect 24510 -16680 24520 -16000
rect 24630 -16680 24640 -16000
rect 24510 -16690 24640 -16680
rect 26110 -16000 26240 -15990
rect 26110 -16680 26120 -16000
rect 26230 -16680 26240 -16000
rect 26110 -16690 26240 -16680
rect 27710 -16000 27840 -15990
rect 27710 -16680 27720 -16000
rect 27830 -16680 27840 -16000
rect 27710 -16690 27840 -16680
rect 29310 -16000 29440 -15990
rect 29310 -16680 29320 -16000
rect 29430 -16680 29440 -16000
rect 29310 -16690 29440 -16680
rect 30910 -16000 31040 -15990
rect 30910 -16680 30920 -16000
rect 31030 -16680 31040 -16000
rect 30910 -16690 31040 -16680
rect -960 -16960 36260 -16760
rect 1200 -17070 1340 -17060
rect 1200 -17190 1210 -17070
rect 1330 -17080 1340 -17070
rect 2800 -17070 2940 -17060
rect 2800 -17080 2810 -17070
rect 1330 -17180 2810 -17080
rect 1330 -17190 1340 -17180
rect 1200 -17200 1340 -17190
rect 2800 -17190 2810 -17180
rect 2930 -17080 2940 -17070
rect 4400 -17070 4540 -17060
rect 4400 -17080 4410 -17070
rect 2930 -17180 4410 -17080
rect 2930 -17190 2940 -17180
rect 2800 -17200 2940 -17190
rect 4400 -17190 4410 -17180
rect 4530 -17080 4540 -17070
rect 6000 -17070 6140 -17060
rect 6000 -17080 6010 -17070
rect 4530 -17180 6010 -17080
rect 4530 -17190 4540 -17180
rect 4400 -17200 4540 -17190
rect 6000 -17190 6010 -17180
rect 6130 -17080 6140 -17070
rect 7600 -17070 7740 -17060
rect 7600 -17080 7610 -17070
rect 6130 -17180 7610 -17080
rect 6130 -17190 6140 -17180
rect 6000 -17200 6140 -17190
rect 7600 -17190 7610 -17180
rect 7730 -17080 7740 -17070
rect 9200 -17070 9340 -17060
rect 15820 -17070 15960 -17060
rect 9200 -17080 9210 -17070
rect 7730 -17180 9210 -17080
rect 7730 -17190 7740 -17180
rect 7600 -17200 7740 -17190
rect 9200 -17190 9210 -17180
rect 9330 -17080 9340 -17070
rect 12620 -17080 12760 -17070
rect 9330 -17180 10700 -17080
rect 9330 -17190 9340 -17180
rect 9200 -17200 9340 -17190
rect 12620 -17200 12630 -17080
rect 12750 -17110 12760 -17080
rect 12750 -17200 15490 -17110
rect 15820 -17190 15830 -17070
rect 15950 -17100 15960 -17070
rect 17420 -17070 17560 -17060
rect 15950 -17190 17090 -17100
rect 15820 -17200 17090 -17190
rect 17420 -17190 17430 -17070
rect 17550 -17100 17560 -17070
rect 19020 -17070 19160 -17060
rect 17550 -17190 18690 -17100
rect 17420 -17200 18690 -17190
rect 19020 -17190 19030 -17070
rect 19150 -17100 19160 -17070
rect 20620 -17070 20760 -17060
rect 19150 -17190 20290 -17100
rect 19020 -17200 20290 -17190
rect 20620 -17190 20630 -17070
rect 20750 -17100 20760 -17070
rect 22220 -17070 22360 -17060
rect 20750 -17190 21890 -17100
rect 20620 -17200 21890 -17190
rect 22220 -17190 22230 -17070
rect 22350 -17100 22360 -17070
rect 23820 -17070 23960 -17060
rect 22350 -17190 23490 -17100
rect 22220 -17200 23490 -17190
rect 23820 -17190 23830 -17070
rect 23950 -17100 23960 -17070
rect 27020 -17070 27160 -17060
rect 27020 -17100 27030 -17070
rect 23950 -17190 25090 -17100
rect 23820 -17200 25090 -17190
rect 25660 -17190 27030 -17100
rect 27150 -17100 27160 -17070
rect 28620 -17070 28760 -17060
rect 27150 -17190 28290 -17100
rect 25660 -17200 28290 -17190
rect 28620 -17190 28630 -17070
rect 28750 -17100 28760 -17070
rect 28750 -17190 31490 -17100
rect 28620 -17200 31490 -17190
rect 12620 -17210 12760 -17200
rect 1560 -17380 33200 -17260
rect 1420 -17510 1560 -17500
rect 1420 -17630 1430 -17510
rect 1550 -17520 1560 -17510
rect 1660 -17520 2060 -17430
rect 2290 -17520 2690 -17430
rect 3020 -17510 3160 -17500
rect 3020 -17520 3030 -17510
rect 1550 -17620 3030 -17520
rect 1550 -17630 1560 -17620
rect 1420 -17640 1560 -17630
rect 1660 -17640 2690 -17620
rect 3020 -17630 3030 -17620
rect 3150 -17520 3160 -17510
rect 3260 -17520 3660 -17430
rect 3890 -17520 4290 -17430
rect 4620 -17510 4760 -17500
rect 4620 -17520 4630 -17510
rect 3150 -17620 4630 -17520
rect 3150 -17630 3160 -17620
rect 3020 -17640 3160 -17630
rect 3260 -17640 4290 -17620
rect 4620 -17630 4630 -17620
rect 4750 -17520 4760 -17510
rect 4860 -17520 5260 -17430
rect 5490 -17520 5890 -17430
rect 6220 -17510 6360 -17500
rect 6220 -17520 6230 -17510
rect 4750 -17620 6230 -17520
rect 4750 -17630 4760 -17620
rect 4620 -17640 4760 -17630
rect 4860 -17640 5890 -17620
rect 6220 -17630 6230 -17620
rect 6350 -17520 6360 -17510
rect 6460 -17520 6860 -17430
rect 7090 -17520 7490 -17430
rect 7820 -17510 7960 -17500
rect 7820 -17520 7830 -17510
rect 6350 -17620 7830 -17520
rect 6350 -17630 6360 -17620
rect 6220 -17640 6360 -17630
rect 6460 -17640 7490 -17620
rect 7820 -17630 7830 -17620
rect 7950 -17520 7960 -17510
rect 8060 -17520 8460 -17430
rect 8690 -17520 9090 -17430
rect 9420 -17510 9560 -17500
rect 9420 -17520 9430 -17510
rect 7950 -17620 9430 -17520
rect 7950 -17630 7960 -17620
rect 7820 -17640 7960 -17630
rect 8060 -17640 9090 -17620
rect 9420 -17630 9430 -17620
rect 9550 -17520 9560 -17510
rect 9660 -17520 10060 -17430
rect 10290 -17520 10690 -17430
rect 9550 -17620 10690 -17520
rect 9550 -17630 9560 -17620
rect 9420 -17640 9560 -17630
rect 9660 -17640 10690 -17620
rect 1660 -17730 2060 -17640
rect 2290 -17730 2690 -17640
rect 3260 -17730 3660 -17640
rect 3890 -17730 4290 -17640
rect 4860 -17730 5260 -17640
rect 5490 -17730 5890 -17640
rect 6460 -17730 6860 -17640
rect 7090 -17730 7490 -17640
rect 8060 -17730 8460 -17640
rect 8690 -17730 9090 -17640
rect 9660 -17730 10060 -17640
rect 10290 -17730 10690 -17640
rect 12860 -17520 13260 -17430
rect 13490 -17520 13890 -17430
rect 14460 -17520 14860 -17430
rect 15090 -17520 15490 -17430
rect 12860 -17640 15490 -17520
rect 12860 -17730 13260 -17640
rect 13490 -17730 13890 -17640
rect 14460 -17730 14860 -17640
rect 15090 -17730 15490 -17640
rect 15600 -17520 15740 -17510
rect 15600 -17640 15610 -17520
rect 15730 -17530 15740 -17520
rect 16060 -17530 16450 -17430
rect 16700 -17530 17090 -17430
rect 15730 -17630 17090 -17530
rect 15730 -17640 15740 -17630
rect 15600 -17650 15740 -17640
rect 16060 -17730 16450 -17630
rect 16700 -17730 17090 -17630
rect 17200 -17520 17340 -17510
rect 17200 -17640 17210 -17520
rect 17330 -17530 17340 -17520
rect 17660 -17530 18050 -17430
rect 18300 -17530 18690 -17430
rect 17330 -17630 18690 -17530
rect 17330 -17640 17340 -17630
rect 17200 -17650 17340 -17640
rect 17660 -17730 18050 -17630
rect 18300 -17730 18690 -17630
rect 18800 -17520 18940 -17510
rect 18800 -17640 18810 -17520
rect 18930 -17530 18940 -17520
rect 19260 -17530 19650 -17430
rect 19900 -17530 20290 -17430
rect 18930 -17630 20290 -17530
rect 18930 -17640 18940 -17630
rect 18800 -17650 18940 -17640
rect 19260 -17730 19650 -17630
rect 19900 -17730 20290 -17630
rect 20400 -17520 20540 -17510
rect 20400 -17640 20410 -17520
rect 20530 -17530 20540 -17520
rect 20860 -17530 21250 -17430
rect 21500 -17530 21890 -17430
rect 20530 -17630 21890 -17530
rect 20530 -17640 20540 -17630
rect 20400 -17650 20540 -17640
rect 20860 -17730 21250 -17630
rect 21500 -17730 21890 -17630
rect 22000 -17520 22140 -17510
rect 22000 -17640 22010 -17520
rect 22130 -17530 22140 -17520
rect 22460 -17530 22850 -17430
rect 23100 -17530 23490 -17430
rect 22130 -17630 23490 -17530
rect 22130 -17640 22140 -17630
rect 22000 -17650 22140 -17640
rect 22460 -17730 22850 -17630
rect 23100 -17730 23490 -17630
rect 23600 -17520 23740 -17510
rect 23600 -17640 23610 -17520
rect 23730 -17530 23740 -17520
rect 24060 -17530 24450 -17430
rect 24700 -17530 25090 -17430
rect 23730 -17630 25090 -17530
rect 23730 -17640 23740 -17630
rect 23600 -17650 23740 -17640
rect 24060 -17730 24450 -17630
rect 24700 -17730 25090 -17630
rect 25660 -17530 26050 -17430
rect 26300 -17530 26690 -17430
rect 27260 -17468 27657 -17430
rect 27893 -17468 28290 -17430
rect 26800 -17520 26940 -17510
rect 26800 -17530 26810 -17520
rect 25660 -17630 26810 -17530
rect 25660 -17730 26050 -17630
rect 26300 -17730 26690 -17630
rect 26800 -17640 26810 -17630
rect 26930 -17530 26940 -17520
rect 27260 -17530 27650 -17468
rect 27900 -17530 28290 -17468
rect 28860 -17468 29257 -17430
rect 29493 -17468 29890 -17430
rect 26930 -17630 28290 -17530
rect 26930 -17640 26940 -17630
rect 26800 -17650 26940 -17640
rect 27260 -17690 27650 -17630
rect 27900 -17690 28290 -17630
rect 28400 -17520 28540 -17510
rect 28400 -17640 28410 -17520
rect 28530 -17530 28540 -17520
rect 28860 -17530 29250 -17468
rect 29500 -17530 29890 -17468
rect 30460 -17468 30857 -17430
rect 31093 -17468 31490 -17430
rect 30460 -17530 30850 -17468
rect 31100 -17530 31490 -17468
rect 28530 -17630 31490 -17530
rect 28530 -17640 28540 -17630
rect 28400 -17650 28540 -17640
rect 27260 -17730 27657 -17690
rect 27893 -17730 28290 -17690
rect 28860 -17690 29250 -17630
rect 29500 -17690 29890 -17630
rect 28860 -17730 29257 -17690
rect 29493 -17730 29890 -17690
rect 30460 -17690 30850 -17630
rect 31100 -17690 31490 -17630
rect 30460 -17730 30857 -17690
rect 31093 -17730 31490 -17690
rect 16510 -17800 16640 -17790
rect 2120 -17810 2240 -17800
rect 2120 -17970 2130 -17810
rect 2120 -18470 2130 -18170
rect 2230 -17970 2240 -17810
rect 3720 -17810 3840 -17800
rect 3720 -17970 3730 -17810
rect 2230 -18470 2240 -18170
rect 2120 -18480 2240 -18470
rect 3720 -18470 3730 -18170
rect 3830 -17970 3840 -17810
rect 5320 -17810 5440 -17800
rect 5320 -17970 5330 -17810
rect 3830 -18470 3840 -18170
rect 3720 -18480 3840 -18470
rect 5320 -18470 5330 -18170
rect 5430 -17970 5440 -17810
rect 6920 -17810 7040 -17800
rect 6920 -17970 6930 -17810
rect 5430 -18470 5440 -18170
rect 5320 -18480 5440 -18470
rect 6920 -18470 6930 -18170
rect 7030 -17970 7040 -17810
rect 8520 -17810 8640 -17800
rect 7030 -18470 7040 -18170
rect 6920 -18480 7040 -18470
rect 8520 -18470 8530 -17810
rect 8630 -18470 8640 -17810
rect 8520 -18480 8640 -18470
rect 10120 -17810 10240 -17800
rect 10120 -18470 10130 -17810
rect 10230 -18470 10240 -17810
rect 10120 -18480 10240 -18470
rect 11710 -17810 11840 -17800
rect 11710 -18470 11720 -17810
rect 11830 -18470 11840 -17810
rect 11710 -18480 11840 -18470
rect 13310 -17810 13440 -17800
rect 13310 -18470 13320 -17810
rect 13430 -18470 13440 -17810
rect 13310 -18480 13440 -18470
rect 14910 -17810 15040 -17800
rect 14910 -18470 14920 -17810
rect 15030 -18470 15040 -17810
rect 14910 -18480 15040 -18470
rect 16510 -18480 16520 -17800
rect 16630 -18480 16640 -17800
rect 16510 -18490 16640 -18480
rect 18110 -17800 18240 -17790
rect 18110 -18480 18120 -17800
rect 18230 -18480 18240 -17800
rect 18110 -18490 18240 -18480
rect 19710 -17800 19840 -17790
rect 19710 -18480 19720 -17800
rect 19830 -18480 19840 -17800
rect 19710 -18490 19840 -18480
rect 21310 -17800 21440 -17790
rect 21310 -18480 21320 -17800
rect 21430 -18480 21440 -17800
rect 21310 -18490 21440 -18480
rect 22910 -17800 23040 -17790
rect 22910 -18480 22920 -17800
rect 23030 -18480 23040 -17800
rect 22910 -18490 23040 -18480
rect 24510 -17800 24640 -17790
rect 24510 -18480 24520 -17800
rect 24630 -18480 24640 -17800
rect 24510 -18490 24640 -18480
rect 26110 -17800 26240 -17790
rect 26110 -18480 26120 -17800
rect 26230 -18480 26240 -17800
rect 26110 -18490 26240 -18480
rect 27710 -17800 27840 -17790
rect 27710 -18480 27720 -17800
rect 27830 -18480 27840 -17800
rect 27710 -18490 27840 -18480
rect 29310 -17800 29440 -17790
rect 29310 -18480 29320 -17800
rect 29430 -18480 29440 -17800
rect 29310 -18490 29440 -18480
rect 30910 -17800 31040 -17790
rect 30910 -18480 30920 -17800
rect 31030 -18480 31040 -17800
rect 30910 -18490 31040 -18480
rect -960 -18760 36260 -18560
rect 1200 -18870 1340 -18860
rect 1200 -18990 1210 -18870
rect 1330 -18880 1340 -18870
rect 2800 -18870 2940 -18860
rect 2800 -18880 2810 -18870
rect 1330 -18980 2810 -18880
rect 1330 -18990 1340 -18980
rect 1200 -19000 1340 -18990
rect 2800 -18990 2810 -18980
rect 2930 -18880 2940 -18870
rect 4400 -18870 4540 -18860
rect 4400 -18880 4410 -18870
rect 2930 -18980 4410 -18880
rect 2930 -18990 2940 -18980
rect 2800 -19000 2940 -18990
rect 4400 -18990 4410 -18980
rect 4530 -18880 4540 -18870
rect 6000 -18870 6140 -18860
rect 6000 -18880 6010 -18870
rect 4530 -18980 6010 -18880
rect 4530 -18990 4540 -18980
rect 4400 -19000 4540 -18990
rect 6000 -18990 6010 -18980
rect 6130 -18880 6140 -18870
rect 7600 -18870 7740 -18860
rect 7600 -18880 7610 -18870
rect 6130 -18980 7610 -18880
rect 6130 -18990 6140 -18980
rect 6000 -19000 6140 -18990
rect 7600 -18990 7610 -18980
rect 7730 -18880 7740 -18870
rect 9200 -18870 9340 -18860
rect 15820 -18870 15960 -18860
rect 9200 -18880 9210 -18870
rect 7730 -18980 9210 -18880
rect 7730 -18990 7740 -18980
rect 7600 -19000 7740 -18990
rect 9200 -18990 9210 -18980
rect 9330 -18880 9340 -18870
rect 12400 -18880 12540 -18870
rect 9330 -18980 10700 -18880
rect 9330 -18990 9340 -18980
rect 9200 -19000 9340 -18990
rect 12400 -19000 12410 -18880
rect 12530 -18910 12540 -18880
rect 12530 -19000 15490 -18910
rect 15820 -18990 15830 -18870
rect 15950 -18900 15960 -18870
rect 17420 -18870 17560 -18860
rect 15950 -18990 17090 -18900
rect 15820 -19000 17090 -18990
rect 17420 -18990 17430 -18870
rect 17550 -18900 17560 -18870
rect 19020 -18870 19160 -18860
rect 17550 -18990 18690 -18900
rect 17420 -19000 18690 -18990
rect 19020 -18990 19030 -18870
rect 19150 -18900 19160 -18870
rect 20620 -18870 20760 -18860
rect 19150 -18990 20290 -18900
rect 19020 -19000 20290 -18990
rect 20620 -18990 20630 -18870
rect 20750 -18900 20760 -18870
rect 22220 -18870 22360 -18860
rect 20750 -18990 21890 -18900
rect 20620 -19000 21890 -18990
rect 22220 -18990 22230 -18870
rect 22350 -18900 22360 -18870
rect 23820 -18870 23960 -18860
rect 22350 -18990 23490 -18900
rect 22220 -19000 23490 -18990
rect 23820 -18990 23830 -18870
rect 23950 -18900 23960 -18870
rect 27020 -18870 27160 -18860
rect 27020 -18900 27030 -18870
rect 23950 -18990 25090 -18900
rect 23820 -19000 25090 -18990
rect 25660 -18990 27030 -18900
rect 27150 -18900 27160 -18870
rect 28620 -18870 28760 -18860
rect 27150 -18990 28290 -18900
rect 25660 -19000 28290 -18990
rect 28620 -18990 28630 -18870
rect 28750 -18900 28760 -18870
rect 28750 -18990 31490 -18900
rect 28620 -19000 31490 -18990
rect 12400 -19010 12540 -19000
rect 1560 -19180 33200 -19060
rect 1420 -19310 1560 -19300
rect 1420 -19430 1430 -19310
rect 1550 -19320 1560 -19310
rect 1660 -19320 2060 -19230
rect 2290 -19320 2690 -19230
rect 3020 -19310 3160 -19300
rect 3020 -19320 3030 -19310
rect 1550 -19420 3030 -19320
rect 1550 -19430 1560 -19420
rect 1420 -19440 1560 -19430
rect 1660 -19440 2690 -19420
rect 3020 -19430 3030 -19420
rect 3150 -19320 3160 -19310
rect 3260 -19320 3660 -19230
rect 3890 -19320 4290 -19230
rect 4620 -19310 4760 -19300
rect 4620 -19320 4630 -19310
rect 3150 -19420 4630 -19320
rect 3150 -19430 3160 -19420
rect 3020 -19440 3160 -19430
rect 3260 -19440 4290 -19420
rect 4620 -19430 4630 -19420
rect 4750 -19320 4760 -19310
rect 4860 -19320 5260 -19230
rect 5490 -19320 5890 -19230
rect 6220 -19310 6360 -19300
rect 6220 -19320 6230 -19310
rect 4750 -19420 6230 -19320
rect 4750 -19430 4760 -19420
rect 4620 -19440 4760 -19430
rect 4860 -19440 5890 -19420
rect 6220 -19430 6230 -19420
rect 6350 -19320 6360 -19310
rect 6460 -19320 6860 -19230
rect 7090 -19320 7490 -19230
rect 7820 -19310 7960 -19300
rect 7820 -19320 7830 -19310
rect 6350 -19420 7830 -19320
rect 6350 -19430 6360 -19420
rect 6220 -19440 6360 -19430
rect 6460 -19440 7490 -19420
rect 7820 -19430 7830 -19420
rect 7950 -19320 7960 -19310
rect 8060 -19320 8460 -19230
rect 8690 -19320 9090 -19230
rect 9420 -19310 9560 -19300
rect 9420 -19320 9430 -19310
rect 7950 -19420 9430 -19320
rect 7950 -19430 7960 -19420
rect 7820 -19440 7960 -19430
rect 8060 -19440 9090 -19420
rect 9420 -19430 9430 -19420
rect 9550 -19320 9560 -19310
rect 9660 -19320 10060 -19230
rect 10290 -19320 10690 -19230
rect 9550 -19420 10690 -19320
rect 9550 -19430 9560 -19420
rect 9420 -19440 9560 -19430
rect 9660 -19440 10690 -19420
rect 1660 -19530 2060 -19440
rect 2290 -19530 2690 -19440
rect 3260 -19530 3660 -19440
rect 3890 -19530 4290 -19440
rect 4860 -19530 5260 -19440
rect 5490 -19530 5890 -19440
rect 6460 -19530 6860 -19440
rect 7090 -19530 7490 -19440
rect 8060 -19530 8460 -19440
rect 8690 -19530 9090 -19440
rect 9660 -19530 10060 -19440
rect 10290 -19530 10690 -19440
rect 12860 -19320 13260 -19230
rect 13490 -19320 13890 -19230
rect 14460 -19320 14860 -19230
rect 15090 -19320 15490 -19230
rect 12860 -19440 15490 -19320
rect 12860 -19530 13260 -19440
rect 13490 -19530 13890 -19440
rect 14460 -19530 14860 -19440
rect 15090 -19530 15490 -19440
rect 15600 -19320 15740 -19310
rect 15600 -19440 15610 -19320
rect 15730 -19330 15740 -19320
rect 16060 -19330 16450 -19230
rect 16700 -19330 17090 -19230
rect 15730 -19430 17090 -19330
rect 15730 -19440 15740 -19430
rect 15600 -19450 15740 -19440
rect 16060 -19530 16450 -19430
rect 16700 -19530 17090 -19430
rect 17200 -19320 17340 -19310
rect 17200 -19440 17210 -19320
rect 17330 -19330 17340 -19320
rect 17660 -19330 18050 -19230
rect 18300 -19330 18690 -19230
rect 17330 -19430 18690 -19330
rect 17330 -19440 17340 -19430
rect 17200 -19450 17340 -19440
rect 17660 -19530 18050 -19430
rect 18300 -19530 18690 -19430
rect 18800 -19320 18940 -19310
rect 18800 -19440 18810 -19320
rect 18930 -19330 18940 -19320
rect 19260 -19330 19650 -19230
rect 19900 -19330 20290 -19230
rect 18930 -19430 20290 -19330
rect 18930 -19440 18940 -19430
rect 18800 -19450 18940 -19440
rect 19260 -19530 19650 -19430
rect 19900 -19530 20290 -19430
rect 20400 -19320 20540 -19310
rect 20400 -19440 20410 -19320
rect 20530 -19330 20540 -19320
rect 20860 -19330 21250 -19230
rect 21500 -19330 21890 -19230
rect 20530 -19430 21890 -19330
rect 20530 -19440 20540 -19430
rect 20400 -19450 20540 -19440
rect 20860 -19530 21250 -19430
rect 21500 -19530 21890 -19430
rect 22000 -19320 22140 -19310
rect 22000 -19440 22010 -19320
rect 22130 -19330 22140 -19320
rect 22460 -19330 22850 -19230
rect 23100 -19330 23490 -19230
rect 22130 -19430 23490 -19330
rect 22130 -19440 22140 -19430
rect 22000 -19450 22140 -19440
rect 22460 -19530 22850 -19430
rect 23100 -19530 23490 -19430
rect 23600 -19320 23740 -19310
rect 23600 -19440 23610 -19320
rect 23730 -19330 23740 -19320
rect 24060 -19330 24450 -19230
rect 24700 -19330 25090 -19230
rect 23730 -19430 25090 -19330
rect 23730 -19440 23740 -19430
rect 23600 -19450 23740 -19440
rect 24060 -19530 24450 -19430
rect 24700 -19530 25090 -19430
rect 25660 -19330 26050 -19230
rect 26300 -19330 26690 -19230
rect 27260 -19268 27657 -19230
rect 27893 -19268 28290 -19230
rect 26800 -19320 26940 -19310
rect 26800 -19330 26810 -19320
rect 25660 -19430 26810 -19330
rect 25660 -19530 26050 -19430
rect 26300 -19530 26690 -19430
rect 26800 -19440 26810 -19430
rect 26930 -19330 26940 -19320
rect 27260 -19330 27650 -19268
rect 27900 -19330 28290 -19268
rect 28860 -19268 29257 -19230
rect 29493 -19268 29890 -19230
rect 26930 -19430 28290 -19330
rect 26930 -19440 26940 -19430
rect 26800 -19450 26940 -19440
rect 27260 -19490 27650 -19430
rect 27900 -19490 28290 -19430
rect 28400 -19320 28540 -19310
rect 28400 -19440 28410 -19320
rect 28530 -19330 28540 -19320
rect 28860 -19330 29250 -19268
rect 29500 -19330 29890 -19268
rect 30460 -19268 30857 -19230
rect 31093 -19268 31490 -19230
rect 30460 -19330 30850 -19268
rect 31100 -19330 31490 -19268
rect 28530 -19430 31490 -19330
rect 28530 -19440 28540 -19430
rect 28400 -19450 28540 -19440
rect 27260 -19530 27657 -19490
rect 27893 -19530 28290 -19490
rect 28860 -19490 29250 -19430
rect 29500 -19490 29890 -19430
rect 28860 -19530 29257 -19490
rect 29493 -19530 29890 -19490
rect 30460 -19490 30850 -19430
rect 31100 -19490 31490 -19430
rect 30460 -19530 30857 -19490
rect 31093 -19530 31490 -19490
rect 16510 -19600 16640 -19590
rect 2120 -19610 2240 -19600
rect 2120 -20170 2130 -19610
rect 2230 -20170 2240 -19610
rect 3720 -19610 3840 -19600
rect 3720 -20170 3730 -19610
rect 3830 -20170 3840 -19610
rect 5320 -19610 5440 -19600
rect 5320 -20170 5330 -19610
rect 5430 -20170 5440 -19610
rect 6920 -19610 7040 -19600
rect 6920 -20170 6930 -19610
rect 7030 -20170 7040 -19610
rect 8520 -19610 8640 -19600
rect 8520 -20270 8530 -19610
rect 8630 -20270 8640 -19610
rect 8520 -20280 8640 -20270
rect 10120 -19610 10240 -19600
rect 10120 -20270 10130 -19610
rect 10230 -20270 10240 -19610
rect 10120 -20280 10240 -20270
rect 11710 -19610 11840 -19600
rect 11710 -20270 11720 -19610
rect 11830 -20270 11840 -19610
rect 11710 -20280 11840 -20270
rect 13310 -19610 13440 -19600
rect 13310 -20270 13320 -19610
rect 13430 -20270 13440 -19610
rect 13310 -20280 13440 -20270
rect 14910 -19610 15040 -19600
rect 14910 -20270 14920 -19610
rect 15030 -20270 15040 -19610
rect 14910 -20280 15040 -20270
rect 16510 -20280 16520 -19600
rect 16630 -20280 16640 -19600
rect 16510 -20290 16640 -20280
rect 18110 -19600 18240 -19590
rect 18110 -20280 18120 -19600
rect 18230 -20280 18240 -19600
rect 18110 -20290 18240 -20280
rect 19710 -19600 19840 -19590
rect 19710 -20280 19720 -19600
rect 19830 -20280 19840 -19600
rect 19710 -20290 19840 -20280
rect 21310 -19600 21440 -19590
rect 21310 -20280 21320 -19600
rect 21430 -20280 21440 -19600
rect 21310 -20290 21440 -20280
rect 22910 -19600 23040 -19590
rect 22910 -20280 22920 -19600
rect 23030 -20280 23040 -19600
rect 22910 -20290 23040 -20280
rect 24510 -19600 24640 -19590
rect 24510 -20280 24520 -19600
rect 24630 -20280 24640 -19600
rect 24510 -20290 24640 -20280
rect 26110 -19600 26240 -19590
rect 26110 -20280 26120 -19600
rect 26230 -20280 26240 -19600
rect 26110 -20290 26240 -20280
rect 27710 -19600 27840 -19590
rect 27710 -20280 27720 -19600
rect 27830 -20280 27840 -19600
rect 27710 -20290 27840 -20280
rect 29310 -19600 29440 -19590
rect 29310 -20280 29320 -19600
rect 29430 -20280 29440 -19600
rect 29310 -20290 29440 -20280
rect 30910 -19600 31040 -19590
rect 30910 -20280 30920 -19600
rect 31030 -20280 31040 -19600
rect 30910 -20290 31040 -20280
rect -960 -20560 36260 -20360
rect 1200 -20670 1340 -20660
rect 1200 -20790 1210 -20670
rect 1330 -20680 1340 -20670
rect 2800 -20670 2940 -20660
rect 2800 -20680 2810 -20670
rect 1330 -20780 2810 -20680
rect 1330 -20790 1340 -20780
rect 1200 -20800 1340 -20790
rect 2800 -20790 2810 -20780
rect 2930 -20680 2940 -20670
rect 4400 -20670 4540 -20660
rect 4400 -20680 4410 -20670
rect 2930 -20780 4410 -20680
rect 2930 -20790 2940 -20780
rect 2800 -20800 2940 -20790
rect 4400 -20790 4410 -20780
rect 4530 -20680 4540 -20670
rect 6000 -20670 6140 -20660
rect 6000 -20680 6010 -20670
rect 4530 -20780 6010 -20680
rect 4530 -20790 4540 -20780
rect 4400 -20800 4540 -20790
rect 6000 -20790 6010 -20780
rect 6130 -20680 6140 -20670
rect 7600 -20670 7740 -20660
rect 7600 -20680 7610 -20670
rect 6130 -20780 7610 -20680
rect 6130 -20790 6140 -20780
rect 6000 -20800 6140 -20790
rect 7600 -20790 7610 -20780
rect 7730 -20680 7740 -20670
rect 9200 -20670 9340 -20660
rect 9200 -20680 9210 -20670
rect 7730 -20780 9210 -20680
rect 7730 -20790 7740 -20780
rect 7600 -20800 7740 -20790
rect 9200 -20790 9210 -20780
rect 9330 -20680 9340 -20670
rect 15820 -20670 15960 -20660
rect 9330 -20780 10700 -20680
rect 9330 -20790 9340 -20780
rect 9200 -20800 9340 -20790
rect 15820 -20790 15830 -20670
rect 15950 -20700 15960 -20670
rect 17420 -20670 17560 -20660
rect 15950 -20790 17090 -20700
rect 15820 -20800 17090 -20790
rect 17420 -20790 17430 -20670
rect 17550 -20700 17560 -20670
rect 19020 -20670 19160 -20660
rect 17550 -20790 18690 -20700
rect 17420 -20800 18690 -20790
rect 19020 -20790 19030 -20670
rect 19150 -20700 19160 -20670
rect 20620 -20670 20760 -20660
rect 19150 -20790 20290 -20700
rect 19020 -20800 20290 -20790
rect 20620 -20790 20630 -20670
rect 20750 -20700 20760 -20670
rect 22220 -20670 22360 -20660
rect 20750 -20790 21890 -20700
rect 20620 -20800 21890 -20790
rect 22220 -20790 22230 -20670
rect 22350 -20700 22360 -20670
rect 23820 -20670 23960 -20660
rect 22350 -20790 23490 -20700
rect 22220 -20800 23490 -20790
rect 23820 -20790 23830 -20670
rect 23950 -20700 23960 -20670
rect 27020 -20670 27160 -20660
rect 27020 -20700 27030 -20670
rect 23950 -20790 25090 -20700
rect 23820 -20800 25090 -20790
rect 25660 -20790 27030 -20700
rect 27150 -20700 27160 -20670
rect 28620 -20670 28760 -20660
rect 27150 -20790 28290 -20700
rect 25660 -20800 28290 -20790
rect 28620 -20790 28630 -20670
rect 28750 -20700 28760 -20670
rect 28750 -20790 31490 -20700
rect 28620 -20800 31490 -20790
rect 1560 -20980 33200 -20860
rect 1420 -21110 1560 -21100
rect 1420 -21230 1430 -21110
rect 1550 -21120 1560 -21110
rect 1660 -21120 2060 -21030
rect 2290 -21120 2690 -21030
rect 3020 -21110 3160 -21100
rect 3020 -21120 3030 -21110
rect 1550 -21220 3030 -21120
rect 1550 -21230 1560 -21220
rect 1420 -21240 1560 -21230
rect 1660 -21240 2690 -21220
rect 3020 -21230 3030 -21220
rect 3150 -21120 3160 -21110
rect 3260 -21120 3660 -21030
rect 3890 -21120 4290 -21030
rect 4620 -21110 4760 -21100
rect 4620 -21120 4630 -21110
rect 3150 -21220 4630 -21120
rect 3150 -21230 3160 -21220
rect 3020 -21240 3160 -21230
rect 3260 -21240 4290 -21220
rect 4620 -21230 4630 -21220
rect 4750 -21120 4760 -21110
rect 4860 -21120 5260 -21030
rect 5490 -21120 5890 -21030
rect 6220 -21110 6360 -21100
rect 6220 -21120 6230 -21110
rect 4750 -21220 6230 -21120
rect 4750 -21230 4760 -21220
rect 4620 -21240 4760 -21230
rect 4860 -21240 5890 -21220
rect 6220 -21230 6230 -21220
rect 6350 -21120 6360 -21110
rect 6460 -21120 6860 -21030
rect 7090 -21120 7490 -21030
rect 7820 -21110 7960 -21100
rect 7820 -21120 7830 -21110
rect 6350 -21220 7830 -21120
rect 6350 -21230 6360 -21220
rect 6220 -21240 6360 -21230
rect 6460 -21240 7490 -21220
rect 7820 -21230 7830 -21220
rect 7950 -21120 7960 -21110
rect 8060 -21120 8460 -21030
rect 8690 -21120 9090 -21030
rect 9420 -21110 9560 -21100
rect 9420 -21120 9430 -21110
rect 7950 -21220 9430 -21120
rect 7950 -21230 7960 -21220
rect 7820 -21240 7960 -21230
rect 8060 -21240 9090 -21220
rect 9420 -21230 9430 -21220
rect 9550 -21120 9560 -21110
rect 9660 -21120 10060 -21030
rect 10290 -21120 10690 -21030
rect 9550 -21220 10690 -21120
rect 9550 -21230 9560 -21220
rect 9420 -21240 9560 -21230
rect 9660 -21240 10690 -21220
rect 1660 -21330 2060 -21240
rect 2290 -21330 2690 -21240
rect 3260 -21330 3660 -21240
rect 3890 -21330 4290 -21240
rect 4860 -21330 5260 -21240
rect 5490 -21330 5890 -21240
rect 6460 -21330 6860 -21240
rect 7090 -21330 7490 -21240
rect 8060 -21330 8460 -21240
rect 8690 -21330 9090 -21240
rect 9660 -21330 10060 -21240
rect 10290 -21330 10690 -21240
rect 15600 -21120 15740 -21110
rect 15600 -21240 15610 -21120
rect 15730 -21130 15740 -21120
rect 16060 -21130 16450 -21030
rect 16700 -21130 17090 -21030
rect 15730 -21230 17090 -21130
rect 15730 -21240 15740 -21230
rect 15600 -21250 15740 -21240
rect 16060 -21330 16450 -21230
rect 16700 -21330 17090 -21230
rect 17200 -21120 17340 -21110
rect 17200 -21240 17210 -21120
rect 17330 -21130 17340 -21120
rect 17660 -21130 18050 -21030
rect 18300 -21130 18690 -21030
rect 17330 -21230 18690 -21130
rect 17330 -21240 17340 -21230
rect 17200 -21250 17340 -21240
rect 17660 -21330 18050 -21230
rect 18300 -21330 18690 -21230
rect 18800 -21120 18940 -21110
rect 18800 -21240 18810 -21120
rect 18930 -21130 18940 -21120
rect 19260 -21130 19650 -21030
rect 19900 -21130 20290 -21030
rect 18930 -21230 20290 -21130
rect 18930 -21240 18940 -21230
rect 18800 -21250 18940 -21240
rect 19260 -21330 19650 -21230
rect 19900 -21330 20290 -21230
rect 20400 -21120 20540 -21110
rect 20400 -21240 20410 -21120
rect 20530 -21130 20540 -21120
rect 20860 -21130 21250 -21030
rect 21500 -21130 21890 -21030
rect 20530 -21230 21890 -21130
rect 20530 -21240 20540 -21230
rect 20400 -21250 20540 -21240
rect 20860 -21330 21250 -21230
rect 21500 -21330 21890 -21230
rect 22000 -21120 22140 -21110
rect 22000 -21240 22010 -21120
rect 22130 -21130 22140 -21120
rect 22460 -21130 22850 -21030
rect 23100 -21130 23490 -21030
rect 22130 -21230 23490 -21130
rect 22130 -21240 22140 -21230
rect 22000 -21250 22140 -21240
rect 22460 -21330 22850 -21230
rect 23100 -21330 23490 -21230
rect 23600 -21120 23740 -21110
rect 23600 -21240 23610 -21120
rect 23730 -21130 23740 -21120
rect 24060 -21130 24450 -21030
rect 24700 -21130 25090 -21030
rect 23730 -21230 25090 -21130
rect 23730 -21240 23740 -21230
rect 23600 -21250 23740 -21240
rect 24060 -21330 24450 -21230
rect 24700 -21330 25090 -21230
rect 25660 -21130 26050 -21030
rect 26300 -21130 26690 -21030
rect 27260 -21068 27657 -21030
rect 27893 -21068 28290 -21030
rect 26800 -21120 26940 -21110
rect 26800 -21130 26810 -21120
rect 25660 -21230 26810 -21130
rect 25660 -21330 26050 -21230
rect 26300 -21330 26690 -21230
rect 26800 -21240 26810 -21230
rect 26930 -21130 26940 -21120
rect 27260 -21130 27650 -21068
rect 27900 -21130 28290 -21068
rect 28860 -21068 29257 -21030
rect 29493 -21068 29890 -21030
rect 26930 -21230 28290 -21130
rect 26930 -21240 26940 -21230
rect 26800 -21250 26940 -21240
rect 27260 -21290 27650 -21230
rect 27900 -21290 28290 -21230
rect 28400 -21120 28540 -21110
rect 28400 -21240 28410 -21120
rect 28530 -21130 28540 -21120
rect 28860 -21130 29250 -21068
rect 29500 -21130 29890 -21068
rect 30460 -21068 30857 -21030
rect 31093 -21068 31490 -21030
rect 30460 -21130 30850 -21068
rect 31100 -21130 31490 -21068
rect 28530 -21230 31490 -21130
rect 28530 -21240 28540 -21230
rect 28400 -21250 28540 -21240
rect 27260 -21330 27657 -21290
rect 27893 -21330 28290 -21290
rect 28860 -21290 29250 -21230
rect 29500 -21290 29890 -21230
rect 28860 -21330 29257 -21290
rect 29493 -21330 29890 -21290
rect 30460 -21290 30850 -21230
rect 31100 -21290 31490 -21230
rect 30460 -21330 30857 -21290
rect 31093 -21330 31490 -21290
rect 16510 -21400 16640 -21390
rect 2120 -21410 2240 -21400
rect 2120 -21490 2130 -21410
rect 2120 -22070 2130 -21690
rect 2230 -21490 2240 -21410
rect 3720 -21410 3840 -21400
rect 3720 -21490 3730 -21410
rect 2230 -22070 2240 -21690
rect 2120 -22080 2240 -22070
rect 3720 -22070 3730 -21690
rect 3830 -21490 3840 -21410
rect 5320 -21410 5440 -21400
rect 5320 -21490 5330 -21410
rect 3830 -22070 3840 -21690
rect 3720 -22080 3840 -22070
rect 5320 -22070 5330 -21690
rect 5430 -21490 5440 -21410
rect 6920 -21410 7040 -21400
rect 6920 -21490 6930 -21410
rect 5430 -22070 5440 -21690
rect 5320 -22080 5440 -22070
rect 6920 -22070 6930 -21690
rect 7030 -21490 7040 -21410
rect 8520 -21410 8640 -21400
rect 7030 -22070 7040 -21690
rect 6920 -22080 7040 -22070
rect 8520 -22070 8530 -21410
rect 8630 -22070 8640 -21410
rect 8520 -22080 8640 -22070
rect 10120 -21410 10240 -21400
rect 10120 -22070 10130 -21410
rect 10230 -22070 10240 -21410
rect 10120 -22080 10240 -22070
rect 16510 -22080 16520 -21400
rect 16630 -22080 16640 -21400
rect 16510 -22090 16640 -22080
rect 18110 -21400 18240 -21390
rect 18110 -22080 18120 -21400
rect 18230 -22080 18240 -21400
rect 18110 -22090 18240 -22080
rect 19710 -21400 19840 -21390
rect 19710 -22080 19720 -21400
rect 19830 -22080 19840 -21400
rect 19710 -22090 19840 -22080
rect 21310 -21400 21440 -21390
rect 21310 -22080 21320 -21400
rect 21430 -22080 21440 -21400
rect 21310 -22090 21440 -22080
rect 22910 -21400 23040 -21390
rect 22910 -22080 22920 -21400
rect 23030 -22080 23040 -21400
rect 22910 -22090 23040 -22080
rect 24510 -21400 24640 -21390
rect 24510 -22080 24520 -21400
rect 24630 -22080 24640 -21400
rect 24510 -22090 24640 -22080
rect 26110 -21400 26240 -21390
rect 26110 -22080 26120 -21400
rect 26230 -22080 26240 -21400
rect 26110 -22090 26240 -22080
rect 27710 -21400 27840 -21390
rect 27710 -22080 27720 -21400
rect 27830 -22080 27840 -21400
rect 27710 -22090 27840 -22080
rect 29310 -21400 29440 -21390
rect 29310 -22080 29320 -21400
rect 29430 -22080 29440 -21400
rect 29310 -22090 29440 -22080
rect 30910 -21400 31040 -21390
rect 30910 -22080 30920 -21400
rect 31030 -22080 31040 -21400
rect 30910 -22090 31040 -22080
rect -960 -22360 36260 -22160
rect 2500 -25070 4020 -25060
rect 2500 -25130 2510 -25070
rect 4010 -25130 4020 -25070
rect 2500 -25142 4020 -25130
rect 4700 -25070 6220 -25060
rect 4700 -25130 4710 -25070
rect 6210 -25130 6220 -25070
rect 4700 -25142 6220 -25130
rect 6900 -25070 8420 -25060
rect 6900 -25130 6910 -25070
rect 8410 -25130 8420 -25070
rect 6900 -25142 8420 -25130
rect 9100 -25070 10620 -25060
rect 9100 -25130 9110 -25070
rect 10610 -25130 10620 -25070
rect 9100 -25142 10620 -25130
rect 11300 -25070 12820 -25060
rect 11300 -25130 11310 -25070
rect 12810 -25130 12820 -25070
rect 11300 -25142 12820 -25130
rect 13500 -25070 15020 -25060
rect 13500 -25130 13510 -25070
rect 15010 -25130 15020 -25070
rect 13500 -25142 15020 -25130
rect 15700 -25070 17220 -25060
rect 15700 -25130 15710 -25070
rect 17210 -25130 17220 -25070
rect 15700 -25142 17220 -25130
rect 17900 -25070 19420 -25060
rect 17900 -25130 17910 -25070
rect 19410 -25130 19420 -25070
rect 17900 -25142 19420 -25130
rect 1900 -25230 2310 -25170
rect 4100 -25230 4440 -25170
rect 4500 -25230 4510 -25170
rect 6300 -25230 6640 -25170
rect 6700 -25230 6710 -25170
rect 8500 -25230 8620 -25170
rect 8680 -25230 8910 -25170
rect 10700 -25230 10820 -25170
rect 10880 -25230 11110 -25170
rect 12900 -25230 13020 -25170
rect 13080 -25230 13310 -25170
rect 15100 -25230 15220 -25170
rect 15280 -25230 15510 -25170
rect 17300 -25230 17640 -25170
rect 17700 -25230 17710 -25170
rect 19500 -25230 19840 -25170
rect 19900 -25230 19910 -25170
rect 2010 -25320 2240 -25260
rect 2300 -25320 2420 -25260
rect 4210 -25340 4440 -25280
rect 4500 -25340 4620 -25280
rect 6410 -25340 6420 -25280
rect 6480 -25340 6820 -25280
rect 8610 -25340 8620 -25280
rect 8680 -25340 9020 -25280
rect 10810 -25340 10820 -25280
rect 10880 -25340 11220 -25280
rect 13010 -25340 13020 -25280
rect 13080 -25340 13420 -25280
rect 15210 -25340 15440 -25280
rect 15500 -25340 15620 -25280
rect 17410 -25340 17640 -25280
rect 17700 -25340 17820 -25280
rect 19610 -25340 20020 -25280
rect -90 -25390 10 -25380
rect -90 -25450 -70 -25390
rect -10 -25450 10 -25390
rect -90 -25460 10 -25450
rect 2110 -25390 2210 -25380
rect 2110 -25450 2130 -25390
rect 2190 -25450 2210 -25390
rect 2110 -25460 2210 -25450
rect 4310 -25390 4410 -25380
rect 4310 -25450 4330 -25390
rect 4390 -25450 4410 -25390
rect 4310 -25460 4410 -25450
rect 6510 -25390 6610 -25380
rect 6510 -25450 6530 -25390
rect 6590 -25450 6610 -25390
rect 6510 -25460 6610 -25450
rect 8710 -25390 8810 -25380
rect 8710 -25450 8730 -25390
rect 8790 -25450 8810 -25390
rect 8710 -25460 8810 -25450
rect 10910 -25390 11010 -25380
rect 10910 -25450 10930 -25390
rect 10990 -25450 11010 -25390
rect 10910 -25460 11010 -25450
rect 13110 -25390 13210 -25380
rect 13110 -25450 13130 -25390
rect 13190 -25450 13210 -25390
rect 13110 -25460 13210 -25450
rect 15310 -25390 15410 -25380
rect 15310 -25450 15330 -25390
rect 15390 -25450 15410 -25390
rect 15310 -25460 15410 -25450
rect 17510 -25390 17610 -25380
rect 17510 -25450 17530 -25390
rect 17590 -25450 17610 -25390
rect 17510 -25460 17610 -25450
rect 19710 -25390 19810 -25380
rect 19710 -25450 19730 -25390
rect 19790 -25450 19810 -25390
rect 19710 -25460 19810 -25450
rect 21910 -25390 22010 -25380
rect 21910 -25450 21930 -25390
rect 21990 -25450 22010 -25390
rect 21910 -25460 22010 -25450
rect 2500 -25700 2700 -25460
rect 2500 -25760 2510 -25700
rect 2690 -25760 2700 -25700
rect 3160 -25700 3360 -25460
rect 3160 -25760 3170 -25700
rect 3350 -25760 3360 -25700
rect 3820 -25700 4020 -25460
rect 3820 -25760 3830 -25700
rect 4010 -25760 4020 -25700
rect 4700 -25700 4900 -25460
rect 4700 -25760 4710 -25700
rect 4890 -25760 4900 -25700
rect 5360 -25700 5560 -25460
rect 5360 -25760 5370 -25700
rect 5550 -25760 5560 -25700
rect 6020 -25700 6220 -25460
rect 6020 -25760 6030 -25700
rect 6210 -25760 6220 -25700
rect 6900 -25560 7100 -25460
rect 6900 -25620 6910 -25560
rect 7090 -25620 7100 -25560
rect 6900 -25760 7100 -25620
rect 7560 -25560 7760 -25460
rect 7560 -25620 7570 -25560
rect 7750 -25620 7760 -25560
rect 7560 -25760 7760 -25620
rect 8220 -25560 8420 -25460
rect 8220 -25620 8230 -25560
rect 8410 -25620 8420 -25560
rect 8220 -25760 8420 -25620
rect 9100 -25560 9300 -25460
rect 9100 -25620 9110 -25560
rect 9290 -25620 9300 -25560
rect 9100 -25760 9300 -25620
rect 9760 -25560 9960 -25460
rect 9760 -25620 9770 -25560
rect 9950 -25620 9960 -25560
rect 9760 -25760 9960 -25620
rect 10420 -25560 10620 -25460
rect 10420 -25620 10430 -25560
rect 10610 -25620 10620 -25560
rect 10420 -25760 10620 -25620
rect 11300 -25560 11500 -25460
rect 11300 -25620 11310 -25560
rect 11490 -25620 11500 -25560
rect 11300 -25760 11500 -25620
rect 11960 -25560 12160 -25460
rect 11960 -25620 11970 -25560
rect 12150 -25620 12160 -25560
rect 11960 -25760 12160 -25620
rect 12620 -25560 12820 -25460
rect 12620 -25620 12630 -25560
rect 12810 -25620 12820 -25560
rect 12620 -25760 12820 -25620
rect 13500 -25560 13700 -25460
rect 13500 -25620 13510 -25560
rect 13690 -25620 13700 -25560
rect 13500 -25760 13700 -25620
rect 14160 -25560 14360 -25460
rect 14160 -25620 14170 -25560
rect 14350 -25620 14360 -25560
rect 14160 -25760 14360 -25620
rect 14820 -25560 15020 -25460
rect 14820 -25620 14830 -25560
rect 15010 -25620 15020 -25560
rect 14820 -25760 15020 -25620
rect 15700 -25700 15900 -25460
rect 15700 -25760 15710 -25700
rect 15890 -25760 15900 -25700
rect 16360 -25700 16560 -25460
rect 16360 -25760 16370 -25700
rect 16550 -25760 16560 -25700
rect 17020 -25700 17220 -25460
rect 17020 -25760 17030 -25700
rect 17210 -25760 17220 -25700
rect 17900 -25700 18100 -25460
rect 17900 -25760 17910 -25700
rect 18090 -25760 18100 -25700
rect 18560 -25700 18760 -25460
rect 18560 -25760 18570 -25700
rect 18750 -25760 18760 -25700
rect 19220 -25700 19420 -25460
rect 19220 -25760 19230 -25700
rect 19410 -25760 19420 -25700
rect 2500 -25870 4020 -25860
rect 2500 -25930 2510 -25870
rect 4010 -25930 4020 -25870
rect 2500 -25942 4020 -25930
rect 4700 -25870 6220 -25860
rect 4700 -25930 4710 -25870
rect 6210 -25930 6220 -25870
rect 4700 -25942 6220 -25930
rect 6900 -25870 8420 -25860
rect 6900 -25930 6910 -25870
rect 8410 -25930 8420 -25870
rect 6900 -25942 8420 -25930
rect 9100 -25870 10620 -25860
rect 9100 -25930 9110 -25870
rect 10610 -25930 10620 -25870
rect 9100 -25942 10620 -25930
rect 11300 -25870 12820 -25860
rect 11300 -25930 11310 -25870
rect 12810 -25930 12820 -25870
rect 11300 -25942 12820 -25930
rect 13500 -25870 15020 -25860
rect 13500 -25930 13510 -25870
rect 15010 -25930 15020 -25870
rect 13500 -25942 15020 -25930
rect 15700 -25870 17220 -25860
rect 15700 -25930 15710 -25870
rect 17210 -25930 17220 -25870
rect 15700 -25942 17220 -25930
rect 17900 -25870 19420 -25860
rect 17900 -25930 17910 -25870
rect 19410 -25930 19420 -25870
rect 17900 -25942 19420 -25930
rect 1900 -26030 2310 -25970
rect 4100 -26030 4220 -25970
rect 4280 -26030 4510 -25970
rect 6300 -26030 6420 -25970
rect 6480 -26030 6710 -25970
rect 8500 -26030 8840 -25970
rect 8900 -26030 8910 -25970
rect 10700 -26030 11040 -25970
rect 11100 -26030 11110 -25970
rect 12900 -26030 13240 -25970
rect 13300 -26030 13310 -25970
rect 15100 -26030 15440 -25970
rect 15500 -26030 15510 -25970
rect 17300 -26030 17420 -25970
rect 17480 -26030 17710 -25970
rect 19500 -26030 19620 -25970
rect 19680 -26030 19910 -25970
rect 2010 -26120 2020 -26060
rect 2080 -26120 2420 -26060
rect 4210 -26140 4220 -26080
rect 4280 -26140 4620 -26080
rect 6410 -26140 6640 -26080
rect 6700 -26140 6820 -26080
rect 8610 -26140 8840 -26080
rect 8900 -26140 9020 -26080
rect 10810 -26140 11040 -26080
rect 11100 -26140 11220 -26080
rect 13010 -26140 13240 -26080
rect 13300 -26140 13420 -26080
rect 15210 -26140 15220 -26080
rect 15280 -26140 15620 -26080
rect 17410 -26140 17420 -26080
rect 17480 -26140 17820 -26080
rect 19610 -26140 20020 -26080
rect -90 -26190 10 -26180
rect -90 -26250 -70 -26190
rect -10 -26250 10 -26190
rect -90 -26260 10 -26250
rect 2110 -26190 2210 -26180
rect 2110 -26250 2130 -26190
rect 2190 -26250 2210 -26190
rect 2110 -26260 2210 -26250
rect 4310 -26190 4410 -26180
rect 4310 -26250 4330 -26190
rect 4390 -26250 4410 -26190
rect 4310 -26260 4410 -26250
rect 6510 -26190 6610 -26180
rect 6510 -26250 6530 -26190
rect 6590 -26250 6610 -26190
rect 6510 -26260 6610 -26250
rect 8710 -26190 8810 -26180
rect 8710 -26250 8730 -26190
rect 8790 -26250 8810 -26190
rect 8710 -26260 8810 -26250
rect 10910 -26190 11010 -26180
rect 10910 -26250 10930 -26190
rect 10990 -26250 11010 -26190
rect 10910 -26260 11010 -26250
rect 13110 -26190 13210 -26180
rect 13110 -26250 13130 -26190
rect 13190 -26250 13210 -26190
rect 13110 -26260 13210 -26250
rect 15310 -26190 15410 -26180
rect 15310 -26250 15330 -26190
rect 15390 -26250 15410 -26190
rect 15310 -26260 15410 -26250
rect 17510 -26190 17610 -26180
rect 17510 -26250 17530 -26190
rect 17590 -26250 17610 -26190
rect 17510 -26260 17610 -26250
rect 19710 -26190 19810 -26180
rect 19710 -26250 19730 -26190
rect 19790 -26250 19810 -26190
rect 19710 -26260 19810 -26250
rect 21910 -26190 22010 -26180
rect 21910 -26250 21930 -26190
rect 21990 -26250 22010 -26190
rect 21910 -26260 22010 -26250
rect 2500 -26360 2700 -26260
rect 2500 -26420 2510 -26360
rect 2690 -26420 2700 -26360
rect 2500 -26560 2700 -26420
rect 3160 -26360 3360 -26260
rect 3160 -26420 3170 -26360
rect 3350 -26420 3360 -26360
rect 3160 -26560 3360 -26420
rect 3820 -26360 4020 -26260
rect 3820 -26420 3830 -26360
rect 4010 -26420 4020 -26360
rect 3820 -26560 4020 -26420
rect 4700 -26360 4900 -26260
rect 4700 -26420 4710 -26360
rect 4890 -26420 4900 -26360
rect 4700 -26560 4900 -26420
rect 5360 -26360 5560 -26260
rect 5360 -26420 5370 -26360
rect 5550 -26420 5560 -26360
rect 5360 -26560 5560 -26420
rect 6020 -26360 6220 -26260
rect 6020 -26420 6030 -26360
rect 6210 -26420 6220 -26360
rect 6020 -26560 6220 -26420
rect 6900 -26500 7100 -26260
rect 6900 -26560 6910 -26500
rect 7090 -26560 7100 -26500
rect 7560 -26500 7760 -26260
rect 7560 -26560 7570 -26500
rect 7750 -26560 7760 -26500
rect 8220 -26500 8420 -26260
rect 8220 -26560 8230 -26500
rect 8410 -26560 8420 -26500
rect 9100 -26500 9300 -26260
rect 9100 -26560 9110 -26500
rect 9290 -26560 9300 -26500
rect 9760 -26500 9960 -26260
rect 9760 -26560 9770 -26500
rect 9950 -26560 9960 -26500
rect 10420 -26500 10620 -26260
rect 10420 -26560 10430 -26500
rect 10610 -26560 10620 -26500
rect 11300 -26500 11500 -26260
rect 11300 -26560 11310 -26500
rect 11490 -26560 11500 -26500
rect 11960 -26500 12160 -26260
rect 11960 -26560 11970 -26500
rect 12150 -26560 12160 -26500
rect 12620 -26500 12820 -26260
rect 12620 -26560 12630 -26500
rect 12810 -26560 12820 -26500
rect 13500 -26500 13700 -26260
rect 13500 -26560 13510 -26500
rect 13690 -26560 13700 -26500
rect 14160 -26500 14360 -26260
rect 14160 -26560 14170 -26500
rect 14350 -26560 14360 -26500
rect 14820 -26500 15020 -26260
rect 14820 -26560 14830 -26500
rect 15010 -26560 15020 -26500
rect 15700 -26360 15900 -26260
rect 15700 -26420 15710 -26360
rect 15890 -26420 15900 -26360
rect 15700 -26560 15900 -26420
rect 16360 -26360 16560 -26260
rect 16360 -26420 16370 -26360
rect 16550 -26420 16560 -26360
rect 16360 -26560 16560 -26420
rect 17020 -26360 17220 -26260
rect 17020 -26420 17030 -26360
rect 17210 -26420 17220 -26360
rect 17020 -26560 17220 -26420
rect 17900 -26360 18100 -26260
rect 17900 -26420 17910 -26360
rect 18090 -26420 18100 -26360
rect 17900 -26560 18100 -26420
rect 18560 -26360 18760 -26260
rect 18560 -26420 18570 -26360
rect 18750 -26420 18760 -26360
rect 18560 -26560 18760 -26420
rect 19220 -26360 19420 -26260
rect 19220 -26420 19230 -26360
rect 19410 -26420 19420 -26360
rect 19220 -26560 19420 -26420
rect 420 -26630 620 -26620
rect 420 -26710 430 -26630
rect 610 -26640 620 -26630
rect 21300 -26630 21500 -26620
rect 21300 -26640 21310 -26630
rect 610 -26700 4040 -26640
rect 4700 -26670 6220 -26660
rect 610 -26710 620 -26700
rect 420 -26720 620 -26710
rect 4700 -26730 4710 -26670
rect 6210 -26730 6220 -26670
rect 4700 -26742 6220 -26730
rect 6900 -26670 8420 -26660
rect 6900 -26730 6910 -26670
rect 8410 -26730 8420 -26670
rect 6900 -26742 8420 -26730
rect 9100 -26670 10620 -26660
rect 9100 -26730 9110 -26670
rect 10610 -26730 10620 -26670
rect 9100 -26742 10620 -26730
rect 11300 -26670 12820 -26660
rect 11300 -26730 11310 -26670
rect 12810 -26730 12820 -26670
rect 11300 -26742 12820 -26730
rect 13500 -26670 15020 -26660
rect 13500 -26730 13510 -26670
rect 15010 -26730 15020 -26670
rect 13500 -26742 15020 -26730
rect 15700 -26670 17220 -26660
rect 15700 -26730 15710 -26670
rect 17210 -26730 17220 -26670
rect 17880 -26700 21310 -26640
rect 21300 -26710 21310 -26700
rect 21490 -26710 21500 -26630
rect 21300 -26720 21500 -26710
rect 15700 -26742 17220 -26730
rect 1900 -26830 2310 -26770
rect 4100 -26830 4510 -26770
rect 6300 -26830 6640 -26770
rect 6700 -26830 6710 -26770
rect 8500 -26830 8620 -26770
rect 8680 -26830 8910 -26770
rect 10700 -26830 10820 -26770
rect 10880 -26830 11110 -26770
rect 12900 -26830 13020 -26770
rect 13080 -26830 13310 -26770
rect 15100 -26830 15220 -26770
rect 15280 -26830 15510 -26770
rect 17300 -26830 17640 -26770
rect 17700 -26830 17710 -26770
rect 19500 -26830 19910 -26770
rect 2010 -26920 2420 -26860
rect 4210 -26940 4440 -26880
rect 4500 -26940 4620 -26880
rect 6410 -26940 6420 -26880
rect 6480 -26940 6820 -26880
rect 8610 -26940 8620 -26880
rect 8680 -26940 9020 -26880
rect 10810 -26940 10820 -26880
rect 10880 -26940 11220 -26880
rect 13010 -26940 13020 -26880
rect 13080 -26940 13420 -26880
rect 15210 -26940 15440 -26880
rect 15500 -26940 15620 -26880
rect 17410 -26940 17820 -26880
rect 19610 -26940 20020 -26880
rect -90 -26990 10 -26980
rect -90 -27050 -70 -26990
rect -10 -27050 10 -26990
rect -90 -27060 10 -27050
rect 2110 -26990 2210 -26980
rect 2110 -27050 2130 -26990
rect 2190 -27050 2210 -26990
rect 2110 -27060 2210 -27050
rect 4310 -26990 4410 -26980
rect 4310 -27050 4330 -26990
rect 4390 -27050 4410 -26990
rect 4310 -27060 4410 -27050
rect 6510 -26990 6610 -26980
rect 6510 -27050 6530 -26990
rect 6590 -27050 6610 -26990
rect 6510 -27060 6610 -27050
rect 8710 -26990 8810 -26980
rect 8710 -27050 8730 -26990
rect 8790 -27050 8810 -26990
rect 8710 -27060 8810 -27050
rect 10910 -26990 11010 -26980
rect 10910 -27050 10930 -26990
rect 10990 -27050 11010 -26990
rect 10910 -27060 11010 -27050
rect 13110 -26990 13210 -26980
rect 13110 -27050 13130 -26990
rect 13190 -27050 13210 -26990
rect 13110 -27060 13210 -27050
rect 15310 -26990 15410 -26980
rect 15310 -27050 15330 -26990
rect 15390 -27050 15410 -26990
rect 15310 -27060 15410 -27050
rect 17510 -26990 17610 -26980
rect 17510 -27050 17530 -26990
rect 17590 -27050 17610 -26990
rect 17510 -27060 17610 -27050
rect 19710 -26990 19810 -26980
rect 19710 -27050 19730 -26990
rect 19790 -27050 19810 -26990
rect 19710 -27060 19810 -27050
rect 21910 -26990 22010 -26980
rect 21910 -27050 21930 -26990
rect 21990 -27050 22010 -26990
rect 21910 -27060 22010 -27050
rect 2500 -27300 2700 -27060
rect 2500 -27360 2510 -27300
rect 2690 -27360 2700 -27300
rect 3160 -27300 3360 -27060
rect 3160 -27360 3170 -27300
rect 3350 -27360 3360 -27300
rect 3820 -27300 4020 -27060
rect 3820 -27360 3830 -27300
rect 4010 -27360 4020 -27300
rect 4700 -27300 4900 -27060
rect 4700 -27360 4710 -27300
rect 4890 -27360 4900 -27300
rect 5360 -27300 5560 -27060
rect 5360 -27360 5370 -27300
rect 5550 -27360 5560 -27300
rect 6020 -27300 6220 -27060
rect 6020 -27360 6030 -27300
rect 6210 -27360 6220 -27300
rect 6900 -27160 7100 -27060
rect 6900 -27220 6910 -27160
rect 7090 -27220 7100 -27160
rect 6900 -27360 7100 -27220
rect 7560 -27160 7760 -27060
rect 7560 -27220 7570 -27160
rect 7750 -27220 7760 -27160
rect 7560 -27360 7760 -27220
rect 8220 -27160 8420 -27060
rect 8220 -27220 8230 -27160
rect 8410 -27220 8420 -27160
rect 8220 -27360 8420 -27220
rect 9100 -27160 9300 -27060
rect 9100 -27220 9110 -27160
rect 9290 -27220 9300 -27160
rect 9100 -27360 9300 -27220
rect 9760 -27160 9960 -27060
rect 9760 -27220 9770 -27160
rect 9950 -27220 9960 -27160
rect 9760 -27360 9960 -27220
rect 10420 -27160 10620 -27060
rect 10420 -27220 10430 -27160
rect 10610 -27220 10620 -27160
rect 10420 -27360 10620 -27220
rect 11300 -27160 11500 -27060
rect 11300 -27220 11310 -27160
rect 11490 -27220 11500 -27160
rect 11300 -27360 11500 -27220
rect 11960 -27160 12160 -27060
rect 11960 -27220 11970 -27160
rect 12150 -27220 12160 -27160
rect 11960 -27360 12160 -27220
rect 12620 -27160 12820 -27060
rect 12620 -27220 12630 -27160
rect 12810 -27220 12820 -27160
rect 12620 -27360 12820 -27220
rect 13500 -27160 13700 -27060
rect 13500 -27220 13510 -27160
rect 13690 -27220 13700 -27160
rect 13500 -27360 13700 -27220
rect 14160 -27160 14360 -27060
rect 14160 -27220 14170 -27160
rect 14350 -27220 14360 -27160
rect 14160 -27360 14360 -27220
rect 14820 -27160 15020 -27060
rect 14820 -27220 14830 -27160
rect 15010 -27220 15020 -27160
rect 14820 -27360 15020 -27220
rect 15700 -27300 15900 -27060
rect 15700 -27360 15710 -27300
rect 15890 -27360 15900 -27300
rect 16360 -27300 16560 -27060
rect 16360 -27360 16370 -27300
rect 16550 -27360 16560 -27300
rect 17020 -27300 17220 -27060
rect 17020 -27360 17030 -27300
rect 17210 -27360 17220 -27300
rect 17900 -27300 18100 -27060
rect 17900 -27360 17910 -27300
rect 18090 -27360 18100 -27300
rect 18560 -27300 18760 -27060
rect 18560 -27360 18570 -27300
rect 18750 -27360 18760 -27300
rect 19220 -27300 19420 -27060
rect 19220 -27360 19230 -27300
rect 19410 -27360 19420 -27300
rect 420 -27430 620 -27420
rect 420 -27510 430 -27430
rect 610 -27440 620 -27430
rect 21300 -27430 21500 -27420
rect 21300 -27440 21310 -27430
rect 610 -27500 4040 -27440
rect 4700 -27470 6220 -27460
rect 610 -27510 620 -27500
rect 420 -27520 620 -27510
rect 4700 -27530 4710 -27470
rect 6210 -27530 6220 -27470
rect 4700 -27542 6220 -27530
rect 6900 -27470 8420 -27460
rect 6900 -27530 6910 -27470
rect 8410 -27530 8420 -27470
rect 6900 -27542 8420 -27530
rect 9100 -27470 10620 -27460
rect 9100 -27530 9110 -27470
rect 10610 -27530 10620 -27470
rect 9100 -27542 10620 -27530
rect 11300 -27470 12820 -27460
rect 11300 -27530 11310 -27470
rect 12810 -27530 12820 -27470
rect 11300 -27542 12820 -27530
rect 13500 -27470 15020 -27460
rect 13500 -27530 13510 -27470
rect 15010 -27530 15020 -27470
rect 13500 -27542 15020 -27530
rect 15700 -27470 17220 -27460
rect 15700 -27530 15710 -27470
rect 17210 -27530 17220 -27470
rect 17880 -27500 21310 -27440
rect 21300 -27510 21310 -27500
rect 21490 -27510 21500 -27430
rect 21300 -27520 21500 -27510
rect 15700 -27542 17220 -27530
rect 1900 -27630 2310 -27570
rect 4100 -27630 4510 -27570
rect 6300 -27630 6420 -27570
rect 6480 -27630 6710 -27570
rect 8500 -27630 8840 -27570
rect 8900 -27630 8910 -27570
rect 10700 -27630 11040 -27570
rect 11100 -27630 11110 -27570
rect 12900 -27630 13240 -27570
rect 13300 -27630 13310 -27570
rect 15100 -27630 15440 -27570
rect 15500 -27630 15510 -27570
rect 17300 -27630 17420 -27570
rect 17480 -27630 17710 -27570
rect 19500 -27630 19910 -27570
rect 2010 -27720 2420 -27660
rect 4210 -27740 4220 -27680
rect 4280 -27740 4620 -27680
rect 6410 -27740 6640 -27680
rect 6700 -27740 6820 -27680
rect 8610 -27740 8840 -27680
rect 8900 -27740 9020 -27680
rect 10810 -27740 11040 -27680
rect 11100 -27740 11220 -27680
rect 13010 -27740 13240 -27680
rect 13300 -27740 13420 -27680
rect 15210 -27740 15220 -27680
rect 15280 -27740 15620 -27680
rect 17410 -27740 17820 -27680
rect 19610 -27740 20020 -27680
rect -90 -27790 10 -27780
rect -90 -27850 -70 -27790
rect -10 -27850 10 -27790
rect -90 -27860 10 -27850
rect 2110 -27790 2210 -27780
rect 2110 -27850 2130 -27790
rect 2190 -27850 2210 -27790
rect 2110 -27860 2210 -27850
rect 4310 -27790 4410 -27780
rect 4310 -27850 4330 -27790
rect 4390 -27850 4410 -27790
rect 4310 -27860 4410 -27850
rect 6510 -27790 6610 -27780
rect 6510 -27850 6530 -27790
rect 6590 -27850 6610 -27790
rect 6510 -27860 6610 -27850
rect 8710 -27790 8810 -27780
rect 8710 -27850 8730 -27790
rect 8790 -27850 8810 -27790
rect 8710 -27860 8810 -27850
rect 10910 -27790 11010 -27780
rect 10910 -27850 10930 -27790
rect 10990 -27850 11010 -27790
rect 10910 -27860 11010 -27850
rect 13110 -27790 13210 -27780
rect 13110 -27850 13130 -27790
rect 13190 -27850 13210 -27790
rect 13110 -27860 13210 -27850
rect 15310 -27790 15410 -27780
rect 15310 -27850 15330 -27790
rect 15390 -27850 15410 -27790
rect 15310 -27860 15410 -27850
rect 17510 -27790 17610 -27780
rect 17510 -27850 17530 -27790
rect 17590 -27850 17610 -27790
rect 17510 -27860 17610 -27850
rect 19710 -27790 19810 -27780
rect 19710 -27850 19730 -27790
rect 19790 -27850 19810 -27790
rect 19710 -27860 19810 -27850
rect 21910 -27790 22010 -27780
rect 21910 -27850 21930 -27790
rect 21990 -27850 22010 -27790
rect 21910 -27860 22010 -27850
rect 2500 -27960 2700 -27860
rect 2500 -28020 2510 -27960
rect 2690 -28020 2700 -27960
rect 2500 -28160 2700 -28020
rect 3160 -27960 3360 -27860
rect 3160 -28020 3170 -27960
rect 3350 -28020 3360 -27960
rect 3160 -28160 3360 -28020
rect 3820 -27960 4020 -27860
rect 3820 -28020 3830 -27960
rect 4010 -28020 4020 -27960
rect 3820 -28160 4020 -28020
rect 4700 -27960 4900 -27860
rect 4700 -28020 4710 -27960
rect 4890 -28020 4900 -27960
rect 4700 -28160 4900 -28020
rect 5360 -27960 5560 -27860
rect 5360 -28020 5370 -27960
rect 5550 -28020 5560 -27960
rect 5360 -28160 5560 -28020
rect 6020 -27960 6220 -27860
rect 6020 -28020 6030 -27960
rect 6210 -28020 6220 -27960
rect 6020 -28160 6220 -28020
rect 6900 -28100 7100 -27860
rect 6900 -28160 6910 -28100
rect 7090 -28160 7100 -28100
rect 7560 -28100 7760 -27860
rect 7560 -28160 7570 -28100
rect 7750 -28160 7760 -28100
rect 8220 -28100 8420 -27860
rect 8220 -28160 8230 -28100
rect 8410 -28160 8420 -28100
rect 9100 -28100 9300 -27860
rect 9100 -28160 9110 -28100
rect 9290 -28160 9300 -28100
rect 9760 -28100 9960 -27860
rect 9760 -28160 9770 -28100
rect 9950 -28160 9960 -28100
rect 10420 -28100 10620 -27860
rect 10420 -28160 10430 -28100
rect 10610 -28160 10620 -28100
rect 11300 -28100 11500 -27860
rect 11300 -28160 11310 -28100
rect 11490 -28160 11500 -28100
rect 11960 -28100 12160 -27860
rect 11960 -28160 11970 -28100
rect 12150 -28160 12160 -28100
rect 12620 -28100 12820 -27860
rect 12620 -28160 12630 -28100
rect 12810 -28160 12820 -28100
rect 13500 -28100 13700 -27860
rect 13500 -28160 13510 -28100
rect 13690 -28160 13700 -28100
rect 14160 -28100 14360 -27860
rect 14160 -28160 14170 -28100
rect 14350 -28160 14360 -28100
rect 14820 -28100 15020 -27860
rect 14820 -28160 14830 -28100
rect 15010 -28160 15020 -28100
rect 15700 -27960 15900 -27860
rect 15700 -28020 15710 -27960
rect 15890 -28020 15900 -27960
rect 15700 -28160 15900 -28020
rect 16360 -27960 16560 -27860
rect 16360 -28020 16370 -27960
rect 16550 -28020 16560 -27960
rect 16360 -28160 16560 -28020
rect 17020 -27960 17220 -27860
rect 17020 -28020 17030 -27960
rect 17210 -28020 17220 -27960
rect 17020 -28160 17220 -28020
rect 17900 -27960 18100 -27860
rect 17900 -28020 17910 -27960
rect 18090 -28020 18100 -27960
rect 17900 -28160 18100 -28020
rect 18560 -27960 18760 -27860
rect 18560 -28020 18570 -27960
rect 18750 -28020 18760 -27960
rect 18560 -28160 18760 -28020
rect 19220 -27960 19420 -27860
rect 19220 -28020 19230 -27960
rect 19410 -28020 19420 -27960
rect 19220 -28160 19420 -28020
rect 420 -28230 620 -28220
rect 420 -28310 430 -28230
rect 610 -28240 620 -28230
rect 21300 -28230 21500 -28220
rect 21300 -28240 21310 -28230
rect 610 -28300 4040 -28240
rect 4700 -28270 6220 -28260
rect 610 -28310 620 -28300
rect 420 -28320 620 -28310
rect 4700 -28330 4710 -28270
rect 6210 -28330 6220 -28270
rect 4700 -28342 6220 -28330
rect 6900 -28270 8420 -28260
rect 6900 -28330 6910 -28270
rect 8410 -28330 8420 -28270
rect 6900 -28342 8420 -28330
rect 9100 -28270 10620 -28260
rect 9100 -28330 9110 -28270
rect 10610 -28330 10620 -28270
rect 9100 -28342 10620 -28330
rect 11300 -28270 12820 -28260
rect 11300 -28330 11310 -28270
rect 12810 -28330 12820 -28270
rect 11300 -28342 12820 -28330
rect 13500 -28270 15020 -28260
rect 13500 -28330 13510 -28270
rect 15010 -28330 15020 -28270
rect 13500 -28342 15020 -28330
rect 15700 -28270 17220 -28260
rect 15700 -28330 15710 -28270
rect 17210 -28330 17220 -28270
rect 17880 -28300 21310 -28240
rect 21300 -28310 21310 -28300
rect 21490 -28310 21500 -28230
rect 21300 -28320 21500 -28310
rect 15700 -28342 17220 -28330
rect 1900 -28430 2310 -28370
rect 4100 -28430 4510 -28370
rect 6300 -28430 6420 -28370
rect 6480 -28430 6710 -28370
rect 8500 -28430 8840 -28370
rect 8900 -28430 8910 -28370
rect 10700 -28430 11040 -28370
rect 11100 -28430 11110 -28370
rect 12900 -28430 13240 -28370
rect 13300 -28430 13310 -28370
rect 15100 -28430 15440 -28370
rect 15500 -28430 15510 -28370
rect 17300 -28430 17420 -28370
rect 17480 -28430 17710 -28370
rect 19500 -28430 19910 -28370
rect 2010 -28520 2420 -28460
rect 4210 -28540 4220 -28480
rect 4280 -28540 4620 -28480
rect 6410 -28540 6640 -28480
rect 6700 -28540 6820 -28480
rect 8610 -28540 8840 -28480
rect 8900 -28540 9020 -28480
rect 10810 -28540 11040 -28480
rect 11100 -28540 11220 -28480
rect 13010 -28540 13240 -28480
rect 13300 -28540 13420 -28480
rect 15210 -28540 15220 -28480
rect 15280 -28540 15620 -28480
rect 17410 -28540 17820 -28480
rect 19610 -28540 20020 -28480
rect -90 -28590 10 -28580
rect -90 -28650 -70 -28590
rect -10 -28650 10 -28590
rect -90 -28660 10 -28650
rect 2110 -28590 2210 -28580
rect 2110 -28650 2130 -28590
rect 2190 -28650 2210 -28590
rect 2110 -28660 2210 -28650
rect 4310 -28590 4410 -28580
rect 4310 -28650 4330 -28590
rect 4390 -28650 4410 -28590
rect 4310 -28660 4410 -28650
rect 6510 -28590 6610 -28580
rect 6510 -28650 6530 -28590
rect 6590 -28650 6610 -28590
rect 6510 -28660 6610 -28650
rect 8710 -28590 8810 -28580
rect 8710 -28650 8730 -28590
rect 8790 -28650 8810 -28590
rect 8710 -28660 8810 -28650
rect 10910 -28590 11010 -28580
rect 10910 -28650 10930 -28590
rect 10990 -28650 11010 -28590
rect 10910 -28660 11010 -28650
rect 13110 -28590 13210 -28580
rect 13110 -28650 13130 -28590
rect 13190 -28650 13210 -28590
rect 13110 -28660 13210 -28650
rect 15310 -28590 15410 -28580
rect 15310 -28650 15330 -28590
rect 15390 -28650 15410 -28590
rect 15310 -28660 15410 -28650
rect 17510 -28590 17610 -28580
rect 17510 -28650 17530 -28590
rect 17590 -28650 17610 -28590
rect 17510 -28660 17610 -28650
rect 19710 -28590 19810 -28580
rect 19710 -28650 19730 -28590
rect 19790 -28650 19810 -28590
rect 19710 -28660 19810 -28650
rect 21910 -28590 22010 -28580
rect 21910 -28650 21930 -28590
rect 21990 -28650 22010 -28590
rect 21910 -28660 22010 -28650
rect 2500 -28760 2700 -28660
rect 2500 -28820 2510 -28760
rect 2690 -28820 2700 -28760
rect 2500 -28960 2700 -28820
rect 3160 -28760 3360 -28660
rect 3160 -28820 3170 -28760
rect 3350 -28820 3360 -28760
rect 3160 -28960 3360 -28820
rect 3820 -28760 4020 -28660
rect 3820 -28820 3830 -28760
rect 4010 -28820 4020 -28760
rect 3820 -28960 4020 -28820
rect 4700 -28760 4900 -28660
rect 4700 -28820 4710 -28760
rect 4890 -28820 4900 -28760
rect 4700 -28960 4900 -28820
rect 5360 -28760 5560 -28660
rect 5360 -28820 5370 -28760
rect 5550 -28820 5560 -28760
rect 5360 -28960 5560 -28820
rect 6020 -28760 6220 -28660
rect 6020 -28820 6030 -28760
rect 6210 -28820 6220 -28760
rect 6020 -28960 6220 -28820
rect 6900 -28900 7100 -28660
rect 6900 -28960 6910 -28900
rect 7090 -28960 7100 -28900
rect 7560 -28900 7760 -28660
rect 7560 -28960 7570 -28900
rect 7750 -28960 7760 -28900
rect 8220 -28900 8420 -28660
rect 8220 -28960 8230 -28900
rect 8410 -28960 8420 -28900
rect 9100 -28900 9300 -28660
rect 9100 -28960 9110 -28900
rect 9290 -28960 9300 -28900
rect 9760 -28900 9960 -28660
rect 9760 -28960 9770 -28900
rect 9950 -28960 9960 -28900
rect 10420 -28900 10620 -28660
rect 10420 -28960 10430 -28900
rect 10610 -28960 10620 -28900
rect 11300 -28900 11500 -28660
rect 11300 -28960 11310 -28900
rect 11490 -28960 11500 -28900
rect 11960 -28900 12160 -28660
rect 11960 -28960 11970 -28900
rect 12150 -28960 12160 -28900
rect 12620 -28900 12820 -28660
rect 12620 -28960 12630 -28900
rect 12810 -28960 12820 -28900
rect 13500 -28900 13700 -28660
rect 13500 -28960 13510 -28900
rect 13690 -28960 13700 -28900
rect 14160 -28900 14360 -28660
rect 14160 -28960 14170 -28900
rect 14350 -28960 14360 -28900
rect 14820 -28900 15020 -28660
rect 14820 -28960 14830 -28900
rect 15010 -28960 15020 -28900
rect 15700 -28760 15900 -28660
rect 15700 -28820 15710 -28760
rect 15890 -28820 15900 -28760
rect 15700 -28960 15900 -28820
rect 16360 -28760 16560 -28660
rect 16360 -28820 16370 -28760
rect 16550 -28820 16560 -28760
rect 16360 -28960 16560 -28820
rect 17020 -28760 17220 -28660
rect 17020 -28820 17030 -28760
rect 17210 -28820 17220 -28760
rect 17020 -28960 17220 -28820
rect 17900 -28760 18100 -28660
rect 17900 -28820 17910 -28760
rect 18090 -28820 18100 -28760
rect 17900 -28960 18100 -28820
rect 18560 -28760 18760 -28660
rect 18560 -28820 18570 -28760
rect 18750 -28820 18760 -28760
rect 18560 -28960 18760 -28820
rect 19220 -28760 19420 -28660
rect 19220 -28820 19230 -28760
rect 19410 -28820 19420 -28760
rect 19220 -28960 19420 -28820
rect 420 -29030 620 -29020
rect 420 -29110 430 -29030
rect 610 -29040 620 -29030
rect 21300 -29030 21500 -29020
rect 21300 -29040 21310 -29030
rect 610 -29100 4040 -29040
rect 4700 -29070 6220 -29060
rect 610 -29110 620 -29100
rect 420 -29120 620 -29110
rect 4700 -29130 4710 -29070
rect 6210 -29130 6220 -29070
rect 4700 -29142 6220 -29130
rect 6900 -29070 8420 -29060
rect 6900 -29130 6910 -29070
rect 8410 -29130 8420 -29070
rect 6900 -29142 8420 -29130
rect 9100 -29070 10620 -29060
rect 9100 -29130 9110 -29070
rect 10610 -29130 10620 -29070
rect 9100 -29142 10620 -29130
rect 11300 -29070 12820 -29060
rect 11300 -29130 11310 -29070
rect 12810 -29130 12820 -29070
rect 11300 -29142 12820 -29130
rect 13500 -29070 15020 -29060
rect 13500 -29130 13510 -29070
rect 15010 -29130 15020 -29070
rect 13500 -29142 15020 -29130
rect 15700 -29070 17220 -29060
rect 15700 -29130 15710 -29070
rect 17210 -29130 17220 -29070
rect 17880 -29100 21310 -29040
rect 21300 -29110 21310 -29100
rect 21490 -29110 21500 -29030
rect 21300 -29120 21500 -29110
rect 15700 -29142 17220 -29130
rect 1900 -29230 2310 -29170
rect 4100 -29230 4510 -29170
rect 6300 -29230 6640 -29170
rect 6700 -29230 6710 -29170
rect 8500 -29230 8620 -29170
rect 8680 -29230 8910 -29170
rect 10700 -29230 10820 -29170
rect 10880 -29230 11110 -29170
rect 12900 -29230 13020 -29170
rect 13080 -29230 13310 -29170
rect 15100 -29230 15220 -29170
rect 15280 -29230 15510 -29170
rect 17300 -29230 17640 -29170
rect 17700 -29230 17710 -29170
rect 19500 -29230 19910 -29170
rect 2010 -29320 2420 -29260
rect 4210 -29340 4440 -29280
rect 4500 -29340 4620 -29280
rect 6410 -29340 6420 -29280
rect 6480 -29340 6820 -29280
rect 8610 -29340 8620 -29280
rect 8680 -29340 9020 -29280
rect 10810 -29340 10820 -29280
rect 10880 -29340 11220 -29280
rect 13010 -29340 13020 -29280
rect 13080 -29340 13420 -29280
rect 15210 -29340 15440 -29280
rect 15500 -29340 15620 -29280
rect 17410 -29340 17820 -29280
rect 19610 -29340 20020 -29280
rect -90 -29390 10 -29380
rect -90 -29450 -70 -29390
rect -10 -29450 10 -29390
rect -90 -29460 10 -29450
rect 2110 -29390 2210 -29380
rect 2110 -29450 2130 -29390
rect 2190 -29450 2210 -29390
rect 2110 -29460 2210 -29450
rect 4310 -29390 4410 -29380
rect 4310 -29450 4330 -29390
rect 4390 -29450 4410 -29390
rect 4310 -29460 4410 -29450
rect 6510 -29390 6610 -29380
rect 6510 -29450 6530 -29390
rect 6590 -29450 6610 -29390
rect 6510 -29460 6610 -29450
rect 8710 -29390 8810 -29380
rect 8710 -29450 8730 -29390
rect 8790 -29450 8810 -29390
rect 8710 -29460 8810 -29450
rect 10910 -29390 11010 -29380
rect 10910 -29450 10930 -29390
rect 10990 -29450 11010 -29390
rect 10910 -29460 11010 -29450
rect 13110 -29390 13210 -29380
rect 13110 -29450 13130 -29390
rect 13190 -29450 13210 -29390
rect 13110 -29460 13210 -29450
rect 15310 -29390 15410 -29380
rect 15310 -29450 15330 -29390
rect 15390 -29450 15410 -29390
rect 15310 -29460 15410 -29450
rect 17510 -29390 17610 -29380
rect 17510 -29450 17530 -29390
rect 17590 -29450 17610 -29390
rect 17510 -29460 17610 -29450
rect 19710 -29390 19810 -29380
rect 19710 -29450 19730 -29390
rect 19790 -29450 19810 -29390
rect 19710 -29460 19810 -29450
rect 21910 -29390 22010 -29380
rect 21910 -29450 21930 -29390
rect 21990 -29450 22010 -29390
rect 21910 -29460 22010 -29450
rect 2500 -29700 2700 -29460
rect 2500 -29760 2510 -29700
rect 2690 -29760 2700 -29700
rect 3160 -29700 3360 -29460
rect 3160 -29760 3170 -29700
rect 3350 -29760 3360 -29700
rect 3820 -29700 4020 -29460
rect 3820 -29760 3830 -29700
rect 4010 -29760 4020 -29700
rect 4700 -29700 4900 -29460
rect 4700 -29760 4710 -29700
rect 4890 -29760 4900 -29700
rect 5360 -29700 5560 -29460
rect 5360 -29760 5370 -29700
rect 5550 -29760 5560 -29700
rect 6020 -29700 6220 -29460
rect 6020 -29760 6030 -29700
rect 6210 -29760 6220 -29700
rect 6900 -29560 7100 -29460
rect 6900 -29620 6910 -29560
rect 7090 -29620 7100 -29560
rect 6900 -29760 7100 -29620
rect 7560 -29560 7760 -29460
rect 7560 -29620 7570 -29560
rect 7750 -29620 7760 -29560
rect 7560 -29760 7760 -29620
rect 8220 -29560 8420 -29460
rect 8220 -29620 8230 -29560
rect 8410 -29620 8420 -29560
rect 8220 -29760 8420 -29620
rect 9100 -29560 9300 -29460
rect 9100 -29620 9110 -29560
rect 9290 -29620 9300 -29560
rect 9100 -29760 9300 -29620
rect 9760 -29560 9960 -29460
rect 9760 -29620 9770 -29560
rect 9950 -29620 9960 -29560
rect 9760 -29760 9960 -29620
rect 10420 -29560 10620 -29460
rect 10420 -29620 10430 -29560
rect 10610 -29620 10620 -29560
rect 10420 -29760 10620 -29620
rect 11300 -29560 11500 -29460
rect 11300 -29620 11310 -29560
rect 11490 -29620 11500 -29560
rect 11300 -29760 11500 -29620
rect 11960 -29560 12160 -29460
rect 11960 -29620 11970 -29560
rect 12150 -29620 12160 -29560
rect 11960 -29760 12160 -29620
rect 12620 -29560 12820 -29460
rect 12620 -29620 12630 -29560
rect 12810 -29620 12820 -29560
rect 12620 -29760 12820 -29620
rect 13500 -29560 13700 -29460
rect 13500 -29620 13510 -29560
rect 13690 -29620 13700 -29560
rect 13500 -29760 13700 -29620
rect 14160 -29560 14360 -29460
rect 14160 -29620 14170 -29560
rect 14350 -29620 14360 -29560
rect 14160 -29760 14360 -29620
rect 14820 -29560 15020 -29460
rect 14820 -29620 14830 -29560
rect 15010 -29620 15020 -29560
rect 14820 -29760 15020 -29620
rect 15700 -29700 15900 -29460
rect 15700 -29760 15710 -29700
rect 15890 -29760 15900 -29700
rect 16360 -29700 16560 -29460
rect 16360 -29760 16370 -29700
rect 16550 -29760 16560 -29700
rect 17020 -29700 17220 -29460
rect 17020 -29760 17030 -29700
rect 17210 -29760 17220 -29700
rect 17900 -29700 18100 -29460
rect 17900 -29760 17910 -29700
rect 18090 -29760 18100 -29700
rect 18560 -29700 18760 -29460
rect 18560 -29760 18570 -29700
rect 18750 -29760 18760 -29700
rect 19220 -29700 19420 -29460
rect 19220 -29760 19230 -29700
rect 19410 -29760 19420 -29700
rect 2500 -29870 4020 -29860
rect 2500 -29930 2510 -29870
rect 4010 -29930 4020 -29870
rect 2500 -29942 4020 -29930
rect 4700 -29870 6220 -29860
rect 4700 -29930 4710 -29870
rect 6210 -29930 6220 -29870
rect 4700 -29942 6220 -29930
rect 6900 -29870 8420 -29860
rect 6900 -29930 6910 -29870
rect 8410 -29930 8420 -29870
rect 6900 -29942 8420 -29930
rect 9100 -29870 10620 -29860
rect 9100 -29930 9110 -29870
rect 10610 -29930 10620 -29870
rect 9100 -29942 10620 -29930
rect 11300 -29870 12820 -29860
rect 11300 -29930 11310 -29870
rect 12810 -29930 12820 -29870
rect 11300 -29942 12820 -29930
rect 13500 -29870 15020 -29860
rect 13500 -29930 13510 -29870
rect 15010 -29930 15020 -29870
rect 13500 -29942 15020 -29930
rect 15700 -29870 17220 -29860
rect 15700 -29930 15710 -29870
rect 17210 -29930 17220 -29870
rect 15700 -29942 17220 -29930
rect 17900 -29870 19420 -29860
rect 17900 -29930 17910 -29870
rect 19410 -29930 19420 -29870
rect 17900 -29942 19420 -29930
rect 1900 -30030 2310 -29970
rect 4100 -30030 4220 -29970
rect 4280 -30030 4510 -29970
rect 6300 -30030 6420 -29970
rect 6480 -30030 6710 -29970
rect 8500 -30030 8840 -29970
rect 8900 -30030 8910 -29970
rect 10700 -30030 11040 -29970
rect 11100 -30030 11110 -29970
rect 12900 -30030 13240 -29970
rect 13300 -30030 13310 -29970
rect 15100 -30030 15440 -29970
rect 15500 -30030 15510 -29970
rect 17300 -30030 17420 -29970
rect 17480 -30030 17710 -29970
rect 19500 -30030 19620 -29970
rect 19680 -30030 19910 -29970
rect 2010 -30120 2020 -30060
rect 2080 -30120 2420 -30060
rect 4210 -30140 4220 -30080
rect 4280 -30140 4620 -30080
rect 6410 -30140 6640 -30080
rect 6700 -30140 6820 -30080
rect 8610 -30140 8840 -30080
rect 8900 -30140 9020 -30080
rect 10810 -30140 11040 -30080
rect 11100 -30140 11220 -30080
rect 13010 -30140 13240 -30080
rect 13300 -30140 13420 -30080
rect 15210 -30140 15220 -30080
rect 15280 -30140 15620 -30080
rect 17410 -30140 17420 -30080
rect 17480 -30140 17820 -30080
rect 19610 -30140 20020 -30080
rect -90 -30190 10 -30180
rect -90 -30250 -70 -30190
rect -10 -30250 10 -30190
rect -90 -30260 10 -30250
rect 2110 -30190 2210 -30180
rect 2110 -30250 2130 -30190
rect 2190 -30250 2210 -30190
rect 2110 -30260 2210 -30250
rect 4310 -30190 4410 -30180
rect 4310 -30250 4330 -30190
rect 4390 -30250 4410 -30190
rect 4310 -30260 4410 -30250
rect 6510 -30190 6610 -30180
rect 6510 -30250 6530 -30190
rect 6590 -30250 6610 -30190
rect 6510 -30260 6610 -30250
rect 8710 -30190 8810 -30180
rect 8710 -30250 8730 -30190
rect 8790 -30250 8810 -30190
rect 8710 -30260 8810 -30250
rect 10910 -30190 11010 -30180
rect 10910 -30250 10930 -30190
rect 10990 -30250 11010 -30190
rect 10910 -30260 11010 -30250
rect 13110 -30190 13210 -30180
rect 13110 -30250 13130 -30190
rect 13190 -30250 13210 -30190
rect 13110 -30260 13210 -30250
rect 15310 -30190 15410 -30180
rect 15310 -30250 15330 -30190
rect 15390 -30250 15410 -30190
rect 15310 -30260 15410 -30250
rect 17510 -30190 17610 -30180
rect 17510 -30250 17530 -30190
rect 17590 -30250 17610 -30190
rect 17510 -30260 17610 -30250
rect 19710 -30190 19810 -30180
rect 19710 -30250 19730 -30190
rect 19790 -30250 19810 -30190
rect 19710 -30260 19810 -30250
rect 21910 -30190 22010 -30180
rect 21910 -30250 21930 -30190
rect 21990 -30250 22010 -30190
rect 21910 -30260 22010 -30250
rect 2500 -30360 2700 -30260
rect 2500 -30420 2510 -30360
rect 2690 -30420 2700 -30360
rect 2500 -30560 2700 -30420
rect 3160 -30360 3360 -30260
rect 3160 -30420 3170 -30360
rect 3350 -30420 3360 -30360
rect 3160 -30560 3360 -30420
rect 3820 -30360 4020 -30260
rect 3820 -30420 3830 -30360
rect 4010 -30420 4020 -30360
rect 3820 -30560 4020 -30420
rect 4700 -30360 4900 -30260
rect 4700 -30420 4710 -30360
rect 4890 -30420 4900 -30360
rect 4700 -30560 4900 -30420
rect 5360 -30360 5560 -30260
rect 5360 -30420 5370 -30360
rect 5550 -30420 5560 -30360
rect 5360 -30560 5560 -30420
rect 6020 -30360 6220 -30260
rect 6020 -30420 6030 -30360
rect 6210 -30420 6220 -30360
rect 6020 -30560 6220 -30420
rect 6900 -30500 7100 -30260
rect 6900 -30560 6910 -30500
rect 7090 -30560 7100 -30500
rect 7560 -30500 7760 -30260
rect 7560 -30560 7570 -30500
rect 7750 -30560 7760 -30500
rect 8220 -30500 8420 -30260
rect 8220 -30560 8230 -30500
rect 8410 -30560 8420 -30500
rect 9100 -30500 9300 -30260
rect 9100 -30560 9110 -30500
rect 9290 -30560 9300 -30500
rect 9760 -30500 9960 -30260
rect 9760 -30560 9770 -30500
rect 9950 -30560 9960 -30500
rect 10420 -30500 10620 -30260
rect 10420 -30560 10430 -30500
rect 10610 -30560 10620 -30500
rect 11300 -30500 11500 -30260
rect 11300 -30560 11310 -30500
rect 11490 -30560 11500 -30500
rect 11960 -30500 12160 -30260
rect 11960 -30560 11970 -30500
rect 12150 -30560 12160 -30500
rect 12620 -30500 12820 -30260
rect 12620 -30560 12630 -30500
rect 12810 -30560 12820 -30500
rect 13500 -30500 13700 -30260
rect 13500 -30560 13510 -30500
rect 13690 -30560 13700 -30500
rect 14160 -30500 14360 -30260
rect 14160 -30560 14170 -30500
rect 14350 -30560 14360 -30500
rect 14820 -30500 15020 -30260
rect 14820 -30560 14830 -30500
rect 15010 -30560 15020 -30500
rect 15700 -30360 15900 -30260
rect 15700 -30420 15710 -30360
rect 15890 -30420 15900 -30360
rect 15700 -30560 15900 -30420
rect 16360 -30360 16560 -30260
rect 16360 -30420 16370 -30360
rect 16550 -30420 16560 -30360
rect 16360 -30560 16560 -30420
rect 17020 -30360 17220 -30260
rect 17020 -30420 17030 -30360
rect 17210 -30420 17220 -30360
rect 17020 -30560 17220 -30420
rect 17900 -30360 18100 -30260
rect 17900 -30420 17910 -30360
rect 18090 -30420 18100 -30360
rect 17900 -30560 18100 -30420
rect 18560 -30360 18760 -30260
rect 18560 -30420 18570 -30360
rect 18750 -30420 18760 -30360
rect 18560 -30560 18760 -30420
rect 19220 -30360 19420 -30260
rect 19220 -30420 19230 -30360
rect 19410 -30420 19420 -30360
rect 19220 -30560 19420 -30420
rect 2500 -30670 4020 -30660
rect 2500 -30730 2510 -30670
rect 4010 -30730 4020 -30670
rect 2500 -30742 4020 -30730
rect 4700 -30670 6220 -30660
rect 4700 -30730 4710 -30670
rect 6210 -30730 6220 -30670
rect 4700 -30742 6220 -30730
rect 6900 -30670 8420 -30660
rect 6900 -30730 6910 -30670
rect 8410 -30730 8420 -30670
rect 6900 -30742 8420 -30730
rect 9100 -30670 10620 -30660
rect 9100 -30730 9110 -30670
rect 10610 -30730 10620 -30670
rect 9100 -30742 10620 -30730
rect 11300 -30670 12820 -30660
rect 11300 -30730 11310 -30670
rect 12810 -30730 12820 -30670
rect 11300 -30742 12820 -30730
rect 13500 -30670 15020 -30660
rect 13500 -30730 13510 -30670
rect 15010 -30730 15020 -30670
rect 13500 -30742 15020 -30730
rect 15700 -30670 17220 -30660
rect 15700 -30730 15710 -30670
rect 17210 -30730 17220 -30670
rect 15700 -30742 17220 -30730
rect 17900 -30670 19420 -30660
rect 17900 -30730 17910 -30670
rect 19410 -30730 19420 -30670
rect 17900 -30740 19420 -30730
rect 1900 -30830 2310 -30770
rect 4100 -30830 4440 -30770
rect 4500 -30830 4510 -30770
rect 6300 -30830 6640 -30770
rect 6700 -30830 6710 -30770
rect 8500 -30830 8620 -30770
rect 8680 -30830 8910 -30770
rect 10700 -30830 10820 -30770
rect 10880 -30830 11110 -30770
rect 12900 -30830 13020 -30770
rect 13080 -30830 13310 -30770
rect 15100 -30830 15220 -30770
rect 15280 -30830 15510 -30770
rect 17300 -30830 17640 -30770
rect 17700 -30830 17710 -30770
rect 19500 -30830 19840 -30770
rect 19900 -30830 19910 -30770
rect 2010 -30920 2240 -30860
rect 2300 -30920 2420 -30860
rect 4210 -30940 4440 -30880
rect 4500 -30940 4620 -30880
rect 6410 -30940 6420 -30880
rect 6480 -30940 6820 -30880
rect 8610 -30940 8620 -30880
rect 8680 -30940 9020 -30880
rect 10810 -30940 10820 -30880
rect 10880 -30940 11220 -30880
rect 13010 -30940 13020 -30880
rect 13080 -30940 13420 -30880
rect 15210 -30940 15440 -30880
rect 15500 -30940 15620 -30880
rect 17410 -30940 17640 -30880
rect 17700 -30940 17820 -30880
rect 19610 -30940 20020 -30880
rect -90 -30990 10 -30980
rect -90 -31050 -70 -30990
rect -10 -31050 10 -30990
rect -90 -31060 10 -31050
rect 2110 -30990 2210 -30980
rect 2110 -31050 2130 -30990
rect 2190 -31050 2210 -30990
rect 2110 -31060 2210 -31050
rect 4310 -30990 4410 -30980
rect 4310 -31050 4330 -30990
rect 4390 -31050 4410 -30990
rect 4310 -31060 4410 -31050
rect 6510 -30990 6610 -30980
rect 6510 -31050 6530 -30990
rect 6590 -31050 6610 -30990
rect 6510 -31060 6610 -31050
rect 8710 -30990 8810 -30980
rect 8710 -31050 8730 -30990
rect 8790 -31050 8810 -30990
rect 8710 -31060 8810 -31050
rect 10910 -30990 11010 -30980
rect 10910 -31050 10930 -30990
rect 10990 -31050 11010 -30990
rect 10910 -31060 11010 -31050
rect 13110 -30990 13210 -30980
rect 13110 -31050 13130 -30990
rect 13190 -31050 13210 -30990
rect 13110 -31060 13210 -31050
rect 15310 -30990 15410 -30980
rect 15310 -31050 15330 -30990
rect 15390 -31050 15410 -30990
rect 15310 -31060 15410 -31050
rect 17510 -30990 17610 -30980
rect 17510 -31050 17530 -30990
rect 17590 -31050 17610 -30990
rect 17510 -31060 17610 -31050
rect 19710 -30990 19810 -30980
rect 19710 -31050 19730 -30990
rect 19790 -31050 19810 -30990
rect 19710 -31060 19810 -31050
rect 21910 -30990 22010 -30980
rect 21910 -31050 21930 -30990
rect 21990 -31050 22010 -30990
rect 21910 -31060 22010 -31050
rect 2500 -31300 2700 -31060
rect 2500 -31360 2510 -31300
rect 2690 -31360 2700 -31300
rect 3160 -31300 3360 -31060
rect 3160 -31360 3170 -31300
rect 3350 -31360 3360 -31300
rect 3820 -31300 4020 -31060
rect 3820 -31360 3830 -31300
rect 4010 -31360 4020 -31300
rect 4700 -31300 4900 -31060
rect 4700 -31360 4710 -31300
rect 4890 -31360 4900 -31300
rect 5360 -31300 5560 -31060
rect 5360 -31360 5370 -31300
rect 5550 -31360 5560 -31300
rect 6020 -31300 6220 -31060
rect 6020 -31360 6030 -31300
rect 6210 -31360 6220 -31300
rect 6900 -31160 7100 -31060
rect 6900 -31220 6910 -31160
rect 7090 -31220 7100 -31160
rect 6900 -31360 7100 -31220
rect 7560 -31160 7760 -31060
rect 7560 -31220 7570 -31160
rect 7750 -31220 7760 -31160
rect 7560 -31360 7760 -31220
rect 8220 -31160 8420 -31060
rect 8220 -31220 8230 -31160
rect 8410 -31220 8420 -31160
rect 8220 -31360 8420 -31220
rect 9100 -31160 9300 -31060
rect 9100 -31220 9110 -31160
rect 9290 -31220 9300 -31160
rect 9100 -31360 9300 -31220
rect 9760 -31160 9960 -31060
rect 9760 -31220 9770 -31160
rect 9950 -31220 9960 -31160
rect 9760 -31360 9960 -31220
rect 10420 -31160 10620 -31060
rect 10420 -31220 10430 -31160
rect 10610 -31220 10620 -31160
rect 10420 -31360 10620 -31220
rect 11300 -31160 11500 -31060
rect 11300 -31220 11310 -31160
rect 11490 -31220 11500 -31160
rect 11300 -31360 11500 -31220
rect 11960 -31160 12160 -31060
rect 11960 -31220 11970 -31160
rect 12150 -31220 12160 -31160
rect 11960 -31360 12160 -31220
rect 12620 -31160 12820 -31060
rect 12620 -31220 12630 -31160
rect 12810 -31220 12820 -31160
rect 12620 -31360 12820 -31220
rect 13500 -31160 13700 -31060
rect 13500 -31220 13510 -31160
rect 13690 -31220 13700 -31160
rect 13500 -31360 13700 -31220
rect 14160 -31160 14360 -31060
rect 14160 -31220 14170 -31160
rect 14350 -31220 14360 -31160
rect 14160 -31360 14360 -31220
rect 14820 -31160 15020 -31060
rect 14820 -31220 14830 -31160
rect 15010 -31220 15020 -31160
rect 14820 -31360 15020 -31220
rect 15700 -31300 15900 -31060
rect 15700 -31360 15710 -31300
rect 15890 -31360 15900 -31300
rect 16360 -31300 16560 -31060
rect 16360 -31360 16370 -31300
rect 16550 -31360 16560 -31300
rect 17020 -31300 17220 -31060
rect 17020 -31360 17030 -31300
rect 17210 -31360 17220 -31300
rect 17900 -31300 18100 -31060
rect 17900 -31360 17910 -31300
rect 18090 -31360 18100 -31300
rect 18560 -31300 18760 -31060
rect 18560 -31360 18570 -31300
rect 18750 -31360 18760 -31300
rect 19220 -31300 19420 -31060
rect 19220 -31360 19230 -31300
rect 19410 -31360 19420 -31300
<< via1 >>
rect 2510 11180 2690 11240
rect 3170 11180 3350 11240
rect 3830 11180 4010 11240
rect 4710 11180 4890 11240
rect 5370 11180 5550 11240
rect 6030 11180 6210 11240
rect 6910 11040 7090 11100
rect 7570 11040 7750 11100
rect 8230 11040 8410 11100
rect 9110 11040 9290 11100
rect 9770 11040 9950 11100
rect 10430 11040 10610 11100
rect 11310 11040 11490 11100
rect 11970 11040 12150 11100
rect 12630 11040 12810 11100
rect 13510 11040 13690 11100
rect 14170 11040 14350 11100
rect 14830 11040 15010 11100
rect 15710 11180 15890 11240
rect 16370 11180 16550 11240
rect 17030 11180 17210 11240
rect 17910 11180 18090 11240
rect 18570 11180 18750 11240
rect 19230 11180 19410 11240
rect -70 10870 -10 10930
rect 2130 10870 2190 10930
rect 4330 10870 4390 10930
rect 6530 10870 6590 10930
rect 8730 10870 8790 10930
rect 10930 10870 10990 10930
rect 13130 10870 13190 10930
rect 15330 10870 15390 10930
rect 17530 10870 17590 10930
rect 19730 10870 19790 10930
rect 21930 10870 21990 10930
rect 4220 10760 4280 10820
rect 6420 10760 6480 10820
rect 8840 10760 8900 10820
rect 11040 10760 11100 10820
rect 13240 10760 13300 10820
rect 15440 10760 15500 10820
rect 17420 10760 17480 10820
rect 19620 10740 19680 10800
rect 2020 10650 2080 10710
rect 4220 10650 4280 10710
rect 6640 10650 6700 10710
rect 8840 10650 8900 10710
rect 11040 10650 11100 10710
rect 13240 10650 13300 10710
rect 15220 10650 15280 10710
rect 17420 10650 17480 10710
rect 2510 10550 4010 10610
rect 4710 10550 6210 10610
rect 6910 10550 8410 10610
rect 9110 10550 10610 10610
rect 11310 10550 12810 10610
rect 13510 10550 15010 10610
rect 15710 10550 17210 10610
rect 17910 10550 19410 10610
rect 2510 10240 2690 10300
rect 3170 10240 3350 10300
rect 3830 10240 4010 10300
rect 4710 10240 4890 10300
rect 5370 10240 5550 10300
rect 6030 10240 6210 10300
rect 6910 10380 7090 10440
rect 7570 10380 7750 10440
rect 8230 10380 8410 10440
rect 9110 10380 9290 10440
rect 9770 10380 9950 10440
rect 10430 10380 10610 10440
rect 11310 10380 11490 10440
rect 11970 10380 12150 10440
rect 12630 10380 12810 10440
rect 13510 10380 13690 10440
rect 14170 10380 14350 10440
rect 14830 10380 15010 10440
rect 15710 10240 15890 10300
rect 16370 10240 16550 10300
rect 17030 10240 17210 10300
rect 17910 10240 18090 10300
rect 18570 10240 18750 10300
rect 19230 10240 19410 10300
rect -70 10070 -10 10130
rect 2130 10070 2190 10130
rect 4330 10070 4390 10130
rect 6530 10070 6590 10130
rect 8730 10070 8790 10130
rect 10930 10070 10990 10130
rect 13130 10070 13190 10130
rect 15330 10070 15390 10130
rect 17530 10070 17590 10130
rect 19730 10070 19790 10130
rect 21930 10070 21990 10130
rect 4440 9960 4500 10020
rect 6640 9960 6700 10020
rect 8620 9960 8680 10020
rect 10820 9960 10880 10020
rect 13020 9960 13080 10020
rect 15220 9960 15280 10020
rect 17640 9960 17700 10020
rect 19840 9940 19900 10000
rect 2240 9850 2300 9910
rect 4440 9850 4500 9910
rect 6420 9850 6480 9910
rect 8620 9850 8680 9910
rect 10820 9850 10880 9910
rect 13020 9850 13080 9910
rect 15440 9850 15500 9910
rect 17640 9850 17700 9910
rect 2510 9750 4010 9810
rect 4710 9750 6210 9810
rect 6910 9750 8410 9810
rect 9110 9750 10610 9810
rect 11310 9750 12810 9810
rect 13510 9750 15010 9810
rect 15710 9750 17210 9810
rect 17910 9750 19410 9810
rect 2510 9580 2690 9640
rect 3170 9580 3350 9640
rect 3830 9580 4010 9640
rect 4710 9580 4890 9640
rect 5370 9580 5550 9640
rect 6030 9580 6210 9640
rect 6910 9440 7090 9500
rect 7570 9440 7750 9500
rect 8230 9440 8410 9500
rect 9110 9440 9290 9500
rect 9770 9440 9950 9500
rect 10430 9440 10610 9500
rect 11310 9440 11490 9500
rect 11970 9440 12150 9500
rect 12630 9440 12810 9500
rect 13510 9440 13690 9500
rect 14170 9440 14350 9500
rect 14830 9440 15010 9500
rect 15710 9580 15890 9640
rect 16370 9580 16550 9640
rect 17030 9580 17210 9640
rect 17910 9580 18090 9640
rect 18570 9580 18750 9640
rect 19230 9580 19410 9640
rect -70 9270 -10 9330
rect 2130 9270 2190 9330
rect 4330 9270 4390 9330
rect 6530 9270 6590 9330
rect 8730 9270 8790 9330
rect 10930 9270 10990 9330
rect 13130 9270 13190 9330
rect 15330 9270 15390 9330
rect 17530 9270 17590 9330
rect 19730 9270 19790 9330
rect 21930 9270 21990 9330
rect 6420 9160 6480 9220
rect 8840 9160 8900 9220
rect 11040 9160 11100 9220
rect 13240 9160 13300 9220
rect 15440 9160 15500 9220
rect 17420 9160 17480 9220
rect 4220 9050 4280 9110
rect 6640 9050 6700 9110
rect 8840 9050 8900 9110
rect 11040 9050 11100 9110
rect 13240 9050 13300 9110
rect 15220 9050 15280 9110
rect 430 8910 610 8990
rect 4710 8950 6210 9010
rect 6910 8950 8410 9010
rect 9110 8950 10610 9010
rect 11310 8950 12810 9010
rect 13510 8950 15010 9010
rect 15710 8950 17210 9010
rect 21310 8910 21490 8990
rect 2510 8640 2690 8700
rect 3170 8640 3350 8700
rect 3830 8640 4010 8700
rect 4710 8640 4890 8700
rect 5370 8640 5550 8700
rect 6030 8640 6210 8700
rect 6910 8780 7090 8840
rect 7570 8780 7750 8840
rect 8230 8780 8410 8840
rect 9110 8780 9290 8840
rect 9770 8780 9950 8840
rect 10430 8780 10610 8840
rect 11310 8780 11490 8840
rect 11970 8780 12150 8840
rect 12630 8780 12810 8840
rect 13510 8780 13690 8840
rect 14170 8780 14350 8840
rect 14830 8780 15010 8840
rect 15710 8640 15890 8700
rect 16370 8640 16550 8700
rect 17030 8640 17210 8700
rect 17910 8640 18090 8700
rect 18570 8640 18750 8700
rect 19230 8640 19410 8700
rect -70 8470 -10 8530
rect 2130 8470 2190 8530
rect 4330 8470 4390 8530
rect 6530 8470 6590 8530
rect 8730 8470 8790 8530
rect 10930 8470 10990 8530
rect 13130 8470 13190 8530
rect 15330 8470 15390 8530
rect 17530 8470 17590 8530
rect 19730 8470 19790 8530
rect 21930 8470 21990 8530
rect 6640 8360 6700 8420
rect 8620 8360 8680 8420
rect 10820 8360 10880 8420
rect 13020 8360 13080 8420
rect 15220 8360 15280 8420
rect 17640 8360 17700 8420
rect 4440 8250 4500 8310
rect 6420 8250 6480 8310
rect 8620 8250 8680 8310
rect 10820 8250 10880 8310
rect 13020 8250 13080 8310
rect 15440 8250 15500 8310
rect 430 8110 610 8190
rect 4710 8150 6210 8210
rect 6910 8150 8410 8210
rect 9110 8150 10610 8210
rect 11310 8150 12810 8210
rect 13510 8150 15010 8210
rect 15710 8150 17210 8210
rect 21310 8110 21490 8190
rect 2510 7840 2690 7900
rect 3170 7840 3350 7900
rect 3830 7840 4010 7900
rect 4710 7840 4890 7900
rect 5370 7840 5550 7900
rect 6030 7840 6210 7900
rect 6910 7980 7090 8040
rect 7570 7980 7750 8040
rect 8230 7980 8410 8040
rect 9110 7980 9290 8040
rect 9770 7980 9950 8040
rect 10430 7980 10610 8040
rect 11310 7980 11490 8040
rect 11970 7980 12150 8040
rect 12630 7980 12810 8040
rect 13510 7980 13690 8040
rect 14170 7980 14350 8040
rect 14830 7980 15010 8040
rect 15710 7840 15890 7900
rect 16370 7840 16550 7900
rect 17030 7840 17210 7900
rect 17910 7840 18090 7900
rect 18570 7840 18750 7900
rect 19230 7840 19410 7900
rect -70 7670 -10 7730
rect 2130 7670 2190 7730
rect 4330 7670 4390 7730
rect 6530 7670 6590 7730
rect 8730 7670 8790 7730
rect 10930 7670 10990 7730
rect 13130 7670 13190 7730
rect 15330 7670 15390 7730
rect 17530 7670 17590 7730
rect 19730 7670 19790 7730
rect 21930 7670 21990 7730
rect 6640 7560 6700 7620
rect 8620 7560 8680 7620
rect 10820 7560 10880 7620
rect 13020 7560 13080 7620
rect 15220 7560 15280 7620
rect 17640 7560 17700 7620
rect 4440 7450 4500 7510
rect 6420 7450 6480 7510
rect 8620 7450 8680 7510
rect 10820 7450 10880 7510
rect 13020 7450 13080 7510
rect 15440 7450 15500 7510
rect 430 7310 610 7390
rect 4710 7350 6210 7410
rect 6910 7350 8410 7410
rect 9110 7350 10610 7410
rect 11310 7350 12810 7410
rect 13510 7350 15010 7410
rect 15710 7350 17210 7410
rect 21310 7310 21490 7390
rect 2510 7180 2690 7240
rect 3170 7180 3350 7240
rect 3830 7180 4010 7240
rect 4710 7180 4890 7240
rect 5370 7180 5550 7240
rect 6030 7180 6210 7240
rect 6910 7040 7090 7100
rect 7570 7040 7750 7100
rect 8230 7040 8410 7100
rect 9110 7040 9290 7100
rect 9770 7040 9950 7100
rect 10430 7040 10610 7100
rect 11310 7040 11490 7100
rect 11970 7040 12150 7100
rect 12630 7040 12810 7100
rect 13510 7040 13690 7100
rect 14170 7040 14350 7100
rect 14830 7040 15010 7100
rect 15710 7180 15890 7240
rect 16370 7180 16550 7240
rect 17030 7180 17210 7240
rect 17910 7180 18090 7240
rect 18570 7180 18750 7240
rect 19230 7180 19410 7240
rect -70 6870 -10 6930
rect 2130 6870 2190 6930
rect 4330 6870 4390 6930
rect 6530 6870 6590 6930
rect 8730 6870 8790 6930
rect 10930 6870 10990 6930
rect 13130 6870 13190 6930
rect 15330 6870 15390 6930
rect 17530 6870 17590 6930
rect 19730 6870 19790 6930
rect 21930 6870 21990 6930
rect 6420 6760 6480 6820
rect 8840 6760 8900 6820
rect 11040 6760 11100 6820
rect 13240 6760 13300 6820
rect 15440 6760 15500 6820
rect 17420 6760 17480 6820
rect 4220 6650 4280 6710
rect 6640 6650 6700 6710
rect 8840 6650 8900 6710
rect 11040 6650 11100 6710
rect 13240 6650 13300 6710
rect 15220 6650 15280 6710
rect 430 6510 610 6590
rect 4710 6550 6210 6610
rect 6910 6550 8410 6610
rect 9110 6550 10610 6610
rect 11310 6550 12810 6610
rect 13510 6550 15010 6610
rect 15710 6550 17210 6610
rect 21310 6510 21490 6590
rect 2510 6240 2690 6300
rect 3170 6240 3350 6300
rect 3830 6240 4010 6300
rect 4710 6240 4890 6300
rect 5370 6240 5550 6300
rect 6030 6240 6210 6300
rect 6910 6380 7090 6440
rect 7570 6380 7750 6440
rect 8230 6380 8410 6440
rect 9110 6380 9290 6440
rect 9770 6380 9950 6440
rect 10430 6380 10610 6440
rect 11310 6380 11490 6440
rect 11970 6380 12150 6440
rect 12630 6380 12810 6440
rect 13510 6380 13690 6440
rect 14170 6380 14350 6440
rect 14830 6380 15010 6440
rect 15710 6240 15890 6300
rect 16370 6240 16550 6300
rect 17030 6240 17210 6300
rect 17910 6240 18090 6300
rect 18570 6240 18750 6300
rect 19230 6240 19410 6300
rect -70 6070 -10 6130
rect 2130 6070 2190 6130
rect 4330 6070 4390 6130
rect 6530 6070 6590 6130
rect 8730 6070 8790 6130
rect 10930 6070 10990 6130
rect 13130 6070 13190 6130
rect 15330 6070 15390 6130
rect 17530 6070 17590 6130
rect 19730 6070 19790 6130
rect 21930 6070 21990 6130
rect 4440 5960 4500 6020
rect 6640 5960 6700 6020
rect 8620 5960 8680 6020
rect 10820 5960 10880 6020
rect 13020 5960 13080 6020
rect 15220 5960 15280 6020
rect 17640 5960 17700 6020
rect 19840 5940 19900 6000
rect 2240 5850 2300 5910
rect 4440 5850 4500 5910
rect 6420 5850 6480 5910
rect 8620 5850 8680 5910
rect 10820 5850 10880 5910
rect 13020 5850 13080 5910
rect 15440 5850 15500 5910
rect 17640 5850 17700 5910
rect 2510 5750 4010 5810
rect 4710 5750 6210 5810
rect 6910 5750 8410 5810
rect 9110 5750 10610 5810
rect 11310 5750 12810 5810
rect 13510 5750 15010 5810
rect 15710 5750 17210 5810
rect 17910 5750 19410 5810
rect 2510 5580 2690 5640
rect 3170 5580 3350 5640
rect 3830 5580 4010 5640
rect 4710 5580 4890 5640
rect 5370 5580 5550 5640
rect 6030 5580 6210 5640
rect 6910 5440 7090 5500
rect 7570 5440 7750 5500
rect 8230 5440 8410 5500
rect 9110 5440 9290 5500
rect 9770 5440 9950 5500
rect 10430 5440 10610 5500
rect 11310 5440 11490 5500
rect 11970 5440 12150 5500
rect 12630 5440 12810 5500
rect 13510 5440 13690 5500
rect 14170 5440 14350 5500
rect 14830 5440 15010 5500
rect 15710 5580 15890 5640
rect 16370 5580 16550 5640
rect 17030 5580 17210 5640
rect 17910 5580 18090 5640
rect 18570 5580 18750 5640
rect 19230 5580 19410 5640
rect -70 5270 -10 5330
rect 2130 5270 2190 5330
rect 4330 5270 4390 5330
rect 6530 5270 6590 5330
rect 8730 5270 8790 5330
rect 10930 5270 10990 5330
rect 13130 5270 13190 5330
rect 15330 5270 15390 5330
rect 17530 5270 17590 5330
rect 19730 5270 19790 5330
rect 21930 5270 21990 5330
rect 4220 5160 4280 5220
rect 6420 5160 6480 5220
rect 8840 5160 8900 5220
rect 11040 5160 11100 5220
rect 13240 5160 13300 5220
rect 15440 5160 15500 5220
rect 17420 5160 17480 5220
rect 19620 5140 19680 5200
rect 2020 5050 2080 5110
rect 4220 5050 4280 5110
rect 6640 5050 6700 5110
rect 8840 5050 8900 5110
rect 11040 5050 11100 5110
rect 13240 5050 13300 5110
rect 15220 5050 15280 5110
rect 17420 5050 17480 5110
rect 2510 4950 4010 5010
rect 4710 4950 6210 5010
rect 6910 4950 8410 5010
rect 9110 4950 10610 5010
rect 11310 4950 12810 5010
rect 13510 4950 15010 5010
rect 15710 4950 17210 5010
rect 17910 4950 19410 5010
rect 2110 1290 2230 1970
rect 3710 1290 3830 1970
rect 5310 1290 5430 1970
rect 6910 1290 7030 1970
rect 8510 1290 8630 1970
rect 10110 1290 10230 1970
rect 11030 1310 11150 1930
rect 12610 1310 12730 1930
rect 13990 1310 14110 1930
rect 14910 1300 15030 1960
rect 16510 1290 16630 1970
rect 18110 1290 18230 1970
rect 19710 1290 19830 1970
rect 21310 1290 21430 1970
rect 22910 1290 23030 1970
rect 24510 1290 24630 1970
rect 26110 1290 26230 1970
rect 27710 1290 27830 1970
rect 29310 1290 29430 1970
rect 30910 1290 31030 1970
rect 32510 1290 32630 1970
rect 34110 1290 34230 1970
rect 35710 1290 35830 1970
rect 1410 1010 1530 1130
rect 3010 1010 3130 1130
rect 4610 1010 4730 1130
rect 6210 1010 6330 1130
rect 7810 1010 7930 1130
rect 9410 1010 9530 1130
rect 11250 1050 11670 1210
rect 15600 1010 15700 1130
rect 17200 1010 17300 1130
rect 18800 1010 18900 1130
rect 20400 1010 20500 1130
rect 22000 1010 22100 1130
rect 23600 1010 23700 1130
rect 26800 1010 26900 1130
rect 28400 1010 28500 1130
rect 12390 750 12510 870
rect 1190 560 1310 680
rect 2790 560 2910 680
rect 4390 560 4510 680
rect 5990 560 6110 680
rect 7590 560 7710 680
rect 9190 560 9310 680
rect 15820 560 15920 680
rect 17420 560 17520 680
rect 19020 560 19120 680
rect 20620 560 20720 680
rect 22220 560 22320 680
rect 23820 560 23920 680
rect 27020 560 27120 680
rect 28620 560 28720 680
rect 31820 560 31920 680
rect 2110 -510 2230 170
rect 3710 -510 3830 170
rect 5310 -510 5430 170
rect 6910 -510 7030 170
rect 8510 -510 8630 170
rect 10110 -510 10230 170
rect 11710 -590 11830 170
rect 13310 -510 13430 170
rect 1410 -790 1530 -670
rect 3010 -790 3130 -670
rect 4610 -790 4730 -670
rect 6210 -790 6330 -670
rect 7810 -790 7930 -670
rect 9410 -790 9530 -670
rect 11270 -750 12270 -590
rect 14910 -590 15030 170
rect 16510 -510 16630 170
rect 18110 -510 18230 170
rect 19710 -510 19830 170
rect 21310 -510 21430 170
rect 22910 -510 23030 170
rect 24510 -510 24630 170
rect 26110 -510 26230 170
rect 27710 -510 27830 170
rect 29310 -510 29430 170
rect 30910 -510 31030 170
rect 32510 -510 32630 170
rect 34110 -510 34230 170
rect 35710 -510 35830 170
rect 12390 -1050 12510 -670
rect 14470 -750 15470 -590
rect 15600 -790 15700 -670
rect 17200 -790 17300 -670
rect 18800 -790 18900 -670
rect 20400 -790 20500 -670
rect 22000 -790 22100 -670
rect 23600 -790 23700 -670
rect 26800 -790 26900 -670
rect 28400 -790 28500 -670
rect 12630 -1070 12750 -930
rect 13970 -1070 14090 -930
rect 1190 -1240 1310 -1120
rect 2790 -1240 2910 -1120
rect 4390 -1240 4510 -1120
rect 5990 -1240 6110 -1120
rect 7590 -1240 7710 -1120
rect 9190 -1240 9310 -1120
rect 10810 -1270 10990 -1210
rect 15820 -1240 15920 -1120
rect 17420 -1240 17520 -1120
rect 19020 -1240 19120 -1120
rect 20620 -1240 20720 -1120
rect 22220 -1240 22320 -1120
rect 23820 -1240 23920 -1120
rect 27020 -1240 27120 -1120
rect 28620 -1240 28720 -1120
rect 31600 -1240 31700 -1120
rect 2110 -2310 2230 -1630
rect 3710 -2310 3830 -1630
rect 5310 -2310 5430 -1630
rect 6910 -2310 7030 -1630
rect 8510 -2310 8630 -1630
rect 10110 -2310 10230 -1630
rect 11710 -2310 11830 -1630
rect 13310 -2310 13430 -1630
rect 14910 -2310 15030 -1630
rect 16510 -2310 16630 -1630
rect 18110 -2310 18230 -1630
rect 19710 -2310 19830 -1630
rect 21310 -2310 21430 -1630
rect 22910 -2310 23030 -1630
rect 24510 -2310 24630 -1630
rect 26110 -2310 26230 -1630
rect 27710 -2310 27830 -1630
rect 29310 -2310 29430 -1630
rect 30910 -2310 31030 -1630
rect 32510 -2310 32630 -1630
rect 34110 -2310 34230 -1630
rect 35710 -2310 35830 -1630
rect 1410 -2590 1530 -2470
rect 3010 -2590 3130 -2470
rect 4610 -2590 4730 -2470
rect 6210 -2590 6330 -2470
rect 7810 -2590 7930 -2470
rect 9410 -2590 9530 -2470
rect 15600 -2590 15700 -2470
rect 17200 -2590 17300 -2470
rect 18800 -2590 18900 -2470
rect 20400 -2590 20500 -2470
rect 22000 -2590 22100 -2470
rect 23600 -2590 23700 -2470
rect 25200 -2590 25300 -2470
rect 26800 -2590 26900 -2470
rect 28400 -2590 28500 -2470
rect 30000 -2590 30100 -2470
rect 12390 -2850 12510 -2730
rect 1190 -3040 1310 -2920
rect 2790 -3040 2910 -2920
rect 4390 -3040 4510 -2920
rect 5990 -3040 6110 -2920
rect 7590 -3040 7710 -2920
rect 9190 -3040 9310 -2920
rect 11010 -3040 11130 -2920
rect 14210 -3040 14330 -2920
rect 14430 -3040 14550 -2920
rect 15820 -3040 15920 -2920
rect 17420 -3040 17520 -2920
rect 19020 -3040 19120 -2920
rect 20620 -3040 20720 -2920
rect 22220 -3040 22320 -2920
rect 23820 -3040 23920 -2920
rect 25420 -3040 25520 -2920
rect 27020 -3040 27120 -2920
rect 28620 -3040 28720 -2920
rect 30220 -3040 30320 -2920
rect 36400 -3030 36500 -2910
rect 12610 -3410 12730 -3310
rect 2110 -4110 2230 -3430
rect 3710 -4110 3830 -3430
rect 5310 -4110 5430 -3430
rect 6910 -4110 7030 -3430
rect 8510 -4110 8630 -3430
rect 10110 -4110 10230 -3430
rect 11710 -4110 11830 -3430
rect 13310 -4110 13430 -3430
rect 14210 -3430 14330 -3310
rect 14910 -4110 15030 -3430
rect 16510 -4110 16630 -3430
rect 18110 -4110 18230 -3430
rect 19710 -4110 19830 -3430
rect 21310 -4110 21430 -3430
rect 22910 -4110 23030 -3430
rect 24510 -4110 24630 -3430
rect 26110 -4110 26230 -3430
rect 27710 -4110 27830 -3430
rect 29310 -4110 29430 -3430
rect 30910 -4110 31030 -3430
rect 32510 -4110 32630 -3430
rect 34110 -4110 34230 -3430
rect 35710 -4110 35830 -3430
rect 1410 -4390 1530 -4270
rect 3010 -4390 3130 -4270
rect 4610 -4390 4730 -4270
rect 6210 -4390 6330 -4270
rect 7810 -4390 7930 -4270
rect 9410 -4390 9530 -4270
rect 15600 -4390 15700 -4270
rect 17200 -4390 17300 -4270
rect 18800 -4390 18900 -4270
rect 20400 -4390 20500 -4270
rect 22000 -4390 22100 -4270
rect 23600 -4390 23700 -4270
rect 25200 -4390 25300 -4270
rect 26800 -4390 26900 -4270
rect 28400 -4390 28500 -4270
rect 30000 -4390 30100 -4270
rect 12390 -4650 12510 -4530
rect 1190 -4840 1310 -4720
rect 2790 -4840 2910 -4720
rect 4390 -4840 4510 -4720
rect 5990 -4840 6110 -4720
rect 7590 -4840 7710 -4720
rect 9190 -4840 9310 -4720
rect 11710 -4930 11830 -4810
rect 12610 -4850 12730 -4730
rect 13630 -4910 13750 -4790
rect 14210 -4850 14330 -4730
rect 15230 -4910 15350 -4790
rect 15820 -4840 15920 -4720
rect 17420 -4840 17520 -4720
rect 19020 -4840 19120 -4720
rect 20620 -4840 20720 -4720
rect 22220 -4840 22320 -4720
rect 23820 -4840 23920 -4720
rect 25420 -4840 25520 -4720
rect 27020 -4840 27120 -4720
rect 28620 -4840 28720 -4720
rect 30220 -4840 30320 -4720
rect 36400 -4830 36500 -4710
rect 11710 -5950 11830 -5830
rect 13310 -5950 13430 -5830
rect 11710 -6170 11830 -6050
rect 13630 -6170 13750 -6050
rect 14230 -6170 14350 -6050
rect 15230 -6170 15350 -6050
rect 12630 -6390 12750 -6270
rect 16510 -6390 16630 -6270
rect 12410 -6610 12530 -6490
rect 14910 -6610 15030 -6490
rect 1210 -8190 1330 -8070
rect 2810 -8190 2930 -8070
rect 4410 -8190 4530 -8070
rect 6010 -8190 6130 -8070
rect 7610 -8190 7730 -8070
rect 9210 -8190 9330 -8070
rect 11710 -8230 11840 -8110
rect 15830 -8190 15950 -8070
rect 17430 -8190 17550 -8070
rect 19030 -8190 19150 -8070
rect 20630 -8190 20750 -8070
rect 22230 -8190 22350 -8070
rect 23830 -8190 23950 -8070
rect 25430 -8190 25550 -8070
rect 27030 -8190 27150 -8070
rect 28630 -8190 28750 -8070
rect 30230 -8190 30350 -8070
rect 1430 -8630 1550 -8510
rect 3030 -8630 3150 -8510
rect 4630 -8630 4750 -8510
rect 6230 -8630 6350 -8510
rect 7830 -8630 7950 -8510
rect 9430 -8630 9550 -8510
rect 2130 -9470 2230 -8810
rect 3730 -9470 3830 -8810
rect 5330 -9470 5430 -8810
rect 6930 -9470 7030 -8810
rect 8530 -9470 8630 -8810
rect 10130 -9470 10230 -8810
rect 11720 -9470 11830 -8810
rect 15610 -8640 15730 -8520
rect 17210 -8640 17330 -8520
rect 18810 -8640 18930 -8520
rect 20410 -8640 20530 -8520
rect 22010 -8640 22130 -8520
rect 23610 -8640 23730 -8520
rect 25210 -8640 25330 -8520
rect 26810 -8640 26930 -8520
rect 28410 -8640 28530 -8520
rect 30010 -8640 30130 -8520
rect 13320 -9470 13430 -8810
rect 14920 -9470 15030 -8810
rect 16520 -9480 16630 -8800
rect 18120 -9480 18230 -8800
rect 19720 -9480 19830 -8800
rect 21320 -9480 21430 -8800
rect 22920 -9480 23030 -8800
rect 24520 -9480 24630 -8800
rect 26120 -9480 26230 -8800
rect 27720 -9480 27830 -8800
rect 29320 -9480 29430 -8800
rect 30920 -9480 31030 -8800
rect 1210 -9990 1330 -9870
rect 2810 -9990 2930 -9870
rect 4410 -9990 4530 -9870
rect 6010 -9990 6130 -9870
rect 7610 -9990 7730 -9870
rect 9210 -9990 9330 -9870
rect 15830 -9990 15950 -9870
rect 17430 -9990 17550 -9870
rect 19030 -9990 19150 -9870
rect 20630 -9990 20750 -9870
rect 22230 -9990 22350 -9870
rect 23830 -9990 23950 -9870
rect 25430 -9990 25550 -9870
rect 27030 -9990 27150 -9870
rect 28630 -9990 28750 -9870
rect 30230 -9990 30350 -9870
rect 1430 -10430 1550 -10310
rect 3030 -10430 3150 -10310
rect 4630 -10430 4750 -10310
rect 6230 -10430 6350 -10310
rect 7830 -10430 7950 -10310
rect 9430 -10430 9550 -10310
rect 11030 -10530 11150 -10410
rect 15610 -10440 15730 -10320
rect 17210 -10440 17330 -10320
rect 18810 -10440 18930 -10320
rect 20410 -10440 20530 -10320
rect 22010 -10440 22130 -10320
rect 23610 -10440 23730 -10320
rect 25210 -10440 25330 -10320
rect 26810 -10440 26930 -10320
rect 28410 -10440 28530 -10320
rect 30010 -10440 30130 -10320
rect 2130 -11270 2230 -10610
rect 3730 -11270 3830 -10610
rect 5330 -11270 5430 -10610
rect 6930 -11270 7030 -10610
rect 8530 -11270 8630 -10610
rect 10130 -11270 10230 -10610
rect 11720 -11270 11830 -10610
rect 13320 -11270 13430 -10610
rect 14920 -11270 15030 -10610
rect 16520 -11280 16630 -10600
rect 18120 -11280 18230 -10600
rect 19720 -11280 19830 -10600
rect 21320 -11280 21430 -10600
rect 22920 -11280 23030 -10600
rect 24520 -11280 24630 -10600
rect 26120 -11280 26230 -10600
rect 27720 -11280 27830 -10600
rect 29320 -11280 29430 -10600
rect 30920 -11280 31030 -10600
rect 1210 -11790 1330 -11670
rect 2810 -11790 2930 -11670
rect 4410 -11790 4530 -11670
rect 6010 -11790 6130 -11670
rect 7610 -11790 7730 -11670
rect 9210 -11790 9330 -11670
rect 13310 -11790 13430 -11670
rect 14230 -11790 14350 -11670
rect 14910 -11790 15030 -11670
rect 15830 -11790 15950 -11670
rect 17430 -11790 17550 -11670
rect 19030 -11790 19150 -11670
rect 20630 -11790 20750 -11670
rect 22230 -11790 22350 -11670
rect 23830 -11790 23950 -11670
rect 25430 -11790 25550 -11670
rect 27030 -11790 27150 -11670
rect 28630 -11790 28750 -11670
rect 30230 -11790 30350 -11670
rect 1430 -12230 1550 -12110
rect 3030 -12230 3150 -12110
rect 4630 -12230 4750 -12110
rect 6230 -12230 6350 -12110
rect 7830 -12230 7950 -12110
rect 9430 -12230 9550 -12110
rect 10810 -12330 10930 -12220
rect 15610 -12240 15730 -12120
rect 17210 -12240 17330 -12120
rect 18810 -12240 18930 -12120
rect 20410 -12240 20530 -12120
rect 22010 -12240 22130 -12120
rect 23610 -12240 23730 -12120
rect 25210 -12240 25330 -12120
rect 26810 -12240 26930 -12120
rect 28410 -12240 28530 -12120
rect 30010 -12240 30130 -12120
rect 2130 -13070 2230 -12410
rect 3730 -13070 3830 -12410
rect 5330 -13070 5430 -12410
rect 6930 -13070 7030 -12410
rect 8530 -13070 8630 -12410
rect 10130 -13070 10230 -12410
rect 11720 -13070 11830 -12410
rect 13320 -13070 13430 -12410
rect 14920 -13070 15030 -12410
rect 16520 -13080 16630 -12400
rect 18120 -13080 18230 -12400
rect 19720 -13080 19830 -12400
rect 21320 -13080 21430 -12400
rect 22920 -13080 23030 -12400
rect 24520 -13080 24630 -12400
rect 26120 -13080 26230 -12400
rect 27720 -13080 27830 -12400
rect 29320 -13080 29430 -12400
rect 30920 -13080 31030 -12400
rect 11270 -13210 11650 -13150
rect 1210 -13590 1330 -13470
rect 2810 -13590 2930 -13470
rect 4410 -13590 4530 -13470
rect 6010 -13590 6130 -13470
rect 7610 -13590 7730 -13470
rect 9210 -13590 9330 -13470
rect 14010 -13600 14130 -13480
rect 15830 -13590 15950 -13470
rect 17430 -13590 17550 -13470
rect 19030 -13590 19150 -13470
rect 20630 -13590 20750 -13470
rect 22230 -13590 22350 -13470
rect 23830 -13590 23950 -13470
rect 25430 -13590 25550 -13470
rect 27030 -13590 27150 -13470
rect 28630 -13590 28750 -13470
rect 30230 -13590 30350 -13470
rect 1430 -14030 1550 -13910
rect 3030 -14030 3150 -13910
rect 4630 -14030 4750 -13910
rect 6230 -14030 6350 -13910
rect 7830 -14030 7950 -13910
rect 9430 -14030 9550 -13910
rect 11270 -14120 11650 -14060
rect 15610 -14040 15730 -13920
rect 17210 -14040 17330 -13920
rect 18810 -14040 18930 -13920
rect 20410 -14040 20530 -13920
rect 22010 -14040 22130 -13920
rect 23610 -14040 23730 -13920
rect 25210 -14040 25330 -13920
rect 26810 -14040 26930 -13920
rect 28410 -14040 28530 -13920
rect 30010 -14040 30130 -13920
rect 2130 -14870 2230 -14210
rect 3730 -14870 3830 -14210
rect 5330 -14870 5430 -14210
rect 6930 -14870 7030 -14210
rect 8530 -14870 8630 -14210
rect 10130 -14870 10230 -14210
rect 11720 -14870 11830 -14210
rect 13320 -14870 13430 -14210
rect 14920 -14870 15030 -14210
rect 16520 -14880 16630 -14200
rect 18120 -14880 18230 -14200
rect 19720 -14880 19830 -14200
rect 21320 -14880 21430 -14200
rect 22920 -14880 23030 -14200
rect 24520 -14880 24630 -14200
rect 26120 -14880 26230 -14200
rect 27720 -14880 27830 -14200
rect 29320 -14880 29430 -14200
rect 30920 -14880 31030 -14200
rect 1210 -15390 1330 -15270
rect 2810 -15390 2930 -15270
rect 4410 -15390 4530 -15270
rect 6010 -15390 6130 -15270
rect 7610 -15390 7730 -15270
rect 9210 -15390 9330 -15270
rect 13330 -15390 13430 -15290
rect 14020 -15410 14120 -15310
rect 14930 -15390 15030 -15290
rect 15830 -15390 15950 -15270
rect 17430 -15390 17550 -15270
rect 19030 -15390 19150 -15270
rect 20630 -15390 20750 -15270
rect 22230 -15390 22350 -15270
rect 23830 -15390 23950 -15270
rect 27030 -15390 27150 -15270
rect 28630 -15390 28750 -15270
rect 1430 -15830 1550 -15710
rect 3030 -15830 3150 -15710
rect 4630 -15830 4750 -15710
rect 6230 -15830 6350 -15710
rect 7830 -15830 7950 -15710
rect 9430 -15830 9550 -15710
rect 15610 -15840 15730 -15720
rect 17210 -15840 17330 -15720
rect 18810 -15840 18930 -15720
rect 20410 -15840 20530 -15720
rect 22010 -15840 22130 -15720
rect 23610 -15840 23730 -15720
rect 26810 -15840 26930 -15720
rect 28410 -15840 28530 -15720
rect 2130 -16670 2230 -16010
rect 3730 -16670 3830 -16010
rect 5330 -16670 5430 -16010
rect 6930 -16670 7030 -16010
rect 8530 -16670 8630 -16010
rect 10130 -16670 10230 -16010
rect 11720 -16670 11830 -16010
rect 13320 -16670 13430 -16010
rect 14920 -16670 15030 -16010
rect 16520 -16680 16630 -16000
rect 18120 -16680 18230 -16000
rect 19720 -16680 19830 -16000
rect 21320 -16680 21430 -16000
rect 22920 -16680 23030 -16000
rect 24520 -16680 24630 -16000
rect 26120 -16680 26230 -16000
rect 27720 -16680 27830 -16000
rect 29320 -16680 29430 -16000
rect 30920 -16680 31030 -16000
rect 1210 -17190 1330 -17070
rect 2810 -17190 2930 -17070
rect 4410 -17190 4530 -17070
rect 6010 -17190 6130 -17070
rect 7610 -17190 7730 -17070
rect 9210 -17190 9330 -17070
rect 12630 -17200 12750 -17080
rect 15830 -17190 15950 -17070
rect 17430 -17190 17550 -17070
rect 19030 -17190 19150 -17070
rect 20630 -17190 20750 -17070
rect 22230 -17190 22350 -17070
rect 23830 -17190 23950 -17070
rect 27030 -17190 27150 -17070
rect 28630 -17190 28750 -17070
rect 1430 -17630 1550 -17510
rect 3030 -17630 3150 -17510
rect 4630 -17630 4750 -17510
rect 6230 -17630 6350 -17510
rect 7830 -17630 7950 -17510
rect 9430 -17630 9550 -17510
rect 15610 -17640 15730 -17520
rect 17210 -17640 17330 -17520
rect 18810 -17640 18930 -17520
rect 20410 -17640 20530 -17520
rect 22010 -17640 22130 -17520
rect 23610 -17640 23730 -17520
rect 26810 -17640 26930 -17520
rect 28410 -17640 28530 -17520
rect 2130 -18470 2230 -17810
rect 3730 -18470 3830 -17810
rect 5330 -18470 5430 -17810
rect 6930 -18470 7030 -17810
rect 8530 -18470 8630 -17810
rect 10130 -18470 10230 -17810
rect 11720 -18470 11830 -17810
rect 13320 -18470 13430 -17810
rect 14920 -18470 15030 -17810
rect 16520 -18480 16630 -17800
rect 18120 -18480 18230 -17800
rect 19720 -18480 19830 -17800
rect 21320 -18480 21430 -17800
rect 22920 -18480 23030 -17800
rect 24520 -18480 24630 -17800
rect 26120 -18480 26230 -17800
rect 27720 -18480 27830 -17800
rect 29320 -18480 29430 -17800
rect 30920 -18480 31030 -17800
rect 1210 -18990 1330 -18870
rect 2810 -18990 2930 -18870
rect 4410 -18990 4530 -18870
rect 6010 -18990 6130 -18870
rect 7610 -18990 7730 -18870
rect 9210 -18990 9330 -18870
rect 12410 -19000 12530 -18880
rect 15830 -18990 15950 -18870
rect 17430 -18990 17550 -18870
rect 19030 -18990 19150 -18870
rect 20630 -18990 20750 -18870
rect 22230 -18990 22350 -18870
rect 23830 -18990 23950 -18870
rect 27030 -18990 27150 -18870
rect 28630 -18990 28750 -18870
rect 1430 -19430 1550 -19310
rect 3030 -19430 3150 -19310
rect 4630 -19430 4750 -19310
rect 6230 -19430 6350 -19310
rect 7830 -19430 7950 -19310
rect 9430 -19430 9550 -19310
rect 15610 -19440 15730 -19320
rect 17210 -19440 17330 -19320
rect 18810 -19440 18930 -19320
rect 20410 -19440 20530 -19320
rect 22010 -19440 22130 -19320
rect 23610 -19440 23730 -19320
rect 26810 -19440 26930 -19320
rect 28410 -19440 28530 -19320
rect 2130 -20270 2230 -19610
rect 3730 -20270 3830 -19610
rect 5330 -20270 5430 -19610
rect 6930 -20270 7030 -19610
rect 8530 -20270 8630 -19610
rect 10130 -20270 10230 -19610
rect 11720 -20270 11830 -19610
rect 13320 -20270 13430 -19610
rect 14920 -20270 15030 -19610
rect 16520 -20280 16630 -19600
rect 18120 -20280 18230 -19600
rect 19720 -20280 19830 -19600
rect 21320 -20280 21430 -19600
rect 22920 -20280 23030 -19600
rect 24520 -20280 24630 -19600
rect 26120 -20280 26230 -19600
rect 27720 -20280 27830 -19600
rect 29320 -20280 29430 -19600
rect 30920 -20280 31030 -19600
rect 1210 -20790 1330 -20670
rect 2810 -20790 2930 -20670
rect 4410 -20790 4530 -20670
rect 6010 -20790 6130 -20670
rect 7610 -20790 7730 -20670
rect 9210 -20790 9330 -20670
rect 15830 -20790 15950 -20670
rect 17430 -20790 17550 -20670
rect 19030 -20790 19150 -20670
rect 20630 -20790 20750 -20670
rect 22230 -20790 22350 -20670
rect 23830 -20790 23950 -20670
rect 27030 -20790 27150 -20670
rect 28630 -20790 28750 -20670
rect 1430 -21230 1550 -21110
rect 3030 -21230 3150 -21110
rect 4630 -21230 4750 -21110
rect 6230 -21230 6350 -21110
rect 7830 -21230 7950 -21110
rect 9430 -21230 9550 -21110
rect 15610 -21240 15730 -21120
rect 17210 -21240 17330 -21120
rect 18810 -21240 18930 -21120
rect 20410 -21240 20530 -21120
rect 22010 -21240 22130 -21120
rect 23610 -21240 23730 -21120
rect 26810 -21240 26930 -21120
rect 28410 -21240 28530 -21120
rect 2130 -22070 2230 -21410
rect 3730 -22070 3830 -21410
rect 5330 -22070 5430 -21410
rect 6930 -22070 7030 -21410
rect 8530 -22070 8630 -21410
rect 10130 -22070 10230 -21410
rect 16520 -22080 16630 -21400
rect 18120 -22080 18230 -21400
rect 19720 -22080 19830 -21400
rect 21320 -22080 21430 -21400
rect 22920 -22080 23030 -21400
rect 24520 -22080 24630 -21400
rect 26120 -22080 26230 -21400
rect 27720 -22080 27830 -21400
rect 29320 -22080 29430 -21400
rect 30920 -22080 31030 -21400
rect 2510 -25130 4010 -25070
rect 4710 -25130 6210 -25070
rect 6910 -25130 8410 -25070
rect 9110 -25130 10610 -25070
rect 11310 -25130 12810 -25070
rect 13510 -25130 15010 -25070
rect 15710 -25130 17210 -25070
rect 17910 -25130 19410 -25070
rect 4440 -25230 4500 -25170
rect 6640 -25230 6700 -25170
rect 8620 -25230 8680 -25170
rect 10820 -25230 10880 -25170
rect 13020 -25230 13080 -25170
rect 15220 -25230 15280 -25170
rect 17640 -25230 17700 -25170
rect 19840 -25230 19900 -25170
rect 2240 -25320 2300 -25260
rect 4440 -25340 4500 -25280
rect 6420 -25340 6480 -25280
rect 8620 -25340 8680 -25280
rect 10820 -25340 10880 -25280
rect 13020 -25340 13080 -25280
rect 15440 -25340 15500 -25280
rect 17640 -25340 17700 -25280
rect -70 -25450 -10 -25390
rect 2130 -25450 2190 -25390
rect 4330 -25450 4390 -25390
rect 6530 -25450 6590 -25390
rect 8730 -25450 8790 -25390
rect 10930 -25450 10990 -25390
rect 13130 -25450 13190 -25390
rect 15330 -25450 15390 -25390
rect 17530 -25450 17590 -25390
rect 19730 -25450 19790 -25390
rect 21930 -25450 21990 -25390
rect 2510 -25760 2690 -25700
rect 3170 -25760 3350 -25700
rect 3830 -25760 4010 -25700
rect 4710 -25760 4890 -25700
rect 5370 -25760 5550 -25700
rect 6030 -25760 6210 -25700
rect 6910 -25620 7090 -25560
rect 7570 -25620 7750 -25560
rect 8230 -25620 8410 -25560
rect 9110 -25620 9290 -25560
rect 9770 -25620 9950 -25560
rect 10430 -25620 10610 -25560
rect 11310 -25620 11490 -25560
rect 11970 -25620 12150 -25560
rect 12630 -25620 12810 -25560
rect 13510 -25620 13690 -25560
rect 14170 -25620 14350 -25560
rect 14830 -25620 15010 -25560
rect 15710 -25760 15890 -25700
rect 16370 -25760 16550 -25700
rect 17030 -25760 17210 -25700
rect 17910 -25760 18090 -25700
rect 18570 -25760 18750 -25700
rect 19230 -25760 19410 -25700
rect 2510 -25930 4010 -25870
rect 4710 -25930 6210 -25870
rect 6910 -25930 8410 -25870
rect 9110 -25930 10610 -25870
rect 11310 -25930 12810 -25870
rect 13510 -25930 15010 -25870
rect 15710 -25930 17210 -25870
rect 17910 -25930 19410 -25870
rect 4220 -26030 4280 -25970
rect 6420 -26030 6480 -25970
rect 8840 -26030 8900 -25970
rect 11040 -26030 11100 -25970
rect 13240 -26030 13300 -25970
rect 15440 -26030 15500 -25970
rect 17420 -26030 17480 -25970
rect 19620 -26030 19680 -25970
rect 2020 -26120 2080 -26060
rect 4220 -26140 4280 -26080
rect 6640 -26140 6700 -26080
rect 8840 -26140 8900 -26080
rect 11040 -26140 11100 -26080
rect 13240 -26140 13300 -26080
rect 15220 -26140 15280 -26080
rect 17420 -26140 17480 -26080
rect -70 -26250 -10 -26190
rect 2130 -26250 2190 -26190
rect 4330 -26250 4390 -26190
rect 6530 -26250 6590 -26190
rect 8730 -26250 8790 -26190
rect 10930 -26250 10990 -26190
rect 13130 -26250 13190 -26190
rect 15330 -26250 15390 -26190
rect 17530 -26250 17590 -26190
rect 19730 -26250 19790 -26190
rect 21930 -26250 21990 -26190
rect 2510 -26420 2690 -26360
rect 3170 -26420 3350 -26360
rect 3830 -26420 4010 -26360
rect 4710 -26420 4890 -26360
rect 5370 -26420 5550 -26360
rect 6030 -26420 6210 -26360
rect 6910 -26560 7090 -26500
rect 7570 -26560 7750 -26500
rect 8230 -26560 8410 -26500
rect 9110 -26560 9290 -26500
rect 9770 -26560 9950 -26500
rect 10430 -26560 10610 -26500
rect 11310 -26560 11490 -26500
rect 11970 -26560 12150 -26500
rect 12630 -26560 12810 -26500
rect 13510 -26560 13690 -26500
rect 14170 -26560 14350 -26500
rect 14830 -26560 15010 -26500
rect 15710 -26420 15890 -26360
rect 16370 -26420 16550 -26360
rect 17030 -26420 17210 -26360
rect 17910 -26420 18090 -26360
rect 18570 -26420 18750 -26360
rect 19230 -26420 19410 -26360
rect 430 -26710 610 -26630
rect 4710 -26730 6210 -26670
rect 6910 -26730 8410 -26670
rect 9110 -26730 10610 -26670
rect 11310 -26730 12810 -26670
rect 13510 -26730 15010 -26670
rect 15710 -26730 17210 -26670
rect 21310 -26710 21490 -26630
rect 6640 -26830 6700 -26770
rect 8620 -26830 8680 -26770
rect 10820 -26830 10880 -26770
rect 13020 -26830 13080 -26770
rect 15220 -26830 15280 -26770
rect 17640 -26830 17700 -26770
rect 4440 -26940 4500 -26880
rect 6420 -26940 6480 -26880
rect 8620 -26940 8680 -26880
rect 10820 -26940 10880 -26880
rect 13020 -26940 13080 -26880
rect 15440 -26940 15500 -26880
rect -70 -27050 -10 -26990
rect 2130 -27050 2190 -26990
rect 4330 -27050 4390 -26990
rect 6530 -27050 6590 -26990
rect 8730 -27050 8790 -26990
rect 10930 -27050 10990 -26990
rect 13130 -27050 13190 -26990
rect 15330 -27050 15390 -26990
rect 17530 -27050 17590 -26990
rect 19730 -27050 19790 -26990
rect 21930 -27050 21990 -26990
rect 2510 -27360 2690 -27300
rect 3170 -27360 3350 -27300
rect 3830 -27360 4010 -27300
rect 4710 -27360 4890 -27300
rect 5370 -27360 5550 -27300
rect 6030 -27360 6210 -27300
rect 6910 -27220 7090 -27160
rect 7570 -27220 7750 -27160
rect 8230 -27220 8410 -27160
rect 9110 -27220 9290 -27160
rect 9770 -27220 9950 -27160
rect 10430 -27220 10610 -27160
rect 11310 -27220 11490 -27160
rect 11970 -27220 12150 -27160
rect 12630 -27220 12810 -27160
rect 13510 -27220 13690 -27160
rect 14170 -27220 14350 -27160
rect 14830 -27220 15010 -27160
rect 15710 -27360 15890 -27300
rect 16370 -27360 16550 -27300
rect 17030 -27360 17210 -27300
rect 17910 -27360 18090 -27300
rect 18570 -27360 18750 -27300
rect 19230 -27360 19410 -27300
rect 430 -27510 610 -27430
rect 4710 -27530 6210 -27470
rect 6910 -27530 8410 -27470
rect 9110 -27530 10610 -27470
rect 11310 -27530 12810 -27470
rect 13510 -27530 15010 -27470
rect 15710 -27530 17210 -27470
rect 21310 -27510 21490 -27430
rect 6420 -27630 6480 -27570
rect 8840 -27630 8900 -27570
rect 11040 -27630 11100 -27570
rect 13240 -27630 13300 -27570
rect 15440 -27630 15500 -27570
rect 17420 -27630 17480 -27570
rect 4220 -27740 4280 -27680
rect 6640 -27740 6700 -27680
rect 8840 -27740 8900 -27680
rect 11040 -27740 11100 -27680
rect 13240 -27740 13300 -27680
rect 15220 -27740 15280 -27680
rect -70 -27850 -10 -27790
rect 2130 -27850 2190 -27790
rect 4330 -27850 4390 -27790
rect 6530 -27850 6590 -27790
rect 8730 -27850 8790 -27790
rect 10930 -27850 10990 -27790
rect 13130 -27850 13190 -27790
rect 15330 -27850 15390 -27790
rect 17530 -27850 17590 -27790
rect 19730 -27850 19790 -27790
rect 21930 -27850 21990 -27790
rect 2510 -28020 2690 -27960
rect 3170 -28020 3350 -27960
rect 3830 -28020 4010 -27960
rect 4710 -28020 4890 -27960
rect 5370 -28020 5550 -27960
rect 6030 -28020 6210 -27960
rect 6910 -28160 7090 -28100
rect 7570 -28160 7750 -28100
rect 8230 -28160 8410 -28100
rect 9110 -28160 9290 -28100
rect 9770 -28160 9950 -28100
rect 10430 -28160 10610 -28100
rect 11310 -28160 11490 -28100
rect 11970 -28160 12150 -28100
rect 12630 -28160 12810 -28100
rect 13510 -28160 13690 -28100
rect 14170 -28160 14350 -28100
rect 14830 -28160 15010 -28100
rect 15710 -28020 15890 -27960
rect 16370 -28020 16550 -27960
rect 17030 -28020 17210 -27960
rect 17910 -28020 18090 -27960
rect 18570 -28020 18750 -27960
rect 19230 -28020 19410 -27960
rect 430 -28310 610 -28230
rect 4710 -28330 6210 -28270
rect 6910 -28330 8410 -28270
rect 9110 -28330 10610 -28270
rect 11310 -28330 12810 -28270
rect 13510 -28330 15010 -28270
rect 15710 -28330 17210 -28270
rect 21310 -28310 21490 -28230
rect 6420 -28430 6480 -28370
rect 8840 -28430 8900 -28370
rect 11040 -28430 11100 -28370
rect 13240 -28430 13300 -28370
rect 15440 -28430 15500 -28370
rect 17420 -28430 17480 -28370
rect 4220 -28540 4280 -28480
rect 6640 -28540 6700 -28480
rect 8840 -28540 8900 -28480
rect 11040 -28540 11100 -28480
rect 13240 -28540 13300 -28480
rect 15220 -28540 15280 -28480
rect -70 -28650 -10 -28590
rect 2130 -28650 2190 -28590
rect 4330 -28650 4390 -28590
rect 6530 -28650 6590 -28590
rect 8730 -28650 8790 -28590
rect 10930 -28650 10990 -28590
rect 13130 -28650 13190 -28590
rect 15330 -28650 15390 -28590
rect 17530 -28650 17590 -28590
rect 19730 -28650 19790 -28590
rect 21930 -28650 21990 -28590
rect 2510 -28820 2690 -28760
rect 3170 -28820 3350 -28760
rect 3830 -28820 4010 -28760
rect 4710 -28820 4890 -28760
rect 5370 -28820 5550 -28760
rect 6030 -28820 6210 -28760
rect 6910 -28960 7090 -28900
rect 7570 -28960 7750 -28900
rect 8230 -28960 8410 -28900
rect 9110 -28960 9290 -28900
rect 9770 -28960 9950 -28900
rect 10430 -28960 10610 -28900
rect 11310 -28960 11490 -28900
rect 11970 -28960 12150 -28900
rect 12630 -28960 12810 -28900
rect 13510 -28960 13690 -28900
rect 14170 -28960 14350 -28900
rect 14830 -28960 15010 -28900
rect 15710 -28820 15890 -28760
rect 16370 -28820 16550 -28760
rect 17030 -28820 17210 -28760
rect 17910 -28820 18090 -28760
rect 18570 -28820 18750 -28760
rect 19230 -28820 19410 -28760
rect 430 -29110 610 -29030
rect 4710 -29130 6210 -29070
rect 6910 -29130 8410 -29070
rect 9110 -29130 10610 -29070
rect 11310 -29130 12810 -29070
rect 13510 -29130 15010 -29070
rect 15710 -29130 17210 -29070
rect 21310 -29110 21490 -29030
rect 6640 -29230 6700 -29170
rect 8620 -29230 8680 -29170
rect 10820 -29230 10880 -29170
rect 13020 -29230 13080 -29170
rect 15220 -29230 15280 -29170
rect 17640 -29230 17700 -29170
rect 4440 -29340 4500 -29280
rect 6420 -29340 6480 -29280
rect 8620 -29340 8680 -29280
rect 10820 -29340 10880 -29280
rect 13020 -29340 13080 -29280
rect 15440 -29340 15500 -29280
rect -70 -29450 -10 -29390
rect 2130 -29450 2190 -29390
rect 4330 -29450 4390 -29390
rect 6530 -29450 6590 -29390
rect 8730 -29450 8790 -29390
rect 10930 -29450 10990 -29390
rect 13130 -29450 13190 -29390
rect 15330 -29450 15390 -29390
rect 17530 -29450 17590 -29390
rect 19730 -29450 19790 -29390
rect 21930 -29450 21990 -29390
rect 2510 -29760 2690 -29700
rect 3170 -29760 3350 -29700
rect 3830 -29760 4010 -29700
rect 4710 -29760 4890 -29700
rect 5370 -29760 5550 -29700
rect 6030 -29760 6210 -29700
rect 6910 -29620 7090 -29560
rect 7570 -29620 7750 -29560
rect 8230 -29620 8410 -29560
rect 9110 -29620 9290 -29560
rect 9770 -29620 9950 -29560
rect 10430 -29620 10610 -29560
rect 11310 -29620 11490 -29560
rect 11970 -29620 12150 -29560
rect 12630 -29620 12810 -29560
rect 13510 -29620 13690 -29560
rect 14170 -29620 14350 -29560
rect 14830 -29620 15010 -29560
rect 15710 -29760 15890 -29700
rect 16370 -29760 16550 -29700
rect 17030 -29760 17210 -29700
rect 17910 -29760 18090 -29700
rect 18570 -29760 18750 -29700
rect 19230 -29760 19410 -29700
rect 2510 -29930 4010 -29870
rect 4710 -29930 6210 -29870
rect 6910 -29930 8410 -29870
rect 9110 -29930 10610 -29870
rect 11310 -29930 12810 -29870
rect 13510 -29930 15010 -29870
rect 15710 -29930 17210 -29870
rect 17910 -29930 19410 -29870
rect 4220 -30030 4280 -29970
rect 6420 -30030 6480 -29970
rect 8840 -30030 8900 -29970
rect 11040 -30030 11100 -29970
rect 13240 -30030 13300 -29970
rect 15440 -30030 15500 -29970
rect 17420 -30030 17480 -29970
rect 19620 -30030 19680 -29970
rect 2020 -30120 2080 -30060
rect 4220 -30140 4280 -30080
rect 6640 -30140 6700 -30080
rect 8840 -30140 8900 -30080
rect 11040 -30140 11100 -30080
rect 13240 -30140 13300 -30080
rect 15220 -30140 15280 -30080
rect 17420 -30140 17480 -30080
rect -70 -30250 -10 -30190
rect 2130 -30250 2190 -30190
rect 4330 -30250 4390 -30190
rect 6530 -30250 6590 -30190
rect 8730 -30250 8790 -30190
rect 10930 -30250 10990 -30190
rect 13130 -30250 13190 -30190
rect 15330 -30250 15390 -30190
rect 17530 -30250 17590 -30190
rect 19730 -30250 19790 -30190
rect 21930 -30250 21990 -30190
rect 2510 -30420 2690 -30360
rect 3170 -30420 3350 -30360
rect 3830 -30420 4010 -30360
rect 4710 -30420 4890 -30360
rect 5370 -30420 5550 -30360
rect 6030 -30420 6210 -30360
rect 6910 -30560 7090 -30500
rect 7570 -30560 7750 -30500
rect 8230 -30560 8410 -30500
rect 9110 -30560 9290 -30500
rect 9770 -30560 9950 -30500
rect 10430 -30560 10610 -30500
rect 11310 -30560 11490 -30500
rect 11970 -30560 12150 -30500
rect 12630 -30560 12810 -30500
rect 13510 -30560 13690 -30500
rect 14170 -30560 14350 -30500
rect 14830 -30560 15010 -30500
rect 15710 -30420 15890 -30360
rect 16370 -30420 16550 -30360
rect 17030 -30420 17210 -30360
rect 17910 -30420 18090 -30360
rect 18570 -30420 18750 -30360
rect 19230 -30420 19410 -30360
rect 2510 -30730 4010 -30670
rect 4710 -30730 6210 -30670
rect 6910 -30730 8410 -30670
rect 9110 -30730 10610 -30670
rect 11310 -30730 12810 -30670
rect 13510 -30730 15010 -30670
rect 15710 -30730 17210 -30670
rect 17910 -30730 19410 -30670
rect 4440 -30830 4500 -30770
rect 6640 -30830 6700 -30770
rect 8620 -30830 8680 -30770
rect 10820 -30830 10880 -30770
rect 13020 -30830 13080 -30770
rect 15220 -30830 15280 -30770
rect 17640 -30830 17700 -30770
rect 19840 -30830 19900 -30770
rect 2240 -30920 2300 -30860
rect 4440 -30940 4500 -30880
rect 6420 -30940 6480 -30880
rect 8620 -30940 8680 -30880
rect 10820 -30940 10880 -30880
rect 13020 -30940 13080 -30880
rect 15440 -30940 15500 -30880
rect 17640 -30940 17700 -30880
rect -70 -31050 -10 -30990
rect 2130 -31050 2190 -30990
rect 4330 -31050 4390 -30990
rect 6530 -31050 6590 -30990
rect 8730 -31050 8790 -30990
rect 10930 -31050 10990 -30990
rect 13130 -31050 13190 -30990
rect 15330 -31050 15390 -30990
rect 17530 -31050 17590 -30990
rect 19730 -31050 19790 -30990
rect 21930 -31050 21990 -30990
rect 2510 -31360 2690 -31300
rect 3170 -31360 3350 -31300
rect 3830 -31360 4010 -31300
rect 4710 -31360 4890 -31300
rect 5370 -31360 5550 -31300
rect 6030 -31360 6210 -31300
rect 6910 -31220 7090 -31160
rect 7570 -31220 7750 -31160
rect 8230 -31220 8410 -31160
rect 9110 -31220 9290 -31160
rect 9770 -31220 9950 -31160
rect 10430 -31220 10610 -31160
rect 11310 -31220 11490 -31160
rect 11970 -31220 12150 -31160
rect 12630 -31220 12810 -31160
rect 13510 -31220 13690 -31160
rect 14170 -31220 14350 -31160
rect 14830 -31220 15010 -31160
rect 15710 -31360 15890 -31300
rect 16370 -31360 16550 -31300
rect 17030 -31360 17210 -31300
rect 17910 -31360 18090 -31300
rect 18570 -31360 18750 -31300
rect 19230 -31360 19410 -31300
<< metal2 >>
rect 2020 11720 2080 12020
rect 2200 12010 2340 12020
rect 2200 11890 2210 12010
rect 2330 11890 2340 12010
rect 2200 11880 2340 11890
rect 1980 11710 2120 11720
rect 1980 11590 1990 11710
rect 2110 11590 2120 11710
rect 1980 11580 2120 11590
rect -70 10930 -10 10940
rect -70 10860 -10 10870
rect 2020 10830 2080 11580
rect 2130 10930 2190 10940
rect 2130 10860 2190 10870
rect 2240 10830 2300 11880
rect 4220 11720 4280 12020
rect 4400 12010 4540 12020
rect 4400 11890 4410 12010
rect 4530 11890 4540 12010
rect 4400 11880 4540 11890
rect 4180 11710 4320 11720
rect 4180 11590 4190 11710
rect 4310 11590 4320 11710
rect 4180 11580 4320 11590
rect 2500 11240 2700 11250
rect 2500 11180 2510 11240
rect 2690 11180 2700 11240
rect 2500 11170 2700 11180
rect 3160 11240 3360 11250
rect 3160 11180 3170 11240
rect 3350 11180 3360 11240
rect 3160 11170 3360 11180
rect 3820 11240 4020 11250
rect 3820 11180 3830 11240
rect 4010 11180 4020 11240
rect 3820 11170 4020 11180
rect 2500 11030 2700 11110
rect 3160 11030 3360 11110
rect 3820 11030 4020 11110
rect 4220 10830 4280 11580
rect 4330 10930 4390 10940
rect 4330 10860 4390 10870
rect 4440 10830 4500 11880
rect 6420 11720 6480 12020
rect 6600 12010 6740 12020
rect 6600 11890 6610 12010
rect 6730 11890 6740 12010
rect 6600 11880 6740 11890
rect 6380 11710 6520 11720
rect 6380 11590 6390 11710
rect 6510 11590 6520 11710
rect 6380 11580 6520 11590
rect 4700 11240 4900 11250
rect 4700 11180 4710 11240
rect 4890 11180 4900 11240
rect 4700 11170 4900 11180
rect 5360 11240 5560 11250
rect 5360 11180 5370 11240
rect 5550 11180 5560 11240
rect 5360 11170 5560 11180
rect 6020 11240 6220 11250
rect 6020 11180 6030 11240
rect 6210 11180 6220 11240
rect 6020 11170 6220 11180
rect 4700 11030 4900 11110
rect 5360 11030 5560 11110
rect 6020 11030 6220 11110
rect 6420 10830 6480 11580
rect 6530 10930 6590 10940
rect 6530 10860 6590 10870
rect 6640 10830 6700 11880
rect 8620 11720 8680 12020
rect 8800 12010 8940 12020
rect 8800 11890 8810 12010
rect 8930 11890 8940 12010
rect 8800 11880 8940 11890
rect 8580 11710 8720 11720
rect 8580 11590 8590 11710
rect 8710 11590 8720 11710
rect 8580 11580 8720 11590
rect 6900 11170 7100 11250
rect 7560 11170 7760 11250
rect 8220 11170 8420 11250
rect 6900 11100 7100 11110
rect 6900 11040 6910 11100
rect 7090 11040 7100 11100
rect 6900 11030 7100 11040
rect 7560 11100 7760 11110
rect 7560 11040 7570 11100
rect 7750 11040 7760 11100
rect 7560 11030 7760 11040
rect 8220 11100 8420 11110
rect 8220 11040 8230 11100
rect 8410 11040 8420 11100
rect 8220 11030 8420 11040
rect 8620 10830 8680 11580
rect 8730 10930 8790 10940
rect 8730 10860 8790 10870
rect 8840 10830 8900 11880
rect 10820 11720 10880 12020
rect 11000 12010 11140 12020
rect 11000 11890 11010 12010
rect 11130 11890 11140 12010
rect 11000 11880 11140 11890
rect 10780 11710 10920 11720
rect 10780 11590 10790 11710
rect 10910 11590 10920 11710
rect 10780 11580 10920 11590
rect 9100 11170 9300 11250
rect 9760 11170 9960 11250
rect 10420 11170 10620 11250
rect 9100 11100 9300 11110
rect 9100 11040 9110 11100
rect 9290 11040 9300 11100
rect 9100 11030 9300 11040
rect 9760 11100 9960 11110
rect 9760 11040 9770 11100
rect 9950 11040 9960 11100
rect 9760 11030 9960 11040
rect 10420 11100 10620 11110
rect 10420 11040 10430 11100
rect 10610 11040 10620 11100
rect 10420 11030 10620 11040
rect 10820 10830 10880 11580
rect 10930 10930 10990 10940
rect 10930 10860 10990 10870
rect 11040 10830 11100 11880
rect 13020 11720 13080 12020
rect 13200 12010 13340 12020
rect 13200 11890 13210 12010
rect 13330 11890 13340 12010
rect 13200 11880 13340 11890
rect 12980 11710 13120 11720
rect 12980 11590 12990 11710
rect 13110 11590 13120 11710
rect 12980 11580 13120 11590
rect 11300 11170 11500 11250
rect 11960 11170 12160 11250
rect 12620 11170 12820 11250
rect 11300 11100 11500 11110
rect 11300 11040 11310 11100
rect 11490 11040 11500 11100
rect 11300 11030 11500 11040
rect 11960 11100 12160 11110
rect 11960 11040 11970 11100
rect 12150 11040 12160 11100
rect 11960 11030 12160 11040
rect 12620 11100 12820 11110
rect 12620 11040 12630 11100
rect 12810 11040 12820 11100
rect 12620 11030 12820 11040
rect 13020 10830 13080 11580
rect 13130 10930 13190 10940
rect 13130 10860 13190 10870
rect 13240 10830 13300 11880
rect 15220 11720 15280 12020
rect 15400 12010 15540 12020
rect 15400 11890 15410 12010
rect 15530 11890 15540 12010
rect 15400 11880 15540 11890
rect 15180 11710 15320 11720
rect 15180 11590 15190 11710
rect 15310 11590 15320 11710
rect 15180 11580 15320 11590
rect 13500 11170 13700 11250
rect 14160 11170 14360 11250
rect 14820 11170 15020 11250
rect 13500 11100 13700 11110
rect 13500 11040 13510 11100
rect 13690 11040 13700 11100
rect 13500 11030 13700 11040
rect 14160 11100 14360 11110
rect 14160 11040 14170 11100
rect 14350 11040 14360 11100
rect 14160 11030 14360 11040
rect 14820 11100 15020 11110
rect 14820 11040 14830 11100
rect 15010 11040 15020 11100
rect 14820 11030 15020 11040
rect 15220 10830 15280 11580
rect 15330 10930 15390 10940
rect 15330 10860 15390 10870
rect 15440 10830 15500 11880
rect 17420 11720 17480 12020
rect 17600 12010 17740 12020
rect 17600 11890 17610 12010
rect 17730 11890 17740 12010
rect 17600 11880 17740 11890
rect 17380 11710 17520 11720
rect 17380 11590 17390 11710
rect 17510 11590 17520 11710
rect 17380 11580 17520 11590
rect 15700 11240 15900 11250
rect 15700 11180 15710 11240
rect 15890 11180 15900 11240
rect 15700 11170 15900 11180
rect 16360 11240 16560 11250
rect 16360 11180 16370 11240
rect 16550 11180 16560 11240
rect 16360 11170 16560 11180
rect 17020 11240 17220 11250
rect 17020 11180 17030 11240
rect 17210 11180 17220 11240
rect 17020 11170 17220 11180
rect 15700 11030 15900 11110
rect 16360 11030 16560 11110
rect 17020 11030 17220 11110
rect 17420 10830 17480 11580
rect 17530 10930 17590 10940
rect 17530 10860 17590 10870
rect 17640 10830 17700 11880
rect 19620 11720 19680 12020
rect 19800 12010 19940 12020
rect 19800 11890 19810 12010
rect 19930 11890 19940 12010
rect 19800 11880 19940 11890
rect 19580 11710 19720 11720
rect 19580 11590 19590 11710
rect 19710 11590 19720 11710
rect 19580 11580 19720 11590
rect 17900 11240 18100 11250
rect 17900 11180 17910 11240
rect 18090 11180 18100 11240
rect 17900 11170 18100 11180
rect 18560 11240 18760 11250
rect 18560 11180 18570 11240
rect 18750 11180 18760 11240
rect 18560 11170 18760 11180
rect 19220 11240 19420 11250
rect 19220 11180 19230 11240
rect 19410 11180 19420 11240
rect 19220 11170 19420 11180
rect 17900 11030 18100 11110
rect 18560 11030 18760 11110
rect 19220 11030 19420 11110
rect 2010 10710 2090 10830
rect 2010 10650 2020 10710
rect 2080 10650 2090 10710
rect 2010 10640 2090 10650
rect 2230 10640 2310 10830
rect 4210 10820 4290 10830
rect 4210 10760 4220 10820
rect 4280 10760 4290 10820
rect 4210 10710 4290 10760
rect 4210 10650 4220 10710
rect 4280 10650 4290 10710
rect 4210 10640 4290 10650
rect 4430 10640 4510 10830
rect 6410 10820 6490 10830
rect 6410 10760 6420 10820
rect 6480 10760 6490 10820
rect 6410 10640 6490 10760
rect 6630 10710 6710 10830
rect 6630 10650 6640 10710
rect 6700 10650 6710 10710
rect 6630 10640 6710 10650
rect 8610 10640 8690 10830
rect 8830 10820 8910 10830
rect 8830 10760 8840 10820
rect 8900 10760 8910 10820
rect 8830 10710 8910 10760
rect 8830 10650 8840 10710
rect 8900 10650 8910 10710
rect 8830 10640 8910 10650
rect 10810 10640 10890 10830
rect 11030 10820 11110 10830
rect 11030 10760 11040 10820
rect 11100 10760 11110 10820
rect 11030 10710 11110 10760
rect 11030 10650 11040 10710
rect 11100 10650 11110 10710
rect 11030 10640 11110 10650
rect 13010 10640 13090 10830
rect 13230 10820 13310 10830
rect 13230 10760 13240 10820
rect 13300 10760 13310 10820
rect 13230 10710 13310 10760
rect 13230 10650 13240 10710
rect 13300 10650 13310 10710
rect 13230 10640 13310 10650
rect 15210 10710 15290 10830
rect 15210 10650 15220 10710
rect 15280 10650 15290 10710
rect 15210 10640 15290 10650
rect 15430 10820 15510 10830
rect 15430 10760 15440 10820
rect 15500 10760 15510 10820
rect 15430 10640 15510 10760
rect 17410 10820 17490 10830
rect 17410 10760 17420 10820
rect 17480 10760 17490 10820
rect 17410 10710 17490 10760
rect 17410 10650 17420 10710
rect 17480 10650 17490 10710
rect 17410 10640 17490 10650
rect 17630 10640 17710 10830
rect 19620 10810 19680 11580
rect 19730 10930 19790 10940
rect 19730 10860 19790 10870
rect 19840 10810 19900 11880
rect 21930 10930 21990 10940
rect 21930 10860 21990 10870
rect 19610 10800 19690 10810
rect 19610 10740 19620 10800
rect 19680 10740 19690 10800
rect 19610 10640 19690 10740
rect 19830 10640 19910 10810
rect -70 10130 -10 10140
rect -70 10060 -10 10070
rect 2020 10030 2080 10640
rect 2130 10130 2190 10140
rect 2130 10060 2190 10070
rect 2240 10030 2300 10640
rect 2500 10610 4020 10620
rect 2500 10550 2510 10610
rect 4010 10550 4020 10610
rect 2500 10540 4020 10550
rect 2500 10370 2700 10450
rect 3160 10370 3360 10450
rect 3820 10370 4020 10450
rect 2500 10300 2700 10310
rect 2500 10240 2510 10300
rect 2690 10240 2700 10300
rect 2500 10230 2700 10240
rect 3160 10300 3360 10310
rect 3160 10240 3170 10300
rect 3350 10240 3360 10300
rect 3160 10230 3360 10240
rect 3820 10300 4020 10310
rect 3820 10240 3830 10300
rect 4010 10240 4020 10300
rect 3820 10230 4020 10240
rect 4220 10030 4280 10640
rect 4330 10130 4390 10140
rect 4330 10060 4390 10070
rect 4440 10030 4500 10640
rect 4700 10610 6220 10620
rect 4700 10550 4710 10610
rect 6210 10550 6220 10610
rect 4700 10540 6220 10550
rect 4700 10370 4900 10450
rect 5360 10370 5560 10450
rect 6020 10370 6220 10450
rect 4700 10300 4900 10310
rect 4700 10240 4710 10300
rect 4890 10240 4900 10300
rect 4700 10230 4900 10240
rect 5360 10300 5560 10310
rect 5360 10240 5370 10300
rect 5550 10240 5560 10300
rect 5360 10230 5560 10240
rect 6020 10300 6220 10310
rect 6020 10240 6030 10300
rect 6210 10240 6220 10300
rect 6020 10230 6220 10240
rect 6420 10030 6480 10640
rect 6530 10130 6590 10140
rect 6530 10060 6590 10070
rect 6640 10030 6700 10640
rect 6900 10610 8420 10620
rect 6900 10550 6910 10610
rect 8410 10550 8420 10610
rect 6900 10540 8420 10550
rect 6900 10440 7100 10450
rect 6900 10380 6910 10440
rect 7090 10380 7100 10440
rect 6900 10370 7100 10380
rect 7560 10440 7760 10450
rect 7560 10380 7570 10440
rect 7750 10380 7760 10440
rect 7560 10370 7760 10380
rect 8220 10440 8420 10450
rect 8220 10380 8230 10440
rect 8410 10380 8420 10440
rect 8220 10370 8420 10380
rect 6900 10230 7100 10310
rect 7560 10230 7760 10310
rect 8220 10230 8420 10310
rect 8620 10030 8680 10640
rect 8730 10130 8790 10140
rect 8730 10060 8790 10070
rect 8840 10030 8900 10640
rect 9100 10610 10620 10620
rect 9100 10550 9110 10610
rect 10610 10550 10620 10610
rect 9100 10540 10620 10550
rect 9100 10440 9300 10450
rect 9100 10380 9110 10440
rect 9290 10380 9300 10440
rect 9100 10370 9300 10380
rect 9760 10440 9960 10450
rect 9760 10380 9770 10440
rect 9950 10380 9960 10440
rect 9760 10370 9960 10380
rect 10420 10440 10620 10450
rect 10420 10380 10430 10440
rect 10610 10380 10620 10440
rect 10420 10370 10620 10380
rect 9100 10230 9300 10310
rect 9760 10230 9960 10310
rect 10420 10230 10620 10310
rect 10820 10030 10880 10640
rect 10930 10130 10990 10140
rect 10930 10060 10990 10070
rect 11040 10030 11100 10640
rect 11300 10610 12820 10620
rect 11300 10550 11310 10610
rect 12810 10550 12820 10610
rect 11300 10540 12820 10550
rect 11300 10440 11500 10450
rect 11300 10380 11310 10440
rect 11490 10380 11500 10440
rect 11300 10370 11500 10380
rect 11960 10440 12160 10450
rect 11960 10380 11970 10440
rect 12150 10380 12160 10440
rect 11960 10370 12160 10380
rect 12620 10440 12820 10450
rect 12620 10380 12630 10440
rect 12810 10380 12820 10440
rect 12620 10370 12820 10380
rect 11300 10230 11500 10310
rect 11960 10230 12160 10310
rect 12620 10230 12820 10310
rect 13020 10030 13080 10640
rect 13130 10130 13190 10140
rect 13130 10060 13190 10070
rect 13240 10030 13300 10640
rect 13500 10610 15020 10620
rect 13500 10550 13510 10610
rect 15010 10550 15020 10610
rect 13500 10540 15020 10550
rect 13500 10440 13700 10450
rect 13500 10380 13510 10440
rect 13690 10380 13700 10440
rect 13500 10370 13700 10380
rect 14160 10440 14360 10450
rect 14160 10380 14170 10440
rect 14350 10380 14360 10440
rect 14160 10370 14360 10380
rect 14820 10440 15020 10450
rect 14820 10380 14830 10440
rect 15010 10380 15020 10440
rect 14820 10370 15020 10380
rect 13500 10230 13700 10310
rect 14160 10230 14360 10310
rect 14820 10230 15020 10310
rect 15220 10030 15280 10640
rect 15330 10130 15390 10140
rect 15330 10060 15390 10070
rect 15440 10030 15500 10640
rect 15700 10610 17220 10620
rect 15700 10550 15710 10610
rect 17210 10550 17220 10610
rect 15700 10540 17220 10550
rect 15700 10370 15900 10450
rect 16360 10370 16560 10450
rect 17020 10370 17220 10450
rect 15700 10300 15900 10310
rect 15700 10240 15710 10300
rect 15890 10240 15900 10300
rect 15700 10230 15900 10240
rect 16360 10300 16560 10310
rect 16360 10240 16370 10300
rect 16550 10240 16560 10300
rect 16360 10230 16560 10240
rect 17020 10300 17220 10310
rect 17020 10240 17030 10300
rect 17210 10240 17220 10300
rect 17020 10230 17220 10240
rect 17420 10030 17480 10640
rect 17530 10130 17590 10140
rect 17530 10060 17590 10070
rect 17640 10030 17700 10640
rect 17900 10610 19420 10620
rect 17900 10550 17910 10610
rect 19410 10550 19420 10610
rect 17900 10540 19420 10550
rect 17900 10370 18100 10450
rect 18560 10370 18760 10450
rect 19220 10370 19420 10450
rect 17900 10300 18100 10310
rect 17900 10240 17910 10300
rect 18090 10240 18100 10300
rect 17900 10230 18100 10240
rect 18560 10300 18760 10310
rect 18560 10240 18570 10300
rect 18750 10240 18760 10300
rect 18560 10230 18760 10240
rect 19220 10300 19420 10310
rect 19220 10240 19230 10300
rect 19410 10240 19420 10300
rect 19220 10230 19420 10240
rect 2010 9840 2090 10030
rect 2230 9910 2310 10030
rect 2230 9850 2240 9910
rect 2300 9850 2310 9910
rect 2230 9840 2310 9850
rect 4210 9840 4290 10030
rect 4430 10020 4510 10030
rect 4430 9960 4440 10020
rect 4500 9960 4510 10020
rect 4430 9910 4510 9960
rect 4430 9850 4440 9910
rect 4500 9850 4510 9910
rect 4430 9840 4510 9850
rect 6410 9910 6490 10030
rect 6410 9850 6420 9910
rect 6480 9850 6490 9910
rect 6410 9840 6490 9850
rect 6630 10020 6710 10030
rect 6630 9960 6640 10020
rect 6700 9960 6710 10020
rect 6630 9840 6710 9960
rect 8610 10020 8690 10030
rect 8610 9960 8620 10020
rect 8680 9960 8690 10020
rect 8610 9910 8690 9960
rect 8610 9850 8620 9910
rect 8680 9850 8690 9910
rect 8610 9840 8690 9850
rect 8830 9840 8910 10030
rect 10810 10020 10890 10030
rect 10810 9960 10820 10020
rect 10880 9960 10890 10020
rect 10810 9910 10890 9960
rect 10810 9850 10820 9910
rect 10880 9850 10890 9910
rect 10810 9840 10890 9850
rect 11030 9840 11110 10030
rect 13010 10020 13090 10030
rect 13010 9960 13020 10020
rect 13080 9960 13090 10020
rect 13010 9910 13090 9960
rect 13010 9850 13020 9910
rect 13080 9850 13090 9910
rect 13010 9840 13090 9850
rect 13230 9840 13310 10030
rect 15210 10020 15290 10030
rect 15210 9960 15220 10020
rect 15280 9960 15290 10020
rect 15210 9840 15290 9960
rect 15430 9910 15510 10030
rect 15430 9850 15440 9910
rect 15500 9850 15510 9910
rect 15430 9840 15510 9850
rect 17410 9840 17490 10030
rect 17630 10020 17710 10030
rect 17630 9960 17640 10020
rect 17700 9960 17710 10020
rect 19620 10010 19680 10640
rect 19730 10130 19790 10140
rect 19730 10060 19790 10070
rect 19840 10010 19900 10640
rect 21930 10130 21990 10140
rect 21930 10060 21990 10070
rect 17630 9910 17710 9960
rect 17630 9850 17640 9910
rect 17700 9850 17710 9910
rect 17630 9840 17710 9850
rect 19610 9840 19690 10010
rect 19830 10000 19910 10010
rect 19830 9940 19840 10000
rect 19900 9940 19910 10000
rect 19830 9840 19910 9940
rect -70 9330 -10 9340
rect -70 9260 -10 9270
rect 2020 9230 2080 9840
rect 2130 9330 2190 9340
rect 2130 9260 2190 9270
rect 2240 9230 2300 9840
rect 2500 9810 4020 9820
rect 2500 9750 2510 9810
rect 4010 9750 4020 9810
rect 2500 9740 4020 9750
rect 2500 9640 2700 9650
rect 2500 9580 2510 9640
rect 2690 9580 2700 9640
rect 2500 9570 2700 9580
rect 3160 9640 3360 9650
rect 3160 9580 3170 9640
rect 3350 9580 3360 9640
rect 3160 9570 3360 9580
rect 3820 9640 4020 9650
rect 3820 9580 3830 9640
rect 4010 9580 4020 9640
rect 3820 9570 4020 9580
rect 2500 9430 2700 9510
rect 3160 9430 3360 9510
rect 3820 9430 4020 9510
rect 4220 9230 4280 9840
rect 4330 9330 4390 9340
rect 4330 9260 4390 9270
rect 4440 9230 4500 9840
rect 4700 9810 6220 9820
rect 4700 9750 4710 9810
rect 6210 9750 6220 9810
rect 4700 9740 6220 9750
rect 4700 9640 4900 9650
rect 4700 9580 4710 9640
rect 4890 9580 4900 9640
rect 4700 9570 4900 9580
rect 5360 9640 5560 9650
rect 5360 9580 5370 9640
rect 5550 9580 5560 9640
rect 5360 9570 5560 9580
rect 6020 9640 6220 9650
rect 6020 9580 6030 9640
rect 6210 9580 6220 9640
rect 6020 9570 6220 9580
rect 4700 9430 4900 9510
rect 5360 9430 5560 9510
rect 6020 9430 6220 9510
rect 6420 9230 6480 9840
rect 6530 9330 6590 9340
rect 6530 9260 6590 9270
rect 6640 9230 6700 9840
rect 6900 9810 8420 9820
rect 6900 9750 6910 9810
rect 8410 9750 8420 9810
rect 6900 9740 8420 9750
rect 6900 9570 7100 9650
rect 7560 9570 7760 9650
rect 8220 9570 8420 9650
rect 6900 9500 7100 9510
rect 6900 9440 6910 9500
rect 7090 9440 7100 9500
rect 6900 9430 7100 9440
rect 7560 9500 7760 9510
rect 7560 9440 7570 9500
rect 7750 9440 7760 9500
rect 7560 9430 7760 9440
rect 8220 9500 8420 9510
rect 8220 9440 8230 9500
rect 8410 9440 8420 9500
rect 8220 9430 8420 9440
rect 8620 9230 8680 9840
rect 8730 9330 8790 9340
rect 8730 9260 8790 9270
rect 8840 9230 8900 9840
rect 9100 9810 10620 9820
rect 9100 9750 9110 9810
rect 10610 9750 10620 9810
rect 9100 9740 10620 9750
rect 9100 9570 9300 9650
rect 9760 9570 9960 9650
rect 10420 9570 10620 9650
rect 9100 9500 9300 9510
rect 9100 9440 9110 9500
rect 9290 9440 9300 9500
rect 9100 9430 9300 9440
rect 9760 9500 9960 9510
rect 9760 9440 9770 9500
rect 9950 9440 9960 9500
rect 9760 9430 9960 9440
rect 10420 9500 10620 9510
rect 10420 9440 10430 9500
rect 10610 9440 10620 9500
rect 10420 9430 10620 9440
rect 10820 9230 10880 9840
rect 10930 9330 10990 9340
rect 10930 9260 10990 9270
rect 11040 9230 11100 9840
rect 11300 9810 12820 9820
rect 11300 9750 11310 9810
rect 12810 9750 12820 9810
rect 11300 9740 12820 9750
rect 11300 9570 11500 9650
rect 11960 9570 12160 9650
rect 12620 9570 12820 9650
rect 11300 9500 11500 9510
rect 11300 9440 11310 9500
rect 11490 9440 11500 9500
rect 11300 9430 11500 9440
rect 11960 9500 12160 9510
rect 11960 9440 11970 9500
rect 12150 9440 12160 9500
rect 11960 9430 12160 9440
rect 12620 9500 12820 9510
rect 12620 9440 12630 9500
rect 12810 9440 12820 9500
rect 12620 9430 12820 9440
rect 13020 9230 13080 9840
rect 13130 9330 13190 9340
rect 13130 9260 13190 9270
rect 13240 9230 13300 9840
rect 13500 9810 15020 9820
rect 13500 9750 13510 9810
rect 15010 9750 15020 9810
rect 13500 9740 15020 9750
rect 13500 9570 13700 9650
rect 14160 9570 14360 9650
rect 14820 9570 15020 9650
rect 13500 9500 13700 9510
rect 13500 9440 13510 9500
rect 13690 9440 13700 9500
rect 13500 9430 13700 9440
rect 14160 9500 14360 9510
rect 14160 9440 14170 9500
rect 14350 9440 14360 9500
rect 14160 9430 14360 9440
rect 14820 9500 15020 9510
rect 14820 9440 14830 9500
rect 15010 9440 15020 9500
rect 14820 9430 15020 9440
rect 15220 9230 15280 9840
rect 15330 9330 15390 9340
rect 15330 9260 15390 9270
rect 15440 9230 15500 9840
rect 15700 9810 17220 9820
rect 15700 9750 15710 9810
rect 17210 9750 17220 9810
rect 15700 9740 17220 9750
rect 15700 9640 15900 9650
rect 15700 9580 15710 9640
rect 15890 9580 15900 9640
rect 15700 9570 15900 9580
rect 16360 9640 16560 9650
rect 16360 9580 16370 9640
rect 16550 9580 16560 9640
rect 16360 9570 16560 9580
rect 17020 9640 17220 9650
rect 17020 9580 17030 9640
rect 17210 9580 17220 9640
rect 17020 9570 17220 9580
rect 15700 9430 15900 9510
rect 16360 9430 16560 9510
rect 17020 9430 17220 9510
rect 17420 9230 17480 9840
rect 17530 9330 17590 9340
rect 17530 9260 17590 9270
rect 17640 9230 17700 9840
rect 17900 9810 19420 9820
rect 17900 9750 17910 9810
rect 19410 9750 19420 9810
rect 17900 9740 19420 9750
rect 17900 9640 18100 9650
rect 17900 9580 17910 9640
rect 18090 9580 18100 9640
rect 17900 9570 18100 9580
rect 18560 9640 18760 9650
rect 18560 9580 18570 9640
rect 18750 9580 18760 9640
rect 18560 9570 18760 9580
rect 19220 9640 19420 9650
rect 19220 9580 19230 9640
rect 19410 9580 19420 9640
rect 19220 9570 19420 9580
rect 17900 9430 18100 9510
rect 18560 9430 18760 9510
rect 19220 9430 19420 9510
rect 2010 9040 2090 9230
rect 2230 9040 2310 9230
rect 4210 9110 4290 9230
rect 4210 9050 4220 9110
rect 4280 9050 4290 9110
rect 4210 9040 4290 9050
rect 4430 9040 4510 9230
rect 6410 9220 6490 9230
rect 6410 9160 6420 9220
rect 6480 9160 6490 9220
rect 6410 9040 6490 9160
rect 6630 9110 6710 9230
rect 6630 9050 6640 9110
rect 6700 9050 6710 9110
rect 6630 9040 6710 9050
rect 8610 9040 8690 9230
rect 8830 9220 8910 9230
rect 8830 9160 8840 9220
rect 8900 9160 8910 9220
rect 8830 9110 8910 9160
rect 8830 9050 8840 9110
rect 8900 9050 8910 9110
rect 8830 9040 8910 9050
rect 10810 9040 10890 9230
rect 11030 9220 11110 9230
rect 11030 9160 11040 9220
rect 11100 9160 11110 9220
rect 11030 9110 11110 9160
rect 11030 9050 11040 9110
rect 11100 9050 11110 9110
rect 11030 9040 11110 9050
rect 13010 9040 13090 9230
rect 13230 9220 13310 9230
rect 13230 9160 13240 9220
rect 13300 9160 13310 9220
rect 13230 9110 13310 9160
rect 13230 9050 13240 9110
rect 13300 9050 13310 9110
rect 13230 9040 13310 9050
rect 15210 9110 15290 9230
rect 15210 9050 15220 9110
rect 15280 9050 15290 9110
rect 15210 9040 15290 9050
rect 15430 9220 15510 9230
rect 15430 9160 15440 9220
rect 15500 9160 15510 9220
rect 15430 9040 15510 9160
rect 17410 9220 17490 9230
rect 17410 9160 17420 9220
rect 17480 9160 17490 9220
rect 17410 9040 17490 9160
rect 17630 9040 17710 9230
rect 19620 9210 19680 9840
rect 19730 9330 19790 9340
rect 19730 9260 19790 9270
rect 19840 9210 19900 9840
rect 21930 9330 21990 9340
rect 21930 9260 21990 9270
rect 19610 9040 19690 9210
rect 19830 9040 19910 9210
rect 420 8990 620 9000
rect 420 8910 430 8990
rect 610 8910 620 8990
rect 420 8900 620 8910
rect -70 8530 -10 8540
rect -70 8460 -10 8470
rect 2020 8430 2080 9040
rect 2130 8530 2190 8540
rect 2130 8460 2190 8470
rect 2240 8430 2300 9040
rect 2500 8770 2700 8850
rect 3160 8770 3360 8850
rect 3820 8770 4020 8850
rect 2500 8700 2700 8710
rect 2500 8640 2510 8700
rect 2690 8640 2700 8700
rect 2500 8630 2700 8640
rect 3160 8700 3360 8710
rect 3160 8640 3170 8700
rect 3350 8640 3360 8700
rect 3160 8630 3360 8640
rect 3820 8700 4020 8710
rect 3820 8640 3830 8700
rect 4010 8640 4020 8700
rect 3820 8630 4020 8640
rect 4220 8430 4280 9040
rect 4330 8530 4390 8540
rect 4330 8460 4390 8470
rect 4440 8430 4500 9040
rect 4700 9010 6220 9020
rect 4700 8950 4710 9010
rect 6210 8950 6220 9010
rect 4700 8940 6220 8950
rect 4700 8770 4900 8850
rect 5360 8770 5560 8850
rect 6020 8770 6220 8850
rect 4700 8700 4900 8710
rect 4700 8640 4710 8700
rect 4890 8640 4900 8700
rect 4700 8630 4900 8640
rect 5360 8700 5560 8710
rect 5360 8640 5370 8700
rect 5550 8640 5560 8700
rect 5360 8630 5560 8640
rect 6020 8700 6220 8710
rect 6020 8640 6030 8700
rect 6210 8640 6220 8700
rect 6020 8630 6220 8640
rect 6420 8430 6480 9040
rect 6530 8530 6590 8540
rect 6530 8460 6590 8470
rect 6640 8430 6700 9040
rect 6900 9010 8420 9020
rect 6900 8950 6910 9010
rect 8410 8950 8420 9010
rect 6900 8940 8420 8950
rect 6900 8840 7100 8850
rect 6900 8780 6910 8840
rect 7090 8780 7100 8840
rect 6900 8770 7100 8780
rect 7560 8840 7760 8850
rect 7560 8780 7570 8840
rect 7750 8780 7760 8840
rect 7560 8770 7760 8780
rect 8220 8840 8420 8850
rect 8220 8780 8230 8840
rect 8410 8780 8420 8840
rect 8220 8770 8420 8780
rect 6900 8630 7100 8710
rect 7560 8630 7760 8710
rect 8220 8630 8420 8710
rect 8620 8430 8680 9040
rect 8730 8530 8790 8540
rect 8730 8460 8790 8470
rect 8840 8430 8900 9040
rect 9100 9010 10620 9020
rect 9100 8950 9110 9010
rect 10610 8950 10620 9010
rect 9100 8940 10620 8950
rect 9100 8840 9300 8850
rect 9100 8780 9110 8840
rect 9290 8780 9300 8840
rect 9100 8770 9300 8780
rect 9760 8840 9960 8850
rect 9760 8780 9770 8840
rect 9950 8780 9960 8840
rect 9760 8770 9960 8780
rect 10420 8840 10620 8850
rect 10420 8780 10430 8840
rect 10610 8780 10620 8840
rect 10420 8770 10620 8780
rect 9100 8630 9300 8710
rect 9760 8630 9960 8710
rect 10420 8630 10620 8710
rect 10820 8430 10880 9040
rect 10930 8530 10990 8540
rect 10930 8460 10990 8470
rect 11040 8430 11100 9040
rect 11300 9010 12820 9020
rect 11300 8950 11310 9010
rect 12810 8950 12820 9010
rect 11300 8940 12820 8950
rect 11300 8840 11500 8850
rect 11300 8780 11310 8840
rect 11490 8780 11500 8840
rect 11300 8770 11500 8780
rect 11960 8840 12160 8850
rect 11960 8780 11970 8840
rect 12150 8780 12160 8840
rect 11960 8770 12160 8780
rect 12620 8840 12820 8850
rect 12620 8780 12630 8840
rect 12810 8780 12820 8840
rect 12620 8770 12820 8780
rect 11300 8630 11500 8710
rect 11960 8630 12160 8710
rect 12620 8630 12820 8710
rect 13020 8430 13080 9040
rect 13130 8530 13190 8540
rect 13130 8460 13190 8470
rect 13240 8430 13300 9040
rect 13500 9010 15020 9020
rect 13500 8950 13510 9010
rect 15010 8950 15020 9010
rect 13500 8940 15020 8950
rect 13500 8840 13700 8850
rect 13500 8780 13510 8840
rect 13690 8780 13700 8840
rect 13500 8770 13700 8780
rect 14160 8840 14360 8850
rect 14160 8780 14170 8840
rect 14350 8780 14360 8840
rect 14160 8770 14360 8780
rect 14820 8840 15020 8850
rect 14820 8780 14830 8840
rect 15010 8780 15020 8840
rect 14820 8770 15020 8780
rect 13500 8630 13700 8710
rect 14160 8630 14360 8710
rect 14820 8630 15020 8710
rect 15220 8430 15280 9040
rect 15330 8530 15390 8540
rect 15330 8460 15390 8470
rect 15440 8430 15500 9040
rect 15700 9010 17220 9020
rect 15700 8950 15710 9010
rect 17210 8950 17220 9010
rect 15700 8940 17220 8950
rect 15700 8770 15900 8850
rect 16360 8770 16560 8850
rect 17020 8770 17220 8850
rect 15700 8700 15900 8710
rect 15700 8640 15710 8700
rect 15890 8640 15900 8700
rect 15700 8630 15900 8640
rect 16360 8700 16560 8710
rect 16360 8640 16370 8700
rect 16550 8640 16560 8700
rect 16360 8630 16560 8640
rect 17020 8700 17220 8710
rect 17020 8640 17030 8700
rect 17210 8640 17220 8700
rect 17020 8630 17220 8640
rect 17420 8430 17480 9040
rect 17530 8530 17590 8540
rect 17530 8460 17590 8470
rect 17640 8430 17700 9040
rect 17900 8770 18100 8850
rect 18560 8770 18760 8850
rect 19220 8770 19420 8850
rect 17900 8700 18100 8710
rect 17900 8640 17910 8700
rect 18090 8640 18100 8700
rect 17900 8630 18100 8640
rect 18560 8700 18760 8710
rect 18560 8640 18570 8700
rect 18750 8640 18760 8700
rect 18560 8630 18760 8640
rect 19220 8700 19420 8710
rect 19220 8640 19230 8700
rect 19410 8640 19420 8700
rect 19220 8630 19420 8640
rect 2010 8240 2090 8430
rect 2230 8240 2310 8430
rect 4210 8240 4290 8430
rect 4430 8310 4510 8430
rect 4430 8250 4440 8310
rect 4500 8250 4510 8310
rect 4430 8240 4510 8250
rect 6410 8310 6490 8430
rect 6410 8250 6420 8310
rect 6480 8250 6490 8310
rect 6410 8240 6490 8250
rect 6630 8420 6710 8430
rect 6630 8360 6640 8420
rect 6700 8360 6710 8420
rect 6630 8240 6710 8360
rect 8610 8420 8690 8430
rect 8610 8360 8620 8420
rect 8680 8360 8690 8420
rect 8610 8310 8690 8360
rect 8610 8250 8620 8310
rect 8680 8250 8690 8310
rect 8610 8240 8690 8250
rect 8830 8240 8910 8430
rect 10810 8420 10890 8430
rect 10810 8360 10820 8420
rect 10880 8360 10890 8420
rect 10810 8310 10890 8360
rect 10810 8250 10820 8310
rect 10880 8250 10890 8310
rect 10810 8240 10890 8250
rect 11030 8240 11110 8430
rect 13010 8420 13090 8430
rect 13010 8360 13020 8420
rect 13080 8360 13090 8420
rect 13010 8310 13090 8360
rect 13010 8250 13020 8310
rect 13080 8250 13090 8310
rect 13010 8240 13090 8250
rect 13230 8240 13310 8430
rect 15210 8420 15290 8430
rect 15210 8360 15220 8420
rect 15280 8360 15290 8420
rect 15210 8240 15290 8360
rect 15430 8310 15510 8430
rect 15430 8250 15440 8310
rect 15500 8250 15510 8310
rect 15430 8240 15510 8250
rect 17410 8240 17490 8430
rect 17630 8420 17710 8430
rect 17630 8360 17640 8420
rect 17700 8360 17710 8420
rect 19620 8410 19680 9040
rect 19730 8530 19790 8540
rect 19730 8460 19790 8470
rect 19840 8410 19900 9040
rect 21300 8990 21500 9000
rect 21300 8910 21310 8990
rect 21490 8910 21500 8990
rect 21300 8900 21500 8910
rect 21930 8530 21990 8540
rect 21930 8460 21990 8470
rect 17630 8240 17710 8360
rect 19610 8240 19690 8410
rect 19830 8240 19910 8410
rect 420 8190 620 8200
rect 420 8110 430 8190
rect 610 8110 620 8190
rect 420 8100 620 8110
rect -70 7730 -10 7740
rect -70 7660 -10 7670
rect 2020 7630 2080 8240
rect 2130 7730 2190 7740
rect 2130 7660 2190 7670
rect 2240 7630 2300 8240
rect 2500 7970 2700 8050
rect 3160 7970 3360 8050
rect 3820 7970 4020 8050
rect 2500 7900 2700 7910
rect 2500 7840 2510 7900
rect 2690 7840 2700 7900
rect 2500 7830 2700 7840
rect 3160 7900 3360 7910
rect 3160 7840 3170 7900
rect 3350 7840 3360 7900
rect 3160 7830 3360 7840
rect 3820 7900 4020 7910
rect 3820 7840 3830 7900
rect 4010 7840 4020 7900
rect 3820 7830 4020 7840
rect 4220 7630 4280 8240
rect 4330 7730 4390 7740
rect 4330 7660 4390 7670
rect 4440 7630 4500 8240
rect 4700 8210 6220 8220
rect 4700 8150 4710 8210
rect 6210 8150 6220 8210
rect 4700 8140 6220 8150
rect 4700 7970 4900 8050
rect 5360 7970 5560 8050
rect 6020 7970 6220 8050
rect 4700 7900 4900 7910
rect 4700 7840 4710 7900
rect 4890 7840 4900 7900
rect 4700 7830 4900 7840
rect 5360 7900 5560 7910
rect 5360 7840 5370 7900
rect 5550 7840 5560 7900
rect 5360 7830 5560 7840
rect 6020 7900 6220 7910
rect 6020 7840 6030 7900
rect 6210 7840 6220 7900
rect 6020 7830 6220 7840
rect 6420 7630 6480 8240
rect 6530 7730 6590 7740
rect 6530 7660 6590 7670
rect 6640 7630 6700 8240
rect 6900 8210 8420 8220
rect 6900 8150 6910 8210
rect 8410 8150 8420 8210
rect 6900 8140 8420 8150
rect 6900 8040 7100 8050
rect 6900 7980 6910 8040
rect 7090 7980 7100 8040
rect 6900 7970 7100 7980
rect 7560 8040 7760 8050
rect 7560 7980 7570 8040
rect 7750 7980 7760 8040
rect 7560 7970 7760 7980
rect 8220 8040 8420 8050
rect 8220 7980 8230 8040
rect 8410 7980 8420 8040
rect 8220 7970 8420 7980
rect 6900 7830 7100 7910
rect 7560 7830 7760 7910
rect 8220 7830 8420 7910
rect 8620 7630 8680 8240
rect 8730 7730 8790 7740
rect 8730 7660 8790 7670
rect 8840 7630 8900 8240
rect 9100 8210 10620 8220
rect 9100 8150 9110 8210
rect 10610 8150 10620 8210
rect 9100 8140 10620 8150
rect 9100 8040 9300 8050
rect 9100 7980 9110 8040
rect 9290 7980 9300 8040
rect 9100 7970 9300 7980
rect 9760 8040 9960 8050
rect 9760 7980 9770 8040
rect 9950 7980 9960 8040
rect 9760 7970 9960 7980
rect 10420 8040 10620 8050
rect 10420 7980 10430 8040
rect 10610 7980 10620 8040
rect 10420 7970 10620 7980
rect 9100 7830 9300 7910
rect 9760 7830 9960 7910
rect 10420 7830 10620 7910
rect 10820 7630 10880 8240
rect 10930 7730 10990 7740
rect 10930 7660 10990 7670
rect 11040 7630 11100 8240
rect 11300 8210 12820 8220
rect 11300 8150 11310 8210
rect 12810 8150 12820 8210
rect 11300 8140 12820 8150
rect 11300 8040 11500 8050
rect 11300 7980 11310 8040
rect 11490 7980 11500 8040
rect 11300 7970 11500 7980
rect 11960 8040 12160 8050
rect 11960 7980 11970 8040
rect 12150 7980 12160 8040
rect 11960 7970 12160 7980
rect 12620 8040 12820 8050
rect 12620 7980 12630 8040
rect 12810 7980 12820 8040
rect 12620 7970 12820 7980
rect 11300 7830 11500 7910
rect 11960 7830 12160 7910
rect 12620 7830 12820 7910
rect 13020 7630 13080 8240
rect 13130 7730 13190 7740
rect 13130 7660 13190 7670
rect 13240 7630 13300 8240
rect 13500 8210 15020 8220
rect 13500 8150 13510 8210
rect 15010 8150 15020 8210
rect 13500 8140 15020 8150
rect 13500 8040 13700 8050
rect 13500 7980 13510 8040
rect 13690 7980 13700 8040
rect 13500 7970 13700 7980
rect 14160 8040 14360 8050
rect 14160 7980 14170 8040
rect 14350 7980 14360 8040
rect 14160 7970 14360 7980
rect 14820 8040 15020 8050
rect 14820 7980 14830 8040
rect 15010 7980 15020 8040
rect 14820 7970 15020 7980
rect 13500 7830 13700 7910
rect 14160 7830 14360 7910
rect 14820 7830 15020 7910
rect 15220 7630 15280 8240
rect 15330 7730 15390 7740
rect 15330 7660 15390 7670
rect 15440 7630 15500 8240
rect 15700 8210 17220 8220
rect 15700 8150 15710 8210
rect 17210 8150 17220 8210
rect 15700 8140 17220 8150
rect 15700 7970 15900 8050
rect 16360 7970 16560 8050
rect 17020 7970 17220 8050
rect 15700 7900 15900 7910
rect 15700 7840 15710 7900
rect 15890 7840 15900 7900
rect 15700 7830 15900 7840
rect 16360 7900 16560 7910
rect 16360 7840 16370 7900
rect 16550 7840 16560 7900
rect 16360 7830 16560 7840
rect 17020 7900 17220 7910
rect 17020 7840 17030 7900
rect 17210 7840 17220 7900
rect 17020 7830 17220 7840
rect 17420 7630 17480 8240
rect 17530 7730 17590 7740
rect 17530 7660 17590 7670
rect 17640 7630 17700 8240
rect 17900 7970 18100 8050
rect 18560 7970 18760 8050
rect 19220 7970 19420 8050
rect 17900 7900 18100 7910
rect 17900 7840 17910 7900
rect 18090 7840 18100 7900
rect 17900 7830 18100 7840
rect 18560 7900 18760 7910
rect 18560 7840 18570 7900
rect 18750 7840 18760 7900
rect 18560 7830 18760 7840
rect 19220 7900 19420 7910
rect 19220 7840 19230 7900
rect 19410 7840 19420 7900
rect 19220 7830 19420 7840
rect 2010 7440 2090 7630
rect 2230 7440 2310 7630
rect 4210 7440 4290 7630
rect 4430 7510 4510 7630
rect 4430 7450 4440 7510
rect 4500 7450 4510 7510
rect 4430 7440 4510 7450
rect 6410 7510 6490 7630
rect 6410 7450 6420 7510
rect 6480 7450 6490 7510
rect 6410 7440 6490 7450
rect 6630 7620 6710 7630
rect 6630 7560 6640 7620
rect 6700 7560 6710 7620
rect 6630 7440 6710 7560
rect 8610 7620 8690 7630
rect 8610 7560 8620 7620
rect 8680 7560 8690 7620
rect 8610 7510 8690 7560
rect 8610 7450 8620 7510
rect 8680 7450 8690 7510
rect 8610 7440 8690 7450
rect 8830 7440 8910 7630
rect 10810 7620 10890 7630
rect 10810 7560 10820 7620
rect 10880 7560 10890 7620
rect 10810 7510 10890 7560
rect 10810 7450 10820 7510
rect 10880 7450 10890 7510
rect 10810 7440 10890 7450
rect 11030 7440 11110 7630
rect 13010 7620 13090 7630
rect 13010 7560 13020 7620
rect 13080 7560 13090 7620
rect 13010 7510 13090 7560
rect 13010 7450 13020 7510
rect 13080 7450 13090 7510
rect 13010 7440 13090 7450
rect 13230 7440 13310 7630
rect 15210 7620 15290 7630
rect 15210 7560 15220 7620
rect 15280 7560 15290 7620
rect 15210 7440 15290 7560
rect 15430 7510 15510 7630
rect 15430 7450 15440 7510
rect 15500 7450 15510 7510
rect 15430 7440 15510 7450
rect 17410 7440 17490 7630
rect 17630 7620 17710 7630
rect 17630 7560 17640 7620
rect 17700 7560 17710 7620
rect 19620 7610 19680 8240
rect 19730 7730 19790 7740
rect 19730 7660 19790 7670
rect 19840 7610 19900 8240
rect 21300 8190 21500 8200
rect 21300 8110 21310 8190
rect 21490 8110 21500 8190
rect 21300 8100 21500 8110
rect 21930 7730 21990 7740
rect 21930 7660 21990 7670
rect 17630 7440 17710 7560
rect 19610 7440 19690 7610
rect 19830 7440 19910 7610
rect 420 7390 620 7400
rect 420 7310 430 7390
rect 610 7310 620 7390
rect 420 7300 620 7310
rect -70 6930 -10 6940
rect -70 6860 -10 6870
rect 2020 6830 2080 7440
rect 2130 6930 2190 6940
rect 2130 6860 2190 6870
rect 2240 6830 2300 7440
rect 2500 7240 2700 7250
rect 2500 7180 2510 7240
rect 2690 7180 2700 7240
rect 2500 7170 2700 7180
rect 3160 7240 3360 7250
rect 3160 7180 3170 7240
rect 3350 7180 3360 7240
rect 3160 7170 3360 7180
rect 3820 7240 4020 7250
rect 3820 7180 3830 7240
rect 4010 7180 4020 7240
rect 3820 7170 4020 7180
rect 2500 7030 2700 7110
rect 3160 7030 3360 7110
rect 3820 7030 4020 7110
rect 4220 6830 4280 7440
rect 4330 6930 4390 6940
rect 4330 6860 4390 6870
rect 4440 6830 4500 7440
rect 4700 7410 6220 7420
rect 4700 7350 4710 7410
rect 6210 7350 6220 7410
rect 4700 7340 6220 7350
rect 4700 7240 4900 7250
rect 4700 7180 4710 7240
rect 4890 7180 4900 7240
rect 4700 7170 4900 7180
rect 5360 7240 5560 7250
rect 5360 7180 5370 7240
rect 5550 7180 5560 7240
rect 5360 7170 5560 7180
rect 6020 7240 6220 7250
rect 6020 7180 6030 7240
rect 6210 7180 6220 7240
rect 6020 7170 6220 7180
rect 4700 7030 4900 7110
rect 5360 7030 5560 7110
rect 6020 7030 6220 7110
rect 6420 6830 6480 7440
rect 6530 6930 6590 6940
rect 6530 6860 6590 6870
rect 6640 6830 6700 7440
rect 6900 7410 8420 7420
rect 6900 7350 6910 7410
rect 8410 7350 8420 7410
rect 6900 7340 8420 7350
rect 6900 7170 7100 7250
rect 7560 7170 7760 7250
rect 8220 7170 8420 7250
rect 6900 7100 7100 7110
rect 6900 7040 6910 7100
rect 7090 7040 7100 7100
rect 6900 7030 7100 7040
rect 7560 7100 7760 7110
rect 7560 7040 7570 7100
rect 7750 7040 7760 7100
rect 7560 7030 7760 7040
rect 8220 7100 8420 7110
rect 8220 7040 8230 7100
rect 8410 7040 8420 7100
rect 8220 7030 8420 7040
rect 8620 6830 8680 7440
rect 8730 6930 8790 6940
rect 8730 6860 8790 6870
rect 8840 6830 8900 7440
rect 9100 7410 10620 7420
rect 9100 7350 9110 7410
rect 10610 7350 10620 7410
rect 9100 7340 10620 7350
rect 9100 7170 9300 7250
rect 9760 7170 9960 7250
rect 10420 7170 10620 7250
rect 9100 7100 9300 7110
rect 9100 7040 9110 7100
rect 9290 7040 9300 7100
rect 9100 7030 9300 7040
rect 9760 7100 9960 7110
rect 9760 7040 9770 7100
rect 9950 7040 9960 7100
rect 9760 7030 9960 7040
rect 10420 7100 10620 7110
rect 10420 7040 10430 7100
rect 10610 7040 10620 7100
rect 10420 7030 10620 7040
rect 10820 6830 10880 7440
rect 10930 6930 10990 6940
rect 10930 6860 10990 6870
rect 11040 6830 11100 7440
rect 11300 7410 12820 7420
rect 11300 7350 11310 7410
rect 12810 7350 12820 7410
rect 11300 7340 12820 7350
rect 11300 7170 11500 7250
rect 11960 7170 12160 7250
rect 12620 7170 12820 7250
rect 11300 7100 11500 7110
rect 11300 7040 11310 7100
rect 11490 7040 11500 7100
rect 11300 7030 11500 7040
rect 11960 7100 12160 7110
rect 11960 7040 11970 7100
rect 12150 7040 12160 7100
rect 11960 7030 12160 7040
rect 12620 7100 12820 7110
rect 12620 7040 12630 7100
rect 12810 7040 12820 7100
rect 12620 7030 12820 7040
rect 13020 6830 13080 7440
rect 13130 6930 13190 6940
rect 13130 6860 13190 6870
rect 13240 6830 13300 7440
rect 13500 7410 15020 7420
rect 13500 7350 13510 7410
rect 15010 7350 15020 7410
rect 13500 7340 15020 7350
rect 13500 7170 13700 7250
rect 14160 7170 14360 7250
rect 14820 7170 15020 7250
rect 13500 7100 13700 7110
rect 13500 7040 13510 7100
rect 13690 7040 13700 7100
rect 13500 7030 13700 7040
rect 14160 7100 14360 7110
rect 14160 7040 14170 7100
rect 14350 7040 14360 7100
rect 14160 7030 14360 7040
rect 14820 7100 15020 7110
rect 14820 7040 14830 7100
rect 15010 7040 15020 7100
rect 14820 7030 15020 7040
rect 15220 6830 15280 7440
rect 15330 6930 15390 6940
rect 15330 6860 15390 6870
rect 15440 6830 15500 7440
rect 15700 7410 17220 7420
rect 15700 7350 15710 7410
rect 17210 7350 17220 7410
rect 15700 7340 17220 7350
rect 15700 7240 15900 7250
rect 15700 7180 15710 7240
rect 15890 7180 15900 7240
rect 15700 7170 15900 7180
rect 16360 7240 16560 7250
rect 16360 7180 16370 7240
rect 16550 7180 16560 7240
rect 16360 7170 16560 7180
rect 17020 7240 17220 7250
rect 17020 7180 17030 7240
rect 17210 7180 17220 7240
rect 17020 7170 17220 7180
rect 15700 7030 15900 7110
rect 16360 7030 16560 7110
rect 17020 7030 17220 7110
rect 17420 6830 17480 7440
rect 17530 6930 17590 6940
rect 17530 6860 17590 6870
rect 17640 6830 17700 7440
rect 17900 7240 18100 7250
rect 17900 7180 17910 7240
rect 18090 7180 18100 7240
rect 17900 7170 18100 7180
rect 18560 7240 18760 7250
rect 18560 7180 18570 7240
rect 18750 7180 18760 7240
rect 18560 7170 18760 7180
rect 19220 7240 19420 7250
rect 19220 7180 19230 7240
rect 19410 7180 19420 7240
rect 19220 7170 19420 7180
rect 17900 7030 18100 7110
rect 18560 7030 18760 7110
rect 19220 7030 19420 7110
rect 2010 6640 2090 6830
rect 2230 6640 2310 6830
rect 4210 6710 4290 6830
rect 4210 6650 4220 6710
rect 4280 6650 4290 6710
rect 4210 6640 4290 6650
rect 4430 6640 4510 6830
rect 6410 6820 6490 6830
rect 6410 6760 6420 6820
rect 6480 6760 6490 6820
rect 6410 6640 6490 6760
rect 6630 6710 6710 6830
rect 6630 6650 6640 6710
rect 6700 6650 6710 6710
rect 6630 6640 6710 6650
rect 8610 6640 8690 6830
rect 8830 6820 8910 6830
rect 8830 6760 8840 6820
rect 8900 6760 8910 6820
rect 8830 6710 8910 6760
rect 8830 6650 8840 6710
rect 8900 6650 8910 6710
rect 8830 6640 8910 6650
rect 10810 6640 10890 6830
rect 11030 6820 11110 6830
rect 11030 6760 11040 6820
rect 11100 6760 11110 6820
rect 11030 6710 11110 6760
rect 11030 6650 11040 6710
rect 11100 6650 11110 6710
rect 11030 6640 11110 6650
rect 13010 6640 13090 6830
rect 13230 6820 13310 6830
rect 13230 6760 13240 6820
rect 13300 6760 13310 6820
rect 13230 6710 13310 6760
rect 13230 6650 13240 6710
rect 13300 6650 13310 6710
rect 13230 6640 13310 6650
rect 15210 6710 15290 6830
rect 15210 6650 15220 6710
rect 15280 6650 15290 6710
rect 15210 6640 15290 6650
rect 15430 6820 15510 6830
rect 15430 6760 15440 6820
rect 15500 6760 15510 6820
rect 15430 6640 15510 6760
rect 17410 6820 17490 6830
rect 17410 6760 17420 6820
rect 17480 6760 17490 6820
rect 17410 6640 17490 6760
rect 17630 6640 17710 6830
rect 19620 6810 19680 7440
rect 19730 6930 19790 6940
rect 19730 6860 19790 6870
rect 19840 6810 19900 7440
rect 21300 7390 21500 7400
rect 21300 7310 21310 7390
rect 21490 7310 21500 7390
rect 21300 7300 21500 7310
rect 21930 6930 21990 6940
rect 21930 6860 21990 6870
rect 19610 6640 19690 6810
rect 19830 6640 19910 6810
rect 420 6590 620 6600
rect 420 6510 430 6590
rect 610 6510 620 6590
rect 420 6500 620 6510
rect -70 6130 -10 6140
rect -70 6060 -10 6070
rect 2020 6030 2080 6640
rect 2130 6130 2190 6140
rect 2130 6060 2190 6070
rect 2240 6030 2300 6640
rect 2500 6370 2700 6450
rect 3160 6370 3360 6450
rect 3820 6370 4020 6450
rect 2500 6300 2700 6310
rect 2500 6240 2510 6300
rect 2690 6240 2700 6300
rect 2500 6230 2700 6240
rect 3160 6300 3360 6310
rect 3160 6240 3170 6300
rect 3350 6240 3360 6300
rect 3160 6230 3360 6240
rect 3820 6300 4020 6310
rect 3820 6240 3830 6300
rect 4010 6240 4020 6300
rect 3820 6230 4020 6240
rect 4220 6030 4280 6640
rect 4330 6130 4390 6140
rect 4330 6060 4390 6070
rect 4440 6030 4500 6640
rect 4700 6610 6220 6620
rect 4700 6550 4710 6610
rect 6210 6550 6220 6610
rect 4700 6540 6220 6550
rect 4700 6370 4900 6450
rect 5360 6370 5560 6450
rect 6020 6370 6220 6450
rect 4700 6300 4900 6310
rect 4700 6240 4710 6300
rect 4890 6240 4900 6300
rect 4700 6230 4900 6240
rect 5360 6300 5560 6310
rect 5360 6240 5370 6300
rect 5550 6240 5560 6300
rect 5360 6230 5560 6240
rect 6020 6300 6220 6310
rect 6020 6240 6030 6300
rect 6210 6240 6220 6300
rect 6020 6230 6220 6240
rect 6420 6030 6480 6640
rect 6530 6130 6590 6140
rect 6530 6060 6590 6070
rect 6640 6030 6700 6640
rect 6900 6610 8420 6620
rect 6900 6550 6910 6610
rect 8410 6550 8420 6610
rect 6900 6540 8420 6550
rect 6900 6440 7100 6450
rect 6900 6380 6910 6440
rect 7090 6380 7100 6440
rect 6900 6370 7100 6380
rect 7560 6440 7760 6450
rect 7560 6380 7570 6440
rect 7750 6380 7760 6440
rect 7560 6370 7760 6380
rect 8220 6440 8420 6450
rect 8220 6380 8230 6440
rect 8410 6380 8420 6440
rect 8220 6370 8420 6380
rect 6900 6230 7100 6310
rect 7560 6230 7760 6310
rect 8220 6230 8420 6310
rect 8620 6030 8680 6640
rect 8730 6130 8790 6140
rect 8730 6060 8790 6070
rect 8840 6030 8900 6640
rect 9100 6610 10620 6620
rect 9100 6550 9110 6610
rect 10610 6550 10620 6610
rect 9100 6540 10620 6550
rect 9100 6440 9300 6450
rect 9100 6380 9110 6440
rect 9290 6380 9300 6440
rect 9100 6370 9300 6380
rect 9760 6440 9960 6450
rect 9760 6380 9770 6440
rect 9950 6380 9960 6440
rect 9760 6370 9960 6380
rect 10420 6440 10620 6450
rect 10420 6380 10430 6440
rect 10610 6380 10620 6440
rect 10420 6370 10620 6380
rect 9100 6230 9300 6310
rect 9760 6230 9960 6310
rect 10420 6230 10620 6310
rect 10820 6030 10880 6640
rect 10930 6130 10990 6140
rect 10930 6060 10990 6070
rect 11040 6030 11100 6640
rect 11300 6610 12820 6620
rect 11300 6550 11310 6610
rect 12810 6550 12820 6610
rect 11300 6540 12820 6550
rect 11300 6440 11500 6450
rect 11300 6380 11310 6440
rect 11490 6380 11500 6440
rect 11300 6370 11500 6380
rect 11960 6440 12160 6450
rect 11960 6380 11970 6440
rect 12150 6380 12160 6440
rect 11960 6370 12160 6380
rect 12620 6440 12820 6450
rect 12620 6380 12630 6440
rect 12810 6380 12820 6440
rect 12620 6370 12820 6380
rect 11300 6230 11500 6310
rect 11960 6230 12160 6310
rect 12620 6230 12820 6310
rect 13020 6030 13080 6640
rect 13130 6130 13190 6140
rect 13130 6060 13190 6070
rect 13240 6030 13300 6640
rect 13500 6610 15020 6620
rect 13500 6550 13510 6610
rect 15010 6550 15020 6610
rect 13500 6540 15020 6550
rect 13500 6440 13700 6450
rect 13500 6380 13510 6440
rect 13690 6380 13700 6440
rect 13500 6370 13700 6380
rect 14160 6440 14360 6450
rect 14160 6380 14170 6440
rect 14350 6380 14360 6440
rect 14160 6370 14360 6380
rect 14820 6440 15020 6450
rect 14820 6380 14830 6440
rect 15010 6380 15020 6440
rect 14820 6370 15020 6380
rect 13500 6230 13700 6310
rect 14160 6230 14360 6310
rect 14820 6230 15020 6310
rect 15220 6030 15280 6640
rect 15330 6130 15390 6140
rect 15330 6060 15390 6070
rect 15440 6030 15500 6640
rect 15700 6610 17220 6620
rect 15700 6550 15710 6610
rect 17210 6550 17220 6610
rect 15700 6540 17220 6550
rect 15700 6370 15900 6450
rect 16360 6370 16560 6450
rect 17020 6370 17220 6450
rect 15700 6300 15900 6310
rect 15700 6240 15710 6300
rect 15890 6240 15900 6300
rect 15700 6230 15900 6240
rect 16360 6300 16560 6310
rect 16360 6240 16370 6300
rect 16550 6240 16560 6300
rect 16360 6230 16560 6240
rect 17020 6300 17220 6310
rect 17020 6240 17030 6300
rect 17210 6240 17220 6300
rect 17020 6230 17220 6240
rect 17420 6030 17480 6640
rect 17530 6130 17590 6140
rect 17530 6060 17590 6070
rect 17640 6030 17700 6640
rect 17900 6370 18100 6450
rect 18560 6370 18760 6450
rect 19220 6370 19420 6450
rect 17900 6300 18100 6310
rect 17900 6240 17910 6300
rect 18090 6240 18100 6300
rect 17900 6230 18100 6240
rect 18560 6300 18760 6310
rect 18560 6240 18570 6300
rect 18750 6240 18760 6300
rect 18560 6230 18760 6240
rect 19220 6300 19420 6310
rect 19220 6240 19230 6300
rect 19410 6240 19420 6300
rect 19220 6230 19420 6240
rect 2010 5840 2090 6030
rect 2230 5910 2310 6030
rect 2230 5850 2240 5910
rect 2300 5850 2310 5910
rect 2230 5840 2310 5850
rect 4210 5840 4290 6030
rect 4430 6020 4510 6030
rect 4430 5960 4440 6020
rect 4500 5960 4510 6020
rect 4430 5910 4510 5960
rect 4430 5850 4440 5910
rect 4500 5850 4510 5910
rect 4430 5840 4510 5850
rect 6410 5910 6490 6030
rect 6410 5850 6420 5910
rect 6480 5850 6490 5910
rect 6410 5840 6490 5850
rect 6630 6020 6710 6030
rect 6630 5960 6640 6020
rect 6700 5960 6710 6020
rect 6630 5840 6710 5960
rect 8610 6020 8690 6030
rect 8610 5960 8620 6020
rect 8680 5960 8690 6020
rect 8610 5910 8690 5960
rect 8610 5850 8620 5910
rect 8680 5850 8690 5910
rect 8610 5840 8690 5850
rect 8830 5840 8910 6030
rect 10810 6020 10890 6030
rect 10810 5960 10820 6020
rect 10880 5960 10890 6020
rect 10810 5910 10890 5960
rect 10810 5850 10820 5910
rect 10880 5850 10890 5910
rect 10810 5840 10890 5850
rect 11030 5840 11110 6030
rect 13010 6020 13090 6030
rect 13010 5960 13020 6020
rect 13080 5960 13090 6020
rect 13010 5910 13090 5960
rect 13010 5850 13020 5910
rect 13080 5850 13090 5910
rect 13010 5840 13090 5850
rect 13230 5840 13310 6030
rect 15210 6020 15290 6030
rect 15210 5960 15220 6020
rect 15280 5960 15290 6020
rect 15210 5840 15290 5960
rect 15430 5910 15510 6030
rect 15430 5850 15440 5910
rect 15500 5850 15510 5910
rect 15430 5840 15510 5850
rect 17410 5840 17490 6030
rect 17630 6020 17710 6030
rect 17630 5960 17640 6020
rect 17700 5960 17710 6020
rect 19620 6010 19680 6640
rect 19730 6130 19790 6140
rect 19730 6060 19790 6070
rect 19840 6010 19900 6640
rect 21300 6590 21500 6600
rect 21300 6510 21310 6590
rect 21490 6510 21500 6590
rect 21300 6500 21500 6510
rect 21930 6130 21990 6140
rect 21930 6060 21990 6070
rect 17630 5910 17710 5960
rect 17630 5850 17640 5910
rect 17700 5850 17710 5910
rect 17630 5840 17710 5850
rect 19610 5840 19690 6010
rect 19830 6000 19910 6010
rect 19830 5940 19840 6000
rect 19900 5940 19910 6000
rect 19830 5840 19910 5940
rect -70 5330 -10 5340
rect -70 5260 -10 5270
rect 2020 5230 2080 5840
rect 2130 5330 2190 5340
rect 2130 5260 2190 5270
rect 2240 5230 2300 5840
rect 2500 5810 4020 5820
rect 2500 5750 2510 5810
rect 4010 5750 4020 5810
rect 2500 5740 4020 5750
rect 2500 5640 2700 5650
rect 2500 5580 2510 5640
rect 2690 5580 2700 5640
rect 2500 5570 2700 5580
rect 3160 5640 3360 5650
rect 3160 5580 3170 5640
rect 3350 5580 3360 5640
rect 3160 5570 3360 5580
rect 3820 5640 4020 5650
rect 3820 5580 3830 5640
rect 4010 5580 4020 5640
rect 3820 5570 4020 5580
rect 2500 5430 2700 5510
rect 3160 5430 3360 5510
rect 3820 5430 4020 5510
rect 4220 5230 4280 5840
rect 4330 5330 4390 5340
rect 4330 5260 4390 5270
rect 4440 5230 4500 5840
rect 4700 5810 6220 5820
rect 4700 5750 4710 5810
rect 6210 5750 6220 5810
rect 4700 5740 6220 5750
rect 4700 5640 4900 5650
rect 4700 5580 4710 5640
rect 4890 5580 4900 5640
rect 4700 5570 4900 5580
rect 5360 5640 5560 5650
rect 5360 5580 5370 5640
rect 5550 5580 5560 5640
rect 5360 5570 5560 5580
rect 6020 5640 6220 5650
rect 6020 5580 6030 5640
rect 6210 5580 6220 5640
rect 6020 5570 6220 5580
rect 4700 5430 4900 5510
rect 5360 5430 5560 5510
rect 6020 5430 6220 5510
rect 6420 5230 6480 5840
rect 6530 5330 6590 5340
rect 6530 5260 6590 5270
rect 6640 5230 6700 5840
rect 6900 5810 8420 5820
rect 6900 5750 6910 5810
rect 8410 5750 8420 5810
rect 6900 5740 8420 5750
rect 6900 5570 7100 5650
rect 7560 5570 7760 5650
rect 8220 5570 8420 5650
rect 6900 5500 7100 5510
rect 6900 5440 6910 5500
rect 7090 5440 7100 5500
rect 6900 5430 7100 5440
rect 7560 5500 7760 5510
rect 7560 5440 7570 5500
rect 7750 5440 7760 5500
rect 7560 5430 7760 5440
rect 8220 5500 8420 5510
rect 8220 5440 8230 5500
rect 8410 5440 8420 5500
rect 8220 5430 8420 5440
rect 8620 5230 8680 5840
rect 8730 5330 8790 5340
rect 8730 5260 8790 5270
rect 8840 5230 8900 5840
rect 9100 5810 10620 5820
rect 9100 5750 9110 5810
rect 10610 5750 10620 5810
rect 9100 5740 10620 5750
rect 9100 5570 9300 5650
rect 9760 5570 9960 5650
rect 10420 5570 10620 5650
rect 9100 5500 9300 5510
rect 9100 5440 9110 5500
rect 9290 5440 9300 5500
rect 9100 5430 9300 5440
rect 9760 5500 9960 5510
rect 9760 5440 9770 5500
rect 9950 5440 9960 5500
rect 9760 5430 9960 5440
rect 10420 5500 10620 5510
rect 10420 5440 10430 5500
rect 10610 5440 10620 5500
rect 10420 5430 10620 5440
rect 10820 5230 10880 5840
rect 10930 5330 10990 5340
rect 10930 5260 10990 5270
rect 11040 5230 11100 5840
rect 11300 5810 12820 5820
rect 11300 5750 11310 5810
rect 12810 5750 12820 5810
rect 11300 5740 12820 5750
rect 11300 5570 11500 5650
rect 11960 5570 12160 5650
rect 12620 5570 12820 5650
rect 11300 5500 11500 5510
rect 11300 5440 11310 5500
rect 11490 5440 11500 5500
rect 11300 5430 11500 5440
rect 11960 5500 12160 5510
rect 11960 5440 11970 5500
rect 12150 5440 12160 5500
rect 11960 5430 12160 5440
rect 12620 5500 12820 5510
rect 12620 5440 12630 5500
rect 12810 5440 12820 5500
rect 12620 5430 12820 5440
rect 13020 5230 13080 5840
rect 13130 5330 13190 5340
rect 13130 5260 13190 5270
rect 13240 5230 13300 5840
rect 13500 5810 15020 5820
rect 13500 5750 13510 5810
rect 15010 5750 15020 5810
rect 13500 5740 15020 5750
rect 13500 5570 13700 5650
rect 14160 5570 14360 5650
rect 14820 5570 15020 5650
rect 13500 5500 13700 5510
rect 13500 5440 13510 5500
rect 13690 5440 13700 5500
rect 13500 5430 13700 5440
rect 14160 5500 14360 5510
rect 14160 5440 14170 5500
rect 14350 5440 14360 5500
rect 14160 5430 14360 5440
rect 14820 5500 15020 5510
rect 14820 5440 14830 5500
rect 15010 5440 15020 5500
rect 14820 5430 15020 5440
rect 15220 5230 15280 5840
rect 15330 5330 15390 5340
rect 15330 5260 15390 5270
rect 15440 5230 15500 5840
rect 15700 5810 17220 5820
rect 15700 5750 15710 5810
rect 17210 5750 17220 5810
rect 15700 5740 17220 5750
rect 15700 5640 15900 5650
rect 15700 5580 15710 5640
rect 15890 5580 15900 5640
rect 15700 5570 15900 5580
rect 16360 5640 16560 5650
rect 16360 5580 16370 5640
rect 16550 5580 16560 5640
rect 16360 5570 16560 5580
rect 17020 5640 17220 5650
rect 17020 5580 17030 5640
rect 17210 5580 17220 5640
rect 17020 5570 17220 5580
rect 15700 5430 15900 5510
rect 16360 5430 16560 5510
rect 17020 5430 17220 5510
rect 17420 5230 17480 5840
rect 17530 5330 17590 5340
rect 17530 5260 17590 5270
rect 17640 5230 17700 5840
rect 17900 5810 19420 5820
rect 17900 5750 17910 5810
rect 19410 5750 19420 5810
rect 17900 5740 19420 5750
rect 17900 5640 18100 5650
rect 17900 5580 17910 5640
rect 18090 5580 18100 5640
rect 17900 5570 18100 5580
rect 18560 5640 18760 5650
rect 18560 5580 18570 5640
rect 18750 5580 18760 5640
rect 18560 5570 18760 5580
rect 19220 5640 19420 5650
rect 19220 5580 19230 5640
rect 19410 5580 19420 5640
rect 19220 5570 19420 5580
rect 17900 5430 18100 5510
rect 18560 5430 18760 5510
rect 19220 5430 19420 5510
rect 2010 5110 2090 5230
rect 2010 5050 2020 5110
rect 2080 5050 2090 5110
rect 2010 5040 2090 5050
rect 2230 5040 2310 5230
rect 4210 5220 4290 5230
rect 4210 5160 4220 5220
rect 4280 5160 4290 5220
rect 4210 5110 4290 5160
rect 4210 5050 4220 5110
rect 4280 5050 4290 5110
rect 4210 5040 4290 5050
rect 4430 5040 4510 5230
rect 6410 5220 6490 5230
rect 6410 5160 6420 5220
rect 6480 5160 6490 5220
rect 6410 5040 6490 5160
rect 6630 5110 6710 5230
rect 6630 5050 6640 5110
rect 6700 5050 6710 5110
rect 6630 5040 6710 5050
rect 8610 5040 8690 5230
rect 8830 5220 8910 5230
rect 8830 5160 8840 5220
rect 8900 5160 8910 5220
rect 8830 5110 8910 5160
rect 8830 5050 8840 5110
rect 8900 5050 8910 5110
rect 8830 5040 8910 5050
rect 10810 5040 10890 5230
rect 11030 5220 11110 5230
rect 11030 5160 11040 5220
rect 11100 5160 11110 5220
rect 11030 5110 11110 5160
rect 11030 5050 11040 5110
rect 11100 5050 11110 5110
rect 11030 5040 11110 5050
rect 13010 5040 13090 5230
rect 13230 5220 13310 5230
rect 13230 5160 13240 5220
rect 13300 5160 13310 5220
rect 13230 5110 13310 5160
rect 13230 5050 13240 5110
rect 13300 5050 13310 5110
rect 13230 5040 13310 5050
rect 15210 5110 15290 5230
rect 15210 5050 15220 5110
rect 15280 5050 15290 5110
rect 15210 5040 15290 5050
rect 15430 5220 15510 5230
rect 15430 5160 15440 5220
rect 15500 5160 15510 5220
rect 15430 5040 15510 5160
rect 17410 5220 17490 5230
rect 17410 5160 17420 5220
rect 17480 5160 17490 5220
rect 17410 5110 17490 5160
rect 17410 5050 17420 5110
rect 17480 5050 17490 5110
rect 17410 5040 17490 5050
rect 17630 5040 17710 5230
rect 19620 5210 19680 5840
rect 19730 5330 19790 5340
rect 19730 5260 19790 5270
rect 19840 5210 19900 5840
rect 21930 5330 21990 5340
rect 21930 5260 21990 5270
rect 19610 5200 19690 5210
rect 19610 5140 19620 5200
rect 19680 5140 19690 5200
rect 19610 5040 19690 5140
rect 19830 5040 19910 5210
rect 2020 4830 2080 5040
rect 2240 4830 2300 5040
rect 2500 5010 4020 5020
rect 2500 4950 2510 5010
rect 4010 4950 4020 5010
rect 2500 4940 4020 4950
rect 4220 4830 4280 5040
rect 4440 4830 4500 5040
rect 4700 5010 6220 5020
rect 4700 4950 4710 5010
rect 6210 4950 6220 5010
rect 4700 4940 6220 4950
rect 6420 4830 6480 5040
rect 6640 4830 6700 5040
rect 6900 5010 8420 5020
rect 6900 4950 6910 5010
rect 8410 4950 8420 5010
rect 6900 4940 8420 4950
rect 8620 4830 8680 5040
rect 8840 4830 8900 5040
rect 9100 5010 10620 5020
rect 9100 4950 9110 5010
rect 10610 4950 10620 5010
rect 9100 4940 10620 4950
rect 10820 4830 10880 5040
rect 11040 4830 11100 5040
rect 11300 5010 12820 5020
rect 11300 4950 11310 5010
rect 12810 4950 12820 5010
rect 11300 4940 12820 4950
rect 13020 4830 13080 5040
rect 13240 4830 13300 5040
rect 13500 5010 15020 5020
rect 13500 4950 13510 5010
rect 15010 4950 15020 5010
rect 13500 4940 15020 4950
rect 15220 4830 15280 5040
rect 15440 4830 15500 5040
rect 15700 5010 17220 5020
rect 15700 4950 15710 5010
rect 17210 4950 17220 5010
rect 15700 4940 17220 4950
rect 17420 4830 17480 5040
rect 17640 4830 17700 5040
rect 17900 5010 19420 5020
rect 17900 4950 17910 5010
rect 19410 4950 19420 5010
rect 17900 4940 19420 4950
rect 19620 4830 19680 5040
rect 19840 4830 19900 5040
rect 31560 3730 31740 3740
rect 31560 3550 31570 3730
rect 31730 3550 31740 3730
rect 31560 3540 31740 3550
rect 1160 3330 1340 3340
rect 1160 3150 1170 3330
rect 1330 3150 1340 3330
rect 1160 3140 1340 3150
rect 2760 3330 2940 3340
rect 2760 3150 2770 3330
rect 2930 3150 2940 3330
rect 2760 3140 2940 3150
rect 4360 3330 4540 3340
rect 4360 3150 4370 3330
rect 4530 3150 4540 3330
rect 4360 3140 4540 3150
rect 5960 3330 6140 3340
rect 5960 3150 5970 3330
rect 6130 3150 6140 3330
rect 5960 3140 6140 3150
rect 7560 3330 7740 3340
rect 7560 3150 7570 3330
rect 7730 3150 7740 3330
rect 7560 3140 7740 3150
rect 9160 3330 9340 3340
rect 9160 3150 9170 3330
rect 9330 3150 9340 3330
rect 9160 3140 9340 3150
rect 1200 690 1300 3140
rect 2100 2230 2240 2240
rect 2100 2070 2110 2230
rect 2230 2070 2240 2230
rect 2100 1970 2240 2070
rect 2100 1290 2110 1970
rect 2230 1290 2240 1970
rect 1420 1140 1520 1160
rect 1400 1130 1540 1140
rect 1400 1010 1410 1130
rect 1530 1010 1540 1130
rect 1400 1000 1540 1010
rect 1180 680 1320 690
rect 1180 560 1190 680
rect 1310 560 1320 680
rect 1180 550 1320 560
rect 1200 -1110 1300 550
rect 1420 -660 1520 1000
rect 2100 430 2240 1290
rect 2800 690 2900 3140
rect 3700 2230 3840 2240
rect 3700 2070 3710 2230
rect 3830 2070 3840 2230
rect 3700 1970 3840 2070
rect 3700 1290 3710 1970
rect 3830 1290 3840 1970
rect 3020 1140 3120 1160
rect 3000 1130 3140 1140
rect 3000 1010 3010 1130
rect 3130 1010 3140 1130
rect 3000 1000 3140 1010
rect 2780 680 2920 690
rect 2780 560 2790 680
rect 2910 560 2920 680
rect 2780 550 2920 560
rect 2100 270 2110 430
rect 2230 270 2240 430
rect 2100 170 2240 270
rect 2100 -510 2110 170
rect 2230 -510 2240 170
rect 1400 -670 1540 -660
rect 1400 -790 1410 -670
rect 1530 -790 1540 -670
rect 1400 -800 1540 -790
rect 1180 -1120 1320 -1110
rect 1180 -1240 1190 -1120
rect 1310 -1240 1320 -1120
rect 1180 -1250 1320 -1240
rect 1200 -2910 1300 -1250
rect 1420 -2460 1520 -800
rect 2100 -1370 2240 -510
rect 2800 -1110 2900 550
rect 3020 -660 3120 1000
rect 3700 430 3840 1290
rect 4400 690 4500 3140
rect 5300 2230 5440 2240
rect 5300 2070 5310 2230
rect 5430 2070 5440 2230
rect 5300 1970 5440 2070
rect 5300 1290 5310 1970
rect 5430 1290 5440 1970
rect 4620 1140 4720 1160
rect 4600 1130 4740 1140
rect 4600 1010 4610 1130
rect 4730 1010 4740 1130
rect 4600 1000 4740 1010
rect 4380 680 4520 690
rect 4380 560 4390 680
rect 4510 560 4520 680
rect 4380 550 4520 560
rect 3700 270 3710 430
rect 3830 270 3840 430
rect 3700 170 3840 270
rect 3700 -510 3710 170
rect 3830 -510 3840 170
rect 3000 -670 3140 -660
rect 3000 -790 3010 -670
rect 3130 -790 3140 -670
rect 3000 -800 3140 -790
rect 2780 -1120 2920 -1110
rect 2780 -1240 2790 -1120
rect 2910 -1240 2920 -1120
rect 2780 -1250 2920 -1240
rect 2100 -1530 2110 -1370
rect 2230 -1530 2240 -1370
rect 2100 -1630 2240 -1530
rect 2100 -2310 2110 -1630
rect 2230 -2310 2240 -1630
rect 1400 -2470 1540 -2460
rect 1400 -2590 1410 -2470
rect 1530 -2590 1540 -2470
rect 1400 -2600 1540 -2590
rect 1180 -2920 1320 -2910
rect 1180 -3040 1190 -2920
rect 1310 -3040 1320 -2920
rect 1180 -3050 1320 -3040
rect 1200 -4710 1300 -3050
rect 1420 -4260 1520 -2600
rect 2100 -3170 2240 -2310
rect 2800 -2910 2900 -1250
rect 3020 -2460 3120 -800
rect 3700 -1370 3840 -510
rect 4400 -1110 4500 550
rect 4620 -660 4720 1000
rect 5300 430 5440 1290
rect 6000 690 6100 3140
rect 6900 2230 7040 2240
rect 6900 2070 6910 2230
rect 7030 2070 7040 2230
rect 6900 1970 7040 2070
rect 6900 1290 6910 1970
rect 7030 1290 7040 1970
rect 6220 1140 6320 1160
rect 6200 1130 6340 1140
rect 6200 1010 6210 1130
rect 6330 1010 6340 1130
rect 6200 1000 6340 1010
rect 5980 680 6120 690
rect 5980 560 5990 680
rect 6110 560 6120 680
rect 5980 550 6120 560
rect 5300 270 5310 430
rect 5430 270 5440 430
rect 5300 170 5440 270
rect 5300 -510 5310 170
rect 5430 -510 5440 170
rect 4600 -670 4740 -660
rect 4600 -790 4610 -670
rect 4730 -790 4740 -670
rect 4600 -800 4740 -790
rect 4380 -1120 4520 -1110
rect 4380 -1240 4390 -1120
rect 4510 -1240 4520 -1120
rect 4380 -1250 4520 -1240
rect 3700 -1530 3710 -1370
rect 3830 -1530 3840 -1370
rect 3700 -1630 3840 -1530
rect 3700 -2310 3710 -1630
rect 3830 -2310 3840 -1630
rect 3000 -2470 3140 -2460
rect 3000 -2590 3010 -2470
rect 3130 -2590 3140 -2470
rect 3000 -2600 3140 -2590
rect 2780 -2920 2920 -2910
rect 2780 -3040 2790 -2920
rect 2910 -3040 2920 -2920
rect 2780 -3050 2920 -3040
rect 2100 -3330 2110 -3170
rect 2230 -3330 2240 -3170
rect 2100 -3430 2240 -3330
rect 2100 -4110 2110 -3430
rect 2230 -4110 2240 -3430
rect 2100 -4120 2240 -4110
rect 1400 -4270 1540 -4260
rect 1400 -4390 1410 -4270
rect 1530 -4390 1540 -4270
rect 1400 -4400 1540 -4390
rect 1420 -4420 1520 -4400
rect 2800 -4710 2900 -3050
rect 3020 -4260 3120 -2600
rect 3700 -3170 3840 -2310
rect 4400 -2910 4500 -1250
rect 4620 -2460 4720 -800
rect 5300 -1370 5440 -510
rect 6000 -1110 6100 550
rect 6220 -660 6320 1000
rect 6900 430 7040 1290
rect 7600 690 7700 3140
rect 8500 2230 8640 2240
rect 8500 2070 8510 2230
rect 8630 2070 8640 2230
rect 8500 1970 8640 2070
rect 8500 1290 8510 1970
rect 8630 1290 8640 1970
rect 7820 1140 7920 1160
rect 7800 1130 7940 1140
rect 7800 1010 7810 1130
rect 7930 1010 7940 1130
rect 7800 1000 7940 1010
rect 7580 680 7720 690
rect 7580 560 7590 680
rect 7710 560 7720 680
rect 7580 550 7720 560
rect 6900 270 6910 430
rect 7030 270 7040 430
rect 6900 170 7040 270
rect 6900 -510 6910 170
rect 7030 -510 7040 170
rect 6200 -670 6340 -660
rect 6200 -790 6210 -670
rect 6330 -790 6340 -670
rect 6200 -800 6340 -790
rect 5980 -1120 6120 -1110
rect 5980 -1240 5990 -1120
rect 6110 -1240 6120 -1120
rect 5980 -1250 6120 -1240
rect 5300 -1530 5310 -1370
rect 5430 -1530 5440 -1370
rect 5300 -1630 5440 -1530
rect 5300 -2310 5310 -1630
rect 5430 -2310 5440 -1630
rect 4600 -2470 4740 -2460
rect 4600 -2590 4610 -2470
rect 4730 -2590 4740 -2470
rect 4600 -2600 4740 -2590
rect 4380 -2920 4520 -2910
rect 4380 -3040 4390 -2920
rect 4510 -3040 4520 -2920
rect 4380 -3050 4520 -3040
rect 3700 -3330 3710 -3170
rect 3830 -3330 3840 -3170
rect 3700 -3430 3840 -3330
rect 3700 -4110 3710 -3430
rect 3830 -4110 3840 -3430
rect 3700 -4120 3840 -4110
rect 3000 -4270 3140 -4260
rect 3000 -4390 3010 -4270
rect 3130 -4390 3140 -4270
rect 3000 -4400 3140 -4390
rect 3020 -4420 3120 -4400
rect 4400 -4710 4500 -3050
rect 4620 -4260 4720 -2600
rect 5300 -3170 5440 -2310
rect 6000 -2910 6100 -1250
rect 6220 -2460 6320 -800
rect 6900 -1370 7040 -510
rect 7600 -1110 7700 550
rect 7820 -660 7920 1000
rect 8500 430 8640 1290
rect 9200 690 9300 3140
rect 11690 2750 11850 2760
rect 11690 2600 11700 2750
rect 11840 2600 11850 2750
rect 11690 2590 11850 2600
rect 10990 2520 11150 2530
rect 10990 2380 11000 2520
rect 11140 2380 11150 2520
rect 10990 2370 11150 2380
rect 10100 2230 10240 2240
rect 10100 2070 10110 2230
rect 10230 2070 10240 2230
rect 10100 1970 10240 2070
rect 10100 1290 10110 1970
rect 10230 1290 10240 1970
rect 11020 1940 11120 2370
rect 11700 2230 11840 2590
rect 12590 2520 12750 2530
rect 12590 2380 12600 2520
rect 12740 2380 12750 2520
rect 12590 2370 12750 2380
rect 13970 2520 14130 2530
rect 13970 2380 13980 2520
rect 14120 2380 14130 2520
rect 13970 2370 14130 2380
rect 11700 2070 11710 2230
rect 11830 2070 11840 2230
rect 11020 1930 11160 1940
rect 11020 1310 11030 1930
rect 11150 1310 11160 1930
rect 11020 1300 11160 1310
rect 9420 1140 9520 1160
rect 9400 1130 9540 1140
rect 9400 1010 9410 1130
rect 9530 1010 9540 1130
rect 9400 1000 9540 1010
rect 9180 680 9320 690
rect 9180 560 9190 680
rect 9310 560 9320 680
rect 9180 550 9320 560
rect 8500 270 8510 430
rect 8630 270 8640 430
rect 8500 170 8640 270
rect 8500 -510 8510 170
rect 8630 -510 8640 170
rect 7800 -670 7940 -660
rect 7800 -790 7810 -670
rect 7930 -790 7940 -670
rect 7800 -800 7940 -790
rect 7580 -1120 7720 -1110
rect 7580 -1240 7590 -1120
rect 7710 -1240 7720 -1120
rect 7580 -1250 7720 -1240
rect 6900 -1530 6910 -1370
rect 7030 -1530 7040 -1370
rect 6900 -1630 7040 -1530
rect 6900 -2310 6910 -1630
rect 7030 -2310 7040 -1630
rect 6200 -2470 6340 -2460
rect 6200 -2590 6210 -2470
rect 6330 -2590 6340 -2470
rect 6200 -2600 6340 -2590
rect 5980 -2920 6120 -2910
rect 5980 -3040 5990 -2920
rect 6110 -3040 6120 -2920
rect 5980 -3050 6120 -3040
rect 5300 -3330 5310 -3170
rect 5430 -3330 5440 -3170
rect 5300 -3430 5440 -3330
rect 5300 -4110 5310 -3430
rect 5430 -4110 5440 -3430
rect 5300 -4120 5440 -4110
rect 4600 -4270 4740 -4260
rect 4600 -4390 4610 -4270
rect 4730 -4390 4740 -4270
rect 4600 -4400 4740 -4390
rect 4620 -4420 4720 -4400
rect 6000 -4710 6100 -3050
rect 6220 -4260 6320 -2600
rect 6900 -3170 7040 -2310
rect 7600 -2910 7700 -1250
rect 7820 -2460 7920 -800
rect 8500 -1370 8640 -510
rect 9200 -1110 9300 550
rect 9420 -660 9520 1000
rect 10100 430 10240 1290
rect 11700 1220 11840 2070
rect 12620 1940 12720 2370
rect 13300 2230 13440 2240
rect 13300 2070 13310 2230
rect 13430 2070 13440 2230
rect 12600 1930 12740 1940
rect 12600 1310 12610 1930
rect 12730 1310 12740 1930
rect 12600 1300 12740 1310
rect 11240 1210 11840 1220
rect 11240 1050 11250 1210
rect 11670 1050 11840 1210
rect 11240 1040 11840 1050
rect 10100 270 10110 430
rect 10230 270 10240 430
rect 10100 170 10240 270
rect 10100 -510 10110 170
rect 10230 -510 10240 170
rect 9400 -670 9540 -660
rect 9400 -790 9410 -670
rect 9530 -790 9540 -670
rect 9400 -800 9540 -790
rect 9180 -1120 9320 -1110
rect 9180 -1240 9190 -1120
rect 9310 -1240 9320 -1120
rect 9180 -1250 9320 -1240
rect 8500 -1530 8510 -1370
rect 8630 -1530 8640 -1370
rect 8500 -1630 8640 -1530
rect 8500 -2310 8510 -1630
rect 8630 -2310 8640 -1630
rect 7800 -2470 7940 -2460
rect 7800 -2590 7810 -2470
rect 7930 -2590 7940 -2470
rect 7800 -2600 7940 -2590
rect 7580 -2920 7720 -2910
rect 7580 -3040 7590 -2920
rect 7710 -3040 7720 -2920
rect 7580 -3050 7720 -3040
rect 6900 -3330 6910 -3170
rect 7030 -3330 7040 -3170
rect 6900 -3430 7040 -3330
rect 6900 -4110 6910 -3430
rect 7030 -4110 7040 -3430
rect 6900 -4120 7040 -4110
rect 6200 -4270 6340 -4260
rect 6200 -4390 6210 -4270
rect 6330 -4390 6340 -4270
rect 6200 -4400 6340 -4390
rect 6220 -4420 6320 -4400
rect 7600 -4710 7700 -3050
rect 7820 -4260 7920 -2600
rect 8500 -3170 8640 -2310
rect 9200 -2910 9300 -1250
rect 9420 -2460 9520 -800
rect 10100 -1370 10240 -510
rect 11700 430 11840 1040
rect 12380 870 12520 880
rect 12380 750 12390 870
rect 12510 750 12520 870
rect 12380 740 12520 750
rect 11700 270 11710 430
rect 11830 270 11840 430
rect 11700 170 11840 270
rect 11700 -580 11710 170
rect 11260 -590 11710 -580
rect 11830 -580 11840 170
rect 11830 -590 12280 -580
rect 11260 -750 11270 -590
rect 12270 -750 12280 -590
rect 12400 -660 12500 740
rect 11260 -760 12280 -750
rect 12380 -670 12520 -660
rect 10100 -1530 10110 -1370
rect 10230 -1530 10240 -1370
rect 10100 -1630 10240 -1530
rect 10100 -2310 10110 -1630
rect 10230 -2310 10240 -1630
rect 9400 -2470 9540 -2460
rect 9400 -2590 9410 -2470
rect 9530 -2590 9540 -2470
rect 9400 -2600 9540 -2590
rect 9180 -2920 9320 -2910
rect 9180 -3040 9190 -2920
rect 9310 -3040 9320 -2920
rect 9180 -3050 9320 -3040
rect 8500 -3330 8510 -3170
rect 8630 -3330 8640 -3170
rect 8500 -3430 8640 -3330
rect 8500 -4110 8510 -3430
rect 8630 -4110 8640 -3430
rect 8500 -4120 8640 -4110
rect 7800 -4270 7940 -4260
rect 7800 -4390 7810 -4270
rect 7930 -4390 7940 -4270
rect 7800 -4400 7940 -4390
rect 7820 -4420 7920 -4400
rect 9200 -4710 9300 -3050
rect 9420 -4260 9520 -2600
rect 10100 -3170 10240 -2310
rect 10100 -3330 10110 -3170
rect 10230 -3330 10240 -3170
rect 10100 -3430 10240 -3330
rect 10100 -4110 10110 -3430
rect 10230 -4110 10240 -3430
rect 10100 -4120 10240 -4110
rect 10800 -1210 11000 -1200
rect 10800 -1270 10810 -1210
rect 10990 -1270 11000 -1210
rect 10800 -1280 11000 -1270
rect 9400 -4270 9540 -4260
rect 9400 -4390 9410 -4270
rect 9530 -4390 9540 -4270
rect 9400 -4400 9540 -4390
rect 9420 -4420 9520 -4400
rect 1180 -4720 1320 -4710
rect 1180 -4840 1190 -4720
rect 1310 -4840 1320 -4720
rect 1180 -4850 1320 -4840
rect 2780 -4720 2920 -4710
rect 2780 -4840 2790 -4720
rect 2910 -4840 2920 -4720
rect 2780 -4850 2920 -4840
rect 4380 -4720 4520 -4710
rect 4380 -4840 4390 -4720
rect 4510 -4840 4520 -4720
rect 4380 -4850 4520 -4840
rect 5980 -4720 6120 -4710
rect 5980 -4840 5990 -4720
rect 6110 -4840 6120 -4720
rect 5980 -4850 6120 -4840
rect 7580 -4720 7720 -4710
rect 7580 -4840 7590 -4720
rect 7710 -4840 7720 -4720
rect 7580 -4850 7720 -4840
rect 9180 -4720 9320 -4710
rect 9180 -4840 9190 -4720
rect 9310 -4840 9320 -4720
rect 9180 -4850 9320 -4840
rect 1200 -4860 1300 -4850
rect 2800 -4880 2900 -4850
rect 4400 -4880 4500 -4850
rect 6000 -4880 6100 -4850
rect 7600 -4880 7700 -4850
rect 9200 -4880 9300 -4850
rect 10800 -5120 10900 -1280
rect 11700 -1370 11840 -760
rect 12380 -1050 12390 -670
rect 12510 -1050 12520 -670
rect 12380 -1060 12520 -1050
rect 12620 -920 12720 1300
rect 13300 430 13440 2070
rect 14000 1940 14100 2370
rect 13980 1930 14120 1940
rect 13980 1310 13990 1930
rect 14110 1310 14120 1930
rect 13980 1300 14120 1310
rect 13300 270 13310 430
rect 13430 270 13440 430
rect 13300 170 13440 270
rect 13300 -510 13310 170
rect 13430 -510 13440 170
rect 12620 -930 12760 -920
rect 11700 -1530 11710 -1370
rect 11830 -1530 11840 -1370
rect 11700 -1630 11840 -1530
rect 11700 -2310 11710 -1630
rect 11830 -2310 11840 -1630
rect 11020 -2910 11120 -2900
rect 11000 -2920 11140 -2910
rect 11000 -3040 11010 -2920
rect 11130 -3040 11140 -2920
rect 11000 -3050 11140 -3040
rect 11020 -4750 11120 -3050
rect 11700 -3170 11840 -2310
rect 12400 -2720 12500 -1060
rect 12620 -1070 12630 -930
rect 12750 -1070 12760 -930
rect 12620 -1100 12760 -1070
rect 13300 -1370 13440 -510
rect 14000 -920 14100 1300
rect 13960 -930 14100 -920
rect 13960 -1070 13970 -930
rect 14090 -1070 14100 -930
rect 13960 -1100 14100 -1070
rect 13300 -1530 13310 -1370
rect 13430 -1530 13440 -1370
rect 13300 -1630 13440 -1530
rect 13300 -2310 13310 -1630
rect 13430 -2310 13440 -1630
rect 12380 -2730 12520 -2720
rect 12380 -2850 12390 -2730
rect 12510 -2850 12520 -2730
rect 12380 -2860 12520 -2850
rect 11700 -3330 11710 -3170
rect 11830 -3330 11840 -3170
rect 11700 -3430 11840 -3330
rect 11700 -4110 11710 -3430
rect 11830 -4110 11840 -3430
rect 11700 -4120 11840 -4110
rect 12400 -4520 12500 -2860
rect 13300 -3170 13440 -2310
rect 14220 -2910 14320 2680
rect 16500 2230 16640 2240
rect 16500 2070 16510 2230
rect 16630 2070 16640 2230
rect 14900 1960 15040 1990
rect 14900 1300 14910 1960
rect 15030 1300 15040 1960
rect 14900 1220 15040 1300
rect 16500 1970 16640 2070
rect 16500 1290 16510 1970
rect 16630 1290 16640 1970
rect 18100 2230 18240 2240
rect 18100 2070 18110 2230
rect 18230 2070 18240 2230
rect 18100 1970 18240 2070
rect 18100 1290 18110 1970
rect 18230 1290 18240 1970
rect 19700 2230 19840 2240
rect 19700 2070 19710 2230
rect 19830 2070 19840 2230
rect 19700 1970 19840 2070
rect 19700 1290 19710 1970
rect 19830 1290 19840 1970
rect 21300 2230 21440 2240
rect 21300 2070 21310 2230
rect 21430 2070 21440 2230
rect 21300 1970 21440 2070
rect 21300 1290 21310 1970
rect 21430 1290 21440 1970
rect 22900 2230 23040 2240
rect 22900 2070 22910 2230
rect 23030 2070 23040 2230
rect 22900 1970 23040 2070
rect 22900 1290 22910 1970
rect 23030 1290 23040 1970
rect 24500 2230 24640 2240
rect 24500 2070 24510 2230
rect 24630 2070 24640 2230
rect 24500 1970 24640 2070
rect 24500 1290 24510 1970
rect 24630 1290 24640 1970
rect 26100 2230 26240 2240
rect 26100 2070 26110 2230
rect 26230 2070 26240 2230
rect 26100 1970 26240 2070
rect 26100 1290 26110 1970
rect 26230 1290 26240 1970
rect 27700 2230 27840 2240
rect 27700 2050 27710 2230
rect 27830 2050 27840 2230
rect 27700 1970 27840 2050
rect 27700 1290 27710 1970
rect 27830 1290 27840 1970
rect 29300 2230 29440 2240
rect 29300 2050 29310 2230
rect 29430 2050 29440 2230
rect 29300 1970 29440 2050
rect 29300 1290 29310 1970
rect 29430 1290 29440 1970
rect 15600 1140 15700 1290
rect 15590 1130 15710 1140
rect 15590 1010 15600 1130
rect 15700 1010 15710 1130
rect 15590 1000 15710 1010
rect 14900 170 15040 440
rect 14900 -580 14910 170
rect 14460 -590 14910 -580
rect 15030 -580 15040 170
rect 15030 -590 15480 -580
rect 14460 -750 14470 -590
rect 15470 -750 15480 -590
rect 15600 -660 15700 1000
rect 15820 690 15920 1290
rect 15810 680 15930 690
rect 15810 560 15820 680
rect 15920 560 15930 680
rect 15810 550 15930 560
rect 14460 -760 15480 -750
rect 15590 -670 15710 -660
rect 14900 -1370 15040 -1360
rect 14900 -1530 14910 -1370
rect 15030 -1530 15040 -1370
rect 14900 -1630 15040 -1530
rect 15240 -1370 15380 -760
rect 15590 -790 15600 -670
rect 15700 -790 15710 -670
rect 15590 -800 15710 -790
rect 15240 -1530 15250 -1370
rect 15370 -1530 15380 -1370
rect 15240 -1540 15380 -1530
rect 14900 -2310 14910 -1630
rect 15030 -2310 15040 -1630
rect 14200 -2920 14340 -2910
rect 14200 -3040 14210 -2920
rect 14330 -3040 14340 -2920
rect 14200 -3050 14340 -3040
rect 14420 -2920 14560 -2910
rect 14420 -3040 14430 -2920
rect 14550 -3040 14560 -2920
rect 14420 -3050 14560 -3040
rect 14440 -3130 14540 -3050
rect 12600 -3310 12740 -3300
rect 12600 -3410 12610 -3310
rect 12730 -3410 12740 -3310
rect 12600 -3420 12740 -3410
rect 13300 -3330 13310 -3170
rect 13430 -3330 13440 -3170
rect 12380 -4530 12520 -4520
rect 12380 -4650 12390 -4530
rect 12510 -4650 12520 -4530
rect 12380 -4660 12520 -4650
rect 12620 -4720 12720 -3420
rect 13300 -3430 13440 -3330
rect 13300 -4110 13310 -3430
rect 13430 -4110 13440 -3430
rect 13300 -4120 13440 -4110
rect 14000 -3240 14540 -3130
rect 14900 -3170 15040 -2310
rect 15600 -2460 15700 -800
rect 15820 -1110 15920 550
rect 16500 430 16640 1290
rect 17200 1140 17300 1290
rect 17190 1130 17310 1140
rect 17190 1010 17200 1130
rect 17300 1010 17310 1130
rect 17190 1000 17310 1010
rect 16500 270 16510 430
rect 16630 270 16640 430
rect 16500 170 16640 270
rect 16500 -510 16510 170
rect 16630 -510 16640 170
rect 15810 -1120 15930 -1110
rect 15810 -1240 15820 -1120
rect 15920 -1240 15930 -1120
rect 15810 -1250 15930 -1240
rect 15590 -2470 15710 -2460
rect 15590 -2590 15600 -2470
rect 15700 -2590 15710 -2470
rect 15590 -2600 15710 -2590
rect 12600 -4730 12740 -4720
rect 11020 -4850 11140 -4750
rect 1220 -8060 1320 -8050
rect 1200 -8070 1340 -8060
rect 1200 -8190 1210 -8070
rect 1330 -8190 1340 -8070
rect 1200 -8200 1340 -8190
rect 1220 -9860 1320 -8200
rect 1440 -8500 1540 -8050
rect 2820 -8060 2920 -8050
rect 2800 -8070 2940 -8060
rect 2800 -8190 2810 -8070
rect 2930 -8190 2940 -8070
rect 2800 -8200 2940 -8190
rect 1420 -8510 1560 -8500
rect 1420 -8630 1430 -8510
rect 1550 -8630 1560 -8510
rect 1420 -8640 1560 -8630
rect 1200 -9870 1340 -9860
rect 1200 -9990 1210 -9870
rect 1330 -9990 1340 -9870
rect 1200 -10000 1340 -9990
rect 1220 -11660 1320 -10000
rect 1440 -10300 1540 -8640
rect 2120 -8810 2240 -8780
rect 2120 -9470 2130 -8810
rect 2230 -9470 2240 -8810
rect 2120 -9590 2240 -9470
rect 2120 -9750 2130 -9590
rect 2230 -9750 2240 -9590
rect 1420 -10310 1560 -10300
rect 1420 -10430 1430 -10310
rect 1550 -10430 1560 -10310
rect 1420 -10440 1560 -10430
rect 1200 -11670 1340 -11660
rect 1200 -11790 1210 -11670
rect 1330 -11790 1340 -11670
rect 1200 -11800 1340 -11790
rect 1220 -13460 1320 -11800
rect 1440 -12100 1540 -10440
rect 2120 -10610 2240 -9750
rect 2820 -9860 2920 -8200
rect 3040 -8500 3140 -8050
rect 4420 -8060 4520 -8050
rect 4400 -8070 4540 -8060
rect 4400 -8190 4410 -8070
rect 4530 -8190 4540 -8070
rect 4400 -8200 4540 -8190
rect 3020 -8510 3160 -8500
rect 3020 -8630 3030 -8510
rect 3150 -8630 3160 -8510
rect 3020 -8640 3160 -8630
rect 2800 -9870 2940 -9860
rect 2800 -9990 2810 -9870
rect 2930 -9990 2940 -9870
rect 2800 -10000 2940 -9990
rect 2120 -11270 2130 -10610
rect 2230 -11270 2240 -10610
rect 2120 -11390 2240 -11270
rect 2120 -11550 2130 -11390
rect 2230 -11550 2240 -11390
rect 1420 -12110 1560 -12100
rect 1420 -12230 1430 -12110
rect 1550 -12230 1560 -12110
rect 1420 -12240 1560 -12230
rect 1200 -13470 1340 -13460
rect 1200 -13590 1210 -13470
rect 1330 -13590 1340 -13470
rect 1200 -13600 1340 -13590
rect 1220 -15260 1320 -13600
rect 1440 -13900 1540 -12240
rect 2120 -12410 2240 -11550
rect 2820 -11660 2920 -10000
rect 3040 -10300 3140 -8640
rect 3720 -8810 3840 -8780
rect 3720 -9470 3730 -8810
rect 3830 -9470 3840 -8810
rect 3720 -9590 3840 -9470
rect 3720 -9750 3730 -9590
rect 3830 -9750 3840 -9590
rect 3020 -10310 3160 -10300
rect 3020 -10430 3030 -10310
rect 3150 -10430 3160 -10310
rect 3020 -10440 3160 -10430
rect 2800 -11670 2940 -11660
rect 2800 -11790 2810 -11670
rect 2930 -11790 2940 -11670
rect 2800 -11800 2940 -11790
rect 2120 -13070 2130 -12410
rect 2230 -13070 2240 -12410
rect 2120 -13190 2240 -13070
rect 2120 -13350 2130 -13190
rect 2230 -13350 2240 -13190
rect 1420 -13910 1560 -13900
rect 1420 -14030 1430 -13910
rect 1550 -14030 1560 -13910
rect 1420 -14040 1560 -14030
rect 1200 -15270 1340 -15260
rect 1200 -15390 1210 -15270
rect 1330 -15390 1340 -15270
rect 1200 -15400 1340 -15390
rect 1220 -17060 1320 -15400
rect 1440 -15700 1540 -14040
rect 2120 -14210 2240 -13350
rect 2820 -13460 2920 -11800
rect 3040 -12100 3140 -10440
rect 3720 -10610 3840 -9750
rect 4420 -9860 4520 -8200
rect 4640 -8500 4740 -8050
rect 6020 -8060 6120 -8050
rect 6000 -8070 6140 -8060
rect 6000 -8190 6010 -8070
rect 6130 -8190 6140 -8070
rect 6000 -8200 6140 -8190
rect 4620 -8510 4760 -8500
rect 4620 -8630 4630 -8510
rect 4750 -8630 4760 -8510
rect 4620 -8640 4760 -8630
rect 4400 -9870 4540 -9860
rect 4400 -9990 4410 -9870
rect 4530 -9990 4540 -9870
rect 4400 -10000 4540 -9990
rect 3720 -11270 3730 -10610
rect 3830 -11270 3840 -10610
rect 3720 -11390 3840 -11270
rect 3720 -11550 3730 -11390
rect 3830 -11550 3840 -11390
rect 3020 -12110 3160 -12100
rect 3020 -12230 3030 -12110
rect 3150 -12230 3160 -12110
rect 3020 -12240 3160 -12230
rect 2800 -13470 2940 -13460
rect 2800 -13590 2810 -13470
rect 2930 -13590 2940 -13470
rect 2800 -13600 2940 -13590
rect 2120 -14870 2130 -14210
rect 2230 -14870 2240 -14210
rect 2120 -14990 2240 -14870
rect 2120 -15150 2130 -14990
rect 2230 -15150 2240 -14990
rect 1420 -15710 1560 -15700
rect 1420 -15830 1430 -15710
rect 1550 -15830 1560 -15710
rect 1420 -15840 1560 -15830
rect 1200 -17070 1340 -17060
rect 1200 -17190 1210 -17070
rect 1330 -17190 1340 -17070
rect 1200 -17200 1340 -17190
rect 1220 -18860 1320 -17200
rect 1440 -17500 1540 -15840
rect 2120 -16010 2240 -15150
rect 2820 -15260 2920 -13600
rect 3040 -13900 3140 -12240
rect 3720 -12410 3840 -11550
rect 4420 -11660 4520 -10000
rect 4640 -10300 4740 -8640
rect 5320 -8810 5440 -8780
rect 5320 -9470 5330 -8810
rect 5430 -9470 5440 -8810
rect 5320 -9590 5440 -9470
rect 5320 -9750 5330 -9590
rect 5430 -9750 5440 -9590
rect 4620 -10310 4760 -10300
rect 4620 -10430 4630 -10310
rect 4750 -10430 4760 -10310
rect 4620 -10440 4760 -10430
rect 4400 -11670 4540 -11660
rect 4400 -11790 4410 -11670
rect 4530 -11790 4540 -11670
rect 4400 -11800 4540 -11790
rect 3720 -13070 3730 -12410
rect 3830 -13070 3840 -12410
rect 3720 -13190 3840 -13070
rect 3720 -13350 3730 -13190
rect 3830 -13350 3840 -13190
rect 3020 -13910 3160 -13900
rect 3020 -14030 3030 -13910
rect 3150 -14030 3160 -13910
rect 3020 -14040 3160 -14030
rect 2800 -15270 2940 -15260
rect 2800 -15390 2810 -15270
rect 2930 -15390 2940 -15270
rect 2800 -15400 2940 -15390
rect 2120 -16670 2130 -16010
rect 2230 -16670 2240 -16010
rect 2120 -16790 2240 -16670
rect 2120 -16950 2130 -16790
rect 2230 -16950 2240 -16790
rect 1420 -17510 1560 -17500
rect 1420 -17630 1430 -17510
rect 1550 -17630 1560 -17510
rect 1420 -17640 1560 -17630
rect 1200 -18870 1340 -18860
rect 1200 -18990 1210 -18870
rect 1330 -18990 1340 -18870
rect 1200 -19000 1340 -18990
rect 1220 -20660 1320 -19000
rect 1440 -19300 1540 -17640
rect 2120 -17810 2240 -16950
rect 2820 -17060 2920 -15400
rect 3040 -15700 3140 -14040
rect 3720 -14210 3840 -13350
rect 4420 -13460 4520 -11800
rect 4640 -12100 4740 -10440
rect 5320 -10610 5440 -9750
rect 6020 -9860 6120 -8200
rect 6240 -8500 6340 -8050
rect 7620 -8060 7720 -8050
rect 7600 -8070 7740 -8060
rect 7600 -8190 7610 -8070
rect 7730 -8190 7740 -8070
rect 7600 -8200 7740 -8190
rect 6220 -8510 6360 -8500
rect 6220 -8630 6230 -8510
rect 6350 -8630 6360 -8510
rect 6220 -8640 6360 -8630
rect 6000 -9870 6140 -9860
rect 6000 -9990 6010 -9870
rect 6130 -9990 6140 -9870
rect 6000 -10000 6140 -9990
rect 5320 -11270 5330 -10610
rect 5430 -11270 5440 -10610
rect 5320 -11390 5440 -11270
rect 5320 -11550 5330 -11390
rect 5430 -11550 5440 -11390
rect 4620 -12110 4760 -12100
rect 4620 -12230 4630 -12110
rect 4750 -12230 4760 -12110
rect 4620 -12240 4760 -12230
rect 4400 -13470 4540 -13460
rect 4400 -13590 4410 -13470
rect 4530 -13590 4540 -13470
rect 4400 -13600 4540 -13590
rect 3720 -14870 3730 -14210
rect 3830 -14870 3840 -14210
rect 3720 -14990 3840 -14870
rect 3720 -15150 3730 -14990
rect 3830 -15150 3840 -14990
rect 3020 -15710 3160 -15700
rect 3020 -15830 3030 -15710
rect 3150 -15830 3160 -15710
rect 3020 -15840 3160 -15830
rect 2800 -17070 2940 -17060
rect 2800 -17190 2810 -17070
rect 2930 -17190 2940 -17070
rect 2800 -17200 2940 -17190
rect 2120 -18470 2130 -17810
rect 2230 -18470 2240 -17810
rect 2120 -18590 2240 -18470
rect 2120 -18750 2130 -18590
rect 2230 -18750 2240 -18590
rect 1420 -19310 1560 -19300
rect 1420 -19430 1430 -19310
rect 1550 -19430 1560 -19310
rect 1420 -19440 1560 -19430
rect 1200 -20670 1340 -20660
rect 1200 -20790 1210 -20670
rect 1330 -20790 1340 -20670
rect 1200 -20800 1340 -20790
rect 1220 -22640 1320 -20800
rect 1440 -21100 1540 -19440
rect 2120 -19610 2240 -18750
rect 2820 -18860 2920 -17200
rect 3040 -17500 3140 -15840
rect 3720 -16010 3840 -15150
rect 4420 -15260 4520 -13600
rect 4640 -13900 4740 -12240
rect 5320 -12410 5440 -11550
rect 6020 -11660 6120 -10000
rect 6240 -10300 6340 -8640
rect 6920 -8810 7040 -8780
rect 6920 -9470 6930 -8810
rect 7030 -9470 7040 -8810
rect 6920 -9590 7040 -9470
rect 6920 -9750 6930 -9590
rect 7030 -9750 7040 -9590
rect 6220 -10310 6360 -10300
rect 6220 -10430 6230 -10310
rect 6350 -10430 6360 -10310
rect 6220 -10440 6360 -10430
rect 6000 -11670 6140 -11660
rect 6000 -11790 6010 -11670
rect 6130 -11790 6140 -11670
rect 6000 -11800 6140 -11790
rect 5320 -13070 5330 -12410
rect 5430 -13070 5440 -12410
rect 5320 -13190 5440 -13070
rect 5320 -13350 5330 -13190
rect 5430 -13350 5440 -13190
rect 4620 -13910 4760 -13900
rect 4620 -14030 4630 -13910
rect 4750 -14030 4760 -13910
rect 4620 -14040 4760 -14030
rect 4400 -15270 4540 -15260
rect 4400 -15390 4410 -15270
rect 4530 -15390 4540 -15270
rect 4400 -15400 4540 -15390
rect 3720 -16670 3730 -16010
rect 3830 -16670 3840 -16010
rect 3720 -16790 3840 -16670
rect 3720 -16950 3730 -16790
rect 3830 -16950 3840 -16790
rect 3020 -17510 3160 -17500
rect 3020 -17630 3030 -17510
rect 3150 -17630 3160 -17510
rect 3020 -17640 3160 -17630
rect 2800 -18870 2940 -18860
rect 2800 -18990 2810 -18870
rect 2930 -18990 2940 -18870
rect 2800 -19000 2940 -18990
rect 2120 -20270 2130 -19610
rect 2230 -20270 2240 -19610
rect 2120 -20390 2240 -20270
rect 2120 -20550 2130 -20390
rect 2230 -20550 2240 -20390
rect 1420 -21110 1560 -21100
rect 1420 -21230 1430 -21110
rect 1550 -21230 1560 -21110
rect 1420 -21240 1560 -21230
rect 2120 -21410 2240 -20550
rect 2820 -20660 2920 -19000
rect 3040 -19300 3140 -17640
rect 3720 -17810 3840 -16950
rect 4420 -17060 4520 -15400
rect 4640 -15700 4740 -14040
rect 5320 -14210 5440 -13350
rect 6020 -13460 6120 -11800
rect 6240 -12100 6340 -10440
rect 6920 -10610 7040 -9750
rect 7620 -9860 7720 -8200
rect 7840 -8500 7940 -8050
rect 9220 -8060 9320 -8050
rect 9200 -8070 9340 -8060
rect 9200 -8190 9210 -8070
rect 9330 -8190 9340 -8070
rect 9200 -8200 9340 -8190
rect 7820 -8510 7960 -8500
rect 7820 -8630 7830 -8510
rect 7950 -8630 7960 -8510
rect 7820 -8640 7960 -8630
rect 7600 -9870 7740 -9860
rect 7600 -9990 7610 -9870
rect 7730 -9990 7740 -9870
rect 7600 -10000 7740 -9990
rect 6920 -11270 6930 -10610
rect 7030 -11270 7040 -10610
rect 6920 -11390 7040 -11270
rect 6920 -11550 6930 -11390
rect 7030 -11550 7040 -11390
rect 6220 -12110 6360 -12100
rect 6220 -12230 6230 -12110
rect 6350 -12230 6360 -12110
rect 6220 -12240 6360 -12230
rect 6000 -13470 6140 -13460
rect 6000 -13590 6010 -13470
rect 6130 -13590 6140 -13470
rect 6000 -13600 6140 -13590
rect 5320 -14870 5330 -14210
rect 5430 -14870 5440 -14210
rect 5320 -14990 5440 -14870
rect 5320 -15150 5330 -14990
rect 5430 -15150 5440 -14990
rect 4620 -15710 4760 -15700
rect 4620 -15830 4630 -15710
rect 4750 -15830 4760 -15710
rect 4620 -15840 4760 -15830
rect 4400 -17070 4540 -17060
rect 4400 -17190 4410 -17070
rect 4530 -17190 4540 -17070
rect 4400 -17200 4540 -17190
rect 3720 -18470 3730 -17810
rect 3830 -18470 3840 -17810
rect 3720 -18590 3840 -18470
rect 3720 -18750 3730 -18590
rect 3830 -18750 3840 -18590
rect 3020 -19310 3160 -19300
rect 3020 -19430 3030 -19310
rect 3150 -19430 3160 -19310
rect 3020 -19440 3160 -19430
rect 2800 -20670 2940 -20660
rect 2800 -20790 2810 -20670
rect 2930 -20790 2940 -20670
rect 2800 -20800 2940 -20790
rect 2120 -22070 2130 -21410
rect 2230 -22070 2240 -21410
rect 2120 -22190 2240 -22070
rect 2120 -22350 2130 -22190
rect 2230 -22350 2240 -22190
rect 2120 -22360 2240 -22350
rect 2820 -23260 2920 -20800
rect 3040 -21100 3140 -19440
rect 3720 -19610 3840 -18750
rect 4420 -18860 4520 -17200
rect 4640 -17500 4740 -15840
rect 5320 -16010 5440 -15150
rect 6020 -15260 6120 -13600
rect 6240 -13900 6340 -12240
rect 6920 -12410 7040 -11550
rect 7620 -11660 7720 -10000
rect 7840 -10300 7940 -8640
rect 8520 -8810 8640 -8780
rect 8520 -9470 8530 -8810
rect 8630 -9470 8640 -8810
rect 8520 -9590 8640 -9470
rect 8520 -9750 8530 -9590
rect 8630 -9750 8640 -9590
rect 7820 -10310 7960 -10300
rect 7820 -10430 7830 -10310
rect 7950 -10430 7960 -10310
rect 7820 -10440 7960 -10430
rect 7600 -11670 7740 -11660
rect 7600 -11790 7610 -11670
rect 7730 -11790 7740 -11670
rect 7600 -11800 7740 -11790
rect 6920 -13070 6930 -12410
rect 7030 -13070 7040 -12410
rect 6920 -13190 7040 -13070
rect 6920 -13350 6930 -13190
rect 7030 -13350 7040 -13190
rect 6220 -13910 6360 -13900
rect 6220 -14030 6230 -13910
rect 6350 -14030 6360 -13910
rect 6220 -14040 6360 -14030
rect 6000 -15270 6140 -15260
rect 6000 -15390 6010 -15270
rect 6130 -15390 6140 -15270
rect 6000 -15400 6140 -15390
rect 5320 -16670 5330 -16010
rect 5430 -16670 5440 -16010
rect 5320 -16790 5440 -16670
rect 5320 -16950 5330 -16790
rect 5430 -16950 5440 -16790
rect 4620 -17510 4760 -17500
rect 4620 -17630 4630 -17510
rect 4750 -17630 4760 -17510
rect 4620 -17640 4760 -17630
rect 4400 -18870 4540 -18860
rect 4400 -18990 4410 -18870
rect 4530 -18990 4540 -18870
rect 4400 -19000 4540 -18990
rect 3720 -20270 3730 -19610
rect 3830 -20270 3840 -19610
rect 3720 -20390 3840 -20270
rect 3720 -20550 3730 -20390
rect 3830 -20550 3840 -20390
rect 3020 -21110 3160 -21100
rect 3020 -21230 3030 -21110
rect 3150 -21230 3160 -21110
rect 3020 -21240 3160 -21230
rect 3720 -21410 3840 -20550
rect 4420 -20660 4520 -19000
rect 4640 -19300 4740 -17640
rect 5320 -17810 5440 -16950
rect 6020 -17060 6120 -15400
rect 6240 -15700 6340 -14040
rect 6920 -14210 7040 -13350
rect 7620 -13460 7720 -11800
rect 7840 -12100 7940 -10440
rect 8520 -10610 8640 -9750
rect 9220 -9860 9320 -8200
rect 9440 -8500 9540 -8050
rect 9420 -8510 9560 -8500
rect 9420 -8630 9430 -8510
rect 9550 -8630 9560 -8510
rect 9420 -8640 9560 -8630
rect 9200 -9870 9340 -9860
rect 9200 -9990 9210 -9870
rect 9330 -9990 9340 -9870
rect 9200 -10000 9340 -9990
rect 8520 -11270 8530 -10610
rect 8630 -11270 8640 -10610
rect 8520 -11390 8640 -11270
rect 8520 -11550 8530 -11390
rect 8630 -11550 8640 -11390
rect 7820 -12110 7960 -12100
rect 7820 -12230 7830 -12110
rect 7950 -12230 7960 -12110
rect 7820 -12240 7960 -12230
rect 7600 -13470 7740 -13460
rect 7600 -13590 7610 -13470
rect 7730 -13590 7740 -13470
rect 7600 -13600 7740 -13590
rect 6920 -14870 6930 -14210
rect 7030 -14870 7040 -14210
rect 6920 -14990 7040 -14870
rect 6920 -15150 6930 -14990
rect 7030 -15150 7040 -14990
rect 6220 -15710 6360 -15700
rect 6220 -15830 6230 -15710
rect 6350 -15830 6360 -15710
rect 6220 -15840 6360 -15830
rect 6000 -17070 6140 -17060
rect 6000 -17190 6010 -17070
rect 6130 -17190 6140 -17070
rect 6000 -17200 6140 -17190
rect 5320 -18470 5330 -17810
rect 5430 -18470 5440 -17810
rect 5320 -18590 5440 -18470
rect 5320 -18750 5330 -18590
rect 5430 -18750 5440 -18590
rect 4620 -19310 4760 -19300
rect 4620 -19430 4630 -19310
rect 4750 -19430 4760 -19310
rect 4620 -19440 4760 -19430
rect 4400 -20670 4540 -20660
rect 4400 -20790 4410 -20670
rect 4530 -20790 4540 -20670
rect 4400 -20800 4540 -20790
rect 3720 -22070 3730 -21410
rect 3830 -22070 3840 -21410
rect 3720 -22190 3840 -22070
rect 3720 -22350 3730 -22190
rect 3830 -22350 3840 -22190
rect 3720 -22360 3840 -22350
rect 4420 -23260 4520 -20800
rect 4640 -21100 4740 -19440
rect 5320 -19610 5440 -18750
rect 6020 -18860 6120 -17200
rect 6240 -17500 6340 -15840
rect 6920 -16010 7040 -15150
rect 7620 -15260 7720 -13600
rect 7840 -13900 7940 -12240
rect 8520 -12410 8640 -11550
rect 9220 -11660 9320 -10000
rect 9440 -10300 9540 -8640
rect 10120 -8810 10240 -8780
rect 10120 -9470 10130 -8810
rect 10230 -9470 10240 -8810
rect 10120 -9590 10240 -9470
rect 10120 -9750 10130 -9590
rect 10230 -9750 10240 -9590
rect 9420 -10310 9560 -10300
rect 9420 -10430 9430 -10310
rect 9550 -10430 9560 -10310
rect 9420 -10440 9560 -10430
rect 9200 -11670 9340 -11660
rect 9200 -11790 9210 -11670
rect 9330 -11790 9340 -11670
rect 9200 -11800 9340 -11790
rect 8520 -13070 8530 -12410
rect 8630 -13070 8640 -12410
rect 8520 -13190 8640 -13070
rect 8520 -13350 8530 -13190
rect 8630 -13350 8640 -13190
rect 7820 -13910 7960 -13900
rect 7820 -14030 7830 -13910
rect 7950 -14030 7960 -13910
rect 7820 -14040 7960 -14030
rect 7600 -15270 7740 -15260
rect 7600 -15390 7610 -15270
rect 7730 -15390 7740 -15270
rect 7600 -15400 7740 -15390
rect 6920 -16670 6930 -16010
rect 7030 -16670 7040 -16010
rect 6920 -16790 7040 -16670
rect 6920 -16950 6930 -16790
rect 7030 -16950 7040 -16790
rect 6220 -17510 6360 -17500
rect 6220 -17630 6230 -17510
rect 6350 -17630 6360 -17510
rect 6220 -17640 6360 -17630
rect 6000 -18870 6140 -18860
rect 6000 -18990 6010 -18870
rect 6130 -18990 6140 -18870
rect 6000 -19000 6140 -18990
rect 5320 -20270 5330 -19610
rect 5430 -20270 5440 -19610
rect 5320 -20390 5440 -20270
rect 5320 -20550 5330 -20390
rect 5430 -20550 5440 -20390
rect 4620 -21110 4760 -21100
rect 4620 -21230 4630 -21110
rect 4750 -21230 4760 -21110
rect 4620 -21240 4760 -21230
rect 5320 -21410 5440 -20550
rect 6020 -20660 6120 -19000
rect 6240 -19300 6340 -17640
rect 6920 -17810 7040 -16950
rect 7620 -17060 7720 -15400
rect 7840 -15700 7940 -14040
rect 8520 -14210 8640 -13350
rect 9220 -13460 9320 -11800
rect 9440 -12100 9540 -10440
rect 10120 -10610 10240 -9750
rect 10120 -11270 10130 -10610
rect 10230 -11270 10240 -10610
rect 10120 -11390 10240 -11270
rect 10120 -11550 10130 -11390
rect 10230 -11550 10240 -11390
rect 9420 -12110 9560 -12100
rect 9420 -12230 9430 -12110
rect 9550 -12230 9560 -12110
rect 9420 -12240 9560 -12230
rect 9200 -13470 9340 -13460
rect 9200 -13590 9210 -13470
rect 9330 -13590 9340 -13470
rect 9200 -13600 9340 -13590
rect 8520 -14870 8530 -14210
rect 8630 -14870 8640 -14210
rect 8520 -14990 8640 -14870
rect 8520 -15150 8530 -14990
rect 8630 -15150 8640 -14990
rect 7820 -15710 7960 -15700
rect 7820 -15830 7830 -15710
rect 7950 -15830 7960 -15710
rect 7820 -15840 7960 -15830
rect 7600 -17070 7740 -17060
rect 7600 -17190 7610 -17070
rect 7730 -17190 7740 -17070
rect 7600 -17200 7740 -17190
rect 6920 -18470 6930 -17810
rect 7030 -18470 7040 -17810
rect 6920 -18590 7040 -18470
rect 6920 -18750 6930 -18590
rect 7030 -18750 7040 -18590
rect 6220 -19310 6360 -19300
rect 6220 -19430 6230 -19310
rect 6350 -19430 6360 -19310
rect 6220 -19440 6360 -19430
rect 6000 -20670 6140 -20660
rect 6000 -20790 6010 -20670
rect 6130 -20790 6140 -20670
rect 6000 -20800 6140 -20790
rect 5320 -22070 5330 -21410
rect 5430 -22070 5440 -21410
rect 5320 -22190 5440 -22070
rect 5320 -22350 5330 -22190
rect 5430 -22350 5440 -22190
rect 5320 -22360 5440 -22350
rect 6020 -23260 6120 -20800
rect 6240 -21100 6340 -19440
rect 6920 -19610 7040 -18750
rect 7620 -18860 7720 -17200
rect 7840 -17500 7940 -15840
rect 8520 -16010 8640 -15150
rect 9220 -15260 9320 -13600
rect 9440 -13900 9540 -12240
rect 10120 -12410 10240 -11550
rect 10820 -12210 10920 -7800
rect 11040 -9580 11140 -4850
rect 11700 -4810 11840 -4800
rect 11700 -4930 11710 -4810
rect 11830 -4930 11840 -4810
rect 12600 -4850 12610 -4730
rect 12730 -4850 12740 -4730
rect 12600 -4860 12740 -4850
rect 13620 -4790 13760 -4780
rect 13620 -4910 13630 -4790
rect 13750 -4910 13760 -4790
rect 13620 -4920 13760 -4910
rect 11700 -4940 11840 -4930
rect 11720 -5820 11820 -4940
rect 11700 -5830 11840 -5820
rect 11700 -5950 11710 -5830
rect 11830 -5950 11840 -5830
rect 11700 -5960 11840 -5950
rect 13300 -5830 13440 -5820
rect 13300 -5950 13310 -5830
rect 13430 -5950 13440 -5830
rect 13300 -5960 13440 -5950
rect 11700 -6050 11840 -6040
rect 11700 -6170 11710 -6050
rect 11830 -6170 11840 -6050
rect 11700 -6180 11840 -6170
rect 11720 -8100 11820 -6180
rect 12620 -6270 12760 -6260
rect 12620 -6390 12630 -6270
rect 12750 -6390 12760 -6270
rect 12620 -6400 12760 -6390
rect 12400 -6490 12540 -6480
rect 12400 -6610 12410 -6490
rect 12530 -6610 12540 -6490
rect 12400 -6620 12540 -6610
rect 11700 -8110 11860 -8100
rect 11700 -8230 11710 -8110
rect 11840 -8140 11860 -8110
rect 11840 -8230 11850 -8140
rect 11700 -8240 11850 -8230
rect 11710 -8810 11840 -8240
rect 11710 -9470 11720 -8810
rect 11830 -9470 11840 -8810
rect 11710 -9480 11840 -9470
rect 11030 -9760 11150 -9580
rect 11040 -10400 11140 -9760
rect 11020 -10410 11160 -10400
rect 11020 -10530 11030 -10410
rect 11150 -10530 11160 -10410
rect 11020 -10540 11160 -10530
rect 11040 -11380 11140 -10540
rect 11710 -10610 11840 -10600
rect 11710 -11270 11720 -10610
rect 11830 -11270 11840 -10610
rect 11030 -11560 11150 -11380
rect 10800 -12220 10940 -12210
rect 10800 -12330 10810 -12220
rect 10930 -12330 10940 -12220
rect 10800 -12340 10940 -12330
rect 10120 -13070 10130 -12410
rect 10230 -13070 10240 -12410
rect 10120 -13190 10240 -13070
rect 11040 -13180 11140 -11560
rect 11710 -12410 11840 -11270
rect 11710 -13070 11720 -12410
rect 11830 -13070 11840 -12410
rect 10120 -13350 10130 -13190
rect 10230 -13350 10240 -13190
rect 9420 -13910 9560 -13900
rect 9420 -14030 9430 -13910
rect 9550 -14030 9560 -13910
rect 9420 -14040 9560 -14030
rect 9200 -15270 9340 -15260
rect 9200 -15390 9210 -15270
rect 9330 -15390 9340 -15270
rect 9200 -15400 9340 -15390
rect 8520 -16670 8530 -16010
rect 8630 -16670 8640 -16010
rect 8520 -16790 8640 -16670
rect 8520 -16950 8530 -16790
rect 8630 -16950 8640 -16790
rect 7820 -17510 7960 -17500
rect 7820 -17630 7830 -17510
rect 7950 -17630 7960 -17510
rect 7820 -17640 7960 -17630
rect 7600 -18870 7740 -18860
rect 7600 -18990 7610 -18870
rect 7730 -18990 7740 -18870
rect 7600 -19000 7740 -18990
rect 6920 -20270 6930 -19610
rect 7030 -20270 7040 -19610
rect 6920 -20390 7040 -20270
rect 6920 -20550 6930 -20390
rect 7030 -20550 7040 -20390
rect 6220 -21110 6360 -21100
rect 6220 -21230 6230 -21110
rect 6350 -21230 6360 -21110
rect 6220 -21240 6360 -21230
rect 6920 -21410 7040 -20550
rect 7620 -20660 7720 -19000
rect 7840 -19300 7940 -17640
rect 8520 -17810 8640 -16950
rect 9220 -17060 9320 -15400
rect 9440 -15700 9540 -14040
rect 10120 -14210 10240 -13350
rect 11030 -13360 11150 -13180
rect 11260 -13210 11270 -13150
rect 11650 -13210 11660 -13150
rect 10120 -14870 10130 -14210
rect 10230 -14870 10240 -14210
rect 10120 -14990 10240 -14870
rect 11040 -14980 11140 -13360
rect 11260 -14060 11660 -13210
rect 11260 -14120 11270 -14060
rect 11650 -14120 11660 -14060
rect 11260 -14130 11660 -14120
rect 11710 -14210 11840 -13070
rect 11710 -14870 11720 -14210
rect 11830 -14870 11840 -14210
rect 11710 -14880 11840 -14870
rect 10120 -15150 10130 -14990
rect 10230 -15150 10240 -14990
rect 9420 -15710 9560 -15700
rect 9420 -15830 9430 -15710
rect 9550 -15830 9560 -15710
rect 9420 -15840 9560 -15830
rect 9200 -17070 9340 -17060
rect 9200 -17190 9210 -17070
rect 9330 -17190 9340 -17070
rect 9200 -17200 9340 -17190
rect 8520 -18470 8530 -17810
rect 8630 -18470 8640 -17810
rect 8520 -18590 8640 -18470
rect 8520 -18750 8530 -18590
rect 8630 -18750 8640 -18590
rect 7820 -19310 7960 -19300
rect 7820 -19430 7830 -19310
rect 7950 -19430 7960 -19310
rect 7820 -19440 7960 -19430
rect 7600 -20670 7740 -20660
rect 7600 -20790 7610 -20670
rect 7730 -20790 7740 -20670
rect 7600 -20800 7740 -20790
rect 6920 -22070 6930 -21410
rect 7030 -22070 7040 -21410
rect 6920 -22190 7040 -22070
rect 6920 -22350 6930 -22190
rect 7030 -22350 7040 -22190
rect 6920 -22360 7040 -22350
rect 7620 -23260 7720 -20800
rect 7840 -21100 7940 -19440
rect 8520 -19610 8640 -18750
rect 9220 -18860 9320 -17200
rect 9440 -17500 9540 -15840
rect 10120 -16010 10240 -15150
rect 11030 -15160 11150 -14980
rect 10120 -16670 10130 -16010
rect 10230 -16670 10240 -16010
rect 10120 -16790 10240 -16670
rect 11040 -16780 11140 -15160
rect 11710 -16010 11840 -16000
rect 11710 -16670 11720 -16010
rect 11830 -16670 11840 -16010
rect 11710 -16680 11840 -16670
rect 10120 -16950 10130 -16790
rect 10230 -16950 10240 -16790
rect 9420 -17510 9560 -17500
rect 9420 -17630 9430 -17510
rect 9550 -17630 9560 -17510
rect 9420 -17640 9560 -17630
rect 9200 -18870 9340 -18860
rect 9200 -18990 9210 -18870
rect 9330 -18990 9340 -18870
rect 9200 -19000 9340 -18990
rect 8520 -20270 8530 -19610
rect 8630 -20270 8640 -19610
rect 8520 -20390 8640 -20270
rect 8520 -20550 8530 -20390
rect 8630 -20550 8640 -20390
rect 7820 -21110 7960 -21100
rect 7820 -21230 7830 -21110
rect 7950 -21230 7960 -21110
rect 7820 -21240 7960 -21230
rect 8520 -21410 8640 -20550
rect 9220 -20660 9320 -19000
rect 9440 -19300 9540 -17640
rect 10120 -17810 10240 -16950
rect 11030 -16960 11150 -16780
rect 10120 -18470 10130 -17810
rect 10230 -18470 10240 -17810
rect 10120 -18590 10240 -18470
rect 11040 -18580 11140 -16960
rect 11710 -17810 11840 -17800
rect 11710 -18470 11720 -17810
rect 11830 -18470 11840 -17810
rect 11710 -18480 11840 -18470
rect 10120 -18750 10130 -18590
rect 10230 -18750 10240 -18590
rect 9420 -19310 9560 -19300
rect 9420 -19430 9430 -19310
rect 9550 -19430 9560 -19310
rect 9420 -19440 9560 -19430
rect 9200 -20670 9340 -20660
rect 9200 -20790 9210 -20670
rect 9330 -20790 9340 -20670
rect 9200 -20800 9340 -20790
rect 8520 -22070 8530 -21410
rect 8630 -22070 8640 -21410
rect 8520 -22190 8640 -22070
rect 8520 -22350 8530 -22190
rect 8630 -22350 8640 -22190
rect 8520 -22360 8640 -22350
rect 9220 -23260 9320 -20800
rect 9440 -21100 9540 -19440
rect 10120 -19610 10240 -18750
rect 11030 -18760 11150 -18580
rect 10120 -20270 10130 -19610
rect 10230 -20270 10240 -19610
rect 10120 -20390 10240 -20270
rect 11040 -20380 11140 -18760
rect 12420 -18870 12520 -6620
rect 12640 -17070 12740 -6400
rect 13310 -8240 13440 -5960
rect 13640 -6040 13740 -4920
rect 14000 -5070 14100 -3240
rect 14200 -3310 14340 -3300
rect 14200 -3430 14210 -3310
rect 14330 -3430 14340 -3310
rect 14200 -3440 14340 -3430
rect 14900 -3330 14910 -3170
rect 15030 -3330 15040 -3170
rect 14900 -3430 15040 -3330
rect 14220 -4720 14320 -3440
rect 14900 -4110 14910 -3430
rect 15030 -4110 15040 -3430
rect 14900 -4120 15040 -4110
rect 15600 -4260 15700 -2600
rect 15820 -2910 15920 -1250
rect 16500 -1370 16640 -510
rect 17200 -660 17300 1000
rect 17420 690 17520 1290
rect 17410 680 17530 690
rect 17410 560 17420 680
rect 17520 560 17530 680
rect 17410 550 17530 560
rect 17190 -670 17310 -660
rect 17190 -790 17200 -670
rect 17300 -790 17310 -670
rect 17190 -800 17310 -790
rect 16500 -1530 16510 -1370
rect 16630 -1530 16640 -1370
rect 16500 -1630 16640 -1530
rect 16500 -2310 16510 -1630
rect 16630 -2310 16640 -1630
rect 15810 -2920 15930 -2910
rect 15810 -3040 15820 -2920
rect 15920 -3040 15930 -2920
rect 15810 -3050 15930 -3040
rect 15590 -4270 15710 -4260
rect 15590 -4390 15600 -4270
rect 15700 -4390 15710 -4270
rect 15590 -4400 15710 -4390
rect 14200 -4730 14340 -4720
rect 14200 -4850 14210 -4730
rect 14330 -4850 14340 -4730
rect 14200 -4860 14340 -4850
rect 15220 -4790 15360 -4780
rect 15220 -4910 15230 -4790
rect 15350 -4910 15360 -4790
rect 15220 -4920 15360 -4910
rect 14000 -5200 14120 -5070
rect 13620 -6050 13760 -6040
rect 13620 -6170 13630 -6050
rect 13750 -6170 13760 -6050
rect 13620 -6180 13760 -6170
rect 13300 -8390 13450 -8240
rect 13310 -8810 13440 -8390
rect 13310 -9470 13320 -8810
rect 13430 -9470 13440 -8810
rect 13310 -9480 13440 -9470
rect 13310 -10610 13440 -10600
rect 13310 -11270 13320 -10610
rect 13430 -11270 13440 -10610
rect 13310 -11280 13440 -11270
rect 13300 -11670 13440 -11660
rect 13300 -11790 13310 -11670
rect 13430 -11790 13440 -11670
rect 13300 -11800 13440 -11790
rect 13310 -12410 13440 -11800
rect 13310 -13070 13320 -12410
rect 13430 -13070 13440 -12410
rect 13310 -13160 13440 -13070
rect 13280 -13170 13470 -13160
rect 13280 -13330 13290 -13170
rect 13460 -13330 13470 -13170
rect 13280 -13340 13470 -13330
rect 13310 -14210 13440 -13340
rect 14020 -13470 14120 -5200
rect 15240 -6040 15340 -4920
rect 15600 -5160 15700 -4400
rect 15820 -4710 15920 -3050
rect 16500 -3170 16640 -2310
rect 17200 -2460 17300 -800
rect 17420 -1110 17520 550
rect 18100 430 18240 1290
rect 18800 1140 18900 1290
rect 18790 1130 18910 1140
rect 18790 1010 18800 1130
rect 18900 1010 18910 1130
rect 18790 1000 18910 1010
rect 18100 270 18110 430
rect 18230 270 18240 430
rect 18100 170 18240 270
rect 18100 -510 18110 170
rect 18230 -510 18240 170
rect 17410 -1120 17530 -1110
rect 17410 -1240 17420 -1120
rect 17520 -1240 17530 -1120
rect 17410 -1250 17530 -1240
rect 17190 -2470 17310 -2460
rect 17190 -2590 17200 -2470
rect 17300 -2590 17310 -2470
rect 17190 -2600 17310 -2590
rect 16500 -3330 16510 -3170
rect 16630 -3330 16640 -3170
rect 16500 -3430 16640 -3330
rect 16500 -4110 16510 -3430
rect 16630 -4110 16640 -3430
rect 15810 -4720 15930 -4710
rect 15810 -4840 15820 -4720
rect 15920 -4840 15930 -4720
rect 15810 -4850 15930 -4840
rect 15560 -5170 15740 -5160
rect 15560 -5350 15570 -5170
rect 15730 -5350 15740 -5170
rect 15560 -5360 15740 -5350
rect 15560 -5570 15740 -5560
rect 15560 -5750 15570 -5570
rect 15730 -5750 15740 -5570
rect 15560 -5760 15740 -5750
rect 14220 -6050 14360 -6040
rect 14220 -6170 14230 -6050
rect 14350 -6170 14360 -6050
rect 14220 -6180 14360 -6170
rect 15220 -6050 15360 -6040
rect 15220 -6170 15230 -6050
rect 15350 -6170 15360 -6050
rect 15220 -6180 15360 -6170
rect 14240 -11660 14340 -6180
rect 14900 -6490 15040 -6480
rect 14900 -6610 14910 -6490
rect 15030 -6610 15040 -6490
rect 14900 -6620 15040 -6610
rect 15620 -8510 15720 -5760
rect 15820 -5960 15920 -4850
rect 15780 -5970 15960 -5960
rect 15780 -6150 15790 -5970
rect 15950 -6150 15960 -5970
rect 15780 -6160 15960 -6150
rect 15840 -8060 15940 -6160
rect 16500 -6270 16640 -4110
rect 17200 -4260 17300 -2600
rect 17420 -2910 17520 -1250
rect 18100 -1370 18240 -510
rect 18800 -660 18900 1000
rect 19020 690 19120 1290
rect 19010 680 19130 690
rect 19010 560 19020 680
rect 19120 560 19130 680
rect 19010 550 19130 560
rect 18790 -670 18910 -660
rect 18790 -790 18800 -670
rect 18900 -790 18910 -670
rect 18790 -800 18910 -790
rect 18100 -1530 18110 -1370
rect 18230 -1530 18240 -1370
rect 18100 -1630 18240 -1530
rect 18100 -2310 18110 -1630
rect 18230 -2310 18240 -1630
rect 17410 -2920 17530 -2910
rect 17410 -3040 17420 -2920
rect 17520 -3040 17530 -2920
rect 17410 -3050 17530 -3040
rect 17190 -4270 17310 -4260
rect 17190 -4390 17200 -4270
rect 17300 -4390 17310 -4270
rect 17190 -4400 17310 -4390
rect 16500 -6390 16510 -6270
rect 16630 -6390 16640 -6270
rect 16500 -6400 16640 -6390
rect 17200 -7160 17300 -4400
rect 17420 -4710 17520 -3050
rect 18100 -3170 18240 -2310
rect 18800 -2460 18900 -800
rect 19020 -1110 19120 550
rect 19700 430 19840 1290
rect 20400 1140 20500 1290
rect 20390 1130 20510 1140
rect 20390 1010 20400 1130
rect 20500 1010 20510 1130
rect 20390 1000 20510 1010
rect 19700 270 19710 430
rect 19830 270 19840 430
rect 19700 170 19840 270
rect 19700 -510 19710 170
rect 19830 -510 19840 170
rect 19010 -1120 19130 -1110
rect 19010 -1240 19020 -1120
rect 19120 -1240 19130 -1120
rect 19010 -1250 19130 -1240
rect 18790 -2470 18910 -2460
rect 18790 -2590 18800 -2470
rect 18900 -2590 18910 -2470
rect 18790 -2600 18910 -2590
rect 18100 -3330 18110 -3170
rect 18230 -3330 18240 -3170
rect 18100 -3430 18240 -3330
rect 18100 -4110 18110 -3430
rect 18230 -4110 18240 -3430
rect 18100 -4120 18240 -4110
rect 18800 -4260 18900 -2600
rect 19020 -2910 19120 -1250
rect 19700 -1370 19840 -510
rect 20400 -660 20500 1000
rect 20620 690 20720 1290
rect 20610 680 20730 690
rect 20610 560 20620 680
rect 20720 560 20730 680
rect 20610 550 20730 560
rect 20390 -670 20510 -660
rect 20390 -790 20400 -670
rect 20500 -790 20510 -670
rect 20390 -800 20510 -790
rect 19700 -1530 19710 -1370
rect 19830 -1530 19840 -1370
rect 19700 -1630 19840 -1530
rect 19700 -2310 19710 -1630
rect 19830 -2310 19840 -1630
rect 19010 -2920 19130 -2910
rect 19010 -3040 19020 -2920
rect 19120 -3040 19130 -2920
rect 19010 -3050 19130 -3040
rect 18790 -4270 18910 -4260
rect 18790 -4390 18800 -4270
rect 18900 -4390 18910 -4270
rect 18790 -4400 18910 -4390
rect 17410 -4720 17530 -4710
rect 17410 -4840 17420 -4720
rect 17520 -4840 17530 -4720
rect 17410 -4850 17530 -4840
rect 17420 -6760 17520 -4850
rect 18800 -5160 18900 -4400
rect 19020 -4710 19120 -3050
rect 19700 -3170 19840 -2310
rect 20400 -2460 20500 -800
rect 20620 -1110 20720 550
rect 21300 430 21440 1290
rect 22000 1140 22100 1290
rect 21990 1130 22110 1140
rect 21990 1010 22000 1130
rect 22100 1010 22110 1130
rect 21990 1000 22110 1010
rect 21300 270 21310 430
rect 21430 270 21440 430
rect 21300 170 21440 270
rect 21300 -510 21310 170
rect 21430 -510 21440 170
rect 20610 -1120 20730 -1110
rect 20610 -1240 20620 -1120
rect 20720 -1240 20730 -1120
rect 20610 -1250 20730 -1240
rect 20390 -2470 20510 -2460
rect 20390 -2590 20400 -2470
rect 20500 -2590 20510 -2470
rect 20390 -2600 20510 -2590
rect 19700 -3330 19710 -3170
rect 19830 -3330 19840 -3170
rect 19700 -3430 19840 -3330
rect 19700 -4110 19710 -3430
rect 19830 -4110 19840 -3430
rect 19700 -4120 19840 -4110
rect 20400 -4260 20500 -2600
rect 20620 -2910 20720 -1250
rect 21300 -1370 21440 -510
rect 22000 -660 22100 1000
rect 22220 690 22320 1290
rect 22210 680 22330 690
rect 22210 560 22220 680
rect 22320 560 22330 680
rect 22210 550 22330 560
rect 21990 -670 22110 -660
rect 21990 -790 22000 -670
rect 22100 -790 22110 -670
rect 21990 -800 22110 -790
rect 21300 -1530 21310 -1370
rect 21430 -1530 21440 -1370
rect 21300 -1630 21440 -1530
rect 21300 -2310 21310 -1630
rect 21430 -2310 21440 -1630
rect 20610 -2920 20730 -2910
rect 20610 -3040 20620 -2920
rect 20720 -3040 20730 -2920
rect 20610 -3050 20730 -3040
rect 20390 -4270 20510 -4260
rect 20390 -4390 20400 -4270
rect 20500 -4390 20510 -4270
rect 20390 -4400 20510 -4390
rect 19010 -4720 19130 -4710
rect 19010 -4840 19020 -4720
rect 19120 -4840 19130 -4720
rect 19010 -4850 19130 -4840
rect 18760 -5170 18940 -5160
rect 18760 -5350 18770 -5170
rect 18930 -5350 18940 -5170
rect 18760 -5360 18940 -5350
rect 18760 -5570 18940 -5560
rect 18760 -5750 18770 -5570
rect 18930 -5750 18940 -5570
rect 18760 -5760 18940 -5750
rect 17380 -6770 17560 -6760
rect 17380 -6950 17390 -6770
rect 17550 -6950 17560 -6770
rect 17380 -6960 17560 -6950
rect 17160 -7170 17340 -7160
rect 17160 -7350 17170 -7170
rect 17330 -7350 17340 -7170
rect 17160 -7360 17340 -7350
rect 17160 -7570 17340 -7560
rect 17160 -7750 17170 -7570
rect 17330 -7750 17340 -7570
rect 17160 -7760 17340 -7750
rect 15820 -8070 15960 -8060
rect 15820 -8190 15830 -8070
rect 15950 -8190 15960 -8070
rect 15820 -8200 15960 -8190
rect 15600 -8520 15740 -8510
rect 15600 -8640 15610 -8520
rect 15730 -8640 15740 -8520
rect 15600 -8650 15740 -8640
rect 14910 -8810 15040 -8800
rect 14910 -9470 14920 -8810
rect 15030 -9470 15040 -8810
rect 14910 -9480 15040 -9470
rect 15620 -10310 15720 -8650
rect 15840 -9860 15940 -8200
rect 17220 -8510 17320 -7760
rect 17440 -8060 17540 -6960
rect 17420 -8070 17560 -8060
rect 17420 -8190 17430 -8070
rect 17550 -8190 17560 -8070
rect 17420 -8200 17560 -8190
rect 17200 -8520 17340 -8510
rect 17200 -8640 17210 -8520
rect 17330 -8640 17340 -8520
rect 17200 -8650 17340 -8640
rect 16510 -8800 16640 -8790
rect 16510 -9480 16520 -8800
rect 16630 -9480 16640 -8800
rect 16510 -9560 16640 -9480
rect 16500 -9570 16650 -9560
rect 16500 -9730 16510 -9570
rect 16640 -9730 16650 -9570
rect 16500 -9740 16650 -9730
rect 15820 -9870 15960 -9860
rect 15820 -9990 15830 -9870
rect 15950 -9990 15960 -9870
rect 15820 -10000 15960 -9990
rect 15600 -10320 15740 -10310
rect 15600 -10440 15610 -10320
rect 15730 -10440 15740 -10320
rect 15600 -10450 15740 -10440
rect 14910 -10610 15040 -10600
rect 14910 -11270 14920 -10610
rect 15030 -11270 15040 -10610
rect 14910 -11280 15040 -11270
rect 14220 -11670 14360 -11660
rect 14220 -11790 14230 -11670
rect 14350 -11790 14360 -11670
rect 14220 -11800 14360 -11790
rect 14900 -11670 15040 -11660
rect 14900 -11790 14910 -11670
rect 15030 -11790 15040 -11670
rect 14900 -11800 15040 -11790
rect 14000 -13480 14140 -13470
rect 14000 -13600 14010 -13480
rect 14130 -13600 14140 -13480
rect 14000 -13610 14140 -13600
rect 13310 -14870 13320 -14210
rect 13430 -14870 13440 -14210
rect 13310 -14960 13440 -14870
rect 13280 -14970 13470 -14960
rect 13280 -15130 13290 -14970
rect 13460 -15130 13470 -14970
rect 13280 -15140 13470 -15130
rect 13310 -15290 13440 -15280
rect 13310 -15390 13330 -15290
rect 13430 -15390 13440 -15290
rect 14020 -15300 14120 -13610
rect 13310 -16010 13440 -15390
rect 14010 -15310 14130 -15300
rect 14010 -15410 14020 -15310
rect 14120 -15410 14130 -15310
rect 14010 -15420 14130 -15410
rect 13310 -16670 13320 -16010
rect 13430 -16670 13440 -16010
rect 13310 -16680 13440 -16670
rect 13310 -16780 13430 -16680
rect 13290 -16790 13460 -16780
rect 13290 -16950 13300 -16790
rect 13450 -16950 13460 -16790
rect 13290 -16960 13460 -16950
rect 12620 -17080 12760 -17070
rect 12620 -17200 12630 -17080
rect 12750 -17200 12760 -17080
rect 12620 -17210 12760 -17200
rect 13310 -17800 13430 -16960
rect 13310 -17810 13440 -17800
rect 13310 -18470 13320 -17810
rect 13430 -18470 13440 -17810
rect 13310 -18580 13440 -18470
rect 13290 -18590 13460 -18580
rect 13290 -18750 13300 -18590
rect 13450 -18750 13460 -18590
rect 13290 -18760 13460 -18750
rect 12400 -18880 12540 -18870
rect 12400 -19000 12410 -18880
rect 12530 -19000 12540 -18880
rect 12400 -19010 12540 -19000
rect 14240 -19320 14340 -11800
rect 14910 -12410 15040 -11800
rect 15620 -12110 15720 -10450
rect 15840 -11660 15940 -10000
rect 16510 -10600 16640 -9740
rect 17220 -10310 17320 -8650
rect 17440 -9860 17540 -8200
rect 18820 -8510 18920 -5760
rect 19020 -5960 19120 -4850
rect 18980 -5970 19160 -5960
rect 18980 -6150 18990 -5970
rect 19150 -6150 19160 -5970
rect 18980 -6160 19160 -6150
rect 19040 -8060 19140 -6160
rect 20400 -7160 20500 -4400
rect 20620 -4710 20720 -3050
rect 21300 -3170 21440 -2310
rect 22000 -2460 22100 -800
rect 22220 -1110 22320 550
rect 22900 430 23040 1290
rect 23600 1140 23700 1290
rect 23590 1130 23710 1140
rect 23590 1010 23600 1130
rect 23700 1010 23710 1130
rect 23590 1000 23710 1010
rect 22900 270 22910 430
rect 23030 270 23040 430
rect 22900 170 23040 270
rect 22900 -510 22910 170
rect 23030 -510 23040 170
rect 22210 -1120 22330 -1110
rect 22210 -1240 22220 -1120
rect 22320 -1240 22330 -1120
rect 22210 -1250 22330 -1240
rect 21990 -2470 22110 -2460
rect 21990 -2590 22000 -2470
rect 22100 -2590 22110 -2470
rect 21990 -2600 22110 -2590
rect 21300 -3330 21310 -3170
rect 21430 -3330 21440 -3170
rect 21300 -3430 21440 -3330
rect 21300 -4110 21310 -3430
rect 21430 -4110 21440 -3430
rect 21300 -4120 21440 -4110
rect 22000 -4260 22100 -2600
rect 22220 -2910 22320 -1250
rect 22900 -1370 23040 -510
rect 23600 -660 23700 1000
rect 23820 690 23920 1290
rect 23810 680 23930 690
rect 23810 560 23820 680
rect 23920 560 23930 680
rect 23810 550 23930 560
rect 23590 -670 23710 -660
rect 23590 -790 23600 -670
rect 23700 -790 23710 -670
rect 23590 -800 23710 -790
rect 22900 -1530 22910 -1370
rect 23030 -1530 23040 -1370
rect 22900 -1630 23040 -1530
rect 22900 -2310 22910 -1630
rect 23030 -2310 23040 -1630
rect 22210 -2920 22330 -2910
rect 22210 -3040 22220 -2920
rect 22320 -3040 22330 -2920
rect 22210 -3050 22330 -3040
rect 21990 -4270 22110 -4260
rect 21990 -4390 22000 -4270
rect 22100 -4390 22110 -4270
rect 21990 -4400 22110 -4390
rect 20610 -4720 20730 -4710
rect 20610 -4840 20620 -4720
rect 20720 -4840 20730 -4720
rect 20610 -4850 20730 -4840
rect 20620 -6760 20720 -4850
rect 22000 -5160 22100 -4400
rect 22220 -4710 22320 -3050
rect 22900 -3170 23040 -2310
rect 23600 -2460 23700 -800
rect 23820 -1110 23920 550
rect 24500 430 24640 1290
rect 24500 270 24510 430
rect 24630 270 24640 430
rect 24500 170 24640 270
rect 24500 -510 24510 170
rect 24630 -510 24640 170
rect 23810 -1120 23930 -1110
rect 23810 -1240 23820 -1120
rect 23920 -1240 23930 -1120
rect 23810 -1250 23930 -1240
rect 23590 -2470 23710 -2460
rect 23590 -2590 23600 -2470
rect 23700 -2590 23710 -2470
rect 23590 -2600 23710 -2590
rect 22900 -3330 22910 -3170
rect 23030 -3330 23040 -3170
rect 22900 -3430 23040 -3330
rect 22900 -4110 22910 -3430
rect 23030 -4110 23040 -3430
rect 22900 -4120 23040 -4110
rect 23600 -4260 23700 -2600
rect 23820 -2910 23920 -1250
rect 24500 -1370 24640 -510
rect 24500 -1530 24510 -1370
rect 24630 -1530 24640 -1370
rect 24500 -1630 24640 -1530
rect 24500 -2310 24510 -1630
rect 24630 -2310 24640 -1630
rect 23810 -2920 23930 -2910
rect 23810 -3040 23820 -2920
rect 23920 -3040 23930 -2920
rect 23810 -3050 23930 -3040
rect 23590 -4270 23710 -4260
rect 23590 -4390 23600 -4270
rect 23700 -4390 23710 -4270
rect 23590 -4400 23710 -4390
rect 22210 -4720 22330 -4710
rect 22210 -4840 22220 -4720
rect 22320 -4840 22330 -4720
rect 22210 -4850 22330 -4840
rect 21960 -5170 22140 -5160
rect 21960 -5350 21970 -5170
rect 22130 -5350 22140 -5170
rect 21960 -5360 22140 -5350
rect 21960 -5570 22140 -5560
rect 21960 -5750 21970 -5570
rect 22130 -5750 22140 -5570
rect 21960 -5760 22140 -5750
rect 20580 -6770 20760 -6760
rect 20580 -6950 20590 -6770
rect 20750 -6950 20760 -6770
rect 20580 -6960 20760 -6950
rect 20360 -7170 20540 -7160
rect 20360 -7350 20370 -7170
rect 20530 -7350 20540 -7170
rect 20360 -7360 20540 -7350
rect 20360 -7570 20540 -7560
rect 20360 -7750 20370 -7570
rect 20530 -7750 20540 -7570
rect 20360 -7760 20540 -7750
rect 19020 -8070 19160 -8060
rect 19020 -8190 19030 -8070
rect 19150 -8190 19160 -8070
rect 19020 -8200 19160 -8190
rect 18800 -8520 18940 -8510
rect 18800 -8640 18810 -8520
rect 18930 -8640 18940 -8520
rect 18800 -8650 18940 -8640
rect 18110 -8800 18240 -8790
rect 18110 -9480 18120 -8800
rect 18230 -9480 18240 -8800
rect 18110 -9560 18240 -9480
rect 18100 -9570 18250 -9560
rect 18100 -9730 18110 -9570
rect 18240 -9730 18250 -9570
rect 18100 -9740 18250 -9730
rect 17420 -9870 17560 -9860
rect 17420 -9990 17430 -9870
rect 17550 -9990 17560 -9870
rect 17420 -10000 17560 -9990
rect 17200 -10320 17340 -10310
rect 17200 -10440 17210 -10320
rect 17330 -10440 17340 -10320
rect 17200 -10450 17340 -10440
rect 16510 -11280 16520 -10600
rect 16630 -11280 16640 -10600
rect 16510 -11360 16640 -11280
rect 16500 -11370 16650 -11360
rect 16500 -11530 16510 -11370
rect 16640 -11530 16650 -11370
rect 16500 -11540 16650 -11530
rect 15820 -11670 15960 -11660
rect 15820 -11790 15830 -11670
rect 15950 -11790 15960 -11670
rect 15820 -11800 15960 -11790
rect 15600 -12120 15740 -12110
rect 15600 -12240 15610 -12120
rect 15730 -12240 15740 -12120
rect 15600 -12250 15740 -12240
rect 14910 -13070 14920 -12410
rect 15030 -13070 15040 -12410
rect 14910 -13160 15040 -13070
rect 14880 -13170 15070 -13160
rect 14880 -13330 14890 -13170
rect 15060 -13330 15070 -13170
rect 14880 -13340 15070 -13330
rect 14910 -14210 15040 -13340
rect 15620 -13910 15720 -12250
rect 15840 -13460 15940 -11800
rect 16510 -12400 16640 -11540
rect 17220 -12110 17320 -10450
rect 17440 -11660 17540 -10000
rect 18110 -10600 18240 -9740
rect 18820 -10310 18920 -8650
rect 19040 -9860 19140 -8200
rect 20420 -8510 20520 -7760
rect 20640 -8060 20740 -6960
rect 20620 -8070 20760 -8060
rect 20620 -8190 20630 -8070
rect 20750 -8190 20760 -8070
rect 20620 -8200 20760 -8190
rect 20400 -8520 20540 -8510
rect 20400 -8640 20410 -8520
rect 20530 -8640 20540 -8520
rect 20400 -8650 20540 -8640
rect 19710 -8800 19840 -8790
rect 19710 -9480 19720 -8800
rect 19830 -9480 19840 -8800
rect 19710 -9560 19840 -9480
rect 19700 -9570 19850 -9560
rect 19700 -9730 19710 -9570
rect 19840 -9730 19850 -9570
rect 19700 -9740 19850 -9730
rect 19020 -9870 19160 -9860
rect 19020 -9990 19030 -9870
rect 19150 -9990 19160 -9870
rect 19020 -10000 19160 -9990
rect 18800 -10320 18940 -10310
rect 18800 -10440 18810 -10320
rect 18930 -10440 18940 -10320
rect 18800 -10450 18940 -10440
rect 18110 -11280 18120 -10600
rect 18230 -11280 18240 -10600
rect 18110 -11360 18240 -11280
rect 18100 -11370 18250 -11360
rect 18100 -11530 18110 -11370
rect 18240 -11530 18250 -11370
rect 18100 -11540 18250 -11530
rect 17420 -11670 17560 -11660
rect 17420 -11790 17430 -11670
rect 17550 -11790 17560 -11670
rect 17420 -11800 17560 -11790
rect 17200 -12120 17340 -12110
rect 17200 -12240 17210 -12120
rect 17330 -12240 17340 -12120
rect 17200 -12250 17340 -12240
rect 16510 -13080 16520 -12400
rect 16630 -13080 16640 -12400
rect 16510 -13160 16640 -13080
rect 16500 -13170 16650 -13160
rect 16500 -13330 16510 -13170
rect 16640 -13330 16650 -13170
rect 16500 -13340 16650 -13330
rect 15820 -13470 15960 -13460
rect 15820 -13590 15830 -13470
rect 15950 -13590 15960 -13470
rect 15820 -13600 15960 -13590
rect 15600 -13920 15740 -13910
rect 15600 -14040 15610 -13920
rect 15730 -14040 15740 -13920
rect 15600 -14050 15740 -14040
rect 14910 -14870 14920 -14210
rect 15030 -14870 15040 -14210
rect 14910 -14960 15040 -14870
rect 14880 -14970 15070 -14960
rect 14880 -15130 14890 -14970
rect 15060 -15130 15070 -14970
rect 14880 -15140 15070 -15130
rect 14910 -15290 15040 -15280
rect 14910 -15390 14930 -15290
rect 15030 -15390 15040 -15290
rect 14910 -16010 15040 -15390
rect 15620 -15710 15720 -14050
rect 15840 -15260 15940 -13600
rect 16510 -14200 16640 -13340
rect 17220 -13910 17320 -12250
rect 17440 -13460 17540 -11800
rect 18110 -12400 18240 -11540
rect 18820 -12110 18920 -10450
rect 19040 -11660 19140 -10000
rect 19710 -10600 19840 -9740
rect 20420 -10310 20520 -8650
rect 20640 -9860 20740 -8200
rect 22020 -8510 22120 -5760
rect 22220 -5960 22320 -4850
rect 22180 -5970 22360 -5960
rect 22180 -6150 22190 -5970
rect 22350 -6150 22360 -5970
rect 22180 -6160 22360 -6150
rect 22240 -8060 22340 -6160
rect 23600 -7160 23700 -4400
rect 23820 -4710 23920 -3050
rect 24500 -3170 24640 -2310
rect 25200 -2460 25300 1290
rect 25190 -2470 25310 -2460
rect 25190 -2590 25200 -2470
rect 25300 -2590 25310 -2470
rect 25190 -2600 25310 -2590
rect 24500 -3330 24510 -3170
rect 24630 -3330 24640 -3170
rect 24500 -3430 24640 -3330
rect 24500 -4110 24510 -3430
rect 24630 -4110 24640 -3430
rect 24500 -4120 24640 -4110
rect 25200 -4260 25300 -2600
rect 25420 -2910 25520 1290
rect 26100 430 26240 1290
rect 26800 1140 26900 1290
rect 26790 1130 26910 1140
rect 26790 1010 26800 1130
rect 26900 1010 26910 1130
rect 26790 1000 26910 1010
rect 26100 270 26110 430
rect 26230 270 26240 430
rect 26100 170 26240 270
rect 26100 -510 26110 170
rect 26230 -510 26240 170
rect 26100 -1370 26240 -510
rect 26800 -660 26900 1000
rect 27020 690 27120 1290
rect 27010 680 27130 690
rect 27010 560 27020 680
rect 27120 560 27130 680
rect 27010 550 27130 560
rect 26790 -670 26910 -660
rect 26790 -790 26800 -670
rect 26900 -790 26910 -670
rect 26790 -800 26910 -790
rect 26100 -1530 26110 -1370
rect 26230 -1530 26240 -1370
rect 26100 -1630 26240 -1530
rect 26100 -2310 26110 -1630
rect 26230 -2310 26240 -1630
rect 25410 -2920 25530 -2910
rect 25410 -3040 25420 -2920
rect 25520 -3040 25530 -2920
rect 25410 -3050 25530 -3040
rect 25190 -4270 25310 -4260
rect 25190 -4390 25200 -4270
rect 25300 -4390 25310 -4270
rect 25190 -4400 25310 -4390
rect 23810 -4720 23930 -4710
rect 23810 -4840 23820 -4720
rect 23920 -4840 23930 -4720
rect 23810 -4850 23930 -4840
rect 23820 -6760 23920 -4850
rect 25200 -5160 25300 -4400
rect 25420 -4710 25520 -3050
rect 26100 -3170 26240 -2310
rect 26800 -2460 26900 -800
rect 27020 -1110 27120 550
rect 27700 430 27840 1290
rect 28400 1140 28500 1290
rect 28391 1130 28510 1140
rect 28391 1010 28400 1130
rect 28500 1010 28510 1130
rect 28391 1000 28510 1010
rect 27700 250 27710 430
rect 27830 250 27840 430
rect 27700 170 27840 250
rect 27700 -510 27710 170
rect 27830 -510 27840 170
rect 27010 -1120 27130 -1110
rect 27010 -1240 27020 -1120
rect 27120 -1240 27130 -1120
rect 27010 -1250 27130 -1240
rect 26791 -2470 26910 -2460
rect 26791 -2590 26800 -2470
rect 26900 -2590 26910 -2470
rect 26791 -2600 26910 -2590
rect 26100 -3330 26110 -3170
rect 26230 -3330 26240 -3170
rect 26100 -3430 26240 -3330
rect 26100 -4110 26110 -3430
rect 26230 -4110 26240 -3430
rect 26100 -4120 26240 -4110
rect 26800 -4260 26900 -2600
rect 27020 -2910 27120 -1250
rect 27700 -1370 27840 -510
rect 28400 -660 28500 1000
rect 28620 690 28720 1290
rect 28611 680 28730 690
rect 28611 560 28620 680
rect 28720 560 28730 680
rect 28611 550 28730 560
rect 28391 -670 28510 -660
rect 28391 -790 28400 -670
rect 28500 -790 28510 -670
rect 28391 -800 28510 -790
rect 27700 -1550 27710 -1370
rect 27830 -1550 27840 -1370
rect 27700 -1630 27840 -1550
rect 27700 -2310 27710 -1630
rect 27830 -2310 27840 -1630
rect 27011 -2920 27130 -2910
rect 27011 -3040 27020 -2920
rect 27120 -3040 27130 -2920
rect 27011 -3050 27130 -3040
rect 26791 -4270 26910 -4260
rect 26791 -4390 26800 -4270
rect 26900 -4390 26910 -4270
rect 26791 -4400 26910 -4390
rect 25410 -4720 25530 -4710
rect 25410 -4840 25420 -4720
rect 25520 -4840 25530 -4720
rect 25410 -4850 25530 -4840
rect 25160 -5170 25340 -5160
rect 25160 -5350 25170 -5170
rect 25330 -5350 25340 -5170
rect 25160 -5360 25340 -5350
rect 25160 -5570 25340 -5560
rect 25160 -5750 25170 -5570
rect 25330 -5750 25340 -5570
rect 25160 -5760 25340 -5750
rect 23780 -6770 23960 -6760
rect 23780 -6950 23790 -6770
rect 23950 -6950 23960 -6770
rect 23780 -6960 23960 -6950
rect 23560 -7170 23740 -7160
rect 23560 -7350 23570 -7170
rect 23730 -7350 23740 -7170
rect 23560 -7360 23740 -7350
rect 23560 -7570 23740 -7560
rect 23560 -7750 23570 -7570
rect 23730 -7750 23740 -7570
rect 23560 -7760 23740 -7750
rect 22220 -8070 22360 -8060
rect 22220 -8190 22230 -8070
rect 22350 -8190 22360 -8070
rect 22220 -8200 22360 -8190
rect 22000 -8520 22140 -8510
rect 22000 -8640 22010 -8520
rect 22130 -8640 22140 -8520
rect 22000 -8650 22140 -8640
rect 21310 -8800 21440 -8790
rect 21310 -9480 21320 -8800
rect 21430 -9480 21440 -8800
rect 21310 -9560 21440 -9480
rect 21300 -9570 21450 -9560
rect 21300 -9730 21310 -9570
rect 21440 -9730 21450 -9570
rect 21300 -9740 21450 -9730
rect 20620 -9870 20760 -9860
rect 20620 -9990 20630 -9870
rect 20750 -9990 20760 -9870
rect 20620 -10000 20760 -9990
rect 20400 -10320 20540 -10310
rect 20400 -10440 20410 -10320
rect 20530 -10440 20540 -10320
rect 20400 -10450 20540 -10440
rect 19710 -11280 19720 -10600
rect 19830 -11280 19840 -10600
rect 19710 -11360 19840 -11280
rect 19700 -11370 19850 -11360
rect 19700 -11530 19710 -11370
rect 19840 -11530 19850 -11370
rect 19700 -11540 19850 -11530
rect 19020 -11670 19160 -11660
rect 19020 -11790 19030 -11670
rect 19150 -11790 19160 -11670
rect 19020 -11800 19160 -11790
rect 18800 -12120 18940 -12110
rect 18800 -12240 18810 -12120
rect 18930 -12240 18940 -12120
rect 18800 -12250 18940 -12240
rect 18110 -13080 18120 -12400
rect 18230 -13080 18240 -12400
rect 18110 -13160 18240 -13080
rect 18100 -13170 18250 -13160
rect 18100 -13330 18110 -13170
rect 18240 -13330 18250 -13170
rect 18100 -13340 18250 -13330
rect 17420 -13470 17560 -13460
rect 17420 -13590 17430 -13470
rect 17550 -13590 17560 -13470
rect 17420 -13600 17560 -13590
rect 17200 -13920 17340 -13910
rect 17200 -14040 17210 -13920
rect 17330 -14040 17340 -13920
rect 17200 -14050 17340 -14040
rect 16510 -14880 16520 -14200
rect 16630 -14880 16640 -14200
rect 16510 -14960 16640 -14880
rect 16500 -14970 16650 -14960
rect 16500 -15130 16510 -14970
rect 16640 -15130 16650 -14970
rect 16500 -15140 16650 -15130
rect 15820 -15270 15960 -15260
rect 15820 -15390 15830 -15270
rect 15950 -15390 15960 -15270
rect 15820 -15400 15960 -15390
rect 15600 -15720 15740 -15710
rect 15600 -15840 15610 -15720
rect 15730 -15840 15740 -15720
rect 15600 -15850 15740 -15840
rect 14910 -16670 14920 -16010
rect 15030 -16670 15040 -16010
rect 14910 -16680 15040 -16670
rect 14910 -16780 15030 -16680
rect 14890 -16790 15060 -16780
rect 14890 -16950 14900 -16790
rect 15050 -16950 15060 -16790
rect 14890 -16960 15060 -16950
rect 14910 -17800 15030 -16960
rect 15620 -17510 15720 -15850
rect 15840 -17060 15940 -15400
rect 16510 -16000 16640 -15140
rect 17220 -15710 17320 -14050
rect 17440 -15260 17540 -13600
rect 18110 -14200 18240 -13340
rect 18820 -13910 18920 -12250
rect 19040 -13460 19140 -11800
rect 19710 -12400 19840 -11540
rect 20420 -12110 20520 -10450
rect 20640 -11660 20740 -10000
rect 21310 -10600 21440 -9740
rect 22020 -10310 22120 -8650
rect 22240 -9860 22340 -8200
rect 23620 -8510 23720 -7760
rect 23840 -8060 23940 -6960
rect 23820 -8070 23960 -8060
rect 23820 -8190 23830 -8070
rect 23950 -8190 23960 -8070
rect 23820 -8200 23960 -8190
rect 23600 -8520 23740 -8510
rect 23600 -8640 23610 -8520
rect 23730 -8640 23740 -8520
rect 23600 -8650 23740 -8640
rect 22910 -8800 23040 -8790
rect 22910 -9480 22920 -8800
rect 23030 -9480 23040 -8800
rect 22910 -9560 23040 -9480
rect 22900 -9570 23050 -9560
rect 22900 -9730 22910 -9570
rect 23040 -9730 23050 -9570
rect 22900 -9740 23050 -9730
rect 22220 -9870 22360 -9860
rect 22220 -9990 22230 -9870
rect 22350 -9990 22360 -9870
rect 22220 -10000 22360 -9990
rect 22000 -10320 22140 -10310
rect 22000 -10440 22010 -10320
rect 22130 -10440 22140 -10320
rect 22000 -10450 22140 -10440
rect 21310 -11280 21320 -10600
rect 21430 -11280 21440 -10600
rect 21310 -11360 21440 -11280
rect 21300 -11370 21450 -11360
rect 21300 -11530 21310 -11370
rect 21440 -11530 21450 -11370
rect 21300 -11540 21450 -11530
rect 20620 -11670 20760 -11660
rect 20620 -11790 20630 -11670
rect 20750 -11790 20760 -11670
rect 20620 -11800 20760 -11790
rect 20400 -12120 20540 -12110
rect 20400 -12240 20410 -12120
rect 20530 -12240 20540 -12120
rect 20400 -12250 20540 -12240
rect 19710 -13080 19720 -12400
rect 19830 -13080 19840 -12400
rect 19710 -13160 19840 -13080
rect 19700 -13170 19850 -13160
rect 19700 -13330 19710 -13170
rect 19840 -13330 19850 -13170
rect 19700 -13340 19850 -13330
rect 19020 -13470 19160 -13460
rect 19020 -13590 19030 -13470
rect 19150 -13590 19160 -13470
rect 19020 -13600 19160 -13590
rect 18800 -13920 18940 -13910
rect 18800 -14040 18810 -13920
rect 18930 -14040 18940 -13920
rect 18800 -14050 18940 -14040
rect 18110 -14880 18120 -14200
rect 18230 -14880 18240 -14200
rect 18110 -14960 18240 -14880
rect 18100 -14970 18250 -14960
rect 18100 -15130 18110 -14970
rect 18240 -15130 18250 -14970
rect 18100 -15140 18250 -15130
rect 17420 -15270 17560 -15260
rect 17420 -15390 17430 -15270
rect 17550 -15390 17560 -15270
rect 17420 -15400 17560 -15390
rect 17200 -15720 17340 -15710
rect 17200 -15840 17210 -15720
rect 17330 -15840 17340 -15720
rect 17200 -15850 17340 -15840
rect 16510 -16680 16520 -16000
rect 16630 -16680 16640 -16000
rect 16510 -16760 16640 -16680
rect 16500 -16770 16650 -16760
rect 16500 -16930 16510 -16770
rect 16640 -16930 16650 -16770
rect 16500 -16940 16650 -16930
rect 15820 -17070 15960 -17060
rect 15820 -17190 15830 -17070
rect 15950 -17190 15960 -17070
rect 15820 -17200 15960 -17190
rect 15600 -17520 15740 -17510
rect 15600 -17640 15610 -17520
rect 15730 -17640 15740 -17520
rect 15600 -17650 15740 -17640
rect 14910 -17810 15040 -17800
rect 14910 -18470 14920 -17810
rect 15030 -18470 15040 -17810
rect 14910 -18580 15040 -18470
rect 14890 -18590 15060 -18580
rect 14890 -18750 14900 -18590
rect 15050 -18750 15060 -18590
rect 14890 -18760 15060 -18750
rect 15620 -19310 15720 -17650
rect 15840 -18860 15940 -17200
rect 16510 -17800 16640 -16940
rect 17220 -17510 17320 -15850
rect 17440 -17060 17540 -15400
rect 18110 -16000 18240 -15140
rect 18820 -15710 18920 -14050
rect 19040 -15260 19140 -13600
rect 19710 -14200 19840 -13340
rect 20420 -13910 20520 -12250
rect 20640 -13460 20740 -11800
rect 21310 -12400 21440 -11540
rect 22020 -12110 22120 -10450
rect 22240 -11660 22340 -10000
rect 22910 -10600 23040 -9740
rect 23620 -10310 23720 -8650
rect 23840 -9860 23940 -8200
rect 25220 -8510 25320 -5760
rect 25420 -5960 25520 -4850
rect 25380 -5970 25560 -5960
rect 25380 -6150 25390 -5970
rect 25550 -6150 25560 -5970
rect 25380 -6160 25560 -6150
rect 25440 -8060 25540 -6160
rect 26800 -7160 26900 -4400
rect 27020 -4710 27120 -3050
rect 27700 -3170 27840 -2310
rect 28400 -2460 28500 -800
rect 28620 -1110 28720 550
rect 29300 430 29440 1290
rect 29300 250 29310 430
rect 29430 250 29440 430
rect 29300 170 29440 250
rect 29300 -510 29310 170
rect 29430 -510 29440 170
rect 28611 -1120 28730 -1110
rect 28611 -1240 28620 -1120
rect 28720 -1240 28730 -1120
rect 28611 -1250 28730 -1240
rect 28390 -2470 28510 -2460
rect 28390 -2590 28400 -2470
rect 28500 -2590 28510 -2470
rect 28390 -2600 28510 -2590
rect 27700 -3350 27710 -3170
rect 27830 -3350 27840 -3170
rect 27700 -3430 27840 -3350
rect 27700 -4110 27710 -3430
rect 27830 -4110 27840 -3430
rect 27011 -4720 27130 -4710
rect 27011 -4840 27020 -4720
rect 27120 -4840 27130 -4720
rect 27011 -4850 27130 -4840
rect 27020 -6760 27120 -4850
rect 27700 -5960 27840 -4110
rect 28400 -4260 28500 -2600
rect 28620 -2910 28720 -1250
rect 29300 -1370 29440 -510
rect 29300 -1550 29310 -1370
rect 29430 -1550 29440 -1370
rect 29300 -1630 29440 -1550
rect 29300 -2310 29310 -1630
rect 29430 -2310 29440 -1630
rect 28610 -2920 28730 -2910
rect 28610 -3040 28620 -2920
rect 28720 -3040 28730 -2920
rect 28610 -3050 28730 -3040
rect 28390 -4270 28510 -4260
rect 28390 -4390 28400 -4270
rect 28500 -4390 28510 -4270
rect 28390 -4400 28510 -4390
rect 28400 -5160 28500 -4400
rect 28620 -4710 28720 -3050
rect 29300 -3170 29440 -2310
rect 30900 2230 31040 2240
rect 30900 2050 30910 2230
rect 31030 2050 31040 2230
rect 30900 1970 31040 2050
rect 30900 1290 30910 1970
rect 31030 1290 31040 1970
rect 30900 430 31040 1290
rect 30900 250 30910 430
rect 31030 250 31040 430
rect 30900 170 31040 250
rect 30900 -510 30910 170
rect 31030 -510 31040 170
rect 30900 -1370 31040 -510
rect 31600 -1110 31700 3540
rect 31820 690 31920 2810
rect 34890 2760 35060 2770
rect 34890 2600 34900 2760
rect 35050 2600 35060 2760
rect 34890 2590 35060 2600
rect 33290 2530 33460 2540
rect 33290 2370 33300 2530
rect 33450 2370 33460 2530
rect 33290 2360 33460 2370
rect 32500 1970 32640 1980
rect 32500 1290 32510 1970
rect 32630 1290 32640 1970
rect 32500 1130 32640 1290
rect 32500 1010 32510 1130
rect 32630 1010 32640 1130
rect 32500 1000 32640 1010
rect 31810 680 31930 690
rect 31810 560 31820 680
rect 31920 560 31930 680
rect 31810 550 31930 560
rect 33310 430 33440 2360
rect 34100 1970 34240 1980
rect 34100 1290 34110 1970
rect 34230 1290 34240 1970
rect 34100 1130 34240 1290
rect 34910 1140 35040 2590
rect 35700 1970 35840 1980
rect 35700 1290 35710 1970
rect 35830 1290 35840 1970
rect 34100 1010 34110 1130
rect 34230 1010 34240 1130
rect 34100 1000 34240 1010
rect 34900 1130 35050 1140
rect 34900 1010 34910 1130
rect 35040 1010 35050 1130
rect 34900 1000 35050 1010
rect 35700 1130 35840 1290
rect 35700 1010 35710 1130
rect 35830 1010 35840 1130
rect 35700 1000 35840 1010
rect 33290 420 33460 430
rect 33290 260 33300 420
rect 33450 260 33460 420
rect 33290 250 33460 260
rect 32500 170 32640 180
rect 32500 -510 32510 170
rect 32630 -510 32640 170
rect 32500 -520 32640 -510
rect 34100 170 34240 180
rect 34100 -510 34110 170
rect 34230 -510 34240 170
rect 34100 -520 34240 -510
rect 31590 -1120 31710 -1110
rect 31590 -1240 31600 -1120
rect 31700 -1240 31710 -1120
rect 31590 -1250 31710 -1240
rect 30900 -1550 30910 -1370
rect 31030 -1550 31040 -1370
rect 30900 -1630 31040 -1550
rect 30900 -2310 30910 -1630
rect 31030 -2310 31040 -1630
rect 29990 -2470 30110 -2460
rect 29990 -2590 30000 -2470
rect 30100 -2590 30110 -2470
rect 29990 -2600 30110 -2590
rect 29300 -3350 29310 -3170
rect 29430 -3350 29440 -3170
rect 29300 -3430 29440 -3350
rect 29300 -4110 29310 -3430
rect 29430 -4110 29440 -3430
rect 28610 -4720 28730 -4710
rect 28610 -4840 28620 -4720
rect 28720 -4840 28730 -4720
rect 28610 -4850 28730 -4840
rect 28360 -5170 28540 -5160
rect 28360 -5350 28370 -5170
rect 28530 -5350 28540 -5170
rect 28360 -5360 28540 -5350
rect 28360 -5570 28540 -5560
rect 28360 -5750 28370 -5570
rect 28530 -5750 28540 -5570
rect 28360 -5760 28540 -5750
rect 27680 -5970 27860 -5960
rect 27680 -6150 27690 -5970
rect 27850 -6150 27860 -5970
rect 27680 -6160 27860 -6150
rect 26980 -6770 27160 -6760
rect 26980 -6950 26990 -6770
rect 27150 -6950 27160 -6770
rect 26980 -6960 27160 -6950
rect 26760 -7170 26940 -7160
rect 26760 -7350 26770 -7170
rect 26930 -7350 26940 -7170
rect 26760 -7360 26940 -7350
rect 26760 -7570 26940 -7560
rect 26760 -7750 26770 -7570
rect 26930 -7750 26940 -7570
rect 26760 -7760 26940 -7750
rect 25420 -8070 25560 -8060
rect 25420 -8190 25430 -8070
rect 25550 -8190 25560 -8070
rect 25420 -8200 25560 -8190
rect 25200 -8520 25340 -8510
rect 25200 -8640 25210 -8520
rect 25330 -8640 25340 -8520
rect 25200 -8650 25340 -8640
rect 24510 -8800 24640 -8790
rect 24510 -9480 24520 -8800
rect 24630 -9480 24640 -8800
rect 24510 -9560 24640 -9480
rect 24500 -9570 24650 -9560
rect 24500 -9730 24510 -9570
rect 24640 -9730 24650 -9570
rect 24500 -9740 24650 -9730
rect 23820 -9870 23960 -9860
rect 23820 -9990 23830 -9870
rect 23950 -9990 23960 -9870
rect 23820 -10000 23960 -9990
rect 23600 -10320 23740 -10310
rect 23600 -10440 23610 -10320
rect 23730 -10440 23740 -10320
rect 23600 -10450 23740 -10440
rect 22910 -11280 22920 -10600
rect 23030 -11280 23040 -10600
rect 22910 -11360 23040 -11280
rect 22900 -11370 23050 -11360
rect 22900 -11530 22910 -11370
rect 23040 -11530 23050 -11370
rect 22900 -11540 23050 -11530
rect 22220 -11670 22360 -11660
rect 22220 -11790 22230 -11670
rect 22350 -11790 22360 -11670
rect 22220 -11800 22360 -11790
rect 22000 -12120 22140 -12110
rect 22000 -12240 22010 -12120
rect 22130 -12240 22140 -12120
rect 22000 -12250 22140 -12240
rect 21310 -13080 21320 -12400
rect 21430 -13080 21440 -12400
rect 21310 -13160 21440 -13080
rect 21300 -13170 21450 -13160
rect 21300 -13330 21310 -13170
rect 21440 -13330 21450 -13170
rect 21300 -13340 21450 -13330
rect 20620 -13470 20760 -13460
rect 20620 -13590 20630 -13470
rect 20750 -13590 20760 -13470
rect 20620 -13600 20760 -13590
rect 20400 -13920 20540 -13910
rect 20400 -14040 20410 -13920
rect 20530 -14040 20540 -13920
rect 20400 -14050 20540 -14040
rect 19710 -14880 19720 -14200
rect 19830 -14880 19840 -14200
rect 19710 -14960 19840 -14880
rect 19700 -14970 19850 -14960
rect 19700 -15130 19710 -14970
rect 19840 -15130 19850 -14970
rect 19700 -15140 19850 -15130
rect 19020 -15270 19160 -15260
rect 19020 -15390 19030 -15270
rect 19150 -15390 19160 -15270
rect 19020 -15400 19160 -15390
rect 18800 -15720 18940 -15710
rect 18800 -15840 18810 -15720
rect 18930 -15840 18940 -15720
rect 18800 -15850 18940 -15840
rect 18110 -16680 18120 -16000
rect 18230 -16680 18240 -16000
rect 18110 -16760 18240 -16680
rect 18100 -16770 18250 -16760
rect 18100 -16930 18110 -16770
rect 18240 -16930 18250 -16770
rect 18100 -16940 18250 -16930
rect 17420 -17070 17560 -17060
rect 17420 -17190 17430 -17070
rect 17550 -17190 17560 -17070
rect 17420 -17200 17560 -17190
rect 17200 -17520 17340 -17510
rect 17200 -17640 17210 -17520
rect 17330 -17640 17340 -17520
rect 17200 -17650 17340 -17640
rect 16510 -18480 16520 -17800
rect 16630 -18480 16640 -17800
rect 16510 -18560 16640 -18480
rect 16500 -18570 16650 -18560
rect 16500 -18730 16510 -18570
rect 16640 -18730 16650 -18570
rect 16500 -18740 16650 -18730
rect 15820 -18870 15960 -18860
rect 15820 -18990 15830 -18870
rect 15950 -18990 15960 -18870
rect 15820 -19000 15960 -18990
rect 15600 -19320 15740 -19310
rect 13310 -19440 15040 -19320
rect 11710 -19610 11840 -19600
rect 11710 -20270 11720 -19610
rect 11830 -20270 11840 -19610
rect 11710 -20280 11840 -20270
rect 13310 -19610 13440 -19440
rect 13310 -20270 13320 -19610
rect 13430 -20270 13440 -19610
rect 13310 -20280 13440 -20270
rect 14910 -19610 15040 -19440
rect 15600 -19440 15610 -19320
rect 15730 -19440 15740 -19320
rect 15600 -19450 15740 -19440
rect 14910 -20270 14920 -19610
rect 15030 -20270 15040 -19610
rect 14910 -20280 15040 -20270
rect 10120 -20550 10130 -20390
rect 10230 -20550 10240 -20390
rect 9420 -21110 9560 -21100
rect 9420 -21230 9430 -21110
rect 9550 -21230 9560 -21110
rect 9420 -21240 9560 -21230
rect 10120 -21410 10240 -20550
rect 11030 -20560 11150 -20380
rect 10120 -22070 10130 -21410
rect 10230 -22070 10240 -21410
rect 10120 -22190 10240 -22070
rect 11040 -22180 11140 -20560
rect 15620 -21110 15720 -19450
rect 15840 -20660 15940 -19000
rect 16510 -19600 16640 -18740
rect 17220 -19310 17320 -17650
rect 17440 -18860 17540 -17200
rect 18110 -17800 18240 -16940
rect 18820 -17510 18920 -15850
rect 19040 -17060 19140 -15400
rect 19710 -16000 19840 -15140
rect 20420 -15710 20520 -14050
rect 20640 -15260 20740 -13600
rect 21310 -14200 21440 -13340
rect 22020 -13910 22120 -12250
rect 22240 -13460 22340 -11800
rect 22910 -12400 23040 -11540
rect 23620 -12110 23720 -10450
rect 23840 -11660 23940 -10000
rect 24510 -10600 24640 -9740
rect 25220 -10310 25320 -8650
rect 25440 -9860 25540 -8200
rect 26820 -8510 26920 -7760
rect 27040 -8060 27140 -6960
rect 27020 -8070 27160 -8060
rect 27020 -8190 27030 -8070
rect 27150 -8190 27160 -8070
rect 27020 -8200 27160 -8190
rect 26800 -8520 26940 -8510
rect 26800 -8640 26810 -8520
rect 26930 -8640 26940 -8520
rect 26800 -8650 26940 -8640
rect 26110 -8800 26240 -8790
rect 26110 -9480 26120 -8800
rect 26230 -9480 26240 -8800
rect 26110 -9560 26240 -9480
rect 26100 -9570 26250 -9560
rect 26100 -9730 26110 -9570
rect 26240 -9730 26250 -9570
rect 26100 -9740 26250 -9730
rect 25420 -9870 25560 -9860
rect 25420 -9990 25430 -9870
rect 25550 -9990 25560 -9870
rect 25420 -10000 25560 -9990
rect 25200 -10320 25340 -10310
rect 25200 -10440 25210 -10320
rect 25330 -10440 25340 -10320
rect 25200 -10450 25340 -10440
rect 24510 -11280 24520 -10600
rect 24630 -11280 24640 -10600
rect 24510 -11360 24640 -11280
rect 24500 -11370 24650 -11360
rect 24500 -11530 24510 -11370
rect 24640 -11530 24650 -11370
rect 24500 -11540 24650 -11530
rect 23820 -11670 23960 -11660
rect 23820 -11790 23830 -11670
rect 23950 -11790 23960 -11670
rect 23820 -11800 23960 -11790
rect 23600 -12120 23740 -12110
rect 23600 -12240 23610 -12120
rect 23730 -12240 23740 -12120
rect 23600 -12250 23740 -12240
rect 22910 -13080 22920 -12400
rect 23030 -13080 23040 -12400
rect 22910 -13160 23040 -13080
rect 22900 -13170 23050 -13160
rect 22900 -13330 22910 -13170
rect 23040 -13330 23050 -13170
rect 22900 -13340 23050 -13330
rect 22220 -13470 22360 -13460
rect 22220 -13590 22230 -13470
rect 22350 -13590 22360 -13470
rect 22220 -13600 22360 -13590
rect 22000 -13920 22140 -13910
rect 22000 -14040 22010 -13920
rect 22130 -14040 22140 -13920
rect 22000 -14050 22140 -14040
rect 21310 -14880 21320 -14200
rect 21430 -14880 21440 -14200
rect 21310 -14960 21440 -14880
rect 21300 -14970 21450 -14960
rect 21300 -15130 21310 -14970
rect 21440 -15130 21450 -14970
rect 21300 -15140 21450 -15130
rect 20620 -15270 20760 -15260
rect 20620 -15390 20630 -15270
rect 20750 -15390 20760 -15270
rect 20620 -15400 20760 -15390
rect 20400 -15720 20540 -15710
rect 20400 -15840 20410 -15720
rect 20530 -15840 20540 -15720
rect 20400 -15850 20540 -15840
rect 19710 -16680 19720 -16000
rect 19830 -16680 19840 -16000
rect 19710 -16760 19840 -16680
rect 19700 -16770 19850 -16760
rect 19700 -16930 19710 -16770
rect 19840 -16930 19850 -16770
rect 19700 -16940 19850 -16930
rect 19020 -17070 19160 -17060
rect 19020 -17190 19030 -17070
rect 19150 -17190 19160 -17070
rect 19020 -17200 19160 -17190
rect 18800 -17520 18940 -17510
rect 18800 -17640 18810 -17520
rect 18930 -17640 18940 -17520
rect 18800 -17650 18940 -17640
rect 18110 -18480 18120 -17800
rect 18230 -18480 18240 -17800
rect 18110 -18560 18240 -18480
rect 18100 -18570 18250 -18560
rect 18100 -18730 18110 -18570
rect 18240 -18730 18250 -18570
rect 18100 -18740 18250 -18730
rect 17420 -18870 17560 -18860
rect 17420 -18990 17430 -18870
rect 17550 -18990 17560 -18870
rect 17420 -19000 17560 -18990
rect 17200 -19320 17340 -19310
rect 17200 -19440 17210 -19320
rect 17330 -19440 17340 -19320
rect 17200 -19450 17340 -19440
rect 16510 -20280 16520 -19600
rect 16630 -20280 16640 -19600
rect 16510 -20360 16640 -20280
rect 16500 -20370 16650 -20360
rect 16500 -20530 16510 -20370
rect 16640 -20530 16650 -20370
rect 16500 -20540 16650 -20530
rect 15820 -20670 15960 -20660
rect 15820 -20790 15830 -20670
rect 15950 -20790 15960 -20670
rect 15820 -20800 15960 -20790
rect 15600 -21120 15740 -21110
rect 15600 -21240 15610 -21120
rect 15730 -21240 15740 -21120
rect 15600 -21250 15740 -21240
rect 15620 -21370 15720 -21250
rect 15840 -21370 15940 -20800
rect 16510 -21400 16640 -20540
rect 17220 -21110 17320 -19450
rect 17440 -20660 17540 -19000
rect 18110 -19600 18240 -18740
rect 18820 -19310 18920 -17650
rect 19040 -18860 19140 -17200
rect 19710 -17800 19840 -16940
rect 20420 -17510 20520 -15850
rect 20640 -17060 20740 -15400
rect 21310 -16000 21440 -15140
rect 22020 -15710 22120 -14050
rect 22240 -15260 22340 -13600
rect 22910 -14200 23040 -13340
rect 23620 -13910 23720 -12250
rect 23840 -13460 23940 -11800
rect 24510 -12400 24640 -11540
rect 25220 -12110 25320 -10450
rect 25440 -11660 25540 -10000
rect 26110 -10600 26240 -9740
rect 26820 -10310 26920 -8650
rect 27040 -9860 27140 -8200
rect 28420 -8510 28520 -5760
rect 28620 -5960 28720 -4850
rect 29300 -5960 29440 -4110
rect 30000 -4260 30100 -2600
rect 30210 -2920 30330 -2910
rect 30210 -3040 30220 -2920
rect 30320 -3040 30330 -2920
rect 30210 -3050 30330 -3040
rect 29990 -4270 30110 -4260
rect 29990 -4390 30000 -4270
rect 30100 -4390 30110 -4270
rect 29990 -4400 30110 -4390
rect 28580 -5970 28760 -5960
rect 28580 -6150 28590 -5970
rect 28750 -6150 28760 -5970
rect 28580 -6160 28760 -6150
rect 29280 -5970 29460 -5960
rect 29280 -6150 29290 -5970
rect 29450 -6150 29460 -5970
rect 29280 -6160 29460 -6150
rect 28640 -8060 28740 -6160
rect 30000 -7160 30100 -4400
rect 30220 -4710 30320 -3050
rect 30900 -3170 31040 -2310
rect 30900 -3350 30910 -3170
rect 31030 -3350 31040 -3170
rect 30900 -3430 31040 -3350
rect 30900 -4110 30910 -3430
rect 31030 -4110 31040 -3430
rect 30210 -4720 30330 -4710
rect 30210 -4840 30220 -4720
rect 30320 -4840 30330 -4720
rect 30210 -4850 30330 -4840
rect 30220 -6760 30320 -4850
rect 30900 -5960 31040 -4110
rect 32500 -1630 32640 -1620
rect 32500 -2310 32510 -1630
rect 32630 -2310 32640 -1630
rect 32500 -2470 32640 -2310
rect 34100 -1630 34240 -1620
rect 34100 -2310 34110 -1630
rect 34230 -2310 34240 -1630
rect 32500 -2590 32510 -2470
rect 32630 -2590 32640 -2470
rect 32500 -3430 32640 -2590
rect 32500 -4110 32510 -3430
rect 32630 -4110 32640 -3430
rect 32500 -4120 32640 -4110
rect 33250 -4400 33390 -2460
rect 34100 -2470 34240 -2310
rect 34910 -2460 35040 1000
rect 35700 170 35840 180
rect 35700 -510 35710 170
rect 35830 -510 35840 170
rect 35700 -520 35840 -510
rect 35700 -1630 35840 -1620
rect 35700 -2310 35710 -1630
rect 35830 -2310 35840 -1630
rect 34100 -2590 34110 -2470
rect 34230 -2590 34240 -2470
rect 34100 -3430 34240 -2590
rect 34900 -2470 35050 -2460
rect 34900 -2590 34910 -2470
rect 35040 -2590 35050 -2470
rect 34900 -2600 35050 -2590
rect 35700 -2470 35840 -2310
rect 35700 -2590 35710 -2470
rect 35830 -2590 35840 -2470
rect 34100 -4110 34110 -3430
rect 34230 -4110 34240 -3430
rect 34100 -4120 34240 -4110
rect 35700 -3430 35840 -2590
rect 36400 -2900 36500 2810
rect 36390 -2910 36510 -2900
rect 36390 -3030 36400 -2910
rect 36500 -3030 36510 -2910
rect 36390 -3040 36510 -3030
rect 35700 -4110 35710 -3430
rect 35830 -4110 35840 -3430
rect 35700 -4120 35840 -4110
rect 36400 -4700 36500 -3040
rect 36390 -4710 36510 -4700
rect 36390 -4830 36400 -4710
rect 36500 -4830 36510 -4710
rect 36390 -4840 36510 -4830
rect 30880 -5970 31060 -5960
rect 30880 -6150 30890 -5970
rect 31050 -6150 31060 -5970
rect 30880 -6160 31060 -6150
rect 30180 -6770 30360 -6760
rect 30180 -6950 30190 -6770
rect 30350 -6950 30360 -6770
rect 30180 -6960 30360 -6950
rect 29960 -7170 30140 -7160
rect 29960 -7350 29970 -7170
rect 30130 -7350 30140 -7170
rect 29960 -7360 30140 -7350
rect 29960 -7570 30140 -7560
rect 29960 -7750 29970 -7570
rect 30130 -7750 30140 -7570
rect 29960 -7760 30140 -7750
rect 28620 -8070 28760 -8060
rect 28620 -8190 28630 -8070
rect 28750 -8190 28760 -8070
rect 28620 -8200 28760 -8190
rect 28400 -8520 28540 -8510
rect 28400 -8640 28410 -8520
rect 28530 -8640 28540 -8520
rect 28400 -8650 28540 -8640
rect 27710 -8800 27840 -8790
rect 27710 -9480 27720 -8800
rect 27830 -9480 27840 -8800
rect 27710 -9560 27840 -9480
rect 27700 -9570 27850 -9560
rect 27700 -9730 27710 -9570
rect 27840 -9730 27850 -9570
rect 27700 -9740 27850 -9730
rect 27020 -9870 27160 -9860
rect 27020 -9990 27030 -9870
rect 27150 -9990 27160 -9870
rect 27020 -10000 27160 -9990
rect 26800 -10320 26940 -10310
rect 26800 -10440 26810 -10320
rect 26930 -10440 26940 -10320
rect 26800 -10450 26940 -10440
rect 26110 -11280 26120 -10600
rect 26230 -11280 26240 -10600
rect 26110 -11360 26240 -11280
rect 26100 -11370 26250 -11360
rect 26100 -11530 26110 -11370
rect 26240 -11530 26250 -11370
rect 26100 -11540 26250 -11530
rect 25420 -11670 25560 -11660
rect 25420 -11790 25430 -11670
rect 25550 -11790 25560 -11670
rect 25420 -11800 25560 -11790
rect 25200 -12120 25340 -12110
rect 25200 -12240 25210 -12120
rect 25330 -12240 25340 -12120
rect 25200 -12250 25340 -12240
rect 24510 -13080 24520 -12400
rect 24630 -13080 24640 -12400
rect 24510 -13160 24640 -13080
rect 24500 -13170 24650 -13160
rect 24500 -13330 24510 -13170
rect 24640 -13330 24650 -13170
rect 24500 -13340 24650 -13330
rect 23820 -13470 23960 -13460
rect 23820 -13590 23830 -13470
rect 23950 -13590 23960 -13470
rect 23820 -13600 23960 -13590
rect 23600 -13920 23740 -13910
rect 23600 -14040 23610 -13920
rect 23730 -14040 23740 -13920
rect 23600 -14050 23740 -14040
rect 22910 -14880 22920 -14200
rect 23030 -14880 23040 -14200
rect 22910 -14960 23040 -14880
rect 22900 -14970 23050 -14960
rect 22900 -15130 22910 -14970
rect 23040 -15130 23050 -14970
rect 22900 -15140 23050 -15130
rect 22220 -15270 22360 -15260
rect 22220 -15390 22230 -15270
rect 22350 -15390 22360 -15270
rect 22220 -15400 22360 -15390
rect 22000 -15720 22140 -15710
rect 22000 -15840 22010 -15720
rect 22130 -15840 22140 -15720
rect 22000 -15850 22140 -15840
rect 21310 -16680 21320 -16000
rect 21430 -16680 21440 -16000
rect 21310 -16760 21440 -16680
rect 21300 -16770 21450 -16760
rect 21300 -16930 21310 -16770
rect 21440 -16930 21450 -16770
rect 21300 -16940 21450 -16930
rect 20620 -17070 20760 -17060
rect 20620 -17190 20630 -17070
rect 20750 -17190 20760 -17070
rect 20620 -17200 20760 -17190
rect 20400 -17520 20540 -17510
rect 20400 -17640 20410 -17520
rect 20530 -17640 20540 -17520
rect 20400 -17650 20540 -17640
rect 19710 -18480 19720 -17800
rect 19830 -18480 19840 -17800
rect 19710 -18560 19840 -18480
rect 19700 -18570 19850 -18560
rect 19700 -18730 19710 -18570
rect 19840 -18730 19850 -18570
rect 19700 -18740 19850 -18730
rect 19020 -18870 19160 -18860
rect 19020 -18990 19030 -18870
rect 19150 -18990 19160 -18870
rect 19020 -19000 19160 -18990
rect 18800 -19320 18940 -19310
rect 18800 -19440 18810 -19320
rect 18930 -19440 18940 -19320
rect 18800 -19450 18940 -19440
rect 18110 -20280 18120 -19600
rect 18230 -20280 18240 -19600
rect 18110 -20360 18240 -20280
rect 18100 -20370 18250 -20360
rect 18100 -20530 18110 -20370
rect 18240 -20530 18250 -20370
rect 18100 -20540 18250 -20530
rect 17420 -20670 17560 -20660
rect 17420 -20790 17430 -20670
rect 17550 -20790 17560 -20670
rect 17420 -20800 17560 -20790
rect 17200 -21120 17340 -21110
rect 17200 -21240 17210 -21120
rect 17330 -21240 17340 -21120
rect 17200 -21250 17340 -21240
rect 17220 -21370 17320 -21250
rect 17440 -21370 17540 -20800
rect 16510 -22080 16520 -21400
rect 16630 -22080 16640 -21400
rect 16510 -22160 16640 -22080
rect 18110 -21400 18240 -20540
rect 18820 -21110 18920 -19450
rect 19040 -20660 19140 -19000
rect 19710 -19600 19840 -18740
rect 20420 -19310 20520 -17650
rect 20640 -18860 20740 -17200
rect 21310 -17800 21440 -16940
rect 22020 -17510 22120 -15850
rect 22240 -17060 22340 -15400
rect 22910 -16000 23040 -15140
rect 23620 -15710 23720 -14050
rect 23840 -15260 23940 -13600
rect 24510 -14200 24640 -13340
rect 25220 -13910 25320 -12250
rect 25440 -13460 25540 -11800
rect 26110 -12400 26240 -11540
rect 26820 -12110 26920 -10450
rect 27040 -11660 27140 -10000
rect 27710 -10600 27840 -9740
rect 28420 -10310 28520 -8650
rect 28640 -9860 28740 -8200
rect 30020 -8510 30120 -7760
rect 30240 -8060 30340 -6960
rect 30220 -8070 30360 -8060
rect 30220 -8190 30230 -8070
rect 30350 -8190 30360 -8070
rect 30220 -8200 30360 -8190
rect 30000 -8520 30140 -8510
rect 30000 -8640 30010 -8520
rect 30130 -8640 30140 -8520
rect 30000 -8650 30140 -8640
rect 29310 -8800 29440 -8790
rect 29310 -9480 29320 -8800
rect 29430 -9480 29440 -8800
rect 29310 -9560 29440 -9480
rect 29300 -9570 29450 -9560
rect 29300 -9730 29310 -9570
rect 29440 -9730 29450 -9570
rect 29300 -9740 29450 -9730
rect 28620 -9870 28760 -9860
rect 28620 -9990 28630 -9870
rect 28750 -9990 28760 -9870
rect 28620 -10000 28760 -9990
rect 28400 -10320 28540 -10310
rect 28400 -10440 28410 -10320
rect 28530 -10440 28540 -10320
rect 28400 -10450 28540 -10440
rect 27710 -11280 27720 -10600
rect 27830 -11280 27840 -10600
rect 27710 -11360 27840 -11280
rect 27700 -11370 27850 -11360
rect 27700 -11530 27710 -11370
rect 27840 -11530 27850 -11370
rect 27700 -11540 27850 -11530
rect 27020 -11670 27160 -11660
rect 27020 -11790 27030 -11670
rect 27150 -11790 27160 -11670
rect 27020 -11800 27160 -11790
rect 26800 -12120 26940 -12110
rect 26800 -12240 26810 -12120
rect 26930 -12240 26940 -12120
rect 26800 -12250 26940 -12240
rect 26110 -13080 26120 -12400
rect 26230 -13080 26240 -12400
rect 26110 -13160 26240 -13080
rect 26100 -13170 26250 -13160
rect 26100 -13330 26110 -13170
rect 26240 -13330 26250 -13170
rect 26100 -13340 26250 -13330
rect 25420 -13470 25560 -13460
rect 25420 -13590 25430 -13470
rect 25550 -13590 25560 -13470
rect 25420 -13600 25560 -13590
rect 25200 -13920 25340 -13910
rect 25200 -14040 25210 -13920
rect 25330 -14040 25340 -13920
rect 25200 -14050 25340 -14040
rect 24510 -14880 24520 -14200
rect 24630 -14880 24640 -14200
rect 24510 -14960 24640 -14880
rect 24500 -14970 24650 -14960
rect 24500 -15130 24510 -14970
rect 24640 -15130 24650 -14970
rect 24500 -15140 24650 -15130
rect 23820 -15270 23960 -15260
rect 23820 -15390 23830 -15270
rect 23950 -15390 23960 -15270
rect 23820 -15400 23960 -15390
rect 23600 -15720 23740 -15710
rect 23600 -15840 23610 -15720
rect 23730 -15840 23740 -15720
rect 23600 -15850 23740 -15840
rect 22910 -16680 22920 -16000
rect 23030 -16680 23040 -16000
rect 22910 -16760 23040 -16680
rect 22900 -16770 23050 -16760
rect 22900 -16930 22910 -16770
rect 23040 -16930 23050 -16770
rect 22900 -16940 23050 -16930
rect 22220 -17070 22360 -17060
rect 22220 -17190 22230 -17070
rect 22350 -17190 22360 -17070
rect 22220 -17200 22360 -17190
rect 22000 -17520 22140 -17510
rect 22000 -17640 22010 -17520
rect 22130 -17640 22140 -17520
rect 22000 -17650 22140 -17640
rect 21310 -18480 21320 -17800
rect 21430 -18480 21440 -17800
rect 21310 -18560 21440 -18480
rect 21300 -18570 21450 -18560
rect 21300 -18730 21310 -18570
rect 21440 -18730 21450 -18570
rect 21300 -18740 21450 -18730
rect 20620 -18870 20760 -18860
rect 20620 -18990 20630 -18870
rect 20750 -18990 20760 -18870
rect 20620 -19000 20760 -18990
rect 20400 -19320 20540 -19310
rect 20400 -19440 20410 -19320
rect 20530 -19440 20540 -19320
rect 20400 -19450 20540 -19440
rect 19710 -20280 19720 -19600
rect 19830 -20280 19840 -19600
rect 19710 -20360 19840 -20280
rect 19700 -20370 19850 -20360
rect 19700 -20530 19710 -20370
rect 19840 -20530 19850 -20370
rect 19700 -20540 19850 -20530
rect 19020 -20670 19160 -20660
rect 19020 -20790 19030 -20670
rect 19150 -20790 19160 -20670
rect 19020 -20800 19160 -20790
rect 18800 -21120 18940 -21110
rect 18800 -21240 18810 -21120
rect 18930 -21240 18940 -21120
rect 18800 -21250 18940 -21240
rect 18820 -21370 18920 -21250
rect 19040 -21370 19140 -20800
rect 18110 -22080 18120 -21400
rect 18230 -22080 18240 -21400
rect 18110 -22160 18240 -22080
rect 19710 -21400 19840 -20540
rect 20420 -21110 20520 -19450
rect 20640 -20660 20740 -19000
rect 21310 -19600 21440 -18740
rect 22020 -19310 22120 -17650
rect 22240 -18860 22340 -17200
rect 22910 -17800 23040 -16940
rect 23620 -17510 23720 -15850
rect 23840 -17060 23940 -15400
rect 24510 -16000 24640 -15140
rect 25220 -15220 25320 -14050
rect 25440 -15220 25540 -13600
rect 26110 -14200 26240 -13340
rect 26820 -13910 26920 -12250
rect 27040 -13460 27140 -11800
rect 27710 -12400 27840 -11540
rect 28420 -12110 28520 -10450
rect 28640 -11660 28740 -10000
rect 29310 -10600 29440 -9740
rect 30020 -10310 30120 -8650
rect 30240 -9860 30340 -8200
rect 30910 -8650 31040 -8030
rect 30910 -8800 31040 -8790
rect 30910 -9480 30920 -8800
rect 31030 -9480 31040 -8800
rect 30910 -9560 31040 -9480
rect 30900 -9570 31050 -9560
rect 30900 -9730 30910 -9570
rect 31040 -9730 31050 -9570
rect 30900 -9740 31050 -9730
rect 30220 -9870 30360 -9860
rect 30220 -9990 30230 -9870
rect 30350 -9990 30360 -9870
rect 30220 -10000 30360 -9990
rect 30000 -10320 30140 -10310
rect 30000 -10440 30010 -10320
rect 30130 -10440 30140 -10320
rect 30000 -10450 30140 -10440
rect 29310 -11280 29320 -10600
rect 29430 -11280 29440 -10600
rect 29310 -11360 29440 -11280
rect 29300 -11370 29450 -11360
rect 29300 -11530 29310 -11370
rect 29440 -11530 29450 -11370
rect 29300 -11540 29450 -11530
rect 28620 -11670 28760 -11660
rect 28620 -11790 28630 -11670
rect 28750 -11790 28760 -11670
rect 28620 -11800 28760 -11790
rect 28400 -12120 28540 -12110
rect 28400 -12240 28410 -12120
rect 28530 -12240 28540 -12120
rect 28400 -12250 28540 -12240
rect 27710 -13080 27720 -12400
rect 27830 -13080 27840 -12400
rect 27710 -13160 27840 -13080
rect 27700 -13170 27850 -13160
rect 27700 -13330 27710 -13170
rect 27840 -13330 27850 -13170
rect 27700 -13340 27850 -13330
rect 27020 -13470 27160 -13460
rect 27020 -13590 27030 -13470
rect 27150 -13590 27160 -13470
rect 27020 -13600 27160 -13590
rect 26800 -13920 26940 -13910
rect 26800 -14040 26810 -13920
rect 26930 -14040 26940 -13920
rect 26800 -14050 26940 -14040
rect 26110 -14880 26120 -14200
rect 26230 -14880 26240 -14200
rect 26110 -14960 26240 -14880
rect 26100 -14970 26250 -14960
rect 26100 -15130 26110 -14970
rect 26240 -15130 26250 -14970
rect 26100 -15140 26250 -15130
rect 24510 -16680 24520 -16000
rect 24630 -16680 24640 -16000
rect 24510 -16760 24640 -16680
rect 26110 -16000 26240 -15140
rect 26820 -15710 26920 -14050
rect 27040 -15260 27140 -13600
rect 27710 -14200 27840 -13340
rect 28420 -13910 28520 -12250
rect 28640 -13460 28740 -11800
rect 29310 -12400 29440 -11540
rect 30020 -12110 30120 -10450
rect 30240 -11660 30340 -10000
rect 30910 -10600 31040 -9740
rect 30910 -11280 30920 -10600
rect 31030 -11280 31040 -10600
rect 30910 -11360 31040 -11280
rect 30900 -11370 31050 -11360
rect 30900 -11530 30910 -11370
rect 31040 -11530 31050 -11370
rect 30900 -11540 31050 -11530
rect 30220 -11670 30360 -11660
rect 30220 -11790 30230 -11670
rect 30350 -11790 30360 -11670
rect 30220 -11800 30360 -11790
rect 30000 -12120 30140 -12110
rect 30000 -12240 30010 -12120
rect 30130 -12240 30140 -12120
rect 30000 -12250 30140 -12240
rect 29310 -13080 29320 -12400
rect 29430 -13080 29440 -12400
rect 29310 -13160 29440 -13080
rect 29300 -13170 29450 -13160
rect 29300 -13330 29310 -13170
rect 29440 -13330 29450 -13170
rect 29300 -13340 29450 -13330
rect 28620 -13470 28760 -13460
rect 28620 -13590 28630 -13470
rect 28750 -13590 28760 -13470
rect 28620 -13600 28760 -13590
rect 28400 -13920 28540 -13910
rect 28400 -14040 28410 -13920
rect 28530 -14040 28540 -13920
rect 28400 -14050 28540 -14040
rect 27710 -14880 27720 -14200
rect 27830 -14880 27840 -14200
rect 27710 -14960 27840 -14880
rect 27700 -14970 27850 -14960
rect 27700 -15130 27710 -14970
rect 27840 -15130 27850 -14970
rect 27700 -15140 27850 -15130
rect 27020 -15270 27160 -15260
rect 27020 -15390 27030 -15270
rect 27150 -15390 27160 -15270
rect 27020 -15400 27160 -15390
rect 26800 -15720 26940 -15710
rect 26800 -15840 26810 -15720
rect 26930 -15840 26940 -15720
rect 26800 -15850 26940 -15840
rect 26110 -16680 26120 -16000
rect 26230 -16680 26240 -16000
rect 26110 -16760 26240 -16680
rect 24500 -16770 24650 -16760
rect 24500 -16930 24510 -16770
rect 24640 -16930 24650 -16770
rect 24500 -16940 24650 -16930
rect 26100 -16770 26250 -16760
rect 26100 -16930 26110 -16770
rect 26240 -16930 26250 -16770
rect 26100 -16940 26250 -16930
rect 23820 -17070 23960 -17060
rect 23820 -17190 23830 -17070
rect 23950 -17190 23960 -17070
rect 23820 -17200 23960 -17190
rect 23600 -17520 23740 -17510
rect 23600 -17640 23610 -17520
rect 23730 -17640 23740 -17520
rect 23600 -17650 23740 -17640
rect 22910 -18480 22920 -17800
rect 23030 -18480 23040 -17800
rect 22910 -18560 23040 -18480
rect 22900 -18570 23050 -18560
rect 22900 -18730 22910 -18570
rect 23040 -18730 23050 -18570
rect 22900 -18740 23050 -18730
rect 22220 -18870 22360 -18860
rect 22220 -18990 22230 -18870
rect 22350 -18990 22360 -18870
rect 22220 -19000 22360 -18990
rect 22000 -19320 22140 -19310
rect 22000 -19440 22010 -19320
rect 22130 -19440 22140 -19320
rect 22000 -19450 22140 -19440
rect 21310 -20280 21320 -19600
rect 21430 -20280 21440 -19600
rect 21310 -20360 21440 -20280
rect 21300 -20370 21450 -20360
rect 21300 -20530 21310 -20370
rect 21440 -20530 21450 -20370
rect 21300 -20540 21450 -20530
rect 20620 -20670 20760 -20660
rect 20620 -20790 20630 -20670
rect 20750 -20790 20760 -20670
rect 20620 -20800 20760 -20790
rect 20400 -21120 20540 -21110
rect 20400 -21240 20410 -21120
rect 20530 -21240 20540 -21120
rect 20400 -21250 20540 -21240
rect 20420 -21370 20520 -21250
rect 20640 -21370 20740 -20800
rect 19710 -22080 19720 -21400
rect 19830 -22080 19840 -21400
rect 19710 -22160 19840 -22080
rect 21310 -21400 21440 -20540
rect 22020 -21110 22120 -19450
rect 22240 -20660 22340 -19000
rect 22910 -19600 23040 -18740
rect 23620 -19310 23720 -17650
rect 23840 -18860 23940 -17200
rect 24510 -17800 24640 -16940
rect 24510 -18480 24520 -17800
rect 24630 -18480 24640 -17800
rect 24510 -18560 24640 -18480
rect 26110 -17800 26240 -16940
rect 26820 -17510 26920 -15850
rect 27040 -17060 27140 -15400
rect 27710 -16000 27840 -15140
rect 28420 -15710 28520 -14050
rect 28640 -15260 28740 -13600
rect 29310 -14200 29440 -13340
rect 30020 -13910 30120 -12250
rect 30240 -13460 30340 -11800
rect 30910 -12400 31040 -11540
rect 30910 -13080 30920 -12400
rect 31030 -13080 31040 -12400
rect 30910 -13160 31040 -13080
rect 30900 -13170 31050 -13160
rect 30900 -13330 30910 -13170
rect 31040 -13330 31050 -13170
rect 30900 -13340 31050 -13330
rect 30220 -13470 30360 -13460
rect 30220 -13590 30230 -13470
rect 30350 -13590 30360 -13470
rect 30220 -13600 30360 -13590
rect 30000 -13920 30140 -13910
rect 30000 -14040 30010 -13920
rect 30130 -14040 30140 -13920
rect 30000 -14050 30140 -14040
rect 29310 -14880 29320 -14200
rect 29430 -14880 29440 -14200
rect 29310 -14960 29440 -14880
rect 29300 -14970 29450 -14960
rect 29300 -15130 29310 -14970
rect 29440 -15130 29450 -14970
rect 29300 -15140 29450 -15130
rect 28620 -15270 28760 -15260
rect 28620 -15390 28630 -15270
rect 28750 -15390 28760 -15270
rect 28620 -15400 28760 -15390
rect 28400 -15720 28540 -15710
rect 28400 -15840 28410 -15720
rect 28530 -15840 28540 -15720
rect 28400 -15850 28540 -15840
rect 27710 -16680 27720 -16000
rect 27830 -16680 27840 -16000
rect 27710 -16760 27840 -16680
rect 27700 -16770 27850 -16760
rect 27700 -16930 27710 -16770
rect 27840 -16930 27850 -16770
rect 27700 -16940 27850 -16930
rect 27020 -17070 27160 -17060
rect 27020 -17190 27030 -17070
rect 27150 -17190 27160 -17070
rect 27020 -17200 27160 -17190
rect 26800 -17520 26940 -17510
rect 26800 -17640 26810 -17520
rect 26930 -17640 26940 -17520
rect 26800 -17650 26940 -17640
rect 26110 -18480 26120 -17800
rect 26230 -18480 26240 -17800
rect 26110 -18560 26240 -18480
rect 24500 -18570 24650 -18560
rect 24500 -18730 24510 -18570
rect 24640 -18730 24650 -18570
rect 24500 -18740 24650 -18730
rect 26100 -18570 26250 -18560
rect 26100 -18730 26110 -18570
rect 26240 -18730 26250 -18570
rect 26100 -18740 26250 -18730
rect 23820 -18870 23960 -18860
rect 23820 -18990 23830 -18870
rect 23950 -18990 23960 -18870
rect 23820 -19000 23960 -18990
rect 23600 -19320 23740 -19310
rect 23600 -19440 23610 -19320
rect 23730 -19440 23740 -19320
rect 23600 -19450 23740 -19440
rect 22910 -20280 22920 -19600
rect 23030 -20280 23040 -19600
rect 22910 -20360 23040 -20280
rect 22900 -20370 23050 -20360
rect 22900 -20530 22910 -20370
rect 23040 -20530 23050 -20370
rect 22900 -20540 23050 -20530
rect 22220 -20670 22360 -20660
rect 22220 -20790 22230 -20670
rect 22350 -20790 22360 -20670
rect 22220 -20800 22360 -20790
rect 22000 -21120 22140 -21110
rect 22000 -21240 22010 -21120
rect 22130 -21240 22140 -21120
rect 22000 -21250 22140 -21240
rect 22020 -21370 22120 -21250
rect 22240 -21370 22340 -20800
rect 21310 -22080 21320 -21400
rect 21430 -22080 21440 -21400
rect 21310 -22160 21440 -22080
rect 22910 -21400 23040 -20540
rect 23620 -21110 23720 -19450
rect 23840 -20660 23940 -19000
rect 24510 -19600 24640 -18740
rect 24510 -20280 24520 -19600
rect 24630 -20280 24640 -19600
rect 24510 -20360 24640 -20280
rect 26110 -19600 26240 -18740
rect 26820 -19310 26920 -17650
rect 27040 -18860 27140 -17200
rect 27710 -17800 27840 -16940
rect 28420 -17510 28520 -15850
rect 28640 -17060 28740 -15400
rect 29310 -16000 29440 -15140
rect 29310 -16680 29320 -16000
rect 29430 -16680 29440 -16000
rect 29310 -16760 29440 -16680
rect 29300 -16770 29450 -16760
rect 29300 -16930 29310 -16770
rect 29440 -16930 29450 -16770
rect 29300 -16940 29450 -16930
rect 28620 -17070 28760 -17060
rect 28620 -17190 28630 -17070
rect 28750 -17190 28760 -17070
rect 28620 -17200 28760 -17190
rect 28400 -17520 28540 -17510
rect 28400 -17640 28410 -17520
rect 28530 -17640 28540 -17520
rect 28400 -17650 28540 -17640
rect 27710 -18480 27720 -17800
rect 27830 -18480 27840 -17800
rect 27710 -18560 27840 -18480
rect 27700 -18570 27850 -18560
rect 27700 -18730 27710 -18570
rect 27840 -18730 27850 -18570
rect 27700 -18740 27850 -18730
rect 27020 -18870 27160 -18860
rect 27020 -18990 27030 -18870
rect 27150 -18990 27160 -18870
rect 27020 -19000 27160 -18990
rect 26800 -19320 26940 -19310
rect 26800 -19440 26810 -19320
rect 26930 -19440 26940 -19320
rect 26800 -19450 26940 -19440
rect 26110 -20280 26120 -19600
rect 26230 -20280 26240 -19600
rect 26110 -20360 26240 -20280
rect 24500 -20370 24650 -20360
rect 24500 -20530 24510 -20370
rect 24640 -20530 24650 -20370
rect 24500 -20540 24650 -20530
rect 26100 -20370 26250 -20360
rect 26100 -20530 26110 -20370
rect 26240 -20530 26250 -20370
rect 26100 -20540 26250 -20530
rect 23820 -20670 23960 -20660
rect 23820 -20790 23830 -20670
rect 23950 -20790 23960 -20670
rect 23820 -20800 23960 -20790
rect 23600 -21120 23740 -21110
rect 23600 -21240 23610 -21120
rect 23730 -21240 23740 -21120
rect 23600 -21250 23740 -21240
rect 23620 -21370 23720 -21250
rect 23840 -21370 23940 -20800
rect 22910 -22080 22920 -21400
rect 23030 -22080 23040 -21400
rect 22910 -22160 23040 -22080
rect 24510 -21400 24640 -20540
rect 24510 -22080 24520 -21400
rect 24630 -22080 24640 -21400
rect 24510 -22160 24640 -22080
rect 26110 -21400 26240 -20540
rect 26820 -21110 26920 -19450
rect 27040 -20660 27140 -19000
rect 27710 -19600 27840 -18740
rect 28420 -19310 28520 -17650
rect 28640 -18860 28740 -17200
rect 29310 -17800 29440 -16940
rect 29310 -18480 29320 -17800
rect 29430 -18480 29440 -17800
rect 29310 -18560 29440 -18480
rect 29300 -18570 29450 -18560
rect 29300 -18730 29310 -18570
rect 29440 -18730 29450 -18570
rect 29300 -18740 29450 -18730
rect 28620 -18870 28760 -18860
rect 28620 -18990 28630 -18870
rect 28750 -18990 28760 -18870
rect 28620 -19000 28760 -18990
rect 28400 -19320 28540 -19310
rect 28400 -19440 28410 -19320
rect 28530 -19440 28540 -19320
rect 28400 -19450 28540 -19440
rect 27710 -20280 27720 -19600
rect 27830 -20280 27840 -19600
rect 27710 -20360 27840 -20280
rect 27700 -20370 27850 -20360
rect 27700 -20530 27710 -20370
rect 27840 -20530 27850 -20370
rect 27700 -20540 27850 -20530
rect 27020 -20670 27160 -20660
rect 27020 -20790 27030 -20670
rect 27150 -20790 27160 -20670
rect 27020 -20800 27160 -20790
rect 26800 -21120 26940 -21110
rect 26800 -21240 26810 -21120
rect 26930 -21240 26940 -21120
rect 26800 -21250 26940 -21240
rect 26820 -21370 26920 -21250
rect 27040 -21370 27140 -20800
rect 26110 -22080 26120 -21400
rect 26230 -22080 26240 -21400
rect 26110 -22160 26240 -22080
rect 27710 -21400 27840 -20540
rect 28420 -21110 28520 -19450
rect 28640 -20660 28740 -19000
rect 29310 -19600 29440 -18740
rect 29310 -20280 29320 -19600
rect 29430 -20280 29440 -19600
rect 29310 -20360 29440 -20280
rect 29300 -20370 29450 -20360
rect 29300 -20530 29310 -20370
rect 29440 -20530 29450 -20370
rect 29300 -20540 29450 -20530
rect 28620 -20670 28760 -20660
rect 28620 -20790 28630 -20670
rect 28750 -20790 28760 -20670
rect 28620 -20800 28760 -20790
rect 28400 -21120 28540 -21110
rect 28400 -21240 28410 -21120
rect 28530 -21240 28540 -21120
rect 28400 -21250 28540 -21240
rect 28420 -21370 28520 -21250
rect 28640 -21370 28740 -20800
rect 27710 -22080 27720 -21400
rect 27830 -22080 27840 -21400
rect 27710 -22160 27840 -22080
rect 29310 -21400 29440 -20540
rect 30020 -21370 30120 -14050
rect 30240 -21370 30340 -13600
rect 30910 -14200 31040 -13340
rect 30910 -14880 30920 -14200
rect 31030 -14880 31040 -14200
rect 30910 -14960 31040 -14880
rect 30900 -14970 31050 -14960
rect 30900 -15130 30910 -14970
rect 31040 -15130 31050 -14970
rect 30900 -15140 31050 -15130
rect 30910 -16000 31040 -15140
rect 30910 -16680 30920 -16000
rect 31030 -16680 31040 -16000
rect 30910 -16760 31040 -16680
rect 30900 -16770 31050 -16760
rect 30900 -16930 30910 -16770
rect 31040 -16930 31050 -16770
rect 30900 -16940 31050 -16930
rect 30910 -17800 31040 -16940
rect 30910 -18480 30920 -17800
rect 31030 -18480 31040 -17800
rect 30910 -18560 31040 -18480
rect 30900 -18570 31050 -18560
rect 30900 -18730 30910 -18570
rect 31040 -18730 31050 -18570
rect 30900 -18740 31050 -18730
rect 30910 -19600 31040 -18740
rect 30910 -20280 30920 -19600
rect 31030 -20280 31040 -19600
rect 30910 -20360 31040 -20280
rect 30900 -20370 31050 -20360
rect 30900 -20530 30910 -20370
rect 31040 -20530 31050 -20370
rect 30900 -20540 31050 -20530
rect 29310 -22080 29320 -21400
rect 29430 -22080 29440 -21400
rect 29310 -22160 29440 -22080
rect 30910 -21400 31040 -20540
rect 30910 -22080 30920 -21400
rect 31030 -22080 31040 -21400
rect 30910 -22160 31040 -22080
rect 16500 -22170 16650 -22160
rect 10120 -22350 10130 -22190
rect 10230 -22350 10240 -22190
rect 10120 -22730 10240 -22350
rect 11030 -22360 11150 -22180
rect 16500 -22330 16510 -22170
rect 16640 -22330 16650 -22170
rect 16500 -22340 16650 -22330
rect 18100 -22170 18250 -22160
rect 18100 -22330 18110 -22170
rect 18240 -22330 18250 -22170
rect 18100 -22340 18250 -22330
rect 19700 -22170 19850 -22160
rect 19700 -22330 19710 -22170
rect 19840 -22330 19850 -22170
rect 19700 -22340 19850 -22330
rect 21300 -22170 21450 -22160
rect 21300 -22330 21310 -22170
rect 21440 -22330 21450 -22170
rect 21300 -22340 21450 -22330
rect 22900 -22170 23050 -22160
rect 22900 -22330 22910 -22170
rect 23040 -22330 23050 -22170
rect 22900 -22340 23050 -22330
rect 24500 -22170 24650 -22160
rect 24500 -22330 24510 -22170
rect 24640 -22330 24650 -22170
rect 24500 -22340 24650 -22330
rect 26100 -22170 26250 -22160
rect 26100 -22330 26110 -22170
rect 26240 -22330 26250 -22170
rect 26100 -22340 26250 -22330
rect 27700 -22170 27850 -22160
rect 27700 -22330 27710 -22170
rect 27840 -22330 27850 -22170
rect 27700 -22340 27850 -22330
rect 29300 -22170 29450 -22160
rect 29300 -22330 29310 -22170
rect 29440 -22330 29450 -22170
rect 29300 -22340 29450 -22330
rect 30900 -22170 31050 -22160
rect 30900 -22330 30910 -22170
rect 31040 -22330 31050 -22170
rect 30900 -22340 31050 -22330
rect 11040 -22730 11150 -22360
rect 11040 -22740 11160 -22730
rect 11040 -22850 11050 -22740
rect 11150 -22850 11160 -22740
rect 11040 -22860 11160 -22850
rect 27710 -22740 27840 -22340
rect 27710 -22850 27720 -22740
rect 27830 -22850 27840 -22740
rect 27710 -22860 27840 -22850
rect 29310 -22740 29440 -22340
rect 29310 -22850 29320 -22740
rect 29430 -22850 29440 -22740
rect 29310 -22860 29440 -22850
rect 30910 -22740 31040 -22340
rect 30910 -22850 30920 -22740
rect 31030 -22850 31040 -22740
rect 30910 -22860 31040 -22850
rect 2780 -23270 2960 -23260
rect 2780 -23450 2790 -23270
rect 2950 -23450 2960 -23270
rect 2780 -23460 2960 -23450
rect 4380 -23270 4560 -23260
rect 4380 -23450 4390 -23270
rect 4550 -23450 4560 -23270
rect 4380 -23460 4560 -23450
rect 5980 -23270 6160 -23260
rect 5980 -23450 5990 -23270
rect 6150 -23450 6160 -23270
rect 5980 -23460 6160 -23450
rect 7580 -23270 7760 -23260
rect 7580 -23450 7590 -23270
rect 7750 -23450 7760 -23270
rect 7580 -23460 7760 -23450
rect 9180 -23270 9360 -23260
rect 9180 -23450 9190 -23270
rect 9350 -23450 9360 -23270
rect 9180 -23460 9360 -23450
rect 2020 -25160 2080 -23820
rect 2240 -25160 2300 -23820
rect 2500 -25070 4020 -25060
rect 2500 -25130 2510 -25070
rect 4010 -25130 4020 -25070
rect 2500 -25140 4020 -25130
rect 4220 -25160 4280 -23820
rect 4440 -25160 4500 -23820
rect 4700 -25070 6220 -25060
rect 4700 -25130 4710 -25070
rect 6210 -25130 6220 -25070
rect 4700 -25140 6220 -25130
rect 6420 -25160 6480 -23820
rect 6640 -25160 6700 -23820
rect 6900 -25070 8420 -25060
rect 6900 -25130 6910 -25070
rect 8410 -25130 8420 -25070
rect 6900 -25140 8420 -25130
rect 8620 -25160 8680 -23820
rect 8840 -25160 8900 -23820
rect 9100 -25070 10620 -25060
rect 9100 -25130 9110 -25070
rect 10610 -25130 10620 -25070
rect 9100 -25140 10620 -25130
rect 10820 -25160 10880 -23820
rect 11040 -25160 11100 -23820
rect 11300 -25070 12820 -25060
rect 11300 -25130 11310 -25070
rect 12810 -25130 12820 -25070
rect 11300 -25140 12820 -25130
rect 13020 -25160 13080 -23820
rect 13240 -25160 13300 -23820
rect 13500 -25070 15020 -25060
rect 13500 -25130 13510 -25070
rect 15010 -25130 15020 -25070
rect 13500 -25140 15020 -25130
rect 15220 -25160 15280 -23820
rect 15440 -25160 15500 -23820
rect 15700 -25070 17220 -25060
rect 15700 -25130 15710 -25070
rect 17210 -25130 17220 -25070
rect 15700 -25140 17220 -25130
rect 17420 -25160 17480 -23820
rect 17640 -25160 17700 -23820
rect 17900 -25070 19420 -25060
rect 17900 -25130 17910 -25070
rect 19410 -25130 19420 -25070
rect 17900 -25140 19420 -25130
rect 19620 -25160 19680 -23820
rect 19840 -25160 19900 -23820
rect 2010 -25330 2090 -25160
rect 2230 -25260 2310 -25160
rect 2230 -25320 2240 -25260
rect 2300 -25320 2310 -25260
rect 2230 -25330 2310 -25320
rect -70 -25390 -10 -25380
rect -70 -25460 -10 -25450
rect 2020 -25960 2080 -25330
rect 2130 -25390 2190 -25380
rect 2130 -25460 2190 -25450
rect 2240 -25960 2300 -25330
rect 4210 -25350 4290 -25160
rect 4430 -25170 4510 -25160
rect 4430 -25230 4440 -25170
rect 4500 -25230 4510 -25170
rect 4430 -25280 4510 -25230
rect 4430 -25340 4440 -25280
rect 4500 -25340 4510 -25280
rect 4430 -25350 4510 -25340
rect 6410 -25280 6490 -25160
rect 6410 -25340 6420 -25280
rect 6480 -25340 6490 -25280
rect 6410 -25350 6490 -25340
rect 6630 -25170 6710 -25160
rect 6630 -25230 6640 -25170
rect 6700 -25230 6710 -25170
rect 6630 -25350 6710 -25230
rect 8610 -25170 8690 -25160
rect 8610 -25230 8620 -25170
rect 8680 -25230 8690 -25170
rect 8610 -25280 8690 -25230
rect 8610 -25340 8620 -25280
rect 8680 -25340 8690 -25280
rect 8610 -25350 8690 -25340
rect 8830 -25350 8910 -25160
rect 10810 -25170 10890 -25160
rect 10810 -25230 10820 -25170
rect 10880 -25230 10890 -25170
rect 10810 -25280 10890 -25230
rect 10810 -25340 10820 -25280
rect 10880 -25340 10890 -25280
rect 10810 -25350 10890 -25340
rect 11030 -25350 11110 -25160
rect 13010 -25170 13090 -25160
rect 13010 -25230 13020 -25170
rect 13080 -25230 13090 -25170
rect 13010 -25280 13090 -25230
rect 13010 -25340 13020 -25280
rect 13080 -25340 13090 -25280
rect 13010 -25350 13090 -25340
rect 13230 -25350 13310 -25160
rect 15210 -25170 15290 -25160
rect 15210 -25230 15220 -25170
rect 15280 -25230 15290 -25170
rect 15210 -25350 15290 -25230
rect 15430 -25280 15510 -25160
rect 15430 -25340 15440 -25280
rect 15500 -25340 15510 -25280
rect 15430 -25350 15510 -25340
rect 17410 -25350 17490 -25160
rect 17630 -25170 17710 -25160
rect 17630 -25230 17640 -25170
rect 17700 -25230 17710 -25170
rect 17630 -25280 17710 -25230
rect 17630 -25340 17640 -25280
rect 17700 -25340 17710 -25280
rect 17630 -25350 17710 -25340
rect 19610 -25350 19690 -25160
rect 19830 -25170 19910 -25160
rect 19830 -25230 19840 -25170
rect 19900 -25230 19910 -25170
rect 19830 -25350 19910 -25230
rect 2500 -25630 2700 -25550
rect 3160 -25630 3360 -25550
rect 3820 -25630 4020 -25550
rect 2500 -25700 2700 -25690
rect 2500 -25760 2510 -25700
rect 2690 -25760 2700 -25700
rect 2500 -25770 2700 -25760
rect 3160 -25700 3360 -25690
rect 3160 -25760 3170 -25700
rect 3350 -25760 3360 -25700
rect 3160 -25770 3360 -25760
rect 3820 -25700 4020 -25690
rect 3820 -25760 3830 -25700
rect 4010 -25760 4020 -25700
rect 3820 -25770 4020 -25760
rect 2500 -25870 4020 -25860
rect 2500 -25930 2510 -25870
rect 4010 -25930 4020 -25870
rect 2500 -25940 4020 -25930
rect 4220 -25960 4280 -25350
rect 4330 -25390 4390 -25380
rect 4330 -25460 4390 -25450
rect 4440 -25960 4500 -25350
rect 4700 -25630 4900 -25550
rect 5360 -25630 5560 -25550
rect 6020 -25630 6220 -25550
rect 4700 -25700 4900 -25690
rect 4700 -25760 4710 -25700
rect 4890 -25760 4900 -25700
rect 4700 -25770 4900 -25760
rect 5360 -25700 5560 -25690
rect 5360 -25760 5370 -25700
rect 5550 -25760 5560 -25700
rect 5360 -25770 5560 -25760
rect 6020 -25700 6220 -25690
rect 6020 -25760 6030 -25700
rect 6210 -25760 6220 -25700
rect 6020 -25770 6220 -25760
rect 4700 -25870 6220 -25860
rect 4700 -25930 4710 -25870
rect 6210 -25930 6220 -25870
rect 4700 -25940 6220 -25930
rect 6420 -25960 6480 -25350
rect 6530 -25390 6590 -25380
rect 6530 -25460 6590 -25450
rect 6640 -25960 6700 -25350
rect 6900 -25560 7100 -25550
rect 6900 -25620 6910 -25560
rect 7090 -25620 7100 -25560
rect 6900 -25630 7100 -25620
rect 7560 -25560 7760 -25550
rect 7560 -25620 7570 -25560
rect 7750 -25620 7760 -25560
rect 7560 -25630 7760 -25620
rect 8220 -25560 8420 -25550
rect 8220 -25620 8230 -25560
rect 8410 -25620 8420 -25560
rect 8220 -25630 8420 -25620
rect 6900 -25770 7100 -25690
rect 7560 -25770 7760 -25690
rect 8220 -25770 8420 -25690
rect 6900 -25870 8420 -25860
rect 6900 -25930 6910 -25870
rect 8410 -25930 8420 -25870
rect 6900 -25940 8420 -25930
rect 8620 -25960 8680 -25350
rect 8730 -25390 8790 -25380
rect 8730 -25460 8790 -25450
rect 8840 -25960 8900 -25350
rect 9100 -25560 9300 -25550
rect 9100 -25620 9110 -25560
rect 9290 -25620 9300 -25560
rect 9100 -25630 9300 -25620
rect 9760 -25560 9960 -25550
rect 9760 -25620 9770 -25560
rect 9950 -25620 9960 -25560
rect 9760 -25630 9960 -25620
rect 10420 -25560 10620 -25550
rect 10420 -25620 10430 -25560
rect 10610 -25620 10620 -25560
rect 10420 -25630 10620 -25620
rect 9100 -25770 9300 -25690
rect 9760 -25770 9960 -25690
rect 10420 -25770 10620 -25690
rect 9100 -25870 10620 -25860
rect 9100 -25930 9110 -25870
rect 10610 -25930 10620 -25870
rect 9100 -25940 10620 -25930
rect 10820 -25960 10880 -25350
rect 10930 -25390 10990 -25380
rect 10930 -25460 10990 -25450
rect 11040 -25960 11100 -25350
rect 11300 -25560 11500 -25550
rect 11300 -25620 11310 -25560
rect 11490 -25620 11500 -25560
rect 11300 -25630 11500 -25620
rect 11960 -25560 12160 -25550
rect 11960 -25620 11970 -25560
rect 12150 -25620 12160 -25560
rect 11960 -25630 12160 -25620
rect 12620 -25560 12820 -25550
rect 12620 -25620 12630 -25560
rect 12810 -25620 12820 -25560
rect 12620 -25630 12820 -25620
rect 11300 -25770 11500 -25690
rect 11960 -25770 12160 -25690
rect 12620 -25770 12820 -25690
rect 11300 -25870 12820 -25860
rect 11300 -25930 11310 -25870
rect 12810 -25930 12820 -25870
rect 11300 -25940 12820 -25930
rect 13020 -25960 13080 -25350
rect 13130 -25390 13190 -25380
rect 13130 -25460 13190 -25450
rect 13240 -25960 13300 -25350
rect 13500 -25560 13700 -25550
rect 13500 -25620 13510 -25560
rect 13690 -25620 13700 -25560
rect 13500 -25630 13700 -25620
rect 14160 -25560 14360 -25550
rect 14160 -25620 14170 -25560
rect 14350 -25620 14360 -25560
rect 14160 -25630 14360 -25620
rect 14820 -25560 15020 -25550
rect 14820 -25620 14830 -25560
rect 15010 -25620 15020 -25560
rect 14820 -25630 15020 -25620
rect 13500 -25770 13700 -25690
rect 14160 -25770 14360 -25690
rect 14820 -25770 15020 -25690
rect 13500 -25870 15020 -25860
rect 13500 -25930 13510 -25870
rect 15010 -25930 15020 -25870
rect 13500 -25940 15020 -25930
rect 15220 -25960 15280 -25350
rect 15330 -25390 15390 -25380
rect 15330 -25460 15390 -25450
rect 15440 -25960 15500 -25350
rect 15700 -25630 15900 -25550
rect 16360 -25630 16560 -25550
rect 17020 -25630 17220 -25550
rect 15700 -25700 15900 -25690
rect 15700 -25760 15710 -25700
rect 15890 -25760 15900 -25700
rect 15700 -25770 15900 -25760
rect 16360 -25700 16560 -25690
rect 16360 -25760 16370 -25700
rect 16550 -25760 16560 -25700
rect 16360 -25770 16560 -25760
rect 17020 -25700 17220 -25690
rect 17020 -25760 17030 -25700
rect 17210 -25760 17220 -25700
rect 17020 -25770 17220 -25760
rect 15700 -25870 17220 -25860
rect 15700 -25930 15710 -25870
rect 17210 -25930 17220 -25870
rect 15700 -25940 17220 -25930
rect 17420 -25960 17480 -25350
rect 17530 -25390 17590 -25380
rect 17530 -25460 17590 -25450
rect 17640 -25960 17700 -25350
rect 17900 -25630 18100 -25550
rect 18560 -25630 18760 -25550
rect 19220 -25630 19420 -25550
rect 17900 -25700 18100 -25690
rect 17900 -25760 17910 -25700
rect 18090 -25760 18100 -25700
rect 17900 -25770 18100 -25760
rect 18560 -25700 18760 -25690
rect 18560 -25760 18570 -25700
rect 18750 -25760 18760 -25700
rect 18560 -25770 18760 -25760
rect 19220 -25700 19420 -25690
rect 19220 -25760 19230 -25700
rect 19410 -25760 19420 -25700
rect 19220 -25770 19420 -25760
rect 17900 -25870 19420 -25860
rect 17900 -25930 17910 -25870
rect 19410 -25930 19420 -25870
rect 17900 -25940 19420 -25930
rect 19620 -25960 19680 -25350
rect 19730 -25390 19790 -25380
rect 19730 -25460 19790 -25450
rect 19840 -25960 19900 -25350
rect 21930 -25390 21990 -25380
rect 21930 -25460 21990 -25450
rect 2010 -26060 2090 -25960
rect 2010 -26120 2020 -26060
rect 2080 -26120 2090 -26060
rect 2010 -26130 2090 -26120
rect 2230 -26130 2310 -25960
rect 4210 -25970 4290 -25960
rect 4210 -26030 4220 -25970
rect 4280 -26030 4290 -25970
rect 4210 -26080 4290 -26030
rect -70 -26190 -10 -26180
rect -70 -26260 -10 -26250
rect 420 -26630 620 -26620
rect 420 -26710 430 -26630
rect 610 -26710 620 -26630
rect 420 -26720 620 -26710
rect 2020 -26760 2080 -26130
rect 2130 -26190 2190 -26180
rect 2130 -26260 2190 -26250
rect 2240 -26760 2300 -26130
rect 4210 -26140 4220 -26080
rect 4280 -26140 4290 -26080
rect 4210 -26150 4290 -26140
rect 4430 -26150 4510 -25960
rect 6410 -25970 6490 -25960
rect 6410 -26030 6420 -25970
rect 6480 -26030 6490 -25970
rect 6410 -26150 6490 -26030
rect 6630 -26080 6710 -25960
rect 6630 -26140 6640 -26080
rect 6700 -26140 6710 -26080
rect 6630 -26150 6710 -26140
rect 8610 -26150 8690 -25960
rect 8830 -25970 8910 -25960
rect 8830 -26030 8840 -25970
rect 8900 -26030 8910 -25970
rect 8830 -26080 8910 -26030
rect 8830 -26140 8840 -26080
rect 8900 -26140 8910 -26080
rect 8830 -26150 8910 -26140
rect 10810 -26150 10890 -25960
rect 11030 -25970 11110 -25960
rect 11030 -26030 11040 -25970
rect 11100 -26030 11110 -25970
rect 11030 -26080 11110 -26030
rect 11030 -26140 11040 -26080
rect 11100 -26140 11110 -26080
rect 11030 -26150 11110 -26140
rect 13010 -26150 13090 -25960
rect 13230 -25970 13310 -25960
rect 13230 -26030 13240 -25970
rect 13300 -26030 13310 -25970
rect 13230 -26080 13310 -26030
rect 13230 -26140 13240 -26080
rect 13300 -26140 13310 -26080
rect 13230 -26150 13310 -26140
rect 15210 -26080 15290 -25960
rect 15210 -26140 15220 -26080
rect 15280 -26140 15290 -26080
rect 15210 -26150 15290 -26140
rect 15430 -25970 15510 -25960
rect 15430 -26030 15440 -25970
rect 15500 -26030 15510 -25970
rect 15430 -26150 15510 -26030
rect 17410 -25970 17490 -25960
rect 17410 -26030 17420 -25970
rect 17480 -26030 17490 -25970
rect 17410 -26080 17490 -26030
rect 17410 -26140 17420 -26080
rect 17480 -26140 17490 -26080
rect 17410 -26150 17490 -26140
rect 17630 -26150 17710 -25960
rect 19610 -25970 19690 -25960
rect 19610 -26030 19620 -25970
rect 19680 -26030 19690 -25970
rect 19610 -26150 19690 -26030
rect 19830 -26150 19910 -25960
rect 2500 -26360 2700 -26350
rect 2500 -26420 2510 -26360
rect 2690 -26420 2700 -26360
rect 2500 -26430 2700 -26420
rect 3160 -26360 3360 -26350
rect 3160 -26420 3170 -26360
rect 3350 -26420 3360 -26360
rect 3160 -26430 3360 -26420
rect 3820 -26360 4020 -26350
rect 3820 -26420 3830 -26360
rect 4010 -26420 4020 -26360
rect 3820 -26430 4020 -26420
rect 2500 -26570 2700 -26490
rect 3160 -26570 3360 -26490
rect 3820 -26570 4020 -26490
rect 4220 -26760 4280 -26150
rect 4330 -26190 4390 -26180
rect 4330 -26260 4390 -26250
rect 4440 -26760 4500 -26150
rect 4700 -26360 4900 -26350
rect 4700 -26420 4710 -26360
rect 4890 -26420 4900 -26360
rect 4700 -26430 4900 -26420
rect 5360 -26360 5560 -26350
rect 5360 -26420 5370 -26360
rect 5550 -26420 5560 -26360
rect 5360 -26430 5560 -26420
rect 6020 -26360 6220 -26350
rect 6020 -26420 6030 -26360
rect 6210 -26420 6220 -26360
rect 6020 -26430 6220 -26420
rect 4700 -26570 4900 -26490
rect 5360 -26570 5560 -26490
rect 6020 -26570 6220 -26490
rect 4700 -26670 6220 -26660
rect 4700 -26730 4710 -26670
rect 6210 -26730 6220 -26670
rect 4700 -26740 6220 -26730
rect 6420 -26760 6480 -26150
rect 6530 -26190 6590 -26180
rect 6530 -26260 6590 -26250
rect 6640 -26760 6700 -26150
rect 6900 -26430 7100 -26350
rect 7560 -26430 7760 -26350
rect 8220 -26430 8420 -26350
rect 6900 -26500 7100 -26490
rect 6900 -26560 6910 -26500
rect 7090 -26560 7100 -26500
rect 6900 -26570 7100 -26560
rect 7560 -26500 7760 -26490
rect 7560 -26560 7570 -26500
rect 7750 -26560 7760 -26500
rect 7560 -26570 7760 -26560
rect 8220 -26500 8420 -26490
rect 8220 -26560 8230 -26500
rect 8410 -26560 8420 -26500
rect 8220 -26570 8420 -26560
rect 6900 -26670 8420 -26660
rect 6900 -26730 6910 -26670
rect 8410 -26730 8420 -26670
rect 6900 -26740 8420 -26730
rect 8620 -26760 8680 -26150
rect 8730 -26190 8790 -26180
rect 8730 -26260 8790 -26250
rect 8840 -26760 8900 -26150
rect 9100 -26430 9300 -26350
rect 9760 -26430 9960 -26350
rect 10420 -26430 10620 -26350
rect 9100 -26500 9300 -26490
rect 9100 -26560 9110 -26500
rect 9290 -26560 9300 -26500
rect 9100 -26570 9300 -26560
rect 9760 -26500 9960 -26490
rect 9760 -26560 9770 -26500
rect 9950 -26560 9960 -26500
rect 9760 -26570 9960 -26560
rect 10420 -26500 10620 -26490
rect 10420 -26560 10430 -26500
rect 10610 -26560 10620 -26500
rect 10420 -26570 10620 -26560
rect 9100 -26670 10620 -26660
rect 9100 -26730 9110 -26670
rect 10610 -26730 10620 -26670
rect 9100 -26740 10620 -26730
rect 10820 -26760 10880 -26150
rect 10930 -26190 10990 -26180
rect 10930 -26260 10990 -26250
rect 11040 -26760 11100 -26150
rect 11300 -26430 11500 -26350
rect 11960 -26430 12160 -26350
rect 12620 -26430 12820 -26350
rect 11300 -26500 11500 -26490
rect 11300 -26560 11310 -26500
rect 11490 -26560 11500 -26500
rect 11300 -26570 11500 -26560
rect 11960 -26500 12160 -26490
rect 11960 -26560 11970 -26500
rect 12150 -26560 12160 -26500
rect 11960 -26570 12160 -26560
rect 12620 -26500 12820 -26490
rect 12620 -26560 12630 -26500
rect 12810 -26560 12820 -26500
rect 12620 -26570 12820 -26560
rect 11300 -26670 12820 -26660
rect 11300 -26730 11310 -26670
rect 12810 -26730 12820 -26670
rect 11300 -26740 12820 -26730
rect 13020 -26760 13080 -26150
rect 13130 -26190 13190 -26180
rect 13130 -26260 13190 -26250
rect 13240 -26760 13300 -26150
rect 13500 -26430 13700 -26350
rect 14160 -26430 14360 -26350
rect 14820 -26430 15020 -26350
rect 13500 -26500 13700 -26490
rect 13500 -26560 13510 -26500
rect 13690 -26560 13700 -26500
rect 13500 -26570 13700 -26560
rect 14160 -26500 14360 -26490
rect 14160 -26560 14170 -26500
rect 14350 -26560 14360 -26500
rect 14160 -26570 14360 -26560
rect 14820 -26500 15020 -26490
rect 14820 -26560 14830 -26500
rect 15010 -26560 15020 -26500
rect 14820 -26570 15020 -26560
rect 13500 -26670 15020 -26660
rect 13500 -26730 13510 -26670
rect 15010 -26730 15020 -26670
rect 13500 -26740 15020 -26730
rect 15220 -26760 15280 -26150
rect 15330 -26190 15390 -26180
rect 15330 -26260 15390 -26250
rect 15440 -26760 15500 -26150
rect 15700 -26360 15900 -26350
rect 15700 -26420 15710 -26360
rect 15890 -26420 15900 -26360
rect 15700 -26430 15900 -26420
rect 16360 -26360 16560 -26350
rect 16360 -26420 16370 -26360
rect 16550 -26420 16560 -26360
rect 16360 -26430 16560 -26420
rect 17020 -26360 17220 -26350
rect 17020 -26420 17030 -26360
rect 17210 -26420 17220 -26360
rect 17020 -26430 17220 -26420
rect 15700 -26570 15900 -26490
rect 16360 -26570 16560 -26490
rect 17020 -26570 17220 -26490
rect 15700 -26670 17220 -26660
rect 15700 -26730 15710 -26670
rect 17210 -26730 17220 -26670
rect 15700 -26740 17220 -26730
rect 17420 -26760 17480 -26150
rect 17530 -26190 17590 -26180
rect 17530 -26260 17590 -26250
rect 17640 -26760 17700 -26150
rect 17900 -26360 18100 -26350
rect 17900 -26420 17910 -26360
rect 18090 -26420 18100 -26360
rect 17900 -26430 18100 -26420
rect 18560 -26360 18760 -26350
rect 18560 -26420 18570 -26360
rect 18750 -26420 18760 -26360
rect 18560 -26430 18760 -26420
rect 19220 -26360 19420 -26350
rect 19220 -26420 19230 -26360
rect 19410 -26420 19420 -26360
rect 19220 -26430 19420 -26420
rect 17900 -26570 18100 -26490
rect 18560 -26570 18760 -26490
rect 19220 -26570 19420 -26490
rect 19620 -26760 19680 -26150
rect 19730 -26190 19790 -26180
rect 19730 -26260 19790 -26250
rect 19840 -26760 19900 -26150
rect 21930 -26190 21990 -26180
rect 21930 -26260 21990 -26250
rect 21300 -26630 21500 -26620
rect 21300 -26710 21310 -26630
rect 21490 -26710 21500 -26630
rect 21300 -26720 21500 -26710
rect 2010 -26930 2090 -26760
rect 2230 -26930 2310 -26760
rect -70 -26990 -10 -26980
rect -70 -27060 -10 -27050
rect 420 -27430 620 -27420
rect 420 -27510 430 -27430
rect 610 -27510 620 -27430
rect 420 -27520 620 -27510
rect 2020 -27560 2080 -26930
rect 2130 -26990 2190 -26980
rect 2130 -27060 2190 -27050
rect 2240 -27560 2300 -26930
rect 4210 -26950 4290 -26760
rect 4430 -26880 4510 -26760
rect 4430 -26940 4440 -26880
rect 4500 -26940 4510 -26880
rect 4430 -26950 4510 -26940
rect 6410 -26880 6490 -26760
rect 6410 -26940 6420 -26880
rect 6480 -26940 6490 -26880
rect 6410 -26950 6490 -26940
rect 6630 -26770 6710 -26760
rect 6630 -26830 6640 -26770
rect 6700 -26830 6710 -26770
rect 6630 -26950 6710 -26830
rect 8610 -26770 8690 -26760
rect 8610 -26830 8620 -26770
rect 8680 -26830 8690 -26770
rect 8610 -26880 8690 -26830
rect 8610 -26940 8620 -26880
rect 8680 -26940 8690 -26880
rect 8610 -26950 8690 -26940
rect 8830 -26950 8910 -26760
rect 10810 -26770 10890 -26760
rect 10810 -26830 10820 -26770
rect 10880 -26830 10890 -26770
rect 10810 -26880 10890 -26830
rect 10810 -26940 10820 -26880
rect 10880 -26940 10890 -26880
rect 10810 -26950 10890 -26940
rect 11030 -26950 11110 -26760
rect 13010 -26770 13090 -26760
rect 13010 -26830 13020 -26770
rect 13080 -26830 13090 -26770
rect 13010 -26880 13090 -26830
rect 13010 -26940 13020 -26880
rect 13080 -26940 13090 -26880
rect 13010 -26950 13090 -26940
rect 13230 -26950 13310 -26760
rect 15210 -26770 15290 -26760
rect 15210 -26830 15220 -26770
rect 15280 -26830 15290 -26770
rect 15210 -26950 15290 -26830
rect 15430 -26880 15510 -26760
rect 15430 -26940 15440 -26880
rect 15500 -26940 15510 -26880
rect 15430 -26950 15510 -26940
rect 17410 -26950 17490 -26760
rect 17630 -26770 17710 -26760
rect 17630 -26830 17640 -26770
rect 17700 -26830 17710 -26770
rect 17630 -26950 17710 -26830
rect 19610 -26950 19690 -26760
rect 19830 -26950 19910 -26760
rect 2500 -27230 2700 -27150
rect 3160 -27230 3360 -27150
rect 3820 -27230 4020 -27150
rect 2500 -27300 2700 -27290
rect 2500 -27360 2510 -27300
rect 2690 -27360 2700 -27300
rect 2500 -27370 2700 -27360
rect 3160 -27300 3360 -27290
rect 3160 -27360 3170 -27300
rect 3350 -27360 3360 -27300
rect 3160 -27370 3360 -27360
rect 3820 -27300 4020 -27290
rect 3820 -27360 3830 -27300
rect 4010 -27360 4020 -27300
rect 3820 -27370 4020 -27360
rect 4220 -27560 4280 -26950
rect 4330 -26990 4390 -26980
rect 4330 -27060 4390 -27050
rect 4440 -27560 4500 -26950
rect 4700 -27230 4900 -27150
rect 5360 -27230 5560 -27150
rect 6020 -27230 6220 -27150
rect 4700 -27300 4900 -27290
rect 4700 -27360 4710 -27300
rect 4890 -27360 4900 -27300
rect 4700 -27370 4900 -27360
rect 5360 -27300 5560 -27290
rect 5360 -27360 5370 -27300
rect 5550 -27360 5560 -27300
rect 5360 -27370 5560 -27360
rect 6020 -27300 6220 -27290
rect 6020 -27360 6030 -27300
rect 6210 -27360 6220 -27300
rect 6020 -27370 6220 -27360
rect 4700 -27470 6220 -27460
rect 4700 -27530 4710 -27470
rect 6210 -27530 6220 -27470
rect 4700 -27540 6220 -27530
rect 6420 -27560 6480 -26950
rect 6530 -26990 6590 -26980
rect 6530 -27060 6590 -27050
rect 6640 -27560 6700 -26950
rect 6900 -27160 7100 -27150
rect 6900 -27220 6910 -27160
rect 7090 -27220 7100 -27160
rect 6900 -27230 7100 -27220
rect 7560 -27160 7760 -27150
rect 7560 -27220 7570 -27160
rect 7750 -27220 7760 -27160
rect 7560 -27230 7760 -27220
rect 8220 -27160 8420 -27150
rect 8220 -27220 8230 -27160
rect 8410 -27220 8420 -27160
rect 8220 -27230 8420 -27220
rect 6900 -27370 7100 -27290
rect 7560 -27370 7760 -27290
rect 8220 -27370 8420 -27290
rect 6900 -27470 8420 -27460
rect 6900 -27530 6910 -27470
rect 8410 -27530 8420 -27470
rect 6900 -27540 8420 -27530
rect 8620 -27560 8680 -26950
rect 8730 -26990 8790 -26980
rect 8730 -27060 8790 -27050
rect 8840 -27560 8900 -26950
rect 9100 -27160 9300 -27150
rect 9100 -27220 9110 -27160
rect 9290 -27220 9300 -27160
rect 9100 -27230 9300 -27220
rect 9760 -27160 9960 -27150
rect 9760 -27220 9770 -27160
rect 9950 -27220 9960 -27160
rect 9760 -27230 9960 -27220
rect 10420 -27160 10620 -27150
rect 10420 -27220 10430 -27160
rect 10610 -27220 10620 -27160
rect 10420 -27230 10620 -27220
rect 9100 -27370 9300 -27290
rect 9760 -27370 9960 -27290
rect 10420 -27370 10620 -27290
rect 9100 -27470 10620 -27460
rect 9100 -27530 9110 -27470
rect 10610 -27530 10620 -27470
rect 9100 -27540 10620 -27530
rect 10820 -27560 10880 -26950
rect 10930 -26990 10990 -26980
rect 10930 -27060 10990 -27050
rect 11040 -27560 11100 -26950
rect 11300 -27160 11500 -27150
rect 11300 -27220 11310 -27160
rect 11490 -27220 11500 -27160
rect 11300 -27230 11500 -27220
rect 11960 -27160 12160 -27150
rect 11960 -27220 11970 -27160
rect 12150 -27220 12160 -27160
rect 11960 -27230 12160 -27220
rect 12620 -27160 12820 -27150
rect 12620 -27220 12630 -27160
rect 12810 -27220 12820 -27160
rect 12620 -27230 12820 -27220
rect 11300 -27370 11500 -27290
rect 11960 -27370 12160 -27290
rect 12620 -27370 12820 -27290
rect 11300 -27470 12820 -27460
rect 11300 -27530 11310 -27470
rect 12810 -27530 12820 -27470
rect 11300 -27540 12820 -27530
rect 13020 -27560 13080 -26950
rect 13130 -26990 13190 -26980
rect 13130 -27060 13190 -27050
rect 13240 -27560 13300 -26950
rect 13500 -27160 13700 -27150
rect 13500 -27220 13510 -27160
rect 13690 -27220 13700 -27160
rect 13500 -27230 13700 -27220
rect 14160 -27160 14360 -27150
rect 14160 -27220 14170 -27160
rect 14350 -27220 14360 -27160
rect 14160 -27230 14360 -27220
rect 14820 -27160 15020 -27150
rect 14820 -27220 14830 -27160
rect 15010 -27220 15020 -27160
rect 14820 -27230 15020 -27220
rect 13500 -27370 13700 -27290
rect 14160 -27370 14360 -27290
rect 14820 -27370 15020 -27290
rect 13500 -27470 15020 -27460
rect 13500 -27530 13510 -27470
rect 15010 -27530 15020 -27470
rect 13500 -27540 15020 -27530
rect 15220 -27560 15280 -26950
rect 15330 -26990 15390 -26980
rect 15330 -27060 15390 -27050
rect 15440 -27560 15500 -26950
rect 15700 -27230 15900 -27150
rect 16360 -27230 16560 -27150
rect 17020 -27230 17220 -27150
rect 15700 -27300 15900 -27290
rect 15700 -27360 15710 -27300
rect 15890 -27360 15900 -27300
rect 15700 -27370 15900 -27360
rect 16360 -27300 16560 -27290
rect 16360 -27360 16370 -27300
rect 16550 -27360 16560 -27300
rect 16360 -27370 16560 -27360
rect 17020 -27300 17220 -27290
rect 17020 -27360 17030 -27300
rect 17210 -27360 17220 -27300
rect 17020 -27370 17220 -27360
rect 15700 -27470 17220 -27460
rect 15700 -27530 15710 -27470
rect 17210 -27530 17220 -27470
rect 15700 -27540 17220 -27530
rect 17420 -27560 17480 -26950
rect 17530 -26990 17590 -26980
rect 17530 -27060 17590 -27050
rect 17640 -27560 17700 -26950
rect 17900 -27230 18100 -27150
rect 18560 -27230 18760 -27150
rect 19220 -27230 19420 -27150
rect 17900 -27300 18100 -27290
rect 17900 -27360 17910 -27300
rect 18090 -27360 18100 -27300
rect 17900 -27370 18100 -27360
rect 18560 -27300 18760 -27290
rect 18560 -27360 18570 -27300
rect 18750 -27360 18760 -27300
rect 18560 -27370 18760 -27360
rect 19220 -27300 19420 -27290
rect 19220 -27360 19230 -27300
rect 19410 -27360 19420 -27300
rect 19220 -27370 19420 -27360
rect 19620 -27560 19680 -26950
rect 19730 -26990 19790 -26980
rect 19730 -27060 19790 -27050
rect 19840 -27560 19900 -26950
rect 21930 -26990 21990 -26980
rect 21930 -27060 21990 -27050
rect 21300 -27430 21500 -27420
rect 21300 -27510 21310 -27430
rect 21490 -27510 21500 -27430
rect 21300 -27520 21500 -27510
rect 2010 -27730 2090 -27560
rect 2230 -27730 2310 -27560
rect 4210 -27680 4290 -27560
rect -70 -27790 -10 -27780
rect -70 -27860 -10 -27850
rect 420 -28230 620 -28220
rect 420 -28310 430 -28230
rect 610 -28310 620 -28230
rect 420 -28320 620 -28310
rect 2020 -28360 2080 -27730
rect 2130 -27790 2190 -27780
rect 2130 -27860 2190 -27850
rect 2240 -28360 2300 -27730
rect 4210 -27740 4220 -27680
rect 4280 -27740 4290 -27680
rect 4210 -27750 4290 -27740
rect 4430 -27750 4510 -27560
rect 6410 -27570 6490 -27560
rect 6410 -27630 6420 -27570
rect 6480 -27630 6490 -27570
rect 6410 -27750 6490 -27630
rect 6630 -27680 6710 -27560
rect 6630 -27740 6640 -27680
rect 6700 -27740 6710 -27680
rect 6630 -27750 6710 -27740
rect 8610 -27750 8690 -27560
rect 8830 -27570 8910 -27560
rect 8830 -27630 8840 -27570
rect 8900 -27630 8910 -27570
rect 8830 -27680 8910 -27630
rect 8830 -27740 8840 -27680
rect 8900 -27740 8910 -27680
rect 8830 -27750 8910 -27740
rect 10810 -27750 10890 -27560
rect 11030 -27570 11110 -27560
rect 11030 -27630 11040 -27570
rect 11100 -27630 11110 -27570
rect 11030 -27680 11110 -27630
rect 11030 -27740 11040 -27680
rect 11100 -27740 11110 -27680
rect 11030 -27750 11110 -27740
rect 13010 -27750 13090 -27560
rect 13230 -27570 13310 -27560
rect 13230 -27630 13240 -27570
rect 13300 -27630 13310 -27570
rect 13230 -27680 13310 -27630
rect 13230 -27740 13240 -27680
rect 13300 -27740 13310 -27680
rect 13230 -27750 13310 -27740
rect 15210 -27680 15290 -27560
rect 15210 -27740 15220 -27680
rect 15280 -27740 15290 -27680
rect 15210 -27750 15290 -27740
rect 15430 -27570 15510 -27560
rect 15430 -27630 15440 -27570
rect 15500 -27630 15510 -27570
rect 15430 -27750 15510 -27630
rect 17410 -27570 17490 -27560
rect 17410 -27630 17420 -27570
rect 17480 -27630 17490 -27570
rect 17410 -27750 17490 -27630
rect 17630 -27750 17710 -27560
rect 19610 -27750 19690 -27560
rect 19830 -27750 19910 -27560
rect 2500 -27960 2700 -27950
rect 2500 -28020 2510 -27960
rect 2690 -28020 2700 -27960
rect 2500 -28030 2700 -28020
rect 3160 -27960 3360 -27950
rect 3160 -28020 3170 -27960
rect 3350 -28020 3360 -27960
rect 3160 -28030 3360 -28020
rect 3820 -27960 4020 -27950
rect 3820 -28020 3830 -27960
rect 4010 -28020 4020 -27960
rect 3820 -28030 4020 -28020
rect 2500 -28170 2700 -28090
rect 3160 -28170 3360 -28090
rect 3820 -28170 4020 -28090
rect 4220 -28360 4280 -27750
rect 4330 -27790 4390 -27780
rect 4330 -27860 4390 -27850
rect 4440 -28360 4500 -27750
rect 4700 -27960 4900 -27950
rect 4700 -28020 4710 -27960
rect 4890 -28020 4900 -27960
rect 4700 -28030 4900 -28020
rect 5360 -27960 5560 -27950
rect 5360 -28020 5370 -27960
rect 5550 -28020 5560 -27960
rect 5360 -28030 5560 -28020
rect 6020 -27960 6220 -27950
rect 6020 -28020 6030 -27960
rect 6210 -28020 6220 -27960
rect 6020 -28030 6220 -28020
rect 4700 -28170 4900 -28090
rect 5360 -28170 5560 -28090
rect 6020 -28170 6220 -28090
rect 4700 -28270 6220 -28260
rect 4700 -28330 4710 -28270
rect 6210 -28330 6220 -28270
rect 4700 -28340 6220 -28330
rect 6420 -28360 6480 -27750
rect 6530 -27790 6590 -27780
rect 6530 -27860 6590 -27850
rect 6640 -28360 6700 -27750
rect 6900 -28030 7100 -27950
rect 7560 -28030 7760 -27950
rect 8220 -28030 8420 -27950
rect 6900 -28100 7100 -28090
rect 6900 -28160 6910 -28100
rect 7090 -28160 7100 -28100
rect 6900 -28170 7100 -28160
rect 7560 -28100 7760 -28090
rect 7560 -28160 7570 -28100
rect 7750 -28160 7760 -28100
rect 7560 -28170 7760 -28160
rect 8220 -28100 8420 -28090
rect 8220 -28160 8230 -28100
rect 8410 -28160 8420 -28100
rect 8220 -28170 8420 -28160
rect 6900 -28270 8420 -28260
rect 6900 -28330 6910 -28270
rect 8410 -28330 8420 -28270
rect 6900 -28340 8420 -28330
rect 8620 -28360 8680 -27750
rect 8730 -27790 8790 -27780
rect 8730 -27860 8790 -27850
rect 8840 -28360 8900 -27750
rect 9100 -28030 9300 -27950
rect 9760 -28030 9960 -27950
rect 10420 -28030 10620 -27950
rect 9100 -28100 9300 -28090
rect 9100 -28160 9110 -28100
rect 9290 -28160 9300 -28100
rect 9100 -28170 9300 -28160
rect 9760 -28100 9960 -28090
rect 9760 -28160 9770 -28100
rect 9950 -28160 9960 -28100
rect 9760 -28170 9960 -28160
rect 10420 -28100 10620 -28090
rect 10420 -28160 10430 -28100
rect 10610 -28160 10620 -28100
rect 10420 -28170 10620 -28160
rect 9100 -28270 10620 -28260
rect 9100 -28330 9110 -28270
rect 10610 -28330 10620 -28270
rect 9100 -28340 10620 -28330
rect 10820 -28360 10880 -27750
rect 10930 -27790 10990 -27780
rect 10930 -27860 10990 -27850
rect 11040 -28360 11100 -27750
rect 11300 -28030 11500 -27950
rect 11960 -28030 12160 -27950
rect 12620 -28030 12820 -27950
rect 11300 -28100 11500 -28090
rect 11300 -28160 11310 -28100
rect 11490 -28160 11500 -28100
rect 11300 -28170 11500 -28160
rect 11960 -28100 12160 -28090
rect 11960 -28160 11970 -28100
rect 12150 -28160 12160 -28100
rect 11960 -28170 12160 -28160
rect 12620 -28100 12820 -28090
rect 12620 -28160 12630 -28100
rect 12810 -28160 12820 -28100
rect 12620 -28170 12820 -28160
rect 11300 -28270 12820 -28260
rect 11300 -28330 11310 -28270
rect 12810 -28330 12820 -28270
rect 11300 -28340 12820 -28330
rect 13020 -28360 13080 -27750
rect 13130 -27790 13190 -27780
rect 13130 -27860 13190 -27850
rect 13240 -28360 13300 -27750
rect 13500 -28030 13700 -27950
rect 14160 -28030 14360 -27950
rect 14820 -28030 15020 -27950
rect 13500 -28100 13700 -28090
rect 13500 -28160 13510 -28100
rect 13690 -28160 13700 -28100
rect 13500 -28170 13700 -28160
rect 14160 -28100 14360 -28090
rect 14160 -28160 14170 -28100
rect 14350 -28160 14360 -28100
rect 14160 -28170 14360 -28160
rect 14820 -28100 15020 -28090
rect 14820 -28160 14830 -28100
rect 15010 -28160 15020 -28100
rect 14820 -28170 15020 -28160
rect 13500 -28270 15020 -28260
rect 13500 -28330 13510 -28270
rect 15010 -28330 15020 -28270
rect 13500 -28340 15020 -28330
rect 15220 -28360 15280 -27750
rect 15330 -27790 15390 -27780
rect 15330 -27860 15390 -27850
rect 15440 -28360 15500 -27750
rect 15700 -27960 15900 -27950
rect 15700 -28020 15710 -27960
rect 15890 -28020 15900 -27960
rect 15700 -28030 15900 -28020
rect 16360 -27960 16560 -27950
rect 16360 -28020 16370 -27960
rect 16550 -28020 16560 -27960
rect 16360 -28030 16560 -28020
rect 17020 -27960 17220 -27950
rect 17020 -28020 17030 -27960
rect 17210 -28020 17220 -27960
rect 17020 -28030 17220 -28020
rect 15700 -28170 15900 -28090
rect 16360 -28170 16560 -28090
rect 17020 -28170 17220 -28090
rect 15700 -28270 17220 -28260
rect 15700 -28330 15710 -28270
rect 17210 -28330 17220 -28270
rect 15700 -28340 17220 -28330
rect 17420 -28360 17480 -27750
rect 17530 -27790 17590 -27780
rect 17530 -27860 17590 -27850
rect 17640 -28360 17700 -27750
rect 17900 -27960 18100 -27950
rect 17900 -28020 17910 -27960
rect 18090 -28020 18100 -27960
rect 17900 -28030 18100 -28020
rect 18560 -27960 18760 -27950
rect 18560 -28020 18570 -27960
rect 18750 -28020 18760 -27960
rect 18560 -28030 18760 -28020
rect 19220 -27960 19420 -27950
rect 19220 -28020 19230 -27960
rect 19410 -28020 19420 -27960
rect 19220 -28030 19420 -28020
rect 17900 -28170 18100 -28090
rect 18560 -28170 18760 -28090
rect 19220 -28170 19420 -28090
rect 19620 -28360 19680 -27750
rect 19730 -27790 19790 -27780
rect 19730 -27860 19790 -27850
rect 19840 -28360 19900 -27750
rect 21930 -27790 21990 -27780
rect 21930 -27860 21990 -27850
rect 21300 -28230 21500 -28220
rect 21300 -28310 21310 -28230
rect 21490 -28310 21500 -28230
rect 21300 -28320 21500 -28310
rect 2010 -28530 2090 -28360
rect 2230 -28530 2310 -28360
rect 4210 -28480 4290 -28360
rect -70 -28590 -10 -28580
rect -70 -28660 -10 -28650
rect 420 -29030 620 -29020
rect 420 -29110 430 -29030
rect 610 -29110 620 -29030
rect 420 -29120 620 -29110
rect 2020 -29160 2080 -28530
rect 2130 -28590 2190 -28580
rect 2130 -28660 2190 -28650
rect 2240 -29160 2300 -28530
rect 4210 -28540 4220 -28480
rect 4280 -28540 4290 -28480
rect 4210 -28550 4290 -28540
rect 4430 -28550 4510 -28360
rect 6410 -28370 6490 -28360
rect 6410 -28430 6420 -28370
rect 6480 -28430 6490 -28370
rect 6410 -28550 6490 -28430
rect 6630 -28480 6710 -28360
rect 6630 -28540 6640 -28480
rect 6700 -28540 6710 -28480
rect 6630 -28550 6710 -28540
rect 8610 -28550 8690 -28360
rect 8830 -28370 8910 -28360
rect 8830 -28430 8840 -28370
rect 8900 -28430 8910 -28370
rect 8830 -28480 8910 -28430
rect 8830 -28540 8840 -28480
rect 8900 -28540 8910 -28480
rect 8830 -28550 8910 -28540
rect 10810 -28550 10890 -28360
rect 11030 -28370 11110 -28360
rect 11030 -28430 11040 -28370
rect 11100 -28430 11110 -28370
rect 11030 -28480 11110 -28430
rect 11030 -28540 11040 -28480
rect 11100 -28540 11110 -28480
rect 11030 -28550 11110 -28540
rect 13010 -28550 13090 -28360
rect 13230 -28370 13310 -28360
rect 13230 -28430 13240 -28370
rect 13300 -28430 13310 -28370
rect 13230 -28480 13310 -28430
rect 13230 -28540 13240 -28480
rect 13300 -28540 13310 -28480
rect 13230 -28550 13310 -28540
rect 15210 -28480 15290 -28360
rect 15210 -28540 15220 -28480
rect 15280 -28540 15290 -28480
rect 15210 -28550 15290 -28540
rect 15430 -28370 15510 -28360
rect 15430 -28430 15440 -28370
rect 15500 -28430 15510 -28370
rect 15430 -28550 15510 -28430
rect 17410 -28370 17490 -28360
rect 17410 -28430 17420 -28370
rect 17480 -28430 17490 -28370
rect 17410 -28550 17490 -28430
rect 17630 -28550 17710 -28360
rect 19610 -28550 19690 -28360
rect 19830 -28550 19910 -28360
rect 2500 -28760 2700 -28750
rect 2500 -28820 2510 -28760
rect 2690 -28820 2700 -28760
rect 2500 -28830 2700 -28820
rect 3160 -28760 3360 -28750
rect 3160 -28820 3170 -28760
rect 3350 -28820 3360 -28760
rect 3160 -28830 3360 -28820
rect 3820 -28760 4020 -28750
rect 3820 -28820 3830 -28760
rect 4010 -28820 4020 -28760
rect 3820 -28830 4020 -28820
rect 2500 -28970 2700 -28890
rect 3160 -28970 3360 -28890
rect 3820 -28970 4020 -28890
rect 4220 -29160 4280 -28550
rect 4330 -28590 4390 -28580
rect 4330 -28660 4390 -28650
rect 4440 -29160 4500 -28550
rect 4700 -28760 4900 -28750
rect 4700 -28820 4710 -28760
rect 4890 -28820 4900 -28760
rect 4700 -28830 4900 -28820
rect 5360 -28760 5560 -28750
rect 5360 -28820 5370 -28760
rect 5550 -28820 5560 -28760
rect 5360 -28830 5560 -28820
rect 6020 -28760 6220 -28750
rect 6020 -28820 6030 -28760
rect 6210 -28820 6220 -28760
rect 6020 -28830 6220 -28820
rect 4700 -28970 4900 -28890
rect 5360 -28970 5560 -28890
rect 6020 -28970 6220 -28890
rect 4700 -29070 6220 -29060
rect 4700 -29130 4710 -29070
rect 6210 -29130 6220 -29070
rect 4700 -29140 6220 -29130
rect 6420 -29160 6480 -28550
rect 6530 -28590 6590 -28580
rect 6530 -28660 6590 -28650
rect 6640 -29160 6700 -28550
rect 6900 -28830 7100 -28750
rect 7560 -28830 7760 -28750
rect 8220 -28830 8420 -28750
rect 6900 -28900 7100 -28890
rect 6900 -28960 6910 -28900
rect 7090 -28960 7100 -28900
rect 6900 -28970 7100 -28960
rect 7560 -28900 7760 -28890
rect 7560 -28960 7570 -28900
rect 7750 -28960 7760 -28900
rect 7560 -28970 7760 -28960
rect 8220 -28900 8420 -28890
rect 8220 -28960 8230 -28900
rect 8410 -28960 8420 -28900
rect 8220 -28970 8420 -28960
rect 6900 -29070 8420 -29060
rect 6900 -29130 6910 -29070
rect 8410 -29130 8420 -29070
rect 6900 -29140 8420 -29130
rect 8620 -29160 8680 -28550
rect 8730 -28590 8790 -28580
rect 8730 -28660 8790 -28650
rect 8840 -29160 8900 -28550
rect 9100 -28830 9300 -28750
rect 9760 -28830 9960 -28750
rect 10420 -28830 10620 -28750
rect 9100 -28900 9300 -28890
rect 9100 -28960 9110 -28900
rect 9290 -28960 9300 -28900
rect 9100 -28970 9300 -28960
rect 9760 -28900 9960 -28890
rect 9760 -28960 9770 -28900
rect 9950 -28960 9960 -28900
rect 9760 -28970 9960 -28960
rect 10420 -28900 10620 -28890
rect 10420 -28960 10430 -28900
rect 10610 -28960 10620 -28900
rect 10420 -28970 10620 -28960
rect 9100 -29070 10620 -29060
rect 9100 -29130 9110 -29070
rect 10610 -29130 10620 -29070
rect 9100 -29140 10620 -29130
rect 10820 -29160 10880 -28550
rect 10930 -28590 10990 -28580
rect 10930 -28660 10990 -28650
rect 11040 -29160 11100 -28550
rect 11300 -28830 11500 -28750
rect 11960 -28830 12160 -28750
rect 12620 -28830 12820 -28750
rect 11300 -28900 11500 -28890
rect 11300 -28960 11310 -28900
rect 11490 -28960 11500 -28900
rect 11300 -28970 11500 -28960
rect 11960 -28900 12160 -28890
rect 11960 -28960 11970 -28900
rect 12150 -28960 12160 -28900
rect 11960 -28970 12160 -28960
rect 12620 -28900 12820 -28890
rect 12620 -28960 12630 -28900
rect 12810 -28960 12820 -28900
rect 12620 -28970 12820 -28960
rect 11300 -29070 12820 -29060
rect 11300 -29130 11310 -29070
rect 12810 -29130 12820 -29070
rect 11300 -29140 12820 -29130
rect 13020 -29160 13080 -28550
rect 13130 -28590 13190 -28580
rect 13130 -28660 13190 -28650
rect 13240 -29160 13300 -28550
rect 13500 -28830 13700 -28750
rect 14160 -28830 14360 -28750
rect 14820 -28830 15020 -28750
rect 13500 -28900 13700 -28890
rect 13500 -28960 13510 -28900
rect 13690 -28960 13700 -28900
rect 13500 -28970 13700 -28960
rect 14160 -28900 14360 -28890
rect 14160 -28960 14170 -28900
rect 14350 -28960 14360 -28900
rect 14160 -28970 14360 -28960
rect 14820 -28900 15020 -28890
rect 14820 -28960 14830 -28900
rect 15010 -28960 15020 -28900
rect 14820 -28970 15020 -28960
rect 13500 -29070 15020 -29060
rect 13500 -29130 13510 -29070
rect 15010 -29130 15020 -29070
rect 13500 -29140 15020 -29130
rect 15220 -29160 15280 -28550
rect 15330 -28590 15390 -28580
rect 15330 -28660 15390 -28650
rect 15440 -29160 15500 -28550
rect 15700 -28760 15900 -28750
rect 15700 -28820 15710 -28760
rect 15890 -28820 15900 -28760
rect 15700 -28830 15900 -28820
rect 16360 -28760 16560 -28750
rect 16360 -28820 16370 -28760
rect 16550 -28820 16560 -28760
rect 16360 -28830 16560 -28820
rect 17020 -28760 17220 -28750
rect 17020 -28820 17030 -28760
rect 17210 -28820 17220 -28760
rect 17020 -28830 17220 -28820
rect 15700 -28970 15900 -28890
rect 16360 -28970 16560 -28890
rect 17020 -28970 17220 -28890
rect 15700 -29070 17220 -29060
rect 15700 -29130 15710 -29070
rect 17210 -29130 17220 -29070
rect 15700 -29140 17220 -29130
rect 17420 -29160 17480 -28550
rect 17530 -28590 17590 -28580
rect 17530 -28660 17590 -28650
rect 17640 -29160 17700 -28550
rect 17900 -28760 18100 -28750
rect 17900 -28820 17910 -28760
rect 18090 -28820 18100 -28760
rect 17900 -28830 18100 -28820
rect 18560 -28760 18760 -28750
rect 18560 -28820 18570 -28760
rect 18750 -28820 18760 -28760
rect 18560 -28830 18760 -28820
rect 19220 -28760 19420 -28750
rect 19220 -28820 19230 -28760
rect 19410 -28820 19420 -28760
rect 19220 -28830 19420 -28820
rect 17900 -28970 18100 -28890
rect 18560 -28970 18760 -28890
rect 19220 -28970 19420 -28890
rect 19620 -29160 19680 -28550
rect 19730 -28590 19790 -28580
rect 19730 -28660 19790 -28650
rect 19840 -29160 19900 -28550
rect 21930 -28590 21990 -28580
rect 21930 -28660 21990 -28650
rect 21300 -29030 21500 -29020
rect 21300 -29110 21310 -29030
rect 21490 -29110 21500 -29030
rect 21300 -29120 21500 -29110
rect 2010 -29330 2090 -29160
rect 2230 -29330 2310 -29160
rect -70 -29390 -10 -29380
rect -70 -29460 -10 -29450
rect 2020 -29960 2080 -29330
rect 2130 -29390 2190 -29380
rect 2130 -29460 2190 -29450
rect 2240 -29960 2300 -29330
rect 4210 -29350 4290 -29160
rect 4430 -29280 4510 -29160
rect 4430 -29340 4440 -29280
rect 4500 -29340 4510 -29280
rect 4430 -29350 4510 -29340
rect 6410 -29280 6490 -29160
rect 6410 -29340 6420 -29280
rect 6480 -29340 6490 -29280
rect 6410 -29350 6490 -29340
rect 6630 -29170 6710 -29160
rect 6630 -29230 6640 -29170
rect 6700 -29230 6710 -29170
rect 6630 -29350 6710 -29230
rect 8610 -29170 8690 -29160
rect 8610 -29230 8620 -29170
rect 8680 -29230 8690 -29170
rect 8610 -29280 8690 -29230
rect 8610 -29340 8620 -29280
rect 8680 -29340 8690 -29280
rect 8610 -29350 8690 -29340
rect 8830 -29350 8910 -29160
rect 10810 -29170 10890 -29160
rect 10810 -29230 10820 -29170
rect 10880 -29230 10890 -29170
rect 10810 -29280 10890 -29230
rect 10810 -29340 10820 -29280
rect 10880 -29340 10890 -29280
rect 10810 -29350 10890 -29340
rect 11030 -29350 11110 -29160
rect 13010 -29170 13090 -29160
rect 13010 -29230 13020 -29170
rect 13080 -29230 13090 -29170
rect 13010 -29280 13090 -29230
rect 13010 -29340 13020 -29280
rect 13080 -29340 13090 -29280
rect 13010 -29350 13090 -29340
rect 13230 -29350 13310 -29160
rect 15210 -29170 15290 -29160
rect 15210 -29230 15220 -29170
rect 15280 -29230 15290 -29170
rect 15210 -29350 15290 -29230
rect 15430 -29280 15510 -29160
rect 15430 -29340 15440 -29280
rect 15500 -29340 15510 -29280
rect 15430 -29350 15510 -29340
rect 17410 -29350 17490 -29160
rect 17630 -29170 17710 -29160
rect 17630 -29230 17640 -29170
rect 17700 -29230 17710 -29170
rect 17630 -29350 17710 -29230
rect 19610 -29350 19690 -29160
rect 19830 -29350 19910 -29160
rect 2500 -29630 2700 -29550
rect 3160 -29630 3360 -29550
rect 3820 -29630 4020 -29550
rect 2500 -29700 2700 -29690
rect 2500 -29760 2510 -29700
rect 2690 -29760 2700 -29700
rect 2500 -29770 2700 -29760
rect 3160 -29700 3360 -29690
rect 3160 -29760 3170 -29700
rect 3350 -29760 3360 -29700
rect 3160 -29770 3360 -29760
rect 3820 -29700 4020 -29690
rect 3820 -29760 3830 -29700
rect 4010 -29760 4020 -29700
rect 3820 -29770 4020 -29760
rect 2500 -29870 4020 -29860
rect 2500 -29930 2510 -29870
rect 4010 -29930 4020 -29870
rect 2500 -29940 4020 -29930
rect 4220 -29960 4280 -29350
rect 4330 -29390 4390 -29380
rect 4330 -29460 4390 -29450
rect 4440 -29960 4500 -29350
rect 4700 -29630 4900 -29550
rect 5360 -29630 5560 -29550
rect 6020 -29630 6220 -29550
rect 4700 -29700 4900 -29690
rect 4700 -29760 4710 -29700
rect 4890 -29760 4900 -29700
rect 4700 -29770 4900 -29760
rect 5360 -29700 5560 -29690
rect 5360 -29760 5370 -29700
rect 5550 -29760 5560 -29700
rect 5360 -29770 5560 -29760
rect 6020 -29700 6220 -29690
rect 6020 -29760 6030 -29700
rect 6210 -29760 6220 -29700
rect 6020 -29770 6220 -29760
rect 4700 -29870 6220 -29860
rect 4700 -29930 4710 -29870
rect 6210 -29930 6220 -29870
rect 4700 -29940 6220 -29930
rect 6420 -29960 6480 -29350
rect 6530 -29390 6590 -29380
rect 6530 -29460 6590 -29450
rect 6640 -29960 6700 -29350
rect 6900 -29560 7100 -29550
rect 6900 -29620 6910 -29560
rect 7090 -29620 7100 -29560
rect 6900 -29630 7100 -29620
rect 7560 -29560 7760 -29550
rect 7560 -29620 7570 -29560
rect 7750 -29620 7760 -29560
rect 7560 -29630 7760 -29620
rect 8220 -29560 8420 -29550
rect 8220 -29620 8230 -29560
rect 8410 -29620 8420 -29560
rect 8220 -29630 8420 -29620
rect 6900 -29770 7100 -29690
rect 7560 -29770 7760 -29690
rect 8220 -29770 8420 -29690
rect 6900 -29870 8420 -29860
rect 6900 -29930 6910 -29870
rect 8410 -29930 8420 -29870
rect 6900 -29940 8420 -29930
rect 8620 -29960 8680 -29350
rect 8730 -29390 8790 -29380
rect 8730 -29460 8790 -29450
rect 8840 -29960 8900 -29350
rect 9100 -29560 9300 -29550
rect 9100 -29620 9110 -29560
rect 9290 -29620 9300 -29560
rect 9100 -29630 9300 -29620
rect 9760 -29560 9960 -29550
rect 9760 -29620 9770 -29560
rect 9950 -29620 9960 -29560
rect 9760 -29630 9960 -29620
rect 10420 -29560 10620 -29550
rect 10420 -29620 10430 -29560
rect 10610 -29620 10620 -29560
rect 10420 -29630 10620 -29620
rect 9100 -29770 9300 -29690
rect 9760 -29770 9960 -29690
rect 10420 -29770 10620 -29690
rect 9100 -29870 10620 -29860
rect 9100 -29930 9110 -29870
rect 10610 -29930 10620 -29870
rect 9100 -29940 10620 -29930
rect 10820 -29960 10880 -29350
rect 10930 -29390 10990 -29380
rect 10930 -29460 10990 -29450
rect 11040 -29960 11100 -29350
rect 11300 -29560 11500 -29550
rect 11300 -29620 11310 -29560
rect 11490 -29620 11500 -29560
rect 11300 -29630 11500 -29620
rect 11960 -29560 12160 -29550
rect 11960 -29620 11970 -29560
rect 12150 -29620 12160 -29560
rect 11960 -29630 12160 -29620
rect 12620 -29560 12820 -29550
rect 12620 -29620 12630 -29560
rect 12810 -29620 12820 -29560
rect 12620 -29630 12820 -29620
rect 11300 -29770 11500 -29690
rect 11960 -29770 12160 -29690
rect 12620 -29770 12820 -29690
rect 11300 -29870 12820 -29860
rect 11300 -29930 11310 -29870
rect 12810 -29930 12820 -29870
rect 11300 -29940 12820 -29930
rect 13020 -29960 13080 -29350
rect 13130 -29390 13190 -29380
rect 13130 -29460 13190 -29450
rect 13240 -29960 13300 -29350
rect 13500 -29560 13700 -29550
rect 13500 -29620 13510 -29560
rect 13690 -29620 13700 -29560
rect 13500 -29630 13700 -29620
rect 14160 -29560 14360 -29550
rect 14160 -29620 14170 -29560
rect 14350 -29620 14360 -29560
rect 14160 -29630 14360 -29620
rect 14820 -29560 15020 -29550
rect 14820 -29620 14830 -29560
rect 15010 -29620 15020 -29560
rect 14820 -29630 15020 -29620
rect 13500 -29770 13700 -29690
rect 14160 -29770 14360 -29690
rect 14820 -29770 15020 -29690
rect 13500 -29870 15020 -29860
rect 13500 -29930 13510 -29870
rect 15010 -29930 15020 -29870
rect 13500 -29940 15020 -29930
rect 15220 -29960 15280 -29350
rect 15330 -29390 15390 -29380
rect 15330 -29460 15390 -29450
rect 15440 -29960 15500 -29350
rect 15700 -29630 15900 -29550
rect 16360 -29630 16560 -29550
rect 17020 -29630 17220 -29550
rect 15700 -29700 15900 -29690
rect 15700 -29760 15710 -29700
rect 15890 -29760 15900 -29700
rect 15700 -29770 15900 -29760
rect 16360 -29700 16560 -29690
rect 16360 -29760 16370 -29700
rect 16550 -29760 16560 -29700
rect 16360 -29770 16560 -29760
rect 17020 -29700 17220 -29690
rect 17020 -29760 17030 -29700
rect 17210 -29760 17220 -29700
rect 17020 -29770 17220 -29760
rect 15700 -29870 17220 -29860
rect 15700 -29930 15710 -29870
rect 17210 -29930 17220 -29870
rect 15700 -29940 17220 -29930
rect 17420 -29960 17480 -29350
rect 17530 -29390 17590 -29380
rect 17530 -29460 17590 -29450
rect 17640 -29960 17700 -29350
rect 17900 -29630 18100 -29550
rect 18560 -29630 18760 -29550
rect 19220 -29630 19420 -29550
rect 17900 -29700 18100 -29690
rect 17900 -29760 17910 -29700
rect 18090 -29760 18100 -29700
rect 17900 -29770 18100 -29760
rect 18560 -29700 18760 -29690
rect 18560 -29760 18570 -29700
rect 18750 -29760 18760 -29700
rect 18560 -29770 18760 -29760
rect 19220 -29700 19420 -29690
rect 19220 -29760 19230 -29700
rect 19410 -29760 19420 -29700
rect 19220 -29770 19420 -29760
rect 17900 -29870 19420 -29860
rect 17900 -29930 17910 -29870
rect 19410 -29930 19420 -29870
rect 17900 -29940 19420 -29930
rect 19620 -29960 19680 -29350
rect 19730 -29390 19790 -29380
rect 19730 -29460 19790 -29450
rect 19840 -29960 19900 -29350
rect 21930 -29390 21990 -29380
rect 21930 -29460 21990 -29450
rect 2010 -30060 2090 -29960
rect 2010 -30120 2020 -30060
rect 2080 -30120 2090 -30060
rect 2010 -30130 2090 -30120
rect 2230 -30130 2310 -29960
rect 4210 -29970 4290 -29960
rect 4210 -30030 4220 -29970
rect 4280 -30030 4290 -29970
rect 4210 -30080 4290 -30030
rect -70 -30190 -10 -30180
rect -70 -30260 -10 -30250
rect 2020 -30760 2080 -30130
rect 2130 -30190 2190 -30180
rect 2130 -30260 2190 -30250
rect 2240 -30760 2300 -30130
rect 4210 -30140 4220 -30080
rect 4280 -30140 4290 -30080
rect 4210 -30150 4290 -30140
rect 4430 -30150 4510 -29960
rect 6410 -29970 6490 -29960
rect 6410 -30030 6420 -29970
rect 6480 -30030 6490 -29970
rect 6410 -30150 6490 -30030
rect 6630 -30080 6710 -29960
rect 6630 -30140 6640 -30080
rect 6700 -30140 6710 -30080
rect 6630 -30150 6710 -30140
rect 8610 -30150 8690 -29960
rect 8830 -29970 8910 -29960
rect 8830 -30030 8840 -29970
rect 8900 -30030 8910 -29970
rect 8830 -30080 8910 -30030
rect 8830 -30140 8840 -30080
rect 8900 -30140 8910 -30080
rect 8830 -30150 8910 -30140
rect 10810 -30150 10890 -29960
rect 11030 -29970 11110 -29960
rect 11030 -30030 11040 -29970
rect 11100 -30030 11110 -29970
rect 11030 -30080 11110 -30030
rect 11030 -30140 11040 -30080
rect 11100 -30140 11110 -30080
rect 11030 -30150 11110 -30140
rect 13010 -30150 13090 -29960
rect 13230 -29970 13310 -29960
rect 13230 -30030 13240 -29970
rect 13300 -30030 13310 -29970
rect 13230 -30080 13310 -30030
rect 13230 -30140 13240 -30080
rect 13300 -30140 13310 -30080
rect 13230 -30150 13310 -30140
rect 15210 -30080 15290 -29960
rect 15210 -30140 15220 -30080
rect 15280 -30140 15290 -30080
rect 15210 -30150 15290 -30140
rect 15430 -29970 15510 -29960
rect 15430 -30030 15440 -29970
rect 15500 -30030 15510 -29970
rect 15430 -30150 15510 -30030
rect 17410 -29970 17490 -29960
rect 17410 -30030 17420 -29970
rect 17480 -30030 17490 -29970
rect 17410 -30080 17490 -30030
rect 17410 -30140 17420 -30080
rect 17480 -30140 17490 -30080
rect 17410 -30150 17490 -30140
rect 17630 -30150 17710 -29960
rect 19610 -29970 19690 -29960
rect 19610 -30030 19620 -29970
rect 19680 -30030 19690 -29970
rect 19610 -30150 19690 -30030
rect 19830 -30150 19910 -29960
rect 2500 -30360 2700 -30350
rect 2500 -30420 2510 -30360
rect 2690 -30420 2700 -30360
rect 2500 -30430 2700 -30420
rect 3160 -30360 3360 -30350
rect 3160 -30420 3170 -30360
rect 3350 -30420 3360 -30360
rect 3160 -30430 3360 -30420
rect 3820 -30360 4020 -30350
rect 3820 -30420 3830 -30360
rect 4010 -30420 4020 -30360
rect 3820 -30430 4020 -30420
rect 2500 -30570 2700 -30490
rect 3160 -30570 3360 -30490
rect 3820 -30570 4020 -30490
rect 2500 -30670 4020 -30660
rect 2500 -30730 2510 -30670
rect 4010 -30730 4020 -30670
rect 2500 -30740 4020 -30730
rect 4220 -30760 4280 -30150
rect 4330 -30190 4390 -30180
rect 4330 -30260 4390 -30250
rect 4440 -30760 4500 -30150
rect 4700 -30360 4900 -30350
rect 4700 -30420 4710 -30360
rect 4890 -30420 4900 -30360
rect 4700 -30430 4900 -30420
rect 5360 -30360 5560 -30350
rect 5360 -30420 5370 -30360
rect 5550 -30420 5560 -30360
rect 5360 -30430 5560 -30420
rect 6020 -30360 6220 -30350
rect 6020 -30420 6030 -30360
rect 6210 -30420 6220 -30360
rect 6020 -30430 6220 -30420
rect 4700 -30570 4900 -30490
rect 5360 -30570 5560 -30490
rect 6020 -30570 6220 -30490
rect 4700 -30670 6220 -30660
rect 4700 -30730 4710 -30670
rect 6210 -30730 6220 -30670
rect 4700 -30740 6220 -30730
rect 6420 -30760 6480 -30150
rect 6530 -30190 6590 -30180
rect 6530 -30260 6590 -30250
rect 6640 -30760 6700 -30150
rect 6900 -30430 7100 -30350
rect 7560 -30430 7760 -30350
rect 8220 -30430 8420 -30350
rect 6900 -30500 7100 -30490
rect 6900 -30560 6910 -30500
rect 7090 -30560 7100 -30500
rect 6900 -30570 7100 -30560
rect 7560 -30500 7760 -30490
rect 7560 -30560 7570 -30500
rect 7750 -30560 7760 -30500
rect 7560 -30570 7760 -30560
rect 8220 -30500 8420 -30490
rect 8220 -30560 8230 -30500
rect 8410 -30560 8420 -30500
rect 8220 -30570 8420 -30560
rect 6900 -30670 8420 -30660
rect 6900 -30730 6910 -30670
rect 8410 -30730 8420 -30670
rect 6900 -30740 8420 -30730
rect 8620 -30760 8680 -30150
rect 8730 -30190 8790 -30180
rect 8730 -30260 8790 -30250
rect 8840 -30760 8900 -30150
rect 9100 -30430 9300 -30350
rect 9760 -30430 9960 -30350
rect 10420 -30430 10620 -30350
rect 9100 -30500 9300 -30490
rect 9100 -30560 9110 -30500
rect 9290 -30560 9300 -30500
rect 9100 -30570 9300 -30560
rect 9760 -30500 9960 -30490
rect 9760 -30560 9770 -30500
rect 9950 -30560 9960 -30500
rect 9760 -30570 9960 -30560
rect 10420 -30500 10620 -30490
rect 10420 -30560 10430 -30500
rect 10610 -30560 10620 -30500
rect 10420 -30570 10620 -30560
rect 9100 -30670 10620 -30660
rect 9100 -30730 9110 -30670
rect 10610 -30730 10620 -30670
rect 9100 -30740 10620 -30730
rect 10820 -30760 10880 -30150
rect 10930 -30190 10990 -30180
rect 10930 -30260 10990 -30250
rect 11040 -30760 11100 -30150
rect 11300 -30430 11500 -30350
rect 11960 -30430 12160 -30350
rect 12620 -30430 12820 -30350
rect 11300 -30500 11500 -30490
rect 11300 -30560 11310 -30500
rect 11490 -30560 11500 -30500
rect 11300 -30570 11500 -30560
rect 11960 -30500 12160 -30490
rect 11960 -30560 11970 -30500
rect 12150 -30560 12160 -30500
rect 11960 -30570 12160 -30560
rect 12620 -30500 12820 -30490
rect 12620 -30560 12630 -30500
rect 12810 -30560 12820 -30500
rect 12620 -30570 12820 -30560
rect 11300 -30670 12820 -30660
rect 11300 -30730 11310 -30670
rect 12810 -30730 12820 -30670
rect 11300 -30740 12820 -30730
rect 13020 -30760 13080 -30150
rect 13130 -30190 13190 -30180
rect 13130 -30260 13190 -30250
rect 13240 -30760 13300 -30150
rect 13500 -30430 13700 -30350
rect 14160 -30430 14360 -30350
rect 14820 -30430 15020 -30350
rect 13500 -30500 13700 -30490
rect 13500 -30560 13510 -30500
rect 13690 -30560 13700 -30500
rect 13500 -30570 13700 -30560
rect 14160 -30500 14360 -30490
rect 14160 -30560 14170 -30500
rect 14350 -30560 14360 -30500
rect 14160 -30570 14360 -30560
rect 14820 -30500 15020 -30490
rect 14820 -30560 14830 -30500
rect 15010 -30560 15020 -30500
rect 14820 -30570 15020 -30560
rect 13500 -30670 15020 -30660
rect 13500 -30730 13510 -30670
rect 15010 -30730 15020 -30670
rect 13500 -30740 15020 -30730
rect 15220 -30760 15280 -30150
rect 15330 -30190 15390 -30180
rect 15330 -30260 15390 -30250
rect 15440 -30760 15500 -30150
rect 15700 -30360 15900 -30350
rect 15700 -30420 15710 -30360
rect 15890 -30420 15900 -30360
rect 15700 -30430 15900 -30420
rect 16360 -30360 16560 -30350
rect 16360 -30420 16370 -30360
rect 16550 -30420 16560 -30360
rect 16360 -30430 16560 -30420
rect 17020 -30360 17220 -30350
rect 17020 -30420 17030 -30360
rect 17210 -30420 17220 -30360
rect 17020 -30430 17220 -30420
rect 15700 -30570 15900 -30490
rect 16360 -30570 16560 -30490
rect 17020 -30570 17220 -30490
rect 15700 -30670 17220 -30660
rect 15700 -30730 15710 -30670
rect 17210 -30730 17220 -30670
rect 15700 -30740 17220 -30730
rect 17420 -30760 17480 -30150
rect 17530 -30190 17590 -30180
rect 17530 -30260 17590 -30250
rect 17640 -30760 17700 -30150
rect 17900 -30360 18100 -30350
rect 17900 -30420 17910 -30360
rect 18090 -30420 18100 -30360
rect 17900 -30430 18100 -30420
rect 18560 -30360 18760 -30350
rect 18560 -30420 18570 -30360
rect 18750 -30420 18760 -30360
rect 18560 -30430 18760 -30420
rect 19220 -30360 19420 -30350
rect 19220 -30420 19230 -30360
rect 19410 -30420 19420 -30360
rect 19220 -30430 19420 -30420
rect 17900 -30570 18100 -30490
rect 18560 -30570 18760 -30490
rect 19220 -30570 19420 -30490
rect 17900 -30670 19420 -30660
rect 17900 -30730 17910 -30670
rect 19410 -30730 19420 -30670
rect 17900 -30740 19420 -30730
rect 19620 -30760 19680 -30150
rect 19730 -30190 19790 -30180
rect 19730 -30260 19790 -30250
rect 19840 -30760 19900 -30150
rect 21930 -30190 21990 -30180
rect 21930 -30260 21990 -30250
rect 2010 -30930 2090 -30760
rect 2230 -30860 2310 -30760
rect 2230 -30920 2240 -30860
rect 2300 -30920 2310 -30860
rect 2230 -30930 2310 -30920
rect -70 -30990 -10 -30980
rect -70 -31060 -10 -31050
rect 2020 -32420 2080 -30930
rect 2130 -30990 2190 -30980
rect 2130 -31060 2190 -31050
rect 2240 -32420 2300 -30930
rect 4210 -30950 4290 -30760
rect 4430 -30770 4510 -30760
rect 4430 -30830 4440 -30770
rect 4500 -30830 4510 -30770
rect 4430 -30880 4510 -30830
rect 4430 -30940 4440 -30880
rect 4500 -30940 4510 -30880
rect 4430 -30950 4510 -30940
rect 6410 -30880 6490 -30760
rect 6410 -30940 6420 -30880
rect 6480 -30940 6490 -30880
rect 6410 -30950 6490 -30940
rect 6630 -30770 6710 -30760
rect 6630 -30830 6640 -30770
rect 6700 -30830 6710 -30770
rect 6630 -30950 6710 -30830
rect 8610 -30770 8690 -30760
rect 8610 -30830 8620 -30770
rect 8680 -30830 8690 -30770
rect 8610 -30880 8690 -30830
rect 8610 -30940 8620 -30880
rect 8680 -30940 8690 -30880
rect 8610 -30950 8690 -30940
rect 8830 -30950 8910 -30760
rect 10810 -30770 10890 -30760
rect 10810 -30830 10820 -30770
rect 10880 -30830 10890 -30770
rect 10810 -30880 10890 -30830
rect 10810 -30940 10820 -30880
rect 10880 -30940 10890 -30880
rect 10810 -30950 10890 -30940
rect 11030 -30950 11110 -30760
rect 13010 -30770 13090 -30760
rect 13010 -30830 13020 -30770
rect 13080 -30830 13090 -30770
rect 13010 -30880 13090 -30830
rect 13010 -30940 13020 -30880
rect 13080 -30940 13090 -30880
rect 13010 -30950 13090 -30940
rect 13230 -30950 13310 -30760
rect 15210 -30770 15290 -30760
rect 15210 -30830 15220 -30770
rect 15280 -30830 15290 -30770
rect 15210 -30950 15290 -30830
rect 15430 -30880 15510 -30760
rect 15430 -30940 15440 -30880
rect 15500 -30940 15510 -30880
rect 15430 -30950 15510 -30940
rect 17410 -30950 17490 -30760
rect 17630 -30770 17710 -30760
rect 17630 -30830 17640 -30770
rect 17700 -30830 17710 -30770
rect 17630 -30880 17710 -30830
rect 17630 -30940 17640 -30880
rect 17700 -30940 17710 -30880
rect 17630 -30950 17710 -30940
rect 19610 -30950 19690 -30760
rect 19830 -30770 19910 -30760
rect 19830 -30830 19840 -30770
rect 19900 -30830 19910 -30770
rect 19830 -30950 19910 -30830
rect 2500 -31230 2700 -31150
rect 3160 -31230 3360 -31150
rect 3820 -31230 4020 -31150
rect 2500 -31300 2700 -31290
rect 2500 -31360 2510 -31300
rect 2690 -31360 2700 -31300
rect 2500 -31370 2700 -31360
rect 3160 -31300 3360 -31290
rect 3160 -31360 3170 -31300
rect 3350 -31360 3360 -31300
rect 3160 -31370 3360 -31360
rect 3820 -31300 4020 -31290
rect 3820 -31360 3830 -31300
rect 4010 -31360 4020 -31300
rect 3820 -31370 4020 -31360
rect 4220 -32420 4280 -30950
rect 4330 -30990 4390 -30980
rect 4330 -31060 4390 -31050
rect 4440 -32420 4500 -30950
rect 4700 -31230 4900 -31150
rect 5360 -31230 5560 -31150
rect 6020 -31230 6220 -31150
rect 4700 -31300 4900 -31290
rect 4700 -31360 4710 -31300
rect 4890 -31360 4900 -31300
rect 4700 -31370 4900 -31360
rect 5360 -31300 5560 -31290
rect 5360 -31360 5370 -31300
rect 5550 -31360 5560 -31300
rect 5360 -31370 5560 -31360
rect 6020 -31300 6220 -31290
rect 6020 -31360 6030 -31300
rect 6210 -31360 6220 -31300
rect 6020 -31370 6220 -31360
rect 6420 -32420 6480 -30950
rect 6530 -30990 6590 -30980
rect 6530 -31060 6590 -31050
rect 6640 -32420 6700 -30950
rect 6900 -31160 7100 -31150
rect 6900 -31220 6910 -31160
rect 7090 -31220 7100 -31160
rect 6900 -31230 7100 -31220
rect 7560 -31160 7760 -31150
rect 7560 -31220 7570 -31160
rect 7750 -31220 7760 -31160
rect 7560 -31230 7760 -31220
rect 8220 -31160 8420 -31150
rect 8220 -31220 8230 -31160
rect 8410 -31220 8420 -31160
rect 8220 -31230 8420 -31220
rect 6900 -31370 7100 -31290
rect 7560 -31370 7760 -31290
rect 8220 -31370 8420 -31290
rect 8620 -32420 8680 -30950
rect 8730 -30990 8790 -30980
rect 8730 -31060 8790 -31050
rect 8840 -32420 8900 -30950
rect 9100 -31160 9300 -31150
rect 9100 -31220 9110 -31160
rect 9290 -31220 9300 -31160
rect 9100 -31230 9300 -31220
rect 9760 -31160 9960 -31150
rect 9760 -31220 9770 -31160
rect 9950 -31220 9960 -31160
rect 9760 -31230 9960 -31220
rect 10420 -31160 10620 -31150
rect 10420 -31220 10430 -31160
rect 10610 -31220 10620 -31160
rect 10420 -31230 10620 -31220
rect 9100 -31370 9300 -31290
rect 9760 -31370 9960 -31290
rect 10420 -31370 10620 -31290
rect 10820 -32420 10880 -30950
rect 10930 -30990 10990 -30980
rect 10930 -31060 10990 -31050
rect 11040 -32420 11100 -30950
rect 11300 -31160 11500 -31150
rect 11300 -31220 11310 -31160
rect 11490 -31220 11500 -31160
rect 11300 -31230 11500 -31220
rect 11960 -31160 12160 -31150
rect 11960 -31220 11970 -31160
rect 12150 -31220 12160 -31160
rect 11960 -31230 12160 -31220
rect 12620 -31160 12820 -31150
rect 12620 -31220 12630 -31160
rect 12810 -31220 12820 -31160
rect 12620 -31230 12820 -31220
rect 11300 -31370 11500 -31290
rect 11960 -31370 12160 -31290
rect 12620 -31370 12820 -31290
rect 13020 -32420 13080 -30950
rect 13130 -30990 13190 -30980
rect 13130 -31060 13190 -31050
rect 13240 -32420 13300 -30950
rect 13500 -31160 13700 -31150
rect 13500 -31220 13510 -31160
rect 13690 -31220 13700 -31160
rect 13500 -31230 13700 -31220
rect 14160 -31160 14360 -31150
rect 14160 -31220 14170 -31160
rect 14350 -31220 14360 -31160
rect 14160 -31230 14360 -31220
rect 14820 -31160 15020 -31150
rect 14820 -31220 14830 -31160
rect 15010 -31220 15020 -31160
rect 14820 -31230 15020 -31220
rect 13500 -31370 13700 -31290
rect 14160 -31370 14360 -31290
rect 14820 -31370 15020 -31290
rect 15220 -32420 15280 -30950
rect 15330 -30990 15390 -30980
rect 15330 -31060 15390 -31050
rect 15440 -32420 15500 -30950
rect 15700 -31230 15900 -31150
rect 16360 -31230 16560 -31150
rect 17020 -31230 17220 -31150
rect 15700 -31300 15900 -31290
rect 15700 -31360 15710 -31300
rect 15890 -31360 15900 -31300
rect 15700 -31370 15900 -31360
rect 16360 -31300 16560 -31290
rect 16360 -31360 16370 -31300
rect 16550 -31360 16560 -31300
rect 16360 -31370 16560 -31360
rect 17020 -31300 17220 -31290
rect 17020 -31360 17030 -31300
rect 17210 -31360 17220 -31300
rect 17020 -31370 17220 -31360
rect 17420 -32420 17480 -30950
rect 17530 -30990 17590 -30980
rect 17530 -31060 17590 -31050
rect 17640 -32420 17700 -30950
rect 17900 -31230 18100 -31150
rect 18560 -31230 18760 -31150
rect 19220 -31230 19420 -31150
rect 17900 -31300 18100 -31290
rect 17900 -31360 17910 -31300
rect 18090 -31360 18100 -31300
rect 17900 -31370 18100 -31360
rect 18560 -31300 18760 -31290
rect 18560 -31360 18570 -31300
rect 18750 -31360 18760 -31300
rect 18560 -31370 18760 -31360
rect 19220 -31300 19420 -31290
rect 19220 -31360 19230 -31300
rect 19410 -31360 19420 -31300
rect 19220 -31370 19420 -31360
rect 19620 -32420 19680 -30950
rect 19730 -30990 19790 -30980
rect 19730 -31060 19790 -31050
rect 19840 -32420 19900 -30950
rect 21930 -30990 21990 -30980
rect 21930 -31060 21990 -31050
<< via2 >>
rect 2210 11890 2330 12010
rect 1990 11590 2110 11710
rect -70 10870 -10 10930
rect 2130 10870 2190 10930
rect 4410 11890 4530 12010
rect 4190 11590 4310 11710
rect 2510 11180 2690 11240
rect 3170 11180 3350 11240
rect 3830 11180 4010 11240
rect 4330 10870 4390 10930
rect 6610 11890 6730 12010
rect 6390 11590 6510 11710
rect 4710 11180 4890 11240
rect 5370 11180 5550 11240
rect 6030 11180 6210 11240
rect 6530 10870 6590 10930
rect 8810 11890 8930 12010
rect 8590 11590 8710 11710
rect 6910 11040 7090 11100
rect 7570 11040 7750 11100
rect 8230 11040 8410 11100
rect 8730 10870 8790 10930
rect 11010 11890 11130 12010
rect 10790 11590 10910 11710
rect 9110 11040 9290 11100
rect 9770 11040 9950 11100
rect 10430 11040 10610 11100
rect 10930 10870 10990 10930
rect 13210 11890 13330 12010
rect 12990 11590 13110 11710
rect 11310 11040 11490 11100
rect 11970 11040 12150 11100
rect 12630 11040 12810 11100
rect 13130 10870 13190 10930
rect 15410 11890 15530 12010
rect 15190 11590 15310 11710
rect 13510 11040 13690 11100
rect 14170 11040 14350 11100
rect 14830 11040 15010 11100
rect 15330 10870 15390 10930
rect 17610 11890 17730 12010
rect 17390 11590 17510 11710
rect 15710 11180 15890 11240
rect 16370 11180 16550 11240
rect 17030 11180 17210 11240
rect 17530 10870 17590 10930
rect 19810 11890 19930 12010
rect 19590 11590 19710 11710
rect 17910 11180 18090 11240
rect 18570 11180 18750 11240
rect 19230 11180 19410 11240
rect 19730 10870 19790 10930
rect 21930 10870 21990 10930
rect -70 10070 -10 10130
rect 2130 10070 2190 10130
rect 2510 10550 4010 10610
rect 2510 10240 2690 10300
rect 3170 10240 3350 10300
rect 3830 10240 4010 10300
rect 4330 10070 4390 10130
rect 4710 10550 6210 10610
rect 4710 10240 4890 10300
rect 5370 10240 5550 10300
rect 6030 10240 6210 10300
rect 6530 10070 6590 10130
rect 6910 10550 8410 10610
rect 6910 10380 7090 10440
rect 7570 10380 7750 10440
rect 8230 10380 8410 10440
rect 8730 10070 8790 10130
rect 9110 10550 10610 10610
rect 9110 10380 9290 10440
rect 9770 10380 9950 10440
rect 10430 10380 10610 10440
rect 10930 10070 10990 10130
rect 11310 10550 12810 10610
rect 11310 10380 11490 10440
rect 11970 10380 12150 10440
rect 12630 10380 12810 10440
rect 13130 10070 13190 10130
rect 13510 10550 15010 10610
rect 13510 10380 13690 10440
rect 14170 10380 14350 10440
rect 14830 10380 15010 10440
rect 15330 10070 15390 10130
rect 15710 10550 17210 10610
rect 15710 10240 15890 10300
rect 16370 10240 16550 10300
rect 17030 10240 17210 10300
rect 17530 10070 17590 10130
rect 17910 10550 19410 10610
rect 17910 10240 18090 10300
rect 18570 10240 18750 10300
rect 19230 10240 19410 10300
rect 19730 10070 19790 10130
rect 21930 10070 21990 10130
rect -70 9270 -10 9330
rect 2130 9270 2190 9330
rect 2510 9750 4010 9810
rect 2510 9580 2690 9640
rect 3170 9580 3350 9640
rect 3830 9580 4010 9640
rect 4330 9270 4390 9330
rect 4710 9750 6210 9810
rect 4710 9580 4890 9640
rect 5370 9580 5550 9640
rect 6030 9580 6210 9640
rect 6530 9270 6590 9330
rect 6910 9750 8410 9810
rect 6910 9440 7090 9500
rect 7570 9440 7750 9500
rect 8230 9440 8410 9500
rect 8730 9270 8790 9330
rect 9110 9750 10610 9810
rect 9110 9440 9290 9500
rect 9770 9440 9950 9500
rect 10430 9440 10610 9500
rect 10930 9270 10990 9330
rect 11310 9750 12810 9810
rect 11310 9440 11490 9500
rect 11970 9440 12150 9500
rect 12630 9440 12810 9500
rect 13130 9270 13190 9330
rect 13510 9750 15010 9810
rect 13510 9440 13690 9500
rect 14170 9440 14350 9500
rect 14830 9440 15010 9500
rect 15330 9270 15390 9330
rect 15710 9750 17210 9810
rect 15710 9580 15890 9640
rect 16370 9580 16550 9640
rect 17030 9580 17210 9640
rect 17530 9270 17590 9330
rect 17910 9750 19410 9810
rect 17910 9580 18090 9640
rect 18570 9580 18750 9640
rect 19230 9580 19410 9640
rect 19730 9270 19790 9330
rect 21930 9270 21990 9330
rect 430 8910 610 8990
rect -70 8470 -10 8530
rect 2130 8470 2190 8530
rect 2510 8640 2690 8700
rect 3170 8640 3350 8700
rect 3830 8640 4010 8700
rect 4330 8470 4390 8530
rect 4710 8950 6210 9010
rect 4710 8640 4890 8700
rect 5370 8640 5550 8700
rect 6030 8640 6210 8700
rect 6530 8470 6590 8530
rect 6910 8950 8410 9010
rect 6910 8780 7090 8840
rect 7570 8780 7750 8840
rect 8230 8780 8410 8840
rect 8730 8470 8790 8530
rect 9110 8950 10610 9010
rect 9110 8780 9290 8840
rect 9770 8780 9950 8840
rect 10430 8780 10610 8840
rect 10930 8470 10990 8530
rect 11310 8950 12810 9010
rect 11310 8780 11490 8840
rect 11970 8780 12150 8840
rect 12630 8780 12810 8840
rect 13130 8470 13190 8530
rect 13510 8950 15010 9010
rect 13510 8780 13690 8840
rect 14170 8780 14350 8840
rect 14830 8780 15010 8840
rect 15330 8470 15390 8530
rect 15710 8950 17210 9010
rect 15710 8640 15890 8700
rect 16370 8640 16550 8700
rect 17030 8640 17210 8700
rect 17530 8470 17590 8530
rect 17910 8640 18090 8700
rect 18570 8640 18750 8700
rect 19230 8640 19410 8700
rect 19730 8470 19790 8530
rect 21310 8910 21490 8990
rect 21930 8470 21990 8530
rect 430 8110 610 8190
rect -70 7670 -10 7730
rect 2130 7670 2190 7730
rect 2510 7840 2690 7900
rect 3170 7840 3350 7900
rect 3830 7840 4010 7900
rect 4330 7670 4390 7730
rect 4710 8150 6210 8210
rect 4710 7840 4890 7900
rect 5370 7840 5550 7900
rect 6030 7840 6210 7900
rect 6530 7670 6590 7730
rect 6910 8150 8410 8210
rect 6910 7980 7090 8040
rect 7570 7980 7750 8040
rect 8230 7980 8410 8040
rect 8730 7670 8790 7730
rect 9110 8150 10610 8210
rect 9110 7980 9290 8040
rect 9770 7980 9950 8040
rect 10430 7980 10610 8040
rect 10930 7670 10990 7730
rect 11310 8150 12810 8210
rect 11310 7980 11490 8040
rect 11970 7980 12150 8040
rect 12630 7980 12810 8040
rect 13130 7670 13190 7730
rect 13510 8150 15010 8210
rect 13510 7980 13690 8040
rect 14170 7980 14350 8040
rect 14830 7980 15010 8040
rect 15330 7670 15390 7730
rect 15710 8150 17210 8210
rect 15710 7840 15890 7900
rect 16370 7840 16550 7900
rect 17030 7840 17210 7900
rect 17530 7670 17590 7730
rect 17910 7840 18090 7900
rect 18570 7840 18750 7900
rect 19230 7840 19410 7900
rect 19730 7670 19790 7730
rect 21310 8110 21490 8190
rect 21930 7670 21990 7730
rect 430 7310 610 7390
rect -70 6870 -10 6930
rect 2130 6870 2190 6930
rect 2510 7180 2690 7240
rect 3170 7180 3350 7240
rect 3830 7180 4010 7240
rect 4330 6870 4390 6930
rect 4710 7350 6210 7410
rect 4710 7180 4890 7240
rect 5370 7180 5550 7240
rect 6030 7180 6210 7240
rect 6530 6870 6590 6930
rect 6910 7350 8410 7410
rect 6910 7040 7090 7100
rect 7570 7040 7750 7100
rect 8230 7040 8410 7100
rect 8730 6870 8790 6930
rect 9110 7350 10610 7410
rect 9110 7040 9290 7100
rect 9770 7040 9950 7100
rect 10430 7040 10610 7100
rect 10930 6870 10990 6930
rect 11310 7350 12810 7410
rect 11310 7040 11490 7100
rect 11970 7040 12150 7100
rect 12630 7040 12810 7100
rect 13130 6870 13190 6930
rect 13510 7350 15010 7410
rect 13510 7040 13690 7100
rect 14170 7040 14350 7100
rect 14830 7040 15010 7100
rect 15330 6870 15390 6930
rect 15710 7350 17210 7410
rect 15710 7180 15890 7240
rect 16370 7180 16550 7240
rect 17030 7180 17210 7240
rect 17530 6870 17590 6930
rect 17910 7180 18090 7240
rect 18570 7180 18750 7240
rect 19230 7180 19410 7240
rect 19730 6870 19790 6930
rect 21310 7310 21490 7390
rect 21930 6870 21990 6930
rect 430 6510 610 6590
rect -70 6070 -10 6130
rect 2130 6070 2190 6130
rect 2510 6240 2690 6300
rect 3170 6240 3350 6300
rect 3830 6240 4010 6300
rect 4330 6070 4390 6130
rect 4710 6550 6210 6610
rect 4710 6240 4890 6300
rect 5370 6240 5550 6300
rect 6030 6240 6210 6300
rect 6530 6070 6590 6130
rect 6910 6550 8410 6610
rect 6910 6380 7090 6440
rect 7570 6380 7750 6440
rect 8230 6380 8410 6440
rect 8730 6070 8790 6130
rect 9110 6550 10610 6610
rect 9110 6380 9290 6440
rect 9770 6380 9950 6440
rect 10430 6380 10610 6440
rect 10930 6070 10990 6130
rect 11310 6550 12810 6610
rect 11310 6380 11490 6440
rect 11970 6380 12150 6440
rect 12630 6380 12810 6440
rect 13130 6070 13190 6130
rect 13510 6550 15010 6610
rect 13510 6380 13690 6440
rect 14170 6380 14350 6440
rect 14830 6380 15010 6440
rect 15330 6070 15390 6130
rect 15710 6550 17210 6610
rect 15710 6240 15890 6300
rect 16370 6240 16550 6300
rect 17030 6240 17210 6300
rect 17530 6070 17590 6130
rect 17910 6240 18090 6300
rect 18570 6240 18750 6300
rect 19230 6240 19410 6300
rect 19730 6070 19790 6130
rect 21310 6510 21490 6590
rect 21930 6070 21990 6130
rect -70 5270 -10 5330
rect 2130 5270 2190 5330
rect 2510 5750 4010 5810
rect 2510 5580 2690 5640
rect 3170 5580 3350 5640
rect 3830 5580 4010 5640
rect 4330 5270 4390 5330
rect 4710 5750 6210 5810
rect 4710 5580 4890 5640
rect 5370 5580 5550 5640
rect 6030 5580 6210 5640
rect 6530 5270 6590 5330
rect 6910 5750 8410 5810
rect 6910 5440 7090 5500
rect 7570 5440 7750 5500
rect 8230 5440 8410 5500
rect 8730 5270 8790 5330
rect 9110 5750 10610 5810
rect 9110 5440 9290 5500
rect 9770 5440 9950 5500
rect 10430 5440 10610 5500
rect 10930 5270 10990 5330
rect 11310 5750 12810 5810
rect 11310 5440 11490 5500
rect 11970 5440 12150 5500
rect 12630 5440 12810 5500
rect 13130 5270 13190 5330
rect 13510 5750 15010 5810
rect 13510 5440 13690 5500
rect 14170 5440 14350 5500
rect 14830 5440 15010 5500
rect 15330 5270 15390 5330
rect 15710 5750 17210 5810
rect 15710 5580 15890 5640
rect 16370 5580 16550 5640
rect 17030 5580 17210 5640
rect 17530 5270 17590 5330
rect 17910 5750 19410 5810
rect 17910 5580 18090 5640
rect 18570 5580 18750 5640
rect 19230 5580 19410 5640
rect 19730 5270 19790 5330
rect 21930 5270 21990 5330
rect 2510 4950 4010 5010
rect 4710 4950 6210 5010
rect 6910 4950 8410 5010
rect 9110 4950 10610 5010
rect 11310 4950 12810 5010
rect 13510 4950 15010 5010
rect 15710 4950 17210 5010
rect 17910 4950 19410 5010
rect 31570 3550 31730 3730
rect 1170 3150 1330 3330
rect 2770 3150 2930 3330
rect 4370 3150 4530 3330
rect 5970 3150 6130 3330
rect 7570 3150 7730 3330
rect 9170 3150 9330 3330
rect 2110 2070 2230 2230
rect 3710 2070 3830 2230
rect 2110 270 2230 430
rect 5310 2070 5430 2230
rect 3710 270 3830 430
rect 2110 -1530 2230 -1370
rect 6910 2070 7030 2230
rect 5310 270 5430 430
rect 3710 -1530 3830 -1370
rect 2110 -3330 2230 -3170
rect 8510 2070 8630 2230
rect 6910 270 7030 430
rect 5310 -1530 5430 -1370
rect 3710 -3330 3830 -3170
rect 11700 2600 11840 2750
rect 11000 2380 11140 2520
rect 10110 2070 10230 2230
rect 12600 2380 12740 2520
rect 13980 2380 14120 2520
rect 11710 2070 11830 2230
rect 8510 270 8630 430
rect 6910 -1530 7030 -1370
rect 5310 -3330 5430 -3170
rect 13310 2070 13430 2230
rect 10110 270 10230 430
rect 8510 -1530 8630 -1370
rect 6910 -3330 7030 -3170
rect 11710 270 11830 430
rect 10110 -1530 10230 -1370
rect 8510 -3330 8630 -3170
rect 10110 -3330 10230 -3170
rect 13310 270 13430 430
rect 11710 -1530 11830 -1370
rect 13310 -1530 13430 -1370
rect 11710 -3330 11830 -3170
rect 16510 2070 16630 2230
rect 14910 1300 15030 1960
rect 18110 2070 18230 2230
rect 19710 2070 19830 2230
rect 21310 2070 21430 2230
rect 22910 2070 23030 2230
rect 24510 2070 24630 2230
rect 26110 2070 26230 2230
rect 27710 2050 27830 2230
rect 29310 2050 29430 2230
rect 14910 -1530 15030 -1370
rect 15250 -1530 15370 -1370
rect 13310 -3330 13430 -3170
rect 16510 270 16630 430
rect 2130 -9750 2230 -9590
rect 2130 -11550 2230 -11390
rect 3730 -9750 3830 -9590
rect 2130 -13350 2230 -13190
rect 3730 -11550 3830 -11390
rect 2130 -15150 2230 -14990
rect 5330 -9750 5430 -9590
rect 3730 -13350 3830 -13190
rect 2130 -16950 2230 -16790
rect 5330 -11550 5430 -11390
rect 3730 -15150 3830 -14990
rect 2130 -18750 2230 -18590
rect 6930 -9750 7030 -9590
rect 5330 -13350 5430 -13190
rect 3730 -16950 3830 -16790
rect 2130 -20550 2230 -20390
rect 6930 -11550 7030 -11390
rect 5330 -15150 5430 -14990
rect 3730 -18750 3830 -18590
rect 2130 -22350 2230 -22190
rect 8530 -9750 8630 -9590
rect 6930 -13350 7030 -13190
rect 5330 -16950 5430 -16790
rect 3730 -20550 3830 -20390
rect 8530 -11550 8630 -11390
rect 6930 -15150 7030 -14990
rect 5330 -18750 5430 -18590
rect 3730 -22350 3830 -22190
rect 10130 -9750 10230 -9590
rect 8530 -13350 8630 -13190
rect 6930 -16950 7030 -16790
rect 5330 -20550 5430 -20390
rect 10130 -11550 10230 -11390
rect 8530 -15150 8630 -14990
rect 6930 -18750 7030 -18590
rect 5330 -22350 5430 -22190
rect 10130 -13350 10230 -13190
rect 8530 -16950 8630 -16790
rect 6930 -20550 7030 -20390
rect 10130 -15150 10230 -14990
rect 8530 -18750 8630 -18590
rect 6930 -22350 7030 -22190
rect 10130 -16950 10230 -16790
rect 8530 -20550 8630 -20390
rect 10130 -18750 10230 -18590
rect 8530 -22350 8630 -22190
rect 14910 -3330 15030 -3170
rect 16510 -1530 16630 -1370
rect 13290 -13330 13460 -13170
rect 18110 270 18230 430
rect 16510 -3330 16630 -3170
rect 15570 -5350 15730 -5170
rect 15570 -5750 15730 -5570
rect 14910 -6610 15030 -6490
rect 15790 -6150 15950 -5970
rect 18110 -1530 18230 -1370
rect 19710 270 19830 430
rect 18110 -3330 18230 -3170
rect 19710 -1530 19830 -1370
rect 21310 270 21430 430
rect 19710 -3330 19830 -3170
rect 21310 -1530 21430 -1370
rect 18770 -5350 18930 -5170
rect 18770 -5750 18930 -5570
rect 17390 -6950 17550 -6770
rect 17170 -7350 17330 -7170
rect 17170 -7750 17330 -7570
rect 16510 -9730 16640 -9570
rect 13290 -15130 13460 -14970
rect 13300 -16950 13450 -16790
rect 13300 -18750 13450 -18590
rect 18990 -6150 19150 -5970
rect 22910 270 23030 430
rect 21310 -3330 21430 -3170
rect 22910 -1530 23030 -1370
rect 24510 270 24630 430
rect 22910 -3330 23030 -3170
rect 24510 -1530 24630 -1370
rect 21970 -5350 22130 -5170
rect 21970 -5750 22130 -5570
rect 20590 -6950 20750 -6770
rect 20370 -7350 20530 -7170
rect 20370 -7750 20530 -7570
rect 18110 -9730 18240 -9570
rect 16510 -11530 16640 -11370
rect 14890 -13330 15060 -13170
rect 19710 -9730 19840 -9570
rect 18110 -11530 18240 -11370
rect 16510 -13330 16640 -13170
rect 14890 -15130 15060 -14970
rect 22190 -6150 22350 -5970
rect 24510 -3330 24630 -3170
rect 26110 270 26230 430
rect 26110 -1530 26230 -1370
rect 27710 250 27830 430
rect 26110 -3330 26230 -3170
rect 27710 -1550 27830 -1370
rect 25170 -5350 25330 -5170
rect 25170 -5750 25330 -5570
rect 23790 -6950 23950 -6770
rect 23570 -7350 23730 -7170
rect 23570 -7750 23730 -7570
rect 21310 -9730 21440 -9570
rect 19710 -11530 19840 -11370
rect 18110 -13330 18240 -13170
rect 16510 -15130 16640 -14970
rect 14900 -16950 15050 -16790
rect 22910 -9730 23040 -9570
rect 21310 -11530 21440 -11370
rect 19710 -13330 19840 -13170
rect 18110 -15130 18240 -14970
rect 16510 -16930 16640 -16770
rect 14900 -18750 15050 -18590
rect 25390 -6150 25550 -5970
rect 29310 250 29430 430
rect 27710 -3350 27830 -3170
rect 29310 -1550 29430 -1370
rect 30910 2050 31030 2230
rect 30910 250 31030 430
rect 34900 2600 35050 2760
rect 33300 2370 33450 2530
rect 32510 1010 32630 1130
rect 34110 1010 34230 1130
rect 34910 1010 35040 1130
rect 35710 1010 35830 1130
rect 33300 260 33450 420
rect 32510 -510 32630 170
rect 34110 -510 34230 170
rect 30910 -1550 31030 -1370
rect 29310 -3350 29430 -3170
rect 28370 -5350 28530 -5170
rect 28370 -5750 28530 -5570
rect 27690 -6150 27850 -5970
rect 26990 -6950 27150 -6770
rect 26770 -7350 26930 -7170
rect 26770 -7750 26930 -7570
rect 24510 -9730 24640 -9570
rect 22910 -11530 23040 -11370
rect 21310 -13330 21440 -13170
rect 19710 -15130 19840 -14970
rect 18110 -16930 18240 -16770
rect 16510 -18730 16640 -18570
rect 10130 -20550 10230 -20390
rect 26110 -9730 26240 -9570
rect 24510 -11530 24640 -11370
rect 22910 -13330 23040 -13170
rect 21310 -15130 21440 -14970
rect 19710 -16930 19840 -16770
rect 18110 -18730 18240 -18570
rect 16510 -20530 16640 -20370
rect 28590 -6150 28750 -5970
rect 29290 -6150 29450 -5970
rect 30910 -3350 31030 -3170
rect 32510 -2590 32630 -2470
rect 35710 -510 35830 170
rect 34110 -2590 34230 -2470
rect 34910 -2590 35040 -2470
rect 35710 -2590 35830 -2470
rect 30890 -6150 31050 -5970
rect 30190 -6950 30350 -6770
rect 29970 -7350 30130 -7170
rect 29970 -7750 30130 -7570
rect 27710 -9730 27840 -9570
rect 26110 -11530 26240 -11370
rect 24510 -13330 24640 -13170
rect 22910 -15130 23040 -14970
rect 21310 -16930 21440 -16770
rect 19710 -18730 19840 -18570
rect 18110 -20530 18240 -20370
rect 29310 -9730 29440 -9570
rect 27710 -11530 27840 -11370
rect 26110 -13330 26240 -13170
rect 24510 -15130 24640 -14970
rect 22910 -16930 23040 -16770
rect 21310 -18730 21440 -18570
rect 19710 -20530 19840 -20370
rect 30910 -9730 31040 -9570
rect 29310 -11530 29440 -11370
rect 27710 -13330 27840 -13170
rect 26110 -15130 26240 -14970
rect 30910 -11530 31040 -11370
rect 29310 -13330 29440 -13170
rect 27710 -15130 27840 -14970
rect 24510 -16930 24640 -16770
rect 26110 -16930 26240 -16770
rect 22910 -18730 23040 -18570
rect 21310 -20530 21440 -20370
rect 30910 -13330 31040 -13170
rect 29310 -15130 29440 -14970
rect 27710 -16930 27840 -16770
rect 24510 -18730 24640 -18570
rect 26110 -18730 26240 -18570
rect 22910 -20530 23040 -20370
rect 29310 -16930 29440 -16770
rect 27710 -18730 27840 -18570
rect 24510 -20530 24640 -20370
rect 26110 -20530 26240 -20370
rect 29310 -18730 29440 -18570
rect 27710 -20530 27840 -20370
rect 29310 -20530 29440 -20370
rect 30910 -15130 31040 -14970
rect 30910 -16930 31040 -16770
rect 30910 -18730 31040 -18570
rect 30910 -20530 31040 -20370
rect 10130 -22350 10230 -22190
rect 16510 -22330 16640 -22170
rect 18110 -22330 18240 -22170
rect 19710 -22330 19840 -22170
rect 21310 -22330 21440 -22170
rect 22910 -22330 23040 -22170
rect 24510 -22330 24640 -22170
rect 26110 -22330 26240 -22170
rect 27710 -22330 27840 -22170
rect 29310 -22330 29440 -22170
rect 30910 -22330 31040 -22170
rect 11050 -22850 11150 -22740
rect 27720 -22850 27830 -22740
rect 29320 -22850 29430 -22740
rect 30920 -22850 31030 -22740
rect 2790 -23450 2950 -23270
rect 4390 -23450 4550 -23270
rect 5990 -23450 6150 -23270
rect 7590 -23450 7750 -23270
rect 9190 -23450 9350 -23270
rect 2510 -25130 4010 -25070
rect 4710 -25130 6210 -25070
rect 6910 -25130 8410 -25070
rect 9110 -25130 10610 -25070
rect 11310 -25130 12810 -25070
rect 13510 -25130 15010 -25070
rect 15710 -25130 17210 -25070
rect 17910 -25130 19410 -25070
rect -70 -25450 -10 -25390
rect 2130 -25450 2190 -25390
rect 2510 -25760 2690 -25700
rect 3170 -25760 3350 -25700
rect 3830 -25760 4010 -25700
rect 2510 -25930 4010 -25870
rect 4330 -25450 4390 -25390
rect 4710 -25760 4890 -25700
rect 5370 -25760 5550 -25700
rect 6030 -25760 6210 -25700
rect 4710 -25930 6210 -25870
rect 6530 -25450 6590 -25390
rect 6910 -25620 7090 -25560
rect 7570 -25620 7750 -25560
rect 8230 -25620 8410 -25560
rect 6910 -25930 8410 -25870
rect 8730 -25450 8790 -25390
rect 9110 -25620 9290 -25560
rect 9770 -25620 9950 -25560
rect 10430 -25620 10610 -25560
rect 9110 -25930 10610 -25870
rect 10930 -25450 10990 -25390
rect 11310 -25620 11490 -25560
rect 11970 -25620 12150 -25560
rect 12630 -25620 12810 -25560
rect 11310 -25930 12810 -25870
rect 13130 -25450 13190 -25390
rect 13510 -25620 13690 -25560
rect 14170 -25620 14350 -25560
rect 14830 -25620 15010 -25560
rect 13510 -25930 15010 -25870
rect 15330 -25450 15390 -25390
rect 15710 -25760 15890 -25700
rect 16370 -25760 16550 -25700
rect 17030 -25760 17210 -25700
rect 15710 -25930 17210 -25870
rect 17530 -25450 17590 -25390
rect 17910 -25760 18090 -25700
rect 18570 -25760 18750 -25700
rect 19230 -25760 19410 -25700
rect 17910 -25930 19410 -25870
rect 19730 -25450 19790 -25390
rect 21930 -25450 21990 -25390
rect -70 -26250 -10 -26190
rect 430 -26710 610 -26630
rect 2130 -26250 2190 -26190
rect 2510 -26420 2690 -26360
rect 3170 -26420 3350 -26360
rect 3830 -26420 4010 -26360
rect 4330 -26250 4390 -26190
rect 4710 -26420 4890 -26360
rect 5370 -26420 5550 -26360
rect 6030 -26420 6210 -26360
rect 4710 -26730 6210 -26670
rect 6530 -26250 6590 -26190
rect 6910 -26560 7090 -26500
rect 7570 -26560 7750 -26500
rect 8230 -26560 8410 -26500
rect 6910 -26730 8410 -26670
rect 8730 -26250 8790 -26190
rect 9110 -26560 9290 -26500
rect 9770 -26560 9950 -26500
rect 10430 -26560 10610 -26500
rect 9110 -26730 10610 -26670
rect 10930 -26250 10990 -26190
rect 11310 -26560 11490 -26500
rect 11970 -26560 12150 -26500
rect 12630 -26560 12810 -26500
rect 11310 -26730 12810 -26670
rect 13130 -26250 13190 -26190
rect 13510 -26560 13690 -26500
rect 14170 -26560 14350 -26500
rect 14830 -26560 15010 -26500
rect 13510 -26730 15010 -26670
rect 15330 -26250 15390 -26190
rect 15710 -26420 15890 -26360
rect 16370 -26420 16550 -26360
rect 17030 -26420 17210 -26360
rect 15710 -26730 17210 -26670
rect 17530 -26250 17590 -26190
rect 17910 -26420 18090 -26360
rect 18570 -26420 18750 -26360
rect 19230 -26420 19410 -26360
rect 19730 -26250 19790 -26190
rect 21930 -26250 21990 -26190
rect 21310 -26710 21490 -26630
rect -70 -27050 -10 -26990
rect 430 -27510 610 -27430
rect 2130 -27050 2190 -26990
rect 2510 -27360 2690 -27300
rect 3170 -27360 3350 -27300
rect 3830 -27360 4010 -27300
rect 4330 -27050 4390 -26990
rect 4710 -27360 4890 -27300
rect 5370 -27360 5550 -27300
rect 6030 -27360 6210 -27300
rect 4710 -27530 6210 -27470
rect 6530 -27050 6590 -26990
rect 6910 -27220 7090 -27160
rect 7570 -27220 7750 -27160
rect 8230 -27220 8410 -27160
rect 6910 -27530 8410 -27470
rect 8730 -27050 8790 -26990
rect 9110 -27220 9290 -27160
rect 9770 -27220 9950 -27160
rect 10430 -27220 10610 -27160
rect 9110 -27530 10610 -27470
rect 10930 -27050 10990 -26990
rect 11310 -27220 11490 -27160
rect 11970 -27220 12150 -27160
rect 12630 -27220 12810 -27160
rect 11310 -27530 12810 -27470
rect 13130 -27050 13190 -26990
rect 13510 -27220 13690 -27160
rect 14170 -27220 14350 -27160
rect 14830 -27220 15010 -27160
rect 13510 -27530 15010 -27470
rect 15330 -27050 15390 -26990
rect 15710 -27360 15890 -27300
rect 16370 -27360 16550 -27300
rect 17030 -27360 17210 -27300
rect 15710 -27530 17210 -27470
rect 17530 -27050 17590 -26990
rect 17910 -27360 18090 -27300
rect 18570 -27360 18750 -27300
rect 19230 -27360 19410 -27300
rect 19730 -27050 19790 -26990
rect 21930 -27050 21990 -26990
rect 21310 -27510 21490 -27430
rect -70 -27850 -10 -27790
rect 430 -28310 610 -28230
rect 2130 -27850 2190 -27790
rect 2510 -28020 2690 -27960
rect 3170 -28020 3350 -27960
rect 3830 -28020 4010 -27960
rect 4330 -27850 4390 -27790
rect 4710 -28020 4890 -27960
rect 5370 -28020 5550 -27960
rect 6030 -28020 6210 -27960
rect 4710 -28330 6210 -28270
rect 6530 -27850 6590 -27790
rect 6910 -28160 7090 -28100
rect 7570 -28160 7750 -28100
rect 8230 -28160 8410 -28100
rect 6910 -28330 8410 -28270
rect 8730 -27850 8790 -27790
rect 9110 -28160 9290 -28100
rect 9770 -28160 9950 -28100
rect 10430 -28160 10610 -28100
rect 9110 -28330 10610 -28270
rect 10930 -27850 10990 -27790
rect 11310 -28160 11490 -28100
rect 11970 -28160 12150 -28100
rect 12630 -28160 12810 -28100
rect 11310 -28330 12810 -28270
rect 13130 -27850 13190 -27790
rect 13510 -28160 13690 -28100
rect 14170 -28160 14350 -28100
rect 14830 -28160 15010 -28100
rect 13510 -28330 15010 -28270
rect 15330 -27850 15390 -27790
rect 15710 -28020 15890 -27960
rect 16370 -28020 16550 -27960
rect 17030 -28020 17210 -27960
rect 15710 -28330 17210 -28270
rect 17530 -27850 17590 -27790
rect 17910 -28020 18090 -27960
rect 18570 -28020 18750 -27960
rect 19230 -28020 19410 -27960
rect 19730 -27850 19790 -27790
rect 21930 -27850 21990 -27790
rect 21310 -28310 21490 -28230
rect -70 -28650 -10 -28590
rect 430 -29110 610 -29030
rect 2130 -28650 2190 -28590
rect 2510 -28820 2690 -28760
rect 3170 -28820 3350 -28760
rect 3830 -28820 4010 -28760
rect 4330 -28650 4390 -28590
rect 4710 -28820 4890 -28760
rect 5370 -28820 5550 -28760
rect 6030 -28820 6210 -28760
rect 4710 -29130 6210 -29070
rect 6530 -28650 6590 -28590
rect 6910 -28960 7090 -28900
rect 7570 -28960 7750 -28900
rect 8230 -28960 8410 -28900
rect 6910 -29130 8410 -29070
rect 8730 -28650 8790 -28590
rect 9110 -28960 9290 -28900
rect 9770 -28960 9950 -28900
rect 10430 -28960 10610 -28900
rect 9110 -29130 10610 -29070
rect 10930 -28650 10990 -28590
rect 11310 -28960 11490 -28900
rect 11970 -28960 12150 -28900
rect 12630 -28960 12810 -28900
rect 11310 -29130 12810 -29070
rect 13130 -28650 13190 -28590
rect 13510 -28960 13690 -28900
rect 14170 -28960 14350 -28900
rect 14830 -28960 15010 -28900
rect 13510 -29130 15010 -29070
rect 15330 -28650 15390 -28590
rect 15710 -28820 15890 -28760
rect 16370 -28820 16550 -28760
rect 17030 -28820 17210 -28760
rect 15710 -29130 17210 -29070
rect 17530 -28650 17590 -28590
rect 17910 -28820 18090 -28760
rect 18570 -28820 18750 -28760
rect 19230 -28820 19410 -28760
rect 19730 -28650 19790 -28590
rect 21930 -28650 21990 -28590
rect 21310 -29110 21490 -29030
rect -70 -29450 -10 -29390
rect 2130 -29450 2190 -29390
rect 2510 -29760 2690 -29700
rect 3170 -29760 3350 -29700
rect 3830 -29760 4010 -29700
rect 2510 -29930 4010 -29870
rect 4330 -29450 4390 -29390
rect 4710 -29760 4890 -29700
rect 5370 -29760 5550 -29700
rect 6030 -29760 6210 -29700
rect 4710 -29930 6210 -29870
rect 6530 -29450 6590 -29390
rect 6910 -29620 7090 -29560
rect 7570 -29620 7750 -29560
rect 8230 -29620 8410 -29560
rect 6910 -29930 8410 -29870
rect 8730 -29450 8790 -29390
rect 9110 -29620 9290 -29560
rect 9770 -29620 9950 -29560
rect 10430 -29620 10610 -29560
rect 9110 -29930 10610 -29870
rect 10930 -29450 10990 -29390
rect 11310 -29620 11490 -29560
rect 11970 -29620 12150 -29560
rect 12630 -29620 12810 -29560
rect 11310 -29930 12810 -29870
rect 13130 -29450 13190 -29390
rect 13510 -29620 13690 -29560
rect 14170 -29620 14350 -29560
rect 14830 -29620 15010 -29560
rect 13510 -29930 15010 -29870
rect 15330 -29450 15390 -29390
rect 15710 -29760 15890 -29700
rect 16370 -29760 16550 -29700
rect 17030 -29760 17210 -29700
rect 15710 -29930 17210 -29870
rect 17530 -29450 17590 -29390
rect 17910 -29760 18090 -29700
rect 18570 -29760 18750 -29700
rect 19230 -29760 19410 -29700
rect 17910 -29930 19410 -29870
rect 19730 -29450 19790 -29390
rect 21930 -29450 21990 -29390
rect -70 -30250 -10 -30190
rect 2130 -30250 2190 -30190
rect 2510 -30420 2690 -30360
rect 3170 -30420 3350 -30360
rect 3830 -30420 4010 -30360
rect 2510 -30730 4010 -30670
rect 4330 -30250 4390 -30190
rect 4710 -30420 4890 -30360
rect 5370 -30420 5550 -30360
rect 6030 -30420 6210 -30360
rect 4710 -30730 6210 -30670
rect 6530 -30250 6590 -30190
rect 6910 -30560 7090 -30500
rect 7570 -30560 7750 -30500
rect 8230 -30560 8410 -30500
rect 6910 -30730 8410 -30670
rect 8730 -30250 8790 -30190
rect 9110 -30560 9290 -30500
rect 9770 -30560 9950 -30500
rect 10430 -30560 10610 -30500
rect 9110 -30730 10610 -30670
rect 10930 -30250 10990 -30190
rect 11310 -30560 11490 -30500
rect 11970 -30560 12150 -30500
rect 12630 -30560 12810 -30500
rect 11310 -30730 12810 -30670
rect 13130 -30250 13190 -30190
rect 13510 -30560 13690 -30500
rect 14170 -30560 14350 -30500
rect 14830 -30560 15010 -30500
rect 13510 -30730 15010 -30670
rect 15330 -30250 15390 -30190
rect 15710 -30420 15890 -30360
rect 16370 -30420 16550 -30360
rect 17030 -30420 17210 -30360
rect 15710 -30730 17210 -30670
rect 17530 -30250 17590 -30190
rect 17910 -30420 18090 -30360
rect 18570 -30420 18750 -30360
rect 19230 -30420 19410 -30360
rect 17910 -30730 19410 -30670
rect 19730 -30250 19790 -30190
rect 21930 -30250 21990 -30190
rect -70 -31050 -10 -30990
rect 2130 -31050 2190 -30990
rect 2510 -31360 2690 -31300
rect 3170 -31360 3350 -31300
rect 3830 -31360 4010 -31300
rect 4330 -31050 4390 -30990
rect 4710 -31360 4890 -31300
rect 5370 -31360 5550 -31300
rect 6030 -31360 6210 -31300
rect 6530 -31050 6590 -30990
rect 6910 -31220 7090 -31160
rect 7570 -31220 7750 -31160
rect 8230 -31220 8410 -31160
rect 8730 -31050 8790 -30990
rect 9110 -31220 9290 -31160
rect 9770 -31220 9950 -31160
rect 10430 -31220 10610 -31160
rect 10930 -31050 10990 -30990
rect 11310 -31220 11490 -31160
rect 11970 -31220 12150 -31160
rect 12630 -31220 12810 -31160
rect 13130 -31050 13190 -30990
rect 13510 -31220 13690 -31160
rect 14170 -31220 14350 -31160
rect 14830 -31220 15010 -31160
rect 15330 -31050 15390 -30990
rect 15710 -31360 15890 -31300
rect 16370 -31360 16550 -31300
rect 17030 -31360 17210 -31300
rect 17530 -31050 17590 -30990
rect 17910 -31360 18090 -31300
rect 18570 -31360 18750 -31300
rect 19230 -31360 19410 -31300
rect 19730 -31050 19790 -30990
rect 21930 -31050 21990 -30990
<< metal3 >>
rect 2200 12010 2340 12020
rect 2200 12000 2210 12010
rect 2000 11900 2210 12000
rect 2200 11890 2210 11900
rect 2330 12000 2340 12010
rect 4400 12010 4540 12020
rect 4400 12000 4410 12010
rect 2330 11900 4410 12000
rect 2330 11890 2340 11900
rect 2200 11880 2340 11890
rect 4400 11890 4410 11900
rect 4530 12000 4540 12010
rect 6600 12010 6740 12020
rect 6600 12000 6610 12010
rect 4530 11900 6610 12000
rect 4530 11890 4540 11900
rect 4400 11880 4540 11890
rect 6600 11890 6610 11900
rect 6730 12000 6740 12010
rect 8800 12010 8940 12020
rect 8800 12000 8810 12010
rect 6730 11900 8810 12000
rect 6730 11890 6740 11900
rect 6600 11880 6740 11890
rect 8800 11890 8810 11900
rect 8930 12000 8940 12010
rect 11000 12010 11140 12020
rect 11000 12000 11010 12010
rect 8930 11900 11010 12000
rect 8930 11890 8940 11900
rect 8800 11880 8940 11890
rect 11000 11890 11010 11900
rect 11130 12000 11140 12010
rect 13200 12010 13340 12020
rect 13200 12000 13210 12010
rect 11130 11900 13210 12000
rect 11130 11890 11140 11900
rect 11000 11880 11140 11890
rect 13200 11890 13210 11900
rect 13330 12000 13340 12010
rect 15400 12010 15540 12020
rect 15400 12000 15410 12010
rect 13330 11900 15410 12000
rect 13330 11890 13340 11900
rect 13200 11880 13340 11890
rect 15400 11890 15410 11900
rect 15530 12000 15540 12010
rect 17600 12010 17740 12020
rect 17600 12000 17610 12010
rect 15530 11900 17610 12000
rect 15530 11890 15540 11900
rect 15400 11880 15540 11890
rect 17600 11890 17610 11900
rect 17730 12000 17740 12010
rect 19800 12010 19940 12020
rect 19800 12000 19810 12010
rect 17730 11900 19810 12000
rect 17730 11890 17740 11900
rect 17600 11880 17740 11890
rect 19800 11890 19810 11900
rect 19930 12000 19940 12010
rect 19930 11900 28700 12000
rect 19930 11890 19940 11900
rect 19800 11880 19940 11890
rect 1980 11710 2120 11720
rect 1980 11590 1990 11710
rect 2110 11700 2120 11710
rect 4180 11710 4320 11720
rect 4180 11700 4190 11710
rect 2110 11600 4190 11700
rect 2110 11590 2120 11600
rect 1980 11580 2120 11590
rect 4180 11590 4190 11600
rect 4310 11700 4320 11710
rect 6380 11710 6520 11720
rect 6380 11700 6390 11710
rect 4310 11600 6390 11700
rect 4310 11590 4320 11600
rect 4180 11580 4320 11590
rect 6380 11590 6390 11600
rect 6510 11700 6520 11710
rect 8580 11710 8720 11720
rect 8580 11700 8590 11710
rect 6510 11600 8590 11700
rect 6510 11590 6520 11600
rect 6380 11580 6520 11590
rect 8580 11590 8590 11600
rect 8710 11700 8720 11710
rect 10780 11710 10920 11720
rect 10780 11700 10790 11710
rect 8710 11600 10790 11700
rect 8710 11590 8720 11600
rect 8580 11580 8720 11590
rect 10780 11590 10790 11600
rect 10910 11700 10920 11710
rect 12980 11710 13120 11720
rect 12980 11700 12990 11710
rect 10910 11600 12990 11700
rect 10910 11590 10920 11600
rect 10780 11580 10920 11590
rect 12980 11590 12990 11600
rect 13110 11700 13120 11710
rect 15180 11710 15320 11720
rect 15180 11700 15190 11710
rect 13110 11600 15190 11700
rect 13110 11590 13120 11600
rect 12980 11580 13120 11590
rect 15180 11590 15190 11600
rect 15310 11700 15320 11710
rect 17380 11710 17520 11720
rect 17380 11700 17390 11710
rect 15310 11600 17390 11700
rect 15310 11590 15320 11600
rect 15180 11580 15320 11590
rect 17380 11590 17390 11600
rect 17510 11700 17520 11710
rect 19580 11710 19720 11720
rect 19580 11700 19590 11710
rect 17510 11600 19590 11700
rect 17510 11590 17520 11600
rect 17380 11580 17520 11590
rect 19580 11590 19590 11600
rect 19710 11700 19720 11710
rect 19710 11600 28700 11700
rect 19710 11590 19720 11600
rect 19580 11580 19720 11590
rect 820 11250 1020 11260
rect 20500 11250 20700 11260
rect 820 11240 830 11250
rect -220 11180 830 11240
rect 820 11170 830 11180
rect 1010 11240 1020 11250
rect 2500 11240 2700 11250
rect 3160 11240 3360 11250
rect 3820 11240 4020 11250
rect 4700 11240 4900 11250
rect 5360 11240 5560 11250
rect 6020 11240 6220 11250
rect 6900 11240 7100 11250
rect 7560 11240 7760 11250
rect 8220 11240 8420 11250
rect 9100 11240 9300 11250
rect 9760 11240 9960 11250
rect 10420 11240 10620 11250
rect 11300 11240 11500 11250
rect 11960 11240 12160 11250
rect 12620 11240 12820 11250
rect 13500 11240 13700 11250
rect 14160 11240 14360 11250
rect 14820 11240 15020 11250
rect 15700 11240 15900 11250
rect 16360 11240 16560 11250
rect 17020 11240 17220 11250
rect 17900 11240 18100 11250
rect 18560 11240 18760 11250
rect 19220 11240 19420 11250
rect 20500 11240 20510 11250
rect 1010 11180 2510 11240
rect 2690 11180 3170 11240
rect 3350 11180 3830 11240
rect 4010 11180 4710 11240
rect 4890 11180 5370 11240
rect 5550 11180 6030 11240
rect 6210 11180 15710 11240
rect 15890 11180 16370 11240
rect 16550 11180 17030 11240
rect 17210 11180 17910 11240
rect 18090 11180 18570 11240
rect 18750 11180 19230 11240
rect 19410 11180 20510 11240
rect 1010 11170 1020 11180
rect 2500 11170 2700 11180
rect 3160 11170 3360 11180
rect 3820 11170 4020 11180
rect 4700 11170 4900 11180
rect 5360 11170 5560 11180
rect 6020 11170 6220 11180
rect 6900 11170 7100 11180
rect 7560 11170 7760 11180
rect 8220 11170 8420 11180
rect 9100 11170 9300 11180
rect 9760 11170 9960 11180
rect 10420 11170 10620 11180
rect 11300 11170 11500 11180
rect 11960 11170 12160 11180
rect 12620 11170 12820 11180
rect 13500 11170 13700 11180
rect 14160 11170 14360 11180
rect 14820 11170 15020 11180
rect 15700 11170 15900 11180
rect 16360 11170 16560 11180
rect 17020 11170 17220 11180
rect 17900 11170 18100 11180
rect 18560 11170 18760 11180
rect 19220 11170 19420 11180
rect 20500 11170 20510 11180
rect 20690 11240 20700 11250
rect 20690 11180 22180 11240
rect 20690 11170 20700 11180
rect 820 11160 1020 11170
rect 20500 11160 20700 11170
rect 1220 11110 1420 11120
rect 20900 11110 21100 11120
rect 1220 11100 1230 11110
rect -220 11040 1230 11100
rect 1220 11030 1230 11040
rect 1410 11100 1420 11110
rect 2500 11100 2700 11110
rect 3160 11100 3360 11110
rect 3820 11100 4020 11110
rect 4700 11100 4900 11110
rect 5360 11100 5560 11110
rect 6020 11100 6220 11110
rect 6900 11100 7100 11110
rect 7560 11100 7760 11110
rect 8220 11100 8420 11110
rect 9100 11100 9300 11110
rect 9760 11100 9960 11110
rect 10420 11100 10620 11110
rect 11300 11100 11500 11110
rect 11960 11100 12160 11110
rect 12620 11100 12820 11110
rect 13500 11100 13700 11110
rect 14160 11100 14360 11110
rect 14820 11100 15020 11110
rect 15700 11100 15900 11110
rect 16360 11100 16560 11110
rect 17020 11100 17220 11110
rect 17900 11100 18100 11110
rect 18560 11100 18760 11110
rect 19220 11100 19420 11110
rect 20900 11100 20910 11110
rect 1410 11040 6910 11100
rect 7090 11040 7570 11100
rect 7750 11040 8230 11100
rect 8410 11040 9110 11100
rect 9290 11040 9770 11100
rect 9950 11040 10430 11100
rect 10610 11040 11310 11100
rect 11490 11040 11970 11100
rect 12150 11040 12630 11100
rect 12810 11040 13510 11100
rect 13690 11040 14170 11100
rect 14350 11040 14830 11100
rect 15010 11040 20910 11100
rect 1410 11030 1420 11040
rect 2500 11030 2700 11040
rect 3160 11030 3360 11040
rect 3820 11030 4020 11040
rect 4700 11030 4900 11040
rect 5360 11030 5560 11040
rect 6020 11030 6220 11040
rect 6900 11030 7100 11040
rect 7560 11030 7760 11040
rect 8220 11030 8420 11040
rect 9100 11030 9300 11040
rect 9760 11030 9960 11040
rect 10420 11030 10620 11040
rect 11300 11030 11500 11040
rect 11960 11030 12160 11040
rect 12620 11030 12820 11040
rect 13500 11030 13700 11040
rect 14160 11030 14360 11040
rect 14820 11030 15020 11040
rect 15700 11030 15900 11040
rect 16360 11030 16560 11040
rect 17020 11030 17220 11040
rect 17900 11030 18100 11040
rect 18560 11030 18760 11040
rect 19220 11030 19420 11040
rect 20900 11030 20910 11040
rect 21090 11100 21100 11110
rect 21090 11040 22180 11100
rect 21090 11030 21100 11040
rect 1220 11020 1420 11030
rect 20900 11020 21100 11030
rect -110 10940 30 10960
rect -110 10690 -80 10940
rect 0 10690 30 10940
rect -110 10660 30 10690
rect 2090 10940 2230 10960
rect 2090 10690 2120 10940
rect 2200 10690 2230 10940
rect 2090 10660 2230 10690
rect 4290 10940 4430 10960
rect 4290 10690 4320 10940
rect 4400 10690 4430 10940
rect 4290 10660 4430 10690
rect 6490 10940 6630 10960
rect 6490 10690 6520 10940
rect 6600 10690 6630 10940
rect 6490 10660 6630 10690
rect 8690 10940 8830 10960
rect 8690 10690 8720 10940
rect 8800 10690 8830 10940
rect 8690 10660 8830 10690
rect 10890 10940 11030 10960
rect 10890 10690 10920 10940
rect 11000 10690 11030 10940
rect 10890 10660 11030 10690
rect 13090 10940 13230 10960
rect 13090 10690 13120 10940
rect 13200 10690 13230 10940
rect 13090 10660 13230 10690
rect 15290 10940 15430 10960
rect 15290 10690 15320 10940
rect 15400 10690 15430 10940
rect 15290 10660 15430 10690
rect 17490 10940 17630 10960
rect 17490 10690 17520 10940
rect 17600 10690 17630 10940
rect 17490 10660 17630 10690
rect 19690 10940 19830 10960
rect 19690 10690 19720 10940
rect 19800 10690 19830 10940
rect 19690 10660 19830 10690
rect 21890 10940 22030 10960
rect 21890 10690 21920 10940
rect 22000 10690 22030 10940
rect 21890 10660 22030 10690
rect 2500 10610 4020 10620
rect 1620 10590 1820 10600
rect 1620 10580 1630 10590
rect 1600 10520 1630 10580
rect 1620 10510 1630 10520
rect 1810 10580 1820 10590
rect 2500 10580 2510 10610
rect 1810 10550 2510 10580
rect 4010 10580 4020 10610
rect 4700 10610 6220 10620
rect 4700 10580 4710 10610
rect 4010 10550 4710 10580
rect 6210 10580 6220 10610
rect 6900 10610 8420 10620
rect 6900 10580 6910 10610
rect 6210 10550 6910 10580
rect 8410 10580 8420 10610
rect 9100 10610 10620 10620
rect 9100 10580 9110 10610
rect 8410 10550 9110 10580
rect 10610 10580 10620 10610
rect 11300 10610 12820 10620
rect 11300 10580 11310 10610
rect 10610 10550 11310 10580
rect 12810 10580 12820 10610
rect 13500 10610 15020 10620
rect 13500 10580 13510 10610
rect 12810 10550 13510 10580
rect 15010 10580 15020 10610
rect 15700 10610 17220 10620
rect 15700 10580 15710 10610
rect 15010 10550 15710 10580
rect 17210 10580 17220 10610
rect 17900 10610 19420 10620
rect 17900 10580 17910 10610
rect 17210 10550 17910 10580
rect 19410 10580 19420 10610
rect 20100 10590 20300 10600
rect 20100 10580 20110 10590
rect 19410 10550 20110 10580
rect 1810 10520 20110 10550
rect 1810 10510 1820 10520
rect 1620 10500 1820 10510
rect 20100 10510 20110 10520
rect 20290 10580 20300 10590
rect 20290 10520 20320 10580
rect 20290 10510 20300 10520
rect 20100 10500 20300 10510
rect 820 10450 1020 10460
rect 20500 10450 20700 10460
rect 820 10440 830 10450
rect -220 10380 830 10440
rect 820 10370 830 10380
rect 1010 10440 1020 10450
rect 2500 10440 2700 10450
rect 3160 10440 3360 10450
rect 3820 10440 4020 10450
rect 4700 10440 4900 10450
rect 5360 10440 5560 10450
rect 6020 10440 6220 10450
rect 6900 10440 7100 10450
rect 7560 10440 7760 10450
rect 8220 10440 8420 10450
rect 9100 10440 9300 10450
rect 9760 10440 9960 10450
rect 10420 10440 10620 10450
rect 11300 10440 11500 10450
rect 11960 10440 12160 10450
rect 12620 10440 12820 10450
rect 13500 10440 13700 10450
rect 14160 10440 14360 10450
rect 14820 10440 15020 10450
rect 15700 10440 15900 10450
rect 16360 10440 16560 10450
rect 17020 10440 17220 10450
rect 17900 10440 18100 10450
rect 18560 10440 18760 10450
rect 19220 10440 19420 10450
rect 20500 10440 20510 10450
rect 1010 10380 6910 10440
rect 7090 10380 7570 10440
rect 7750 10380 8230 10440
rect 8410 10380 9110 10440
rect 9290 10380 9770 10440
rect 9950 10380 10430 10440
rect 10610 10380 11310 10440
rect 11490 10380 11970 10440
rect 12150 10380 12630 10440
rect 12810 10380 13510 10440
rect 13690 10380 14170 10440
rect 14350 10380 14830 10440
rect 15010 10380 20510 10440
rect 1010 10370 1020 10380
rect 2500 10370 2700 10380
rect 3160 10370 3360 10380
rect 3820 10370 4020 10380
rect 4700 10370 4900 10380
rect 5360 10370 5560 10380
rect 6020 10370 6220 10380
rect 6900 10370 7100 10380
rect 7560 10370 7760 10380
rect 8220 10370 8420 10380
rect 9100 10370 9300 10380
rect 9760 10370 9960 10380
rect 10420 10370 10620 10380
rect 11300 10370 11500 10380
rect 11960 10370 12160 10380
rect 12620 10370 12820 10380
rect 13500 10370 13700 10380
rect 14160 10370 14360 10380
rect 14820 10370 15020 10380
rect 15700 10370 15900 10380
rect 16360 10370 16560 10380
rect 17020 10370 17220 10380
rect 17900 10370 18100 10380
rect 18560 10370 18760 10380
rect 19220 10370 19420 10380
rect 20500 10370 20510 10380
rect 20690 10440 20700 10450
rect 20690 10380 22180 10440
rect 20690 10370 20700 10380
rect 820 10360 1020 10370
rect 20500 10360 20700 10370
rect 1220 10310 1420 10320
rect 20900 10310 21100 10320
rect 1220 10300 1230 10310
rect -220 10240 1230 10300
rect 1220 10230 1230 10240
rect 1410 10300 1420 10310
rect 2500 10300 2700 10310
rect 3160 10300 3360 10310
rect 3820 10300 4020 10310
rect 4700 10300 4900 10310
rect 5360 10300 5560 10310
rect 6020 10300 6220 10310
rect 6900 10300 7100 10310
rect 7560 10300 7760 10310
rect 8220 10300 8420 10310
rect 9100 10300 9300 10310
rect 9760 10300 9960 10310
rect 10420 10300 10620 10310
rect 11300 10300 11500 10310
rect 11960 10300 12160 10310
rect 12620 10300 12820 10310
rect 13500 10300 13700 10310
rect 14160 10300 14360 10310
rect 14820 10300 15020 10310
rect 15700 10300 15900 10310
rect 16360 10300 16560 10310
rect 17020 10300 17220 10310
rect 17900 10300 18100 10310
rect 18560 10300 18760 10310
rect 19220 10300 19420 10310
rect 20900 10300 20910 10310
rect 1410 10240 2510 10300
rect 2690 10240 3170 10300
rect 3350 10240 3830 10300
rect 4010 10240 4710 10300
rect 4890 10240 5370 10300
rect 5550 10240 6030 10300
rect 6210 10240 15710 10300
rect 15890 10240 16370 10300
rect 16550 10240 17030 10300
rect 17210 10240 17910 10300
rect 18090 10240 18570 10300
rect 18750 10240 19230 10300
rect 19410 10240 20910 10300
rect 1410 10230 1420 10240
rect 2500 10230 2700 10240
rect 3160 10230 3360 10240
rect 3820 10230 4020 10240
rect 4700 10230 4900 10240
rect 5360 10230 5560 10240
rect 6020 10230 6220 10240
rect 6900 10230 7100 10240
rect 7560 10230 7760 10240
rect 8220 10230 8420 10240
rect 9100 10230 9300 10240
rect 9760 10230 9960 10240
rect 10420 10230 10620 10240
rect 11300 10230 11500 10240
rect 11960 10230 12160 10240
rect 12620 10230 12820 10240
rect 13500 10230 13700 10240
rect 14160 10230 14360 10240
rect 14820 10230 15020 10240
rect 15700 10230 15900 10240
rect 16360 10230 16560 10240
rect 17020 10230 17220 10240
rect 17900 10230 18100 10240
rect 18560 10230 18760 10240
rect 19220 10230 19420 10240
rect 20900 10230 20910 10240
rect 21090 10300 21100 10310
rect 21090 10240 22180 10300
rect 21090 10230 21100 10240
rect 1220 10220 1420 10230
rect 20900 10220 21100 10230
rect -110 10140 30 10160
rect -110 9890 -80 10140
rect 0 9890 30 10140
rect -110 9860 30 9890
rect 2090 10140 2230 10160
rect 2090 9890 2120 10140
rect 2200 9890 2230 10140
rect 2090 9860 2230 9890
rect 4290 10140 4430 10160
rect 4290 9890 4320 10140
rect 4400 9890 4430 10140
rect 4290 9860 4430 9890
rect 6490 10140 6630 10160
rect 6490 9890 6520 10140
rect 6600 9890 6630 10140
rect 6490 9860 6630 9890
rect 8690 10140 8830 10160
rect 8690 9890 8720 10140
rect 8800 9890 8830 10140
rect 8690 9860 8830 9890
rect 10890 10140 11030 10160
rect 10890 9890 10920 10140
rect 11000 9890 11030 10140
rect 10890 9860 11030 9890
rect 13090 10140 13230 10160
rect 13090 9890 13120 10140
rect 13200 9890 13230 10140
rect 13090 9860 13230 9890
rect 15290 10140 15430 10160
rect 15290 9890 15320 10140
rect 15400 9890 15430 10140
rect 15290 9860 15430 9890
rect 17490 10140 17630 10160
rect 17490 9890 17520 10140
rect 17600 9890 17630 10140
rect 17490 9860 17630 9890
rect 19690 10140 19830 10160
rect 19690 9890 19720 10140
rect 19800 9890 19830 10140
rect 19690 9860 19830 9890
rect 21890 10140 22030 10160
rect 21890 9890 21920 10140
rect 22000 9890 22030 10140
rect 21890 9860 22030 9890
rect 2500 9810 4020 9820
rect 1620 9790 1820 9800
rect 1620 9780 1630 9790
rect 1600 9720 1630 9780
rect 1620 9710 1630 9720
rect 1810 9780 1820 9790
rect 2500 9780 2510 9810
rect 1810 9750 2510 9780
rect 4010 9780 4020 9810
rect 4700 9810 6220 9820
rect 4700 9780 4710 9810
rect 4010 9750 4710 9780
rect 6210 9780 6220 9810
rect 6900 9810 8420 9820
rect 6900 9780 6910 9810
rect 6210 9750 6910 9780
rect 8410 9780 8420 9810
rect 9100 9810 10620 9820
rect 9100 9780 9110 9810
rect 8410 9750 9110 9780
rect 10610 9780 10620 9810
rect 11300 9810 12820 9820
rect 11300 9780 11310 9810
rect 10610 9750 11310 9780
rect 12810 9780 12820 9810
rect 13500 9810 15020 9820
rect 13500 9780 13510 9810
rect 12810 9750 13510 9780
rect 15010 9780 15020 9810
rect 15700 9810 17220 9820
rect 15700 9780 15710 9810
rect 15010 9750 15710 9780
rect 17210 9780 17220 9810
rect 17900 9810 19420 9820
rect 17900 9780 17910 9810
rect 17210 9750 17910 9780
rect 19410 9780 19420 9810
rect 20100 9790 20300 9800
rect 20100 9780 20110 9790
rect 19410 9750 20110 9780
rect 1810 9720 20110 9750
rect 1810 9710 1820 9720
rect 1620 9700 1820 9710
rect 20100 9710 20110 9720
rect 20290 9780 20300 9790
rect 20290 9720 20320 9780
rect 20290 9710 20300 9720
rect 20100 9700 20300 9710
rect 820 9650 1020 9660
rect 20500 9650 20700 9660
rect 820 9640 830 9650
rect -220 9580 830 9640
rect 820 9570 830 9580
rect 1010 9640 1020 9650
rect 2500 9640 2700 9650
rect 3160 9640 3360 9650
rect 3820 9640 4020 9650
rect 4700 9640 4900 9650
rect 5360 9640 5560 9650
rect 6020 9640 6220 9650
rect 6900 9640 7100 9650
rect 7560 9640 7760 9650
rect 8220 9640 8420 9650
rect 9100 9640 9300 9650
rect 9760 9640 9960 9650
rect 10420 9640 10620 9650
rect 11300 9640 11500 9650
rect 11960 9640 12160 9650
rect 12620 9640 12820 9650
rect 13500 9640 13700 9650
rect 14160 9640 14360 9650
rect 14820 9640 15020 9650
rect 15700 9640 15900 9650
rect 16360 9640 16560 9650
rect 17020 9640 17220 9650
rect 17900 9640 18100 9650
rect 18560 9640 18760 9650
rect 19220 9640 19420 9650
rect 20500 9640 20510 9650
rect 1010 9580 2510 9640
rect 2690 9580 3170 9640
rect 3350 9580 3830 9640
rect 4010 9580 4710 9640
rect 4890 9580 5370 9640
rect 5550 9580 6030 9640
rect 6210 9580 15710 9640
rect 15890 9580 16370 9640
rect 16550 9580 17030 9640
rect 17210 9580 17910 9640
rect 18090 9580 18570 9640
rect 18750 9580 19230 9640
rect 19410 9580 20510 9640
rect 1010 9570 1020 9580
rect 2500 9570 2700 9580
rect 3160 9570 3360 9580
rect 3820 9570 4020 9580
rect 4700 9570 4900 9580
rect 5360 9570 5560 9580
rect 6020 9570 6220 9580
rect 6900 9570 7100 9580
rect 7560 9570 7760 9580
rect 8220 9570 8420 9580
rect 9100 9570 9300 9580
rect 9760 9570 9960 9580
rect 10420 9570 10620 9580
rect 11300 9570 11500 9580
rect 11960 9570 12160 9580
rect 12620 9570 12820 9580
rect 13500 9570 13700 9580
rect 14160 9570 14360 9580
rect 14820 9570 15020 9580
rect 15700 9570 15900 9580
rect 16360 9570 16560 9580
rect 17020 9570 17220 9580
rect 17900 9570 18100 9580
rect 18560 9570 18760 9580
rect 19220 9570 19420 9580
rect 20500 9570 20510 9580
rect 20690 9640 20700 9650
rect 20690 9580 22180 9640
rect 20690 9570 20700 9580
rect 820 9560 1020 9570
rect 20500 9560 20700 9570
rect 1220 9510 1420 9520
rect 20900 9510 21100 9520
rect 1220 9500 1230 9510
rect -220 9440 1230 9500
rect 1220 9430 1230 9440
rect 1410 9500 1420 9510
rect 2500 9500 2700 9510
rect 3160 9500 3360 9510
rect 3820 9500 4020 9510
rect 4700 9500 4900 9510
rect 5360 9500 5560 9510
rect 6020 9500 6220 9510
rect 6900 9500 7100 9510
rect 7560 9500 7760 9510
rect 8220 9500 8420 9510
rect 9100 9500 9300 9510
rect 9760 9500 9960 9510
rect 10420 9500 10620 9510
rect 11300 9500 11500 9510
rect 11960 9500 12160 9510
rect 12620 9500 12820 9510
rect 13500 9500 13700 9510
rect 14160 9500 14360 9510
rect 14820 9500 15020 9510
rect 15700 9500 15900 9510
rect 16360 9500 16560 9510
rect 17020 9500 17220 9510
rect 17900 9500 18100 9510
rect 18560 9500 18760 9510
rect 19220 9500 19420 9510
rect 20900 9500 20910 9510
rect 1410 9440 6910 9500
rect 7090 9440 7570 9500
rect 7750 9440 8230 9500
rect 8410 9440 9110 9500
rect 9290 9440 9770 9500
rect 9950 9440 10430 9500
rect 10610 9440 11310 9500
rect 11490 9440 11970 9500
rect 12150 9440 12630 9500
rect 12810 9440 13510 9500
rect 13690 9440 14170 9500
rect 14350 9440 14830 9500
rect 15010 9440 20910 9500
rect 1410 9430 1420 9440
rect 2500 9430 2700 9440
rect 3160 9430 3360 9440
rect 3820 9430 4020 9440
rect 4700 9430 4900 9440
rect 5360 9430 5560 9440
rect 6020 9430 6220 9440
rect 6900 9430 7100 9440
rect 7560 9430 7760 9440
rect 8220 9430 8420 9440
rect 9100 9430 9300 9440
rect 9760 9430 9960 9440
rect 10420 9430 10620 9440
rect 11300 9430 11500 9440
rect 11960 9430 12160 9440
rect 12620 9430 12820 9440
rect 13500 9430 13700 9440
rect 14160 9430 14360 9440
rect 14820 9430 15020 9440
rect 15700 9430 15900 9440
rect 16360 9430 16560 9440
rect 17020 9430 17220 9440
rect 17900 9430 18100 9440
rect 18560 9430 18760 9440
rect 19220 9430 19420 9440
rect 20900 9430 20910 9440
rect 21090 9500 21100 9510
rect 21090 9440 22180 9500
rect 21090 9430 21100 9440
rect 1220 9420 1420 9430
rect 20900 9420 21100 9430
rect -110 9340 30 9360
rect -110 9090 -80 9340
rect 0 9090 30 9340
rect -110 9060 30 9090
rect 2090 9340 2230 9360
rect 2090 9090 2120 9340
rect 2200 9090 2230 9340
rect 2090 9060 2230 9090
rect 4290 9340 4430 9360
rect 4290 9090 4320 9340
rect 4400 9090 4430 9340
rect 4290 9060 4430 9090
rect 6490 9340 6630 9360
rect 6490 9090 6520 9340
rect 6600 9090 6630 9340
rect 6490 9060 6630 9090
rect 8690 9340 8830 9360
rect 8690 9090 8720 9340
rect 8800 9090 8830 9340
rect 8690 9060 8830 9090
rect 10890 9340 11030 9360
rect 10890 9090 10920 9340
rect 11000 9090 11030 9340
rect 10890 9060 11030 9090
rect 13090 9340 13230 9360
rect 13090 9090 13120 9340
rect 13200 9090 13230 9340
rect 13090 9060 13230 9090
rect 15290 9340 15430 9360
rect 15290 9090 15320 9340
rect 15400 9090 15430 9340
rect 15290 9060 15430 9090
rect 17490 9340 17630 9360
rect 17490 9090 17520 9340
rect 17600 9090 17630 9340
rect 17490 9060 17630 9090
rect 19690 9340 19830 9360
rect 19690 9090 19720 9340
rect 19800 9090 19830 9340
rect 19690 9060 19830 9090
rect 21890 9340 22030 9360
rect 21890 9090 21920 9340
rect 22000 9090 22030 9340
rect 21890 9060 22030 9090
rect 4700 9010 6220 9020
rect 420 8990 620 9000
rect 420 8910 430 8990
rect 610 8910 620 8990
rect 1620 8990 1820 9000
rect 1620 8980 1630 8990
rect 1600 8920 1630 8980
rect 420 8900 620 8910
rect 1620 8910 1630 8920
rect 1810 8980 1820 8990
rect 4700 8980 4710 9010
rect 1810 8950 4710 8980
rect 6210 8980 6220 9010
rect 6900 9010 8420 9020
rect 6900 8980 6910 9010
rect 6210 8950 6910 8980
rect 8410 8980 8420 9010
rect 9100 9010 10620 9020
rect 9100 8980 9110 9010
rect 8410 8950 9110 8980
rect 10610 8980 10620 9010
rect 11300 9010 12820 9020
rect 11300 8980 11310 9010
rect 10610 8950 11310 8980
rect 12810 8980 12820 9010
rect 13500 9010 15020 9020
rect 13500 8980 13510 9010
rect 12810 8950 13510 8980
rect 15010 8980 15020 9010
rect 15700 9010 17220 9020
rect 15700 8980 15710 9010
rect 15010 8950 15710 8980
rect 17210 8980 17220 9010
rect 20100 8990 20300 9000
rect 20100 8980 20110 8990
rect 17210 8950 20110 8980
rect 1810 8920 20110 8950
rect 1810 8910 1820 8920
rect 1620 8900 1820 8910
rect 20100 8910 20110 8920
rect 20290 8980 20300 8990
rect 21300 8990 21500 9000
rect 20290 8920 20320 8980
rect 20290 8910 20300 8920
rect 20100 8900 20300 8910
rect 21300 8910 21310 8990
rect 21490 8910 21500 8990
rect 21300 8900 21500 8910
rect 820 8850 1020 8860
rect 20500 8850 20700 8860
rect 820 8840 830 8850
rect -220 8780 830 8840
rect 820 8770 830 8780
rect 1010 8840 1020 8850
rect 2500 8840 2700 8850
rect 3160 8840 3360 8850
rect 3820 8840 4020 8850
rect 4700 8840 4900 8850
rect 5360 8840 5560 8850
rect 6020 8840 6220 8850
rect 6900 8840 7100 8850
rect 7560 8840 7760 8850
rect 8220 8840 8420 8850
rect 9100 8840 9300 8850
rect 9760 8840 9960 8850
rect 10420 8840 10620 8850
rect 11300 8840 11500 8850
rect 11960 8840 12160 8850
rect 12620 8840 12820 8850
rect 13500 8840 13700 8850
rect 14160 8840 14360 8850
rect 14820 8840 15020 8850
rect 15700 8840 15900 8850
rect 16360 8840 16560 8850
rect 17020 8840 17220 8850
rect 17900 8840 18100 8850
rect 18560 8840 18760 8850
rect 19220 8840 19420 8850
rect 20500 8840 20510 8850
rect 1010 8780 6910 8840
rect 7090 8780 7570 8840
rect 7750 8780 8230 8840
rect 8410 8780 9110 8840
rect 9290 8780 9770 8840
rect 9950 8780 10430 8840
rect 10610 8780 11310 8840
rect 11490 8780 11970 8840
rect 12150 8780 12630 8840
rect 12810 8780 13510 8840
rect 13690 8780 14170 8840
rect 14350 8780 14830 8840
rect 15010 8780 20510 8840
rect 1010 8770 1020 8780
rect 2500 8770 2700 8780
rect 3160 8770 3360 8780
rect 3820 8770 4020 8780
rect 4700 8770 4900 8780
rect 5360 8770 5560 8780
rect 6020 8770 6220 8780
rect 6900 8770 7100 8780
rect 7560 8770 7760 8780
rect 8220 8770 8420 8780
rect 9100 8770 9300 8780
rect 9760 8770 9960 8780
rect 10420 8770 10620 8780
rect 11300 8770 11500 8780
rect 11960 8770 12160 8780
rect 12620 8770 12820 8780
rect 13500 8770 13700 8780
rect 14160 8770 14360 8780
rect 14820 8770 15020 8780
rect 15700 8770 15900 8780
rect 16360 8770 16560 8780
rect 17020 8770 17220 8780
rect 17900 8770 18100 8780
rect 18560 8770 18760 8780
rect 19220 8770 19420 8780
rect 20500 8770 20510 8780
rect 20690 8840 20700 8850
rect 20690 8780 22180 8840
rect 20690 8770 20700 8780
rect 820 8760 1020 8770
rect 20500 8760 20700 8770
rect 1220 8710 1420 8720
rect 20900 8710 21100 8720
rect 1220 8700 1230 8710
rect -220 8640 1230 8700
rect 1220 8630 1230 8640
rect 1410 8700 1420 8710
rect 2500 8700 2700 8710
rect 3160 8700 3360 8710
rect 3820 8700 4020 8710
rect 4700 8700 4900 8710
rect 5360 8700 5560 8710
rect 6020 8700 6220 8710
rect 6900 8700 7100 8710
rect 7560 8700 7760 8710
rect 8220 8700 8420 8710
rect 9100 8700 9300 8710
rect 9760 8700 9960 8710
rect 10420 8700 10620 8710
rect 11300 8700 11500 8710
rect 11960 8700 12160 8710
rect 12620 8700 12820 8710
rect 13500 8700 13700 8710
rect 14160 8700 14360 8710
rect 14820 8700 15020 8710
rect 15700 8700 15900 8710
rect 16360 8700 16560 8710
rect 17020 8700 17220 8710
rect 17900 8700 18100 8710
rect 18560 8700 18760 8710
rect 19220 8700 19420 8710
rect 20900 8700 20910 8710
rect 1410 8640 2510 8700
rect 2690 8640 3170 8700
rect 3350 8640 3830 8700
rect 4010 8640 4710 8700
rect 4890 8640 5370 8700
rect 5550 8640 6030 8700
rect 6210 8640 15710 8700
rect 15890 8640 16370 8700
rect 16550 8640 17030 8700
rect 17210 8640 17910 8700
rect 18090 8640 18570 8700
rect 18750 8640 19230 8700
rect 19410 8640 20910 8700
rect 1410 8630 1420 8640
rect 2500 8630 2700 8640
rect 3160 8630 3360 8640
rect 3820 8630 4020 8640
rect 4700 8630 4900 8640
rect 5360 8630 5560 8640
rect 6020 8630 6220 8640
rect 6900 8630 7100 8640
rect 7560 8630 7760 8640
rect 8220 8630 8420 8640
rect 9100 8630 9300 8640
rect 9760 8630 9960 8640
rect 10420 8630 10620 8640
rect 11300 8630 11500 8640
rect 11960 8630 12160 8640
rect 12620 8630 12820 8640
rect 13500 8630 13700 8640
rect 14160 8630 14360 8640
rect 14820 8630 15020 8640
rect 15700 8630 15900 8640
rect 16360 8630 16560 8640
rect 17020 8630 17220 8640
rect 17900 8630 18100 8640
rect 18560 8630 18760 8640
rect 19220 8630 19420 8640
rect 20900 8630 20910 8640
rect 21090 8700 21100 8710
rect 21090 8640 22180 8700
rect 21090 8630 21100 8640
rect 1220 8620 1420 8630
rect 20900 8620 21100 8630
rect -110 8540 30 8560
rect -110 8290 -80 8540
rect 0 8290 30 8540
rect -110 8260 30 8290
rect 2090 8540 2230 8560
rect 2090 8290 2120 8540
rect 2200 8290 2230 8540
rect 2090 8260 2230 8290
rect 4290 8540 4430 8560
rect 4290 8290 4320 8540
rect 4400 8290 4430 8540
rect 4290 8260 4430 8290
rect 6490 8540 6630 8560
rect 6490 8290 6520 8540
rect 6600 8290 6630 8540
rect 6490 8260 6630 8290
rect 8690 8540 8830 8560
rect 8690 8290 8720 8540
rect 8800 8290 8830 8540
rect 8690 8260 8830 8290
rect 10890 8540 11030 8560
rect 10890 8290 10920 8540
rect 11000 8290 11030 8540
rect 10890 8260 11030 8290
rect 13090 8540 13230 8560
rect 13090 8290 13120 8540
rect 13200 8290 13230 8540
rect 13090 8260 13230 8290
rect 15290 8540 15430 8560
rect 15290 8290 15320 8540
rect 15400 8290 15430 8540
rect 15290 8260 15430 8290
rect 17490 8540 17630 8560
rect 17490 8290 17520 8540
rect 17600 8290 17630 8540
rect 17490 8260 17630 8290
rect 19690 8540 19830 8560
rect 19690 8290 19720 8540
rect 19800 8290 19830 8540
rect 19690 8260 19830 8290
rect 21890 8540 22030 8560
rect 21890 8290 21920 8540
rect 22000 8290 22030 8540
rect 21890 8260 22030 8290
rect 4700 8210 6220 8220
rect 420 8190 620 8200
rect 420 8110 430 8190
rect 610 8110 620 8190
rect 1620 8190 1820 8200
rect 1620 8180 1630 8190
rect 1600 8120 1630 8180
rect 420 8100 620 8110
rect 1620 8110 1630 8120
rect 1810 8180 1820 8190
rect 4700 8180 4710 8210
rect 1810 8150 4710 8180
rect 6210 8180 6220 8210
rect 6900 8210 8420 8220
rect 6900 8180 6910 8210
rect 6210 8150 6910 8180
rect 8410 8180 8420 8210
rect 9100 8210 10620 8220
rect 9100 8180 9110 8210
rect 8410 8150 9110 8180
rect 10610 8180 10620 8210
rect 11300 8210 12820 8220
rect 11300 8180 11310 8210
rect 10610 8150 11310 8180
rect 12810 8180 12820 8210
rect 13500 8210 15020 8220
rect 13500 8180 13510 8210
rect 12810 8150 13510 8180
rect 15010 8180 15020 8210
rect 15700 8210 17220 8220
rect 15700 8180 15710 8210
rect 15010 8150 15710 8180
rect 17210 8180 17220 8210
rect 20100 8190 20300 8200
rect 20100 8180 20110 8190
rect 17210 8150 20110 8180
rect 1810 8120 20110 8150
rect 1810 8110 1820 8120
rect 1620 8100 1820 8110
rect 20100 8110 20110 8120
rect 20290 8180 20300 8190
rect 21300 8190 21500 8200
rect 20290 8120 20320 8180
rect 20290 8110 20300 8120
rect 20100 8100 20300 8110
rect 21300 8110 21310 8190
rect 21490 8110 21500 8190
rect 21300 8100 21500 8110
rect 820 8050 1020 8060
rect 20500 8050 20700 8060
rect 820 8040 830 8050
rect -220 7980 830 8040
rect 820 7970 830 7980
rect 1010 8040 1020 8050
rect 2500 8040 2700 8050
rect 3160 8040 3360 8050
rect 3820 8040 4020 8050
rect 4700 8040 4900 8050
rect 5360 8040 5560 8050
rect 6020 8040 6220 8050
rect 6900 8040 7100 8050
rect 7560 8040 7760 8050
rect 8220 8040 8420 8050
rect 9100 8040 9300 8050
rect 9760 8040 9960 8050
rect 10420 8040 10620 8050
rect 11300 8040 11500 8050
rect 11960 8040 12160 8050
rect 12620 8040 12820 8050
rect 13500 8040 13700 8050
rect 14160 8040 14360 8050
rect 14820 8040 15020 8050
rect 15700 8040 15900 8050
rect 16360 8040 16560 8050
rect 17020 8040 17220 8050
rect 17900 8040 18100 8050
rect 18560 8040 18760 8050
rect 19220 8040 19420 8050
rect 20500 8040 20510 8050
rect 1010 7980 6910 8040
rect 7090 7980 7570 8040
rect 7750 7980 8230 8040
rect 8410 7980 9110 8040
rect 9290 7980 9770 8040
rect 9950 7980 10430 8040
rect 10610 7980 11310 8040
rect 11490 7980 11970 8040
rect 12150 7980 12630 8040
rect 12810 7980 13510 8040
rect 13690 7980 14170 8040
rect 14350 7980 14830 8040
rect 15010 7980 20510 8040
rect 1010 7970 1020 7980
rect 2500 7970 2700 7980
rect 3160 7970 3360 7980
rect 3820 7970 4020 7980
rect 4700 7970 4900 7980
rect 5360 7970 5560 7980
rect 6020 7970 6220 7980
rect 6900 7970 7100 7980
rect 7560 7970 7760 7980
rect 8220 7970 8420 7980
rect 9100 7970 9300 7980
rect 9760 7970 9960 7980
rect 10420 7970 10620 7980
rect 11300 7970 11500 7980
rect 11960 7970 12160 7980
rect 12620 7970 12820 7980
rect 13500 7970 13700 7980
rect 14160 7970 14360 7980
rect 14820 7970 15020 7980
rect 15700 7970 15900 7980
rect 16360 7970 16560 7980
rect 17020 7970 17220 7980
rect 17900 7970 18100 7980
rect 18560 7970 18760 7980
rect 19220 7970 19420 7980
rect 20500 7970 20510 7980
rect 20690 8040 20700 8050
rect 20690 7980 22180 8040
rect 20690 7970 20700 7980
rect 820 7960 1020 7970
rect 20500 7960 20700 7970
rect 1220 7910 1420 7920
rect 20900 7910 21100 7920
rect 1220 7900 1230 7910
rect -220 7840 1230 7900
rect 1220 7830 1230 7840
rect 1410 7900 1420 7910
rect 2500 7900 2700 7910
rect 3160 7900 3360 7910
rect 3820 7900 4020 7910
rect 4700 7900 4900 7910
rect 5360 7900 5560 7910
rect 6020 7900 6220 7910
rect 6900 7900 7100 7910
rect 7560 7900 7760 7910
rect 8220 7900 8420 7910
rect 9100 7900 9300 7910
rect 9760 7900 9960 7910
rect 10420 7900 10620 7910
rect 11300 7900 11500 7910
rect 11960 7900 12160 7910
rect 12620 7900 12820 7910
rect 13500 7900 13700 7910
rect 14160 7900 14360 7910
rect 14820 7900 15020 7910
rect 15700 7900 15900 7910
rect 16360 7900 16560 7910
rect 17020 7900 17220 7910
rect 17900 7900 18100 7910
rect 18560 7900 18760 7910
rect 19220 7900 19420 7910
rect 20900 7900 20910 7910
rect 1410 7840 2510 7900
rect 2690 7840 3170 7900
rect 3350 7840 3830 7900
rect 4010 7840 4710 7900
rect 4890 7840 5370 7900
rect 5550 7840 6030 7900
rect 6210 7840 15710 7900
rect 15890 7840 16370 7900
rect 16550 7840 17030 7900
rect 17210 7840 17910 7900
rect 18090 7840 18570 7900
rect 18750 7840 19230 7900
rect 19410 7840 20910 7900
rect 1410 7830 1420 7840
rect 2500 7830 2700 7840
rect 3160 7830 3360 7840
rect 3820 7830 4020 7840
rect 4700 7830 4900 7840
rect 5360 7830 5560 7840
rect 6020 7830 6220 7840
rect 6900 7830 7100 7840
rect 7560 7830 7760 7840
rect 8220 7830 8420 7840
rect 9100 7830 9300 7840
rect 9760 7830 9960 7840
rect 10420 7830 10620 7840
rect 11300 7830 11500 7840
rect 11960 7830 12160 7840
rect 12620 7830 12820 7840
rect 13500 7830 13700 7840
rect 14160 7830 14360 7840
rect 14820 7830 15020 7840
rect 15700 7830 15900 7840
rect 16360 7830 16560 7840
rect 17020 7830 17220 7840
rect 17900 7830 18100 7840
rect 18560 7830 18760 7840
rect 19220 7830 19420 7840
rect 20900 7830 20910 7840
rect 21090 7900 21100 7910
rect 21090 7840 22180 7900
rect 21090 7830 21100 7840
rect 1220 7820 1420 7830
rect 20900 7820 21100 7830
rect -110 7740 30 7760
rect -110 7490 -80 7740
rect 0 7490 30 7740
rect -110 7460 30 7490
rect 2090 7740 2230 7760
rect 2090 7490 2120 7740
rect 2200 7490 2230 7740
rect 2090 7460 2230 7490
rect 4290 7740 4430 7760
rect 4290 7490 4320 7740
rect 4400 7490 4430 7740
rect 4290 7460 4430 7490
rect 6490 7740 6630 7760
rect 6490 7490 6520 7740
rect 6600 7490 6630 7740
rect 6490 7460 6630 7490
rect 8690 7740 8830 7760
rect 8690 7490 8720 7740
rect 8800 7490 8830 7740
rect 8690 7460 8830 7490
rect 10890 7740 11030 7760
rect 10890 7490 10920 7740
rect 11000 7490 11030 7740
rect 10890 7460 11030 7490
rect 13090 7740 13230 7760
rect 13090 7490 13120 7740
rect 13200 7490 13230 7740
rect 13090 7460 13230 7490
rect 15290 7740 15430 7760
rect 15290 7490 15320 7740
rect 15400 7490 15430 7740
rect 15290 7460 15430 7490
rect 17490 7740 17630 7760
rect 17490 7490 17520 7740
rect 17600 7490 17630 7740
rect 17490 7460 17630 7490
rect 19690 7740 19830 7760
rect 19690 7490 19720 7740
rect 19800 7490 19830 7740
rect 19690 7460 19830 7490
rect 21890 7740 22030 7760
rect 21890 7490 21920 7740
rect 22000 7490 22030 7740
rect 21890 7460 22030 7490
rect 4700 7410 6220 7420
rect 420 7390 620 7400
rect 420 7310 430 7390
rect 610 7310 620 7390
rect 1620 7390 1820 7400
rect 1620 7380 1630 7390
rect 1600 7320 1630 7380
rect 420 7300 620 7310
rect 1620 7310 1630 7320
rect 1810 7380 1820 7390
rect 4700 7380 4710 7410
rect 1810 7350 4710 7380
rect 6210 7380 6220 7410
rect 6900 7410 8420 7420
rect 6900 7380 6910 7410
rect 6210 7350 6910 7380
rect 8410 7380 8420 7410
rect 9100 7410 10620 7420
rect 9100 7380 9110 7410
rect 8410 7350 9110 7380
rect 10610 7380 10620 7410
rect 11300 7410 12820 7420
rect 11300 7380 11310 7410
rect 10610 7350 11310 7380
rect 12810 7380 12820 7410
rect 13500 7410 15020 7420
rect 13500 7380 13510 7410
rect 12810 7350 13510 7380
rect 15010 7380 15020 7410
rect 15700 7410 17220 7420
rect 15700 7380 15710 7410
rect 15010 7350 15710 7380
rect 17210 7380 17220 7410
rect 20100 7390 20300 7400
rect 20100 7380 20110 7390
rect 17210 7350 20110 7380
rect 1810 7320 20110 7350
rect 1810 7310 1820 7320
rect 1620 7300 1820 7310
rect 20100 7310 20110 7320
rect 20290 7380 20300 7390
rect 21300 7390 21500 7400
rect 20290 7320 20320 7380
rect 20290 7310 20300 7320
rect 20100 7300 20300 7310
rect 21300 7310 21310 7390
rect 21490 7310 21500 7390
rect 21300 7300 21500 7310
rect 820 7250 1020 7260
rect 20500 7250 20700 7260
rect 820 7240 830 7250
rect -220 7180 830 7240
rect 820 7170 830 7180
rect 1010 7240 1020 7250
rect 2500 7240 2700 7250
rect 3160 7240 3360 7250
rect 3820 7240 4020 7250
rect 4700 7240 4900 7250
rect 5360 7240 5560 7250
rect 6020 7240 6220 7250
rect 6900 7240 7100 7250
rect 7560 7240 7760 7250
rect 8220 7240 8420 7250
rect 9100 7240 9300 7250
rect 9760 7240 9960 7250
rect 10420 7240 10620 7250
rect 11300 7240 11500 7250
rect 11960 7240 12160 7250
rect 12620 7240 12820 7250
rect 13500 7240 13700 7250
rect 14160 7240 14360 7250
rect 14820 7240 15020 7250
rect 15700 7240 15900 7250
rect 16360 7240 16560 7250
rect 17020 7240 17220 7250
rect 17900 7240 18100 7250
rect 18560 7240 18760 7250
rect 19220 7240 19420 7250
rect 20500 7240 20510 7250
rect 1010 7180 2510 7240
rect 2690 7180 3170 7240
rect 3350 7180 3830 7240
rect 4010 7180 4710 7240
rect 4890 7180 5370 7240
rect 5550 7180 6030 7240
rect 6210 7180 15710 7240
rect 15890 7180 16370 7240
rect 16550 7180 17030 7240
rect 17210 7180 17910 7240
rect 18090 7180 18570 7240
rect 18750 7180 19230 7240
rect 19410 7180 20510 7240
rect 1010 7170 1020 7180
rect 2500 7170 2700 7180
rect 3160 7170 3360 7180
rect 3820 7170 4020 7180
rect 4700 7170 4900 7180
rect 5360 7170 5560 7180
rect 6020 7170 6220 7180
rect 6900 7170 7100 7180
rect 7560 7170 7760 7180
rect 8220 7170 8420 7180
rect 9100 7170 9300 7180
rect 9760 7170 9960 7180
rect 10420 7170 10620 7180
rect 11300 7170 11500 7180
rect 11960 7170 12160 7180
rect 12620 7170 12820 7180
rect 13500 7170 13700 7180
rect 14160 7170 14360 7180
rect 14820 7170 15020 7180
rect 15700 7170 15900 7180
rect 16360 7170 16560 7180
rect 17020 7170 17220 7180
rect 17900 7170 18100 7180
rect 18560 7170 18760 7180
rect 19220 7170 19420 7180
rect 20500 7170 20510 7180
rect 20690 7240 20700 7250
rect 20690 7180 22180 7240
rect 20690 7170 20700 7180
rect 820 7160 1020 7170
rect 20500 7160 20700 7170
rect 1220 7110 1420 7120
rect 20900 7110 21100 7120
rect 1220 7100 1230 7110
rect -220 7040 1230 7100
rect 1220 7030 1230 7040
rect 1410 7100 1420 7110
rect 2500 7100 2700 7110
rect 3160 7100 3360 7110
rect 3820 7100 4020 7110
rect 4700 7100 4900 7110
rect 5360 7100 5560 7110
rect 6020 7100 6220 7110
rect 6900 7100 7100 7110
rect 7560 7100 7760 7110
rect 8220 7100 8420 7110
rect 9100 7100 9300 7110
rect 9760 7100 9960 7110
rect 10420 7100 10620 7110
rect 11300 7100 11500 7110
rect 11960 7100 12160 7110
rect 12620 7100 12820 7110
rect 13500 7100 13700 7110
rect 14160 7100 14360 7110
rect 14820 7100 15020 7110
rect 15700 7100 15900 7110
rect 16360 7100 16560 7110
rect 17020 7100 17220 7110
rect 17900 7100 18100 7110
rect 18560 7100 18760 7110
rect 19220 7100 19420 7110
rect 20900 7100 20910 7110
rect 1410 7040 6910 7100
rect 7090 7040 7570 7100
rect 7750 7040 8230 7100
rect 8410 7040 9110 7100
rect 9290 7040 9770 7100
rect 9950 7040 10430 7100
rect 10610 7040 11310 7100
rect 11490 7040 11970 7100
rect 12150 7040 12630 7100
rect 12810 7040 13510 7100
rect 13690 7040 14170 7100
rect 14350 7040 14830 7100
rect 15010 7040 20910 7100
rect 1410 7030 1420 7040
rect 2500 7030 2700 7040
rect 3160 7030 3360 7040
rect 3820 7030 4020 7040
rect 4700 7030 4900 7040
rect 5360 7030 5560 7040
rect 6020 7030 6220 7040
rect 6900 7030 7100 7040
rect 7560 7030 7760 7040
rect 8220 7030 8420 7040
rect 9100 7030 9300 7040
rect 9760 7030 9960 7040
rect 10420 7030 10620 7040
rect 11300 7030 11500 7040
rect 11960 7030 12160 7040
rect 12620 7030 12820 7040
rect 13500 7030 13700 7040
rect 14160 7030 14360 7040
rect 14820 7030 15020 7040
rect 15700 7030 15900 7040
rect 16360 7030 16560 7040
rect 17020 7030 17220 7040
rect 17900 7030 18100 7040
rect 18560 7030 18760 7040
rect 19220 7030 19420 7040
rect 20900 7030 20910 7040
rect 21090 7100 21100 7110
rect 21090 7040 22180 7100
rect 21090 7030 21100 7040
rect 1220 7020 1420 7030
rect 20900 7020 21100 7030
rect -110 6940 30 6960
rect -110 6690 -80 6940
rect 0 6690 30 6940
rect -110 6660 30 6690
rect 2090 6940 2230 6960
rect 2090 6690 2120 6940
rect 2200 6690 2230 6940
rect 2090 6660 2230 6690
rect 4290 6940 4430 6960
rect 4290 6690 4320 6940
rect 4400 6690 4430 6940
rect 4290 6660 4430 6690
rect 6490 6940 6630 6960
rect 6490 6690 6520 6940
rect 6600 6690 6630 6940
rect 6490 6660 6630 6690
rect 8690 6940 8830 6960
rect 8690 6690 8720 6940
rect 8800 6690 8830 6940
rect 8690 6660 8830 6690
rect 10890 6940 11030 6960
rect 10890 6690 10920 6940
rect 11000 6690 11030 6940
rect 10890 6660 11030 6690
rect 13090 6940 13230 6960
rect 13090 6690 13120 6940
rect 13200 6690 13230 6940
rect 13090 6660 13230 6690
rect 15290 6940 15430 6960
rect 15290 6690 15320 6940
rect 15400 6690 15430 6940
rect 15290 6660 15430 6690
rect 17490 6940 17630 6960
rect 17490 6690 17520 6940
rect 17600 6690 17630 6940
rect 17490 6660 17630 6690
rect 19690 6940 19830 6960
rect 19690 6690 19720 6940
rect 19800 6690 19830 6940
rect 19690 6660 19830 6690
rect 21890 6940 22030 6960
rect 21890 6690 21920 6940
rect 22000 6690 22030 6940
rect 21890 6660 22030 6690
rect 4700 6610 6220 6620
rect 420 6590 620 6600
rect 420 6510 430 6590
rect 610 6510 620 6590
rect 1620 6590 1820 6600
rect 1620 6580 1630 6590
rect 1600 6520 1630 6580
rect 420 6500 620 6510
rect 1620 6510 1630 6520
rect 1810 6580 1820 6590
rect 4700 6580 4710 6610
rect 1810 6550 4710 6580
rect 6210 6580 6220 6610
rect 6900 6610 8420 6620
rect 6900 6580 6910 6610
rect 6210 6550 6910 6580
rect 8410 6580 8420 6610
rect 9100 6610 10620 6620
rect 9100 6580 9110 6610
rect 8410 6550 9110 6580
rect 10610 6580 10620 6610
rect 11300 6610 12820 6620
rect 11300 6580 11310 6610
rect 10610 6550 11310 6580
rect 12810 6580 12820 6610
rect 13500 6610 15020 6620
rect 13500 6580 13510 6610
rect 12810 6550 13510 6580
rect 15010 6580 15020 6610
rect 15700 6610 17220 6620
rect 15700 6580 15710 6610
rect 15010 6550 15710 6580
rect 17210 6580 17220 6610
rect 20100 6590 20300 6600
rect 20100 6580 20110 6590
rect 17210 6550 20110 6580
rect 1810 6520 20110 6550
rect 1810 6510 1820 6520
rect 1620 6500 1820 6510
rect 20100 6510 20110 6520
rect 20290 6580 20300 6590
rect 21300 6590 21500 6600
rect 20290 6520 20320 6580
rect 20290 6510 20300 6520
rect 20100 6500 20300 6510
rect 21300 6510 21310 6590
rect 21490 6510 21500 6590
rect 21300 6500 21500 6510
rect 820 6450 1020 6460
rect 20500 6450 20700 6460
rect 820 6440 830 6450
rect -220 6380 830 6440
rect 820 6370 830 6380
rect 1010 6440 1020 6450
rect 2500 6440 2700 6450
rect 3160 6440 3360 6450
rect 3820 6440 4020 6450
rect 4700 6440 4900 6450
rect 5360 6440 5560 6450
rect 6020 6440 6220 6450
rect 6900 6440 7100 6450
rect 7560 6440 7760 6450
rect 8220 6440 8420 6450
rect 9100 6440 9300 6450
rect 9760 6440 9960 6450
rect 10420 6440 10620 6450
rect 11300 6440 11500 6450
rect 11960 6440 12160 6450
rect 12620 6440 12820 6450
rect 13500 6440 13700 6450
rect 14160 6440 14360 6450
rect 14820 6440 15020 6450
rect 15700 6440 15900 6450
rect 16360 6440 16560 6450
rect 17020 6440 17220 6450
rect 17900 6440 18100 6450
rect 18560 6440 18760 6450
rect 19220 6440 19420 6450
rect 20500 6440 20510 6450
rect 1010 6380 6910 6440
rect 7090 6380 7570 6440
rect 7750 6380 8230 6440
rect 8410 6380 9110 6440
rect 9290 6380 9770 6440
rect 9950 6380 10430 6440
rect 10610 6380 11310 6440
rect 11490 6380 11970 6440
rect 12150 6380 12630 6440
rect 12810 6380 13510 6440
rect 13690 6380 14170 6440
rect 14350 6380 14830 6440
rect 15010 6380 20510 6440
rect 1010 6370 1020 6380
rect 2500 6370 2700 6380
rect 3160 6370 3360 6380
rect 3820 6370 4020 6380
rect 4700 6370 4900 6380
rect 5360 6370 5560 6380
rect 6020 6370 6220 6380
rect 6900 6370 7100 6380
rect 7560 6370 7760 6380
rect 8220 6370 8420 6380
rect 9100 6370 9300 6380
rect 9760 6370 9960 6380
rect 10420 6370 10620 6380
rect 11300 6370 11500 6380
rect 11960 6370 12160 6380
rect 12620 6370 12820 6380
rect 13500 6370 13700 6380
rect 14160 6370 14360 6380
rect 14820 6370 15020 6380
rect 15700 6370 15900 6380
rect 16360 6370 16560 6380
rect 17020 6370 17220 6380
rect 17900 6370 18100 6380
rect 18560 6370 18760 6380
rect 19220 6370 19420 6380
rect 20500 6370 20510 6380
rect 20690 6440 20700 6450
rect 20690 6380 22180 6440
rect 20690 6370 20700 6380
rect 820 6360 1020 6370
rect 20500 6360 20700 6370
rect 1220 6310 1420 6320
rect 20900 6310 21100 6320
rect 1220 6300 1230 6310
rect -220 6240 1230 6300
rect 1220 6230 1230 6240
rect 1410 6300 1420 6310
rect 2500 6300 2700 6310
rect 3160 6300 3360 6310
rect 3820 6300 4020 6310
rect 4700 6300 4900 6310
rect 5360 6300 5560 6310
rect 6020 6300 6220 6310
rect 6900 6300 7100 6310
rect 7560 6300 7760 6310
rect 8220 6300 8420 6310
rect 9100 6300 9300 6310
rect 9760 6300 9960 6310
rect 10420 6300 10620 6310
rect 11300 6300 11500 6310
rect 11960 6300 12160 6310
rect 12620 6300 12820 6310
rect 13500 6300 13700 6310
rect 14160 6300 14360 6310
rect 14820 6300 15020 6310
rect 15700 6300 15900 6310
rect 16360 6300 16560 6310
rect 17020 6300 17220 6310
rect 17900 6300 18100 6310
rect 18560 6300 18760 6310
rect 19220 6300 19420 6310
rect 20900 6300 20910 6310
rect 1410 6240 2510 6300
rect 2690 6240 3170 6300
rect 3350 6240 3830 6300
rect 4010 6240 4710 6300
rect 4890 6240 5370 6300
rect 5550 6240 6030 6300
rect 6210 6240 15710 6300
rect 15890 6240 16370 6300
rect 16550 6240 17030 6300
rect 17210 6240 17910 6300
rect 18090 6240 18570 6300
rect 18750 6240 19230 6300
rect 19410 6240 20910 6300
rect 1410 6230 1420 6240
rect 2500 6230 2700 6240
rect 3160 6230 3360 6240
rect 3820 6230 4020 6240
rect 4700 6230 4900 6240
rect 5360 6230 5560 6240
rect 6020 6230 6220 6240
rect 6900 6230 7100 6240
rect 7560 6230 7760 6240
rect 8220 6230 8420 6240
rect 9100 6230 9300 6240
rect 9760 6230 9960 6240
rect 10420 6230 10620 6240
rect 11300 6230 11500 6240
rect 11960 6230 12160 6240
rect 12620 6230 12820 6240
rect 13500 6230 13700 6240
rect 14160 6230 14360 6240
rect 14820 6230 15020 6240
rect 15700 6230 15900 6240
rect 16360 6230 16560 6240
rect 17020 6230 17220 6240
rect 17900 6230 18100 6240
rect 18560 6230 18760 6240
rect 19220 6230 19420 6240
rect 20900 6230 20910 6240
rect 21090 6300 21100 6310
rect 21090 6240 22180 6300
rect 21090 6230 21100 6240
rect 1220 6220 1420 6230
rect 20900 6220 21100 6230
rect -110 6140 30 6160
rect -110 5890 -80 6140
rect 0 5890 30 6140
rect -110 5860 30 5890
rect 2090 6140 2230 6160
rect 2090 5890 2120 6140
rect 2200 5890 2230 6140
rect 2090 5860 2230 5890
rect 4290 6140 4430 6160
rect 4290 5890 4320 6140
rect 4400 5890 4430 6140
rect 4290 5860 4430 5890
rect 6490 6140 6630 6160
rect 6490 5890 6520 6140
rect 6600 5890 6630 6140
rect 6490 5860 6630 5890
rect 8690 6140 8830 6160
rect 8690 5890 8720 6140
rect 8800 5890 8830 6140
rect 8690 5860 8830 5890
rect 10890 6140 11030 6160
rect 10890 5890 10920 6140
rect 11000 5890 11030 6140
rect 10890 5860 11030 5890
rect 13090 6140 13230 6160
rect 13090 5890 13120 6140
rect 13200 5890 13230 6140
rect 13090 5860 13230 5890
rect 15290 6140 15430 6160
rect 15290 5890 15320 6140
rect 15400 5890 15430 6140
rect 15290 5860 15430 5890
rect 17490 6140 17630 6160
rect 17490 5890 17520 6140
rect 17600 5890 17630 6140
rect 17490 5860 17630 5890
rect 19690 6140 19830 6160
rect 19690 5890 19720 6140
rect 19800 5890 19830 6140
rect 19690 5860 19830 5890
rect 21890 6140 22030 6160
rect 21890 5890 21920 6140
rect 22000 5890 22030 6140
rect 21890 5860 22030 5890
rect 2500 5810 4020 5820
rect 1620 5790 1820 5800
rect 1620 5780 1630 5790
rect 1600 5720 1630 5780
rect 1620 5710 1630 5720
rect 1810 5780 1820 5790
rect 2500 5780 2510 5810
rect 1810 5750 2510 5780
rect 4010 5780 4020 5810
rect 4700 5810 6220 5820
rect 4700 5780 4710 5810
rect 4010 5750 4710 5780
rect 6210 5780 6220 5810
rect 6900 5810 8420 5820
rect 6900 5780 6910 5810
rect 6210 5750 6910 5780
rect 8410 5780 8420 5810
rect 9100 5810 10620 5820
rect 9100 5780 9110 5810
rect 8410 5750 9110 5780
rect 10610 5780 10620 5810
rect 11300 5810 12820 5820
rect 11300 5780 11310 5810
rect 10610 5750 11310 5780
rect 12810 5780 12820 5810
rect 13500 5810 15020 5820
rect 13500 5780 13510 5810
rect 12810 5750 13510 5780
rect 15010 5780 15020 5810
rect 15700 5810 17220 5820
rect 15700 5780 15710 5810
rect 15010 5750 15710 5780
rect 17210 5780 17220 5810
rect 17900 5810 19420 5820
rect 17900 5780 17910 5810
rect 17210 5750 17910 5780
rect 19410 5780 19420 5810
rect 20100 5790 20300 5800
rect 20100 5780 20110 5790
rect 19410 5750 20110 5780
rect 1810 5720 20110 5750
rect 1810 5710 1820 5720
rect 1620 5700 1820 5710
rect 20100 5710 20110 5720
rect 20290 5780 20300 5790
rect 20290 5720 20320 5780
rect 20290 5710 20300 5720
rect 20100 5700 20300 5710
rect 820 5650 1020 5660
rect 20500 5650 20700 5660
rect 820 5640 830 5650
rect -220 5580 830 5640
rect 820 5570 830 5580
rect 1010 5640 1020 5650
rect 2500 5640 2700 5650
rect 3160 5640 3360 5650
rect 3820 5640 4020 5650
rect 4700 5640 4900 5650
rect 5360 5640 5560 5650
rect 6020 5640 6220 5650
rect 6900 5640 7100 5650
rect 7560 5640 7760 5650
rect 8220 5640 8420 5650
rect 9100 5640 9300 5650
rect 9760 5640 9960 5650
rect 10420 5640 10620 5650
rect 11300 5640 11500 5650
rect 11960 5640 12160 5650
rect 12620 5640 12820 5650
rect 13500 5640 13700 5650
rect 14160 5640 14360 5650
rect 14820 5640 15020 5650
rect 15700 5640 15900 5650
rect 16360 5640 16560 5650
rect 17020 5640 17220 5650
rect 17900 5640 18100 5650
rect 18560 5640 18760 5650
rect 19220 5640 19420 5650
rect 20500 5640 20510 5650
rect 1010 5580 2510 5640
rect 2690 5580 3170 5640
rect 3350 5580 3830 5640
rect 4010 5580 4710 5640
rect 4890 5580 5370 5640
rect 5550 5580 6030 5640
rect 6210 5580 15710 5640
rect 15890 5580 16370 5640
rect 16550 5580 17030 5640
rect 17210 5580 17910 5640
rect 18090 5580 18570 5640
rect 18750 5580 19230 5640
rect 19410 5580 20510 5640
rect 1010 5570 1020 5580
rect 2500 5570 2700 5580
rect 3160 5570 3360 5580
rect 3820 5570 4020 5580
rect 4700 5570 4900 5580
rect 5360 5570 5560 5580
rect 6020 5570 6220 5580
rect 6900 5570 7100 5580
rect 7560 5570 7760 5580
rect 8220 5570 8420 5580
rect 9100 5570 9300 5580
rect 9760 5570 9960 5580
rect 10420 5570 10620 5580
rect 11300 5570 11500 5580
rect 11960 5570 12160 5580
rect 12620 5570 12820 5580
rect 13500 5570 13700 5580
rect 14160 5570 14360 5580
rect 14820 5570 15020 5580
rect 15700 5570 15900 5580
rect 16360 5570 16560 5580
rect 17020 5570 17220 5580
rect 17900 5570 18100 5580
rect 18560 5570 18760 5580
rect 19220 5570 19420 5580
rect 20500 5570 20510 5580
rect 20690 5640 20700 5650
rect 20690 5580 22180 5640
rect 20690 5570 20700 5580
rect 820 5560 1020 5570
rect 20500 5560 20700 5570
rect 1220 5510 1420 5520
rect 20900 5510 21100 5520
rect 1220 5500 1230 5510
rect -220 5440 1230 5500
rect 1220 5430 1230 5440
rect 1410 5500 1420 5510
rect 2500 5500 2700 5510
rect 3160 5500 3360 5510
rect 3820 5500 4020 5510
rect 4700 5500 4900 5510
rect 5360 5500 5560 5510
rect 6020 5500 6220 5510
rect 6900 5500 7100 5510
rect 7560 5500 7760 5510
rect 8220 5500 8420 5510
rect 9100 5500 9300 5510
rect 9760 5500 9960 5510
rect 10420 5500 10620 5510
rect 11300 5500 11500 5510
rect 11960 5500 12160 5510
rect 12620 5500 12820 5510
rect 13500 5500 13700 5510
rect 14160 5500 14360 5510
rect 14820 5500 15020 5510
rect 15700 5500 15900 5510
rect 16360 5500 16560 5510
rect 17020 5500 17220 5510
rect 17900 5500 18100 5510
rect 18560 5500 18760 5510
rect 19220 5500 19420 5510
rect 20900 5500 20910 5510
rect 1410 5440 6910 5500
rect 7090 5440 7570 5500
rect 7750 5440 8230 5500
rect 8410 5440 9110 5500
rect 9290 5440 9770 5500
rect 9950 5440 10430 5500
rect 10610 5440 11310 5500
rect 11490 5440 11970 5500
rect 12150 5440 12630 5500
rect 12810 5440 13510 5500
rect 13690 5440 14170 5500
rect 14350 5440 14830 5500
rect 15010 5440 20910 5500
rect 1410 5430 1420 5440
rect 2500 5430 2700 5440
rect 3160 5430 3360 5440
rect 3820 5430 4020 5440
rect 4700 5430 4900 5440
rect 5360 5430 5560 5440
rect 6020 5430 6220 5440
rect 6900 5430 7100 5440
rect 7560 5430 7760 5440
rect 8220 5430 8420 5440
rect 9100 5430 9300 5440
rect 9760 5430 9960 5440
rect 10420 5430 10620 5440
rect 11300 5430 11500 5440
rect 11960 5430 12160 5440
rect 12620 5430 12820 5440
rect 13500 5430 13700 5440
rect 14160 5430 14360 5440
rect 14820 5430 15020 5440
rect 15700 5430 15900 5440
rect 16360 5430 16560 5440
rect 17020 5430 17220 5440
rect 17900 5430 18100 5440
rect 18560 5430 18760 5440
rect 19220 5430 19420 5440
rect 20900 5430 20910 5440
rect 21090 5500 21100 5510
rect 21090 5440 22180 5500
rect 21090 5430 21100 5440
rect 1220 5420 1420 5430
rect 20900 5420 21100 5430
rect -110 5340 30 5360
rect -110 5090 -80 5340
rect 0 5090 30 5340
rect -110 5060 30 5090
rect 2090 5340 2230 5360
rect 2090 5090 2120 5340
rect 2200 5090 2230 5340
rect 2090 5060 2230 5090
rect 4290 5340 4430 5360
rect 4290 5090 4320 5340
rect 4400 5090 4430 5340
rect 4290 5060 4430 5090
rect 6490 5340 6630 5360
rect 6490 5090 6520 5340
rect 6600 5090 6630 5340
rect 6490 5060 6630 5090
rect 8690 5340 8830 5360
rect 8690 5090 8720 5340
rect 8800 5090 8830 5340
rect 8690 5060 8830 5090
rect 10890 5340 11030 5360
rect 10890 5090 10920 5340
rect 11000 5090 11030 5340
rect 10890 5060 11030 5090
rect 13090 5340 13230 5360
rect 13090 5090 13120 5340
rect 13200 5090 13230 5340
rect 13090 5060 13230 5090
rect 15290 5340 15430 5360
rect 15290 5090 15320 5340
rect 15400 5090 15430 5340
rect 15290 5060 15430 5090
rect 17490 5340 17630 5360
rect 17490 5090 17520 5340
rect 17600 5090 17630 5340
rect 17490 5060 17630 5090
rect 19690 5340 19830 5360
rect 19690 5090 19720 5340
rect 19800 5090 19830 5340
rect 19690 5060 19830 5090
rect 21890 5340 22030 5360
rect 21890 5090 21920 5340
rect 22000 5090 22030 5340
rect 21890 5060 22030 5090
rect 2500 5010 4020 5020
rect 1620 4990 1820 5000
rect 1620 4980 1630 4990
rect 1600 4920 1630 4980
rect 1620 4910 1630 4920
rect 1810 4980 1820 4990
rect 2500 4980 2510 5010
rect 1810 4950 2510 4980
rect 4010 4980 4020 5010
rect 4700 5010 6220 5020
rect 4700 4980 4710 5010
rect 4010 4950 4710 4980
rect 6210 4980 6220 5010
rect 6900 5010 8420 5020
rect 6900 4980 6910 5010
rect 6210 4950 6910 4980
rect 8410 4980 8420 5010
rect 9100 5010 10620 5020
rect 9100 4980 9110 5010
rect 8410 4950 9110 4980
rect 10610 4980 10620 5010
rect 11300 5010 12820 5020
rect 11300 4980 11310 5010
rect 10610 4950 11310 4980
rect 12810 4980 12820 5010
rect 13500 5010 15020 5020
rect 13500 4980 13510 5010
rect 12810 4950 13510 4980
rect 15010 4980 15020 5010
rect 15700 5010 17220 5020
rect 15700 4980 15710 5010
rect 15010 4950 15710 4980
rect 17210 4980 17220 5010
rect 17900 5010 19420 5020
rect 17900 4980 17910 5010
rect 17210 4950 17910 4980
rect 19410 4980 19420 5010
rect 20100 4990 20300 5000
rect 20100 4980 20110 4990
rect 19410 4950 20110 4980
rect 1810 4920 20110 4950
rect 1810 4910 1820 4920
rect 1620 4900 1820 4910
rect 20100 4910 20110 4920
rect 20290 4980 20300 4990
rect 20290 4920 20320 4980
rect 20290 4910 20300 4920
rect 20100 4900 20300 4910
rect -300 4340 32680 4540
rect -300 3940 32680 4140
rect -300 3730 31740 3740
rect -300 3550 430 3730
rect 610 3550 21310 3730
rect 21490 3550 31570 3730
rect 31730 3550 31740 3730
rect -300 3540 31740 3550
rect 1160 3330 20300 3340
rect 1160 3150 1170 3330
rect 1330 3150 1630 3330
rect 1810 3150 2770 3330
rect 2930 3150 4370 3330
rect 4530 3150 5970 3330
rect 6130 3150 7570 3330
rect 7730 3150 9170 3330
rect 9330 3150 20110 3330
rect 20290 3150 20300 3330
rect 1160 3140 20300 3150
rect 34890 2760 35060 2770
rect 11690 2750 11850 2760
rect 11690 2600 11700 2750
rect 11840 2740 11850 2750
rect 34890 2740 34900 2760
rect 11840 2610 34900 2740
rect 11840 2600 11850 2610
rect 11690 2590 11850 2600
rect 34890 2600 34900 2610
rect 35050 2600 35060 2760
rect 34890 2590 35060 2600
rect 33290 2530 33460 2540
rect 10990 2520 11150 2530
rect 10990 2380 11000 2520
rect 11140 2510 11150 2520
rect 12590 2520 12750 2530
rect 12590 2510 12600 2520
rect 11140 2380 12600 2510
rect 12740 2510 12750 2520
rect 13970 2520 14130 2530
rect 13970 2510 13980 2520
rect 12740 2380 13980 2510
rect 14120 2380 14130 2520
rect 33290 2510 33300 2530
rect 10990 2370 11150 2380
rect 12590 2370 12750 2380
rect 13970 2370 14130 2380
rect 14900 2380 33300 2510
rect 2090 2230 13440 2240
rect 2090 2070 2110 2230
rect 2230 2070 3710 2230
rect 3830 2070 5310 2230
rect 5430 2070 6910 2230
rect 7030 2070 8510 2230
rect 8630 2070 10110 2230
rect 10230 2070 11710 2230
rect 11830 2070 13310 2230
rect 13430 2070 13440 2230
rect 2090 2060 13440 2070
rect 14900 1960 15040 2380
rect 33290 2370 33300 2380
rect 33450 2370 33460 2530
rect 33290 2360 33460 2370
rect 16500 2230 26240 2240
rect 16500 2070 16510 2230
rect 16630 2070 18110 2230
rect 18230 2070 19710 2230
rect 19830 2070 21310 2230
rect 21430 2070 22910 2230
rect 23030 2070 24510 2230
rect 24630 2070 26110 2230
rect 26230 2070 26240 2230
rect 16500 2060 26240 2070
rect 27700 2230 31040 2240
rect 27700 2050 27710 2230
rect 27830 2050 29310 2230
rect 29430 2050 30910 2230
rect 31030 2050 31040 2230
rect 27700 2040 31040 2050
rect 14900 1300 14910 1960
rect 15030 1300 15040 1960
rect 14900 1270 15040 1300
rect 32500 1130 32640 1140
rect 34100 1130 34240 1140
rect 34900 1130 35050 1140
rect 35700 1130 35840 1140
rect 32500 1010 32510 1130
rect 32630 1010 34110 1130
rect 34230 1010 34910 1130
rect 35040 1010 35710 1130
rect 35830 1010 35840 1130
rect 32500 1000 32640 1010
rect 34100 1000 34240 1010
rect 34900 1000 35050 1010
rect 35700 1000 35840 1010
rect 2090 430 13440 440
rect 2090 270 2110 430
rect 2230 270 3710 430
rect 3830 270 5310 430
rect 5430 270 6910 430
rect 7030 270 8510 430
rect 8630 270 10110 430
rect 10230 270 11710 430
rect 11830 270 13310 430
rect 13430 270 13440 430
rect 2090 260 13440 270
rect 16500 430 26240 440
rect 16500 270 16510 430
rect 16630 270 18110 430
rect 18230 270 19710 430
rect 19830 270 21310 430
rect 21430 270 22910 430
rect 23030 270 24510 430
rect 24630 270 26110 430
rect 26230 270 26240 430
rect 16500 260 26240 270
rect 27700 430 31040 440
rect 27700 250 27710 430
rect 27830 250 29310 430
rect 29430 250 30910 430
rect 31030 250 31040 430
rect 27700 240 31040 250
rect 32500 420 35840 430
rect 32500 260 33300 420
rect 33450 260 35840 420
rect 32500 250 35840 260
rect 32500 170 32640 250
rect 32500 -510 32510 170
rect 32630 -510 32640 170
rect 32500 -520 32640 -510
rect 34100 170 34240 250
rect 34100 -510 34110 170
rect 34230 -510 34240 170
rect 34100 -520 34240 -510
rect 35700 170 35840 250
rect 35700 -510 35710 170
rect 35830 -510 35840 170
rect 35700 -520 35840 -510
rect 2090 -1370 15040 -1360
rect 2090 -1530 2110 -1370
rect 2230 -1530 3710 -1370
rect 3830 -1530 5310 -1370
rect 5430 -1530 6910 -1370
rect 7030 -1530 8510 -1370
rect 8630 -1530 10110 -1370
rect 10230 -1530 11710 -1370
rect 11830 -1530 13310 -1370
rect 13430 -1530 14910 -1370
rect 15030 -1530 15040 -1370
rect 2090 -1540 15040 -1530
rect 15240 -1370 26270 -1360
rect 15240 -1530 15250 -1370
rect 15370 -1530 16510 -1370
rect 16630 -1530 18110 -1370
rect 18230 -1530 19710 -1370
rect 19830 -1530 21310 -1370
rect 21430 -1530 22910 -1370
rect 23030 -1530 24510 -1370
rect 24630 -1530 26110 -1370
rect 26230 -1530 26270 -1370
rect 15240 -1540 26270 -1530
rect 27700 -1370 31040 -1360
rect 27700 -1550 27710 -1370
rect 27830 -1550 29310 -1370
rect 29430 -1550 30910 -1370
rect 31030 -1550 31040 -1370
rect 27700 -1560 31040 -1550
rect 32500 -2470 32640 -2460
rect 34100 -2470 34240 -2460
rect 34900 -2470 35050 -2460
rect 35700 -2470 35840 -2460
rect 32500 -2590 32510 -2470
rect 32630 -2590 34110 -2470
rect 34230 -2590 34910 -2470
rect 35040 -2590 35710 -2470
rect 35830 -2590 35840 -2470
rect 32500 -2600 32640 -2590
rect 34100 -2600 34240 -2590
rect 34900 -2600 35050 -2590
rect 35700 -2600 35840 -2590
rect 2090 -3170 15040 -3160
rect 2090 -3330 2110 -3170
rect 2230 -3330 3710 -3170
rect 3830 -3330 5310 -3170
rect 5430 -3330 6910 -3170
rect 7030 -3330 8510 -3170
rect 8630 -3330 10110 -3170
rect 10230 -3330 11710 -3170
rect 11830 -3330 13310 -3170
rect 13430 -3330 14910 -3170
rect 15030 -3330 15040 -3170
rect 2090 -3340 15040 -3330
rect 16500 -3170 26240 -3160
rect 16500 -3330 16510 -3170
rect 16630 -3330 18110 -3170
rect 18230 -3330 19710 -3170
rect 19830 -3330 21310 -3170
rect 21430 -3330 22910 -3170
rect 23030 -3330 24510 -3170
rect 24630 -3330 26110 -3170
rect 26230 -3330 26240 -3170
rect 16500 -3340 26240 -3330
rect 27700 -3170 31040 -3160
rect 27700 -3350 27710 -3170
rect 27830 -3350 29310 -3170
rect 29430 -3350 30910 -3170
rect 31030 -3350 31040 -3170
rect 27700 -3360 31040 -3350
rect -20 -5170 37760 -5160
rect -20 -5350 1630 -5170
rect 1810 -5350 15570 -5170
rect 15730 -5350 18770 -5170
rect 18930 -5350 20910 -5170
rect 21090 -5350 21970 -5170
rect 22130 -5350 25170 -5170
rect 25330 -5350 28370 -5170
rect 28530 -5350 37760 -5170
rect -20 -5360 37760 -5350
rect -20 -5570 37760 -5560
rect -20 -5750 830 -5570
rect 1010 -5750 15570 -5570
rect 15730 -5750 18770 -5570
rect 18930 -5750 20510 -5570
rect 20690 -5750 21970 -5570
rect 22130 -5750 25170 -5570
rect 25330 -5750 28370 -5570
rect 28530 -5750 37760 -5570
rect -20 -5760 37760 -5750
rect -20 -5970 37760 -5960
rect -20 -6150 15790 -5970
rect 15950 -6150 18990 -5970
rect 19150 -6150 22190 -5970
rect 22350 -6150 25390 -5970
rect 25550 -6150 27690 -5970
rect 27850 -6150 28590 -5970
rect 28750 -6150 29290 -5970
rect 29450 -6150 30890 -5970
rect 31050 -6150 37760 -5970
rect -20 -6160 37760 -6150
rect 14900 -6490 15040 -6480
rect 14900 -6610 14910 -6490
rect 15030 -6610 15040 -6490
rect 14900 -6620 15040 -6610
rect -20 -6770 37760 -6760
rect -20 -6950 17390 -6770
rect 17550 -6950 20590 -6770
rect 20750 -6950 23790 -6770
rect 23950 -6950 26990 -6770
rect 27150 -6950 30190 -6770
rect 30350 -6950 37760 -6770
rect -20 -6960 37760 -6950
rect -20 -7170 37760 -7160
rect -20 -7350 830 -7170
rect 1010 -7350 17170 -7170
rect 17330 -7350 20370 -7170
rect 20690 -7350 23570 -7170
rect 23730 -7350 26770 -7170
rect 26930 -7350 29970 -7170
rect 30130 -7350 37760 -7170
rect -20 -7360 37760 -7350
rect -20 -7570 37760 -7560
rect -20 -7750 1230 -7570
rect 1410 -7750 17170 -7570
rect 17330 -7750 20370 -7570
rect 20530 -7750 22070 -7570
rect 22250 -7750 23570 -7570
rect 23730 -7750 26770 -7570
rect 26930 -7750 29970 -7570
rect 30130 -7750 37760 -7570
rect -20 -7760 37760 -7750
rect 16500 -9570 26250 -9560
rect 2120 -9590 10240 -9580
rect 2120 -9750 2130 -9590
rect 2230 -9750 3730 -9590
rect 3830 -9750 5330 -9590
rect 5430 -9750 6930 -9590
rect 7030 -9750 8530 -9590
rect 8630 -9750 10130 -9590
rect 10230 -9750 10240 -9590
rect 16500 -9730 16510 -9570
rect 16640 -9730 18110 -9570
rect 18240 -9730 19710 -9570
rect 19840 -9730 21310 -9570
rect 21440 -9730 22910 -9570
rect 23040 -9730 24510 -9570
rect 24640 -9730 26110 -9570
rect 26240 -9730 26250 -9570
rect 16500 -9740 26250 -9730
rect 27700 -9570 31050 -9560
rect 27700 -9730 27710 -9570
rect 27840 -9730 29310 -9570
rect 29440 -9730 30910 -9570
rect 31040 -9730 31050 -9570
rect 27700 -9740 31050 -9730
rect 2120 -9760 10240 -9750
rect 16500 -11370 26250 -11360
rect 2120 -11390 10240 -11380
rect 2120 -11550 2130 -11390
rect 2230 -11550 3730 -11390
rect 3830 -11550 5330 -11390
rect 5430 -11550 6930 -11390
rect 7030 -11550 8530 -11390
rect 8630 -11550 10130 -11390
rect 10230 -11550 10240 -11390
rect 16500 -11530 16510 -11370
rect 16640 -11530 18110 -11370
rect 18240 -11530 19710 -11370
rect 19840 -11530 21310 -11370
rect 21440 -11530 22910 -11370
rect 23040 -11530 24510 -11370
rect 24640 -11530 26110 -11370
rect 26240 -11530 26250 -11370
rect 16500 -11540 26250 -11530
rect 27700 -11370 31050 -11360
rect 27700 -11530 27710 -11370
rect 27840 -11530 29310 -11370
rect 29440 -11530 30910 -11370
rect 31040 -11530 31050 -11370
rect 27700 -11540 31050 -11530
rect 2120 -11560 10240 -11550
rect 13280 -13170 26250 -13160
rect 2120 -13190 10240 -13180
rect 2120 -13350 2130 -13190
rect 2230 -13350 3730 -13190
rect 3830 -13350 5330 -13190
rect 5430 -13350 6930 -13190
rect 7030 -13350 8530 -13190
rect 8630 -13350 10130 -13190
rect 10230 -13350 10240 -13190
rect 2120 -13360 10240 -13350
rect 13280 -13330 13290 -13170
rect 13460 -13330 14890 -13170
rect 15060 -13330 16510 -13170
rect 16640 -13330 18110 -13170
rect 18240 -13330 19710 -13170
rect 19840 -13330 21310 -13170
rect 21440 -13330 22910 -13170
rect 23040 -13330 24510 -13170
rect 24640 -13330 26110 -13170
rect 26240 -13330 26250 -13170
rect 13280 -13340 26250 -13330
rect 27700 -13170 31050 -13160
rect 27700 -13330 27710 -13170
rect 27840 -13330 29310 -13170
rect 29440 -13330 30910 -13170
rect 31040 -13330 31050 -13170
rect 27700 -13340 31050 -13330
rect 13280 -13360 15070 -13340
rect 13280 -14970 26250 -14960
rect 2120 -14990 10240 -14980
rect 2120 -15150 2130 -14990
rect 2230 -15150 3730 -14990
rect 3830 -15150 5330 -14990
rect 5430 -15150 6930 -14990
rect 7030 -15150 8530 -14990
rect 8630 -15150 10130 -14990
rect 10230 -15150 10240 -14990
rect 2120 -15160 10240 -15150
rect 13280 -15130 13290 -14970
rect 13460 -15130 14890 -14970
rect 15060 -15130 16510 -14970
rect 16640 -15130 18110 -14970
rect 18240 -15130 19710 -14970
rect 19840 -15130 21310 -14970
rect 21440 -15130 22910 -14970
rect 23040 -15130 24510 -14970
rect 24640 -15130 26110 -14970
rect 26240 -15130 26250 -14970
rect 13280 -15140 26250 -15130
rect 27700 -14970 31050 -14960
rect 27700 -15130 27710 -14970
rect 27840 -15130 29310 -14970
rect 29440 -15130 30910 -14970
rect 31040 -15130 31050 -14970
rect 27700 -15140 31050 -15130
rect 13280 -15160 15070 -15140
rect 16500 -16770 26250 -16760
rect 2120 -16790 15090 -16780
rect 2120 -16950 2130 -16790
rect 2230 -16950 3730 -16790
rect 3830 -16950 5330 -16790
rect 5430 -16950 6930 -16790
rect 7030 -16950 8530 -16790
rect 8630 -16950 10130 -16790
rect 10230 -16950 13300 -16790
rect 13450 -16950 14900 -16790
rect 15050 -16950 15090 -16790
rect 16500 -16930 16510 -16770
rect 16640 -16930 18110 -16770
rect 18240 -16930 19710 -16770
rect 19840 -16930 21310 -16770
rect 21440 -16930 22910 -16770
rect 23040 -16930 24510 -16770
rect 24640 -16930 26110 -16770
rect 26240 -16930 26250 -16770
rect 16500 -16940 26250 -16930
rect 27700 -16770 31050 -16760
rect 27700 -16930 27710 -16770
rect 27840 -16930 29310 -16770
rect 29440 -16930 30910 -16770
rect 31040 -16930 31050 -16770
rect 27700 -16940 31050 -16930
rect 2120 -16960 15090 -16950
rect 16500 -18570 26250 -18560
rect 2120 -18590 15060 -18580
rect 2120 -18750 2130 -18590
rect 2230 -18750 3730 -18590
rect 3830 -18750 5330 -18590
rect 5430 -18750 6930 -18590
rect 7030 -18750 8530 -18590
rect 8630 -18750 10130 -18590
rect 10230 -18750 13300 -18590
rect 13450 -18750 14900 -18590
rect 15050 -18750 15060 -18590
rect 16500 -18730 16510 -18570
rect 16640 -18730 18110 -18570
rect 18240 -18730 19710 -18570
rect 19840 -18730 21310 -18570
rect 21440 -18730 22910 -18570
rect 23040 -18730 24510 -18570
rect 24640 -18730 26110 -18570
rect 26240 -18730 26250 -18570
rect 16500 -18740 26250 -18730
rect 27700 -18570 31050 -18560
rect 27700 -18730 27710 -18570
rect 27840 -18730 29310 -18570
rect 29440 -18730 30910 -18570
rect 31040 -18730 31050 -18570
rect 27700 -18740 31050 -18730
rect 2120 -18760 15060 -18750
rect 16500 -20370 26250 -20360
rect 2120 -20390 10240 -20380
rect 2120 -20550 2130 -20390
rect 2230 -20550 3730 -20390
rect 3830 -20550 5330 -20390
rect 5430 -20550 6930 -20390
rect 7030 -20550 8530 -20390
rect 8630 -20550 10130 -20390
rect 10230 -20550 10240 -20390
rect 16500 -20530 16510 -20370
rect 16640 -20530 18110 -20370
rect 18240 -20530 19710 -20370
rect 19840 -20530 21310 -20370
rect 21440 -20530 22910 -20370
rect 23040 -20530 24510 -20370
rect 24640 -20530 26110 -20370
rect 26240 -20530 26250 -20370
rect 16500 -20540 26250 -20530
rect 27700 -20370 31050 -20360
rect 27700 -20530 27710 -20370
rect 27840 -20530 29310 -20370
rect 29440 -20530 30910 -20370
rect 31040 -20530 31050 -20370
rect 27700 -20540 31050 -20530
rect 2120 -20560 10240 -20550
rect 16500 -22170 26250 -22160
rect 2120 -22190 10240 -22180
rect 2120 -22350 2130 -22190
rect 2230 -22350 3730 -22190
rect 3830 -22350 5330 -22190
rect 5430 -22350 6930 -22190
rect 7030 -22350 8530 -22190
rect 8630 -22350 10130 -22190
rect 10230 -22350 10240 -22190
rect 16500 -22330 16510 -22170
rect 16640 -22330 18110 -22170
rect 18240 -22330 19710 -22170
rect 19840 -22330 21310 -22170
rect 21440 -22330 22910 -22170
rect 23040 -22330 24510 -22170
rect 24640 -22330 26110 -22170
rect 26240 -22330 26250 -22170
rect 16500 -22340 26250 -22330
rect 27700 -22170 31050 -22160
rect 27700 -22330 27710 -22170
rect 27840 -22330 29310 -22170
rect 29440 -22330 30910 -22170
rect 31040 -22330 31050 -22170
rect 27700 -22340 31050 -22330
rect 2120 -22360 10240 -22350
rect 11040 -22740 31040 -22730
rect 11040 -22850 11050 -22740
rect 11150 -22850 27720 -22740
rect 27830 -22850 29320 -22740
rect 29430 -22850 30920 -22740
rect 31030 -22850 31040 -22740
rect 11040 -22860 31040 -22850
rect -300 -23270 36260 -23260
rect -300 -23450 1630 -23270
rect 1810 -23450 2790 -23270
rect 2950 -23450 4390 -23270
rect 4550 -23450 5990 -23270
rect 6150 -23450 7590 -23270
rect 7750 -23450 9190 -23270
rect 9350 -23450 20110 -23270
rect 20290 -23450 36260 -23270
rect -300 -23460 36260 -23450
rect -300 -23670 36260 -23660
rect -300 -23850 430 -23670
rect 610 -23850 21310 -23670
rect 21490 -23850 36260 -23670
rect -300 -23860 36260 -23850
rect -300 -24260 36260 -24060
rect -300 -24660 36260 -24460
rect 1620 -25030 1820 -25020
rect 1620 -25040 1630 -25030
rect 1600 -25100 1630 -25040
rect 1620 -25110 1630 -25100
rect 1810 -25040 1820 -25030
rect 20100 -25030 20300 -25020
rect 20100 -25040 20110 -25030
rect 1810 -25070 20110 -25040
rect 1810 -25100 2510 -25070
rect 1810 -25110 1820 -25100
rect 1620 -25120 1820 -25110
rect 2500 -25130 2510 -25100
rect 4010 -25100 4710 -25070
rect 4010 -25130 4020 -25100
rect 2500 -25140 4020 -25130
rect 4700 -25130 4710 -25100
rect 6210 -25100 6910 -25070
rect 6210 -25130 6220 -25100
rect 4700 -25140 6220 -25130
rect 6900 -25130 6910 -25100
rect 8410 -25100 9110 -25070
rect 8410 -25130 8420 -25100
rect 6900 -25140 8420 -25130
rect 9100 -25130 9110 -25100
rect 10610 -25100 11310 -25070
rect 10610 -25130 10620 -25100
rect 9100 -25140 10620 -25130
rect 11300 -25130 11310 -25100
rect 12810 -25100 13510 -25070
rect 12810 -25130 12820 -25100
rect 11300 -25140 12820 -25130
rect 13500 -25130 13510 -25100
rect 15010 -25100 15710 -25070
rect 15010 -25130 15020 -25100
rect 13500 -25140 15020 -25130
rect 15700 -25130 15710 -25100
rect 17210 -25100 17910 -25070
rect 17210 -25130 17220 -25100
rect 15700 -25140 17220 -25130
rect 17900 -25130 17910 -25100
rect 19410 -25100 20110 -25070
rect 19410 -25130 19420 -25100
rect 20100 -25110 20110 -25100
rect 20290 -25040 20300 -25030
rect 20290 -25100 20320 -25040
rect 20290 -25110 20300 -25100
rect 20100 -25120 20300 -25110
rect 17900 -25140 19420 -25130
rect -110 -25210 30 -25180
rect -110 -25460 -80 -25210
rect 0 -25460 30 -25210
rect -110 -25480 30 -25460
rect 2090 -25210 2230 -25180
rect 2090 -25460 2120 -25210
rect 2200 -25460 2230 -25210
rect 2090 -25480 2230 -25460
rect 4290 -25210 4430 -25180
rect 4290 -25460 4320 -25210
rect 4400 -25460 4430 -25210
rect 4290 -25480 4430 -25460
rect 6490 -25210 6630 -25180
rect 6490 -25460 6520 -25210
rect 6600 -25460 6630 -25210
rect 6490 -25480 6630 -25460
rect 8690 -25210 8830 -25180
rect 8690 -25460 8720 -25210
rect 8800 -25460 8830 -25210
rect 8690 -25480 8830 -25460
rect 10890 -25210 11030 -25180
rect 10890 -25460 10920 -25210
rect 11000 -25460 11030 -25210
rect 10890 -25480 11030 -25460
rect 13090 -25210 13230 -25180
rect 13090 -25460 13120 -25210
rect 13200 -25460 13230 -25210
rect 13090 -25480 13230 -25460
rect 15290 -25210 15430 -25180
rect 15290 -25460 15320 -25210
rect 15400 -25460 15430 -25210
rect 15290 -25480 15430 -25460
rect 17490 -25210 17630 -25180
rect 17490 -25460 17520 -25210
rect 17600 -25460 17630 -25210
rect 17490 -25480 17630 -25460
rect 19690 -25210 19830 -25180
rect 19690 -25460 19720 -25210
rect 19800 -25460 19830 -25210
rect 19690 -25480 19830 -25460
rect 21890 -25210 22030 -25180
rect 21890 -25460 21920 -25210
rect 22000 -25460 22030 -25210
rect 21890 -25480 22030 -25460
rect 820 -25550 1020 -25540
rect 20500 -25550 20700 -25540
rect 820 -25560 830 -25550
rect -260 -25620 830 -25560
rect 820 -25630 830 -25620
rect 1010 -25560 1020 -25550
rect 2500 -25560 2700 -25550
rect 3160 -25560 3360 -25550
rect 3820 -25560 4020 -25550
rect 4700 -25560 4900 -25550
rect 5360 -25560 5560 -25550
rect 6020 -25560 6220 -25550
rect 6900 -25560 7100 -25550
rect 7560 -25560 7760 -25550
rect 8220 -25560 8420 -25550
rect 9100 -25560 9300 -25550
rect 9760 -25560 9960 -25550
rect 10420 -25560 10620 -25550
rect 11300 -25560 11500 -25550
rect 11960 -25560 12160 -25550
rect 12620 -25560 12820 -25550
rect 13500 -25560 13700 -25550
rect 14160 -25560 14360 -25550
rect 14820 -25560 15020 -25550
rect 15700 -25560 15900 -25550
rect 16360 -25560 16560 -25550
rect 17020 -25560 17220 -25550
rect 17900 -25560 18100 -25550
rect 18560 -25560 18760 -25550
rect 19220 -25560 19420 -25550
rect 20500 -25560 20510 -25550
rect 1010 -25620 6910 -25560
rect 7090 -25620 7570 -25560
rect 7750 -25620 8230 -25560
rect 8410 -25620 9110 -25560
rect 9290 -25620 9770 -25560
rect 9950 -25620 10430 -25560
rect 10610 -25620 11310 -25560
rect 11490 -25620 11970 -25560
rect 12150 -25620 12630 -25560
rect 12810 -25620 13510 -25560
rect 13690 -25620 14170 -25560
rect 14350 -25620 14830 -25560
rect 15010 -25620 20510 -25560
rect 1010 -25630 1020 -25620
rect 2500 -25630 2700 -25620
rect 3160 -25630 3360 -25620
rect 3820 -25630 4020 -25620
rect 4700 -25630 4900 -25620
rect 5360 -25630 5560 -25620
rect 6020 -25630 6220 -25620
rect 6900 -25630 7100 -25620
rect 7560 -25630 7760 -25620
rect 8220 -25630 8420 -25620
rect 9100 -25630 9300 -25620
rect 9760 -25630 9960 -25620
rect 10420 -25630 10620 -25620
rect 11300 -25630 11500 -25620
rect 11960 -25630 12160 -25620
rect 12620 -25630 12820 -25620
rect 13500 -25630 13700 -25620
rect 14160 -25630 14360 -25620
rect 14820 -25630 15020 -25620
rect 15700 -25630 15900 -25620
rect 16360 -25630 16560 -25620
rect 17020 -25630 17220 -25620
rect 17900 -25630 18100 -25620
rect 18560 -25630 18760 -25620
rect 19220 -25630 19420 -25620
rect 20500 -25630 20510 -25620
rect 20690 -25560 20700 -25550
rect 20690 -25620 22140 -25560
rect 20690 -25630 20700 -25620
rect 820 -25640 1020 -25630
rect 20500 -25640 20700 -25630
rect 1220 -25690 1420 -25680
rect 20900 -25690 21100 -25680
rect 1220 -25700 1230 -25690
rect -260 -25760 1230 -25700
rect 1220 -25770 1230 -25760
rect 1410 -25700 1420 -25690
rect 2500 -25700 2700 -25690
rect 3160 -25700 3360 -25690
rect 3820 -25700 4020 -25690
rect 4700 -25700 4900 -25690
rect 5360 -25700 5560 -25690
rect 6020 -25700 6220 -25690
rect 6900 -25700 7100 -25690
rect 7560 -25700 7760 -25690
rect 8220 -25700 8420 -25690
rect 9100 -25700 9300 -25690
rect 9760 -25700 9960 -25690
rect 10420 -25700 10620 -25690
rect 11300 -25700 11500 -25690
rect 11960 -25700 12160 -25690
rect 12620 -25700 12820 -25690
rect 13500 -25700 13700 -25690
rect 14160 -25700 14360 -25690
rect 14820 -25700 15020 -25690
rect 15700 -25700 15900 -25690
rect 16360 -25700 16560 -25690
rect 17020 -25700 17220 -25690
rect 17900 -25700 18100 -25690
rect 18560 -25700 18760 -25690
rect 19220 -25700 19420 -25690
rect 20900 -25700 20910 -25690
rect 1410 -25760 2510 -25700
rect 2690 -25760 3170 -25700
rect 3350 -25760 3830 -25700
rect 4010 -25760 4710 -25700
rect 4890 -25760 5370 -25700
rect 5550 -25760 6030 -25700
rect 6210 -25760 15710 -25700
rect 15890 -25760 16370 -25700
rect 16550 -25760 17030 -25700
rect 17210 -25760 17910 -25700
rect 18090 -25760 18570 -25700
rect 18750 -25760 19230 -25700
rect 19410 -25760 20910 -25700
rect 1410 -25770 1420 -25760
rect 2500 -25770 2700 -25760
rect 3160 -25770 3360 -25760
rect 3820 -25770 4020 -25760
rect 4700 -25770 4900 -25760
rect 5360 -25770 5560 -25760
rect 6020 -25770 6220 -25760
rect 6900 -25770 7100 -25760
rect 7560 -25770 7760 -25760
rect 8220 -25770 8420 -25760
rect 9100 -25770 9300 -25760
rect 9760 -25770 9960 -25760
rect 10420 -25770 10620 -25760
rect 11300 -25770 11500 -25760
rect 11960 -25770 12160 -25760
rect 12620 -25770 12820 -25760
rect 13500 -25770 13700 -25760
rect 14160 -25770 14360 -25760
rect 14820 -25770 15020 -25760
rect 15700 -25770 15900 -25760
rect 16360 -25770 16560 -25760
rect 17020 -25770 17220 -25760
rect 17900 -25770 18100 -25760
rect 18560 -25770 18760 -25760
rect 19220 -25770 19420 -25760
rect 20900 -25770 20910 -25760
rect 21090 -25700 21100 -25690
rect 21090 -25760 22140 -25700
rect 21090 -25770 21100 -25760
rect 1220 -25780 1420 -25770
rect 20900 -25780 21100 -25770
rect 1620 -25830 1820 -25820
rect 1620 -25840 1630 -25830
rect 1600 -25900 1630 -25840
rect 1620 -25910 1630 -25900
rect 1810 -25840 1820 -25830
rect 20100 -25830 20300 -25820
rect 20100 -25840 20110 -25830
rect 1810 -25870 20110 -25840
rect 1810 -25900 2510 -25870
rect 1810 -25910 1820 -25900
rect 1620 -25920 1820 -25910
rect 2500 -25930 2510 -25900
rect 4010 -25900 4710 -25870
rect 4010 -25930 4020 -25900
rect 2500 -25940 4020 -25930
rect 4700 -25930 4710 -25900
rect 6210 -25900 6910 -25870
rect 6210 -25930 6220 -25900
rect 4700 -25940 6220 -25930
rect 6900 -25930 6910 -25900
rect 8410 -25900 9110 -25870
rect 8410 -25930 8420 -25900
rect 6900 -25940 8420 -25930
rect 9100 -25930 9110 -25900
rect 10610 -25900 11310 -25870
rect 10610 -25930 10620 -25900
rect 9100 -25940 10620 -25930
rect 11300 -25930 11310 -25900
rect 12810 -25900 13510 -25870
rect 12810 -25930 12820 -25900
rect 11300 -25940 12820 -25930
rect 13500 -25930 13510 -25900
rect 15010 -25900 15710 -25870
rect 15010 -25930 15020 -25900
rect 13500 -25940 15020 -25930
rect 15700 -25930 15710 -25900
rect 17210 -25900 17910 -25870
rect 17210 -25930 17220 -25900
rect 15700 -25940 17220 -25930
rect 17900 -25930 17910 -25900
rect 19410 -25900 20110 -25870
rect 19410 -25930 19420 -25900
rect 20100 -25910 20110 -25900
rect 20290 -25840 20300 -25830
rect 20290 -25900 20320 -25840
rect 20290 -25910 20300 -25900
rect 20100 -25920 20300 -25910
rect 17900 -25940 19420 -25930
rect -110 -26010 30 -25980
rect -110 -26260 -80 -26010
rect 0 -26260 30 -26010
rect -110 -26280 30 -26260
rect 2090 -26010 2230 -25980
rect 2090 -26260 2120 -26010
rect 2200 -26260 2230 -26010
rect 2090 -26280 2230 -26260
rect 4290 -26010 4430 -25980
rect 4290 -26260 4320 -26010
rect 4400 -26260 4430 -26010
rect 4290 -26280 4430 -26260
rect 6490 -26010 6630 -25980
rect 6490 -26260 6520 -26010
rect 6600 -26260 6630 -26010
rect 6490 -26280 6630 -26260
rect 8690 -26010 8830 -25980
rect 8690 -26260 8720 -26010
rect 8800 -26260 8830 -26010
rect 8690 -26280 8830 -26260
rect 10890 -26010 11030 -25980
rect 10890 -26260 10920 -26010
rect 11000 -26260 11030 -26010
rect 10890 -26280 11030 -26260
rect 13090 -26010 13230 -25980
rect 13090 -26260 13120 -26010
rect 13200 -26260 13230 -26010
rect 13090 -26280 13230 -26260
rect 15290 -26010 15430 -25980
rect 15290 -26260 15320 -26010
rect 15400 -26260 15430 -26010
rect 15290 -26280 15430 -26260
rect 17490 -26010 17630 -25980
rect 17490 -26260 17520 -26010
rect 17600 -26260 17630 -26010
rect 17490 -26280 17630 -26260
rect 19690 -26010 19830 -25980
rect 19690 -26260 19720 -26010
rect 19800 -26260 19830 -26010
rect 19690 -26280 19830 -26260
rect 21890 -26010 22030 -25980
rect 21890 -26260 21920 -26010
rect 22000 -26260 22030 -26010
rect 21890 -26280 22030 -26260
rect 820 -26350 1020 -26340
rect 20500 -26350 20700 -26340
rect 820 -26360 830 -26350
rect -260 -26420 830 -26360
rect 820 -26430 830 -26420
rect 1010 -26360 1020 -26350
rect 2500 -26360 2700 -26350
rect 3160 -26360 3360 -26350
rect 3820 -26360 4020 -26350
rect 4700 -26360 4900 -26350
rect 5360 -26360 5560 -26350
rect 6020 -26360 6220 -26350
rect 6900 -26360 7100 -26350
rect 7560 -26360 7760 -26350
rect 8220 -26360 8420 -26350
rect 9100 -26360 9300 -26350
rect 9760 -26360 9960 -26350
rect 10420 -26360 10620 -26350
rect 11300 -26360 11500 -26350
rect 11960 -26360 12160 -26350
rect 12620 -26360 12820 -26350
rect 13500 -26360 13700 -26350
rect 14160 -26360 14360 -26350
rect 14820 -26360 15020 -26350
rect 15700 -26360 15900 -26350
rect 16360 -26360 16560 -26350
rect 17020 -26360 17220 -26350
rect 17900 -26360 18100 -26350
rect 18560 -26360 18760 -26350
rect 19220 -26360 19420 -26350
rect 20500 -26360 20510 -26350
rect 1010 -26420 2510 -26360
rect 2690 -26420 3170 -26360
rect 3350 -26420 3830 -26360
rect 4010 -26420 4710 -26360
rect 4890 -26420 5370 -26360
rect 5550 -26420 6030 -26360
rect 6210 -26420 15710 -26360
rect 15890 -26420 16370 -26360
rect 16550 -26420 17030 -26360
rect 17210 -26420 17910 -26360
rect 18090 -26420 18570 -26360
rect 18750 -26420 19230 -26360
rect 19410 -26420 20510 -26360
rect 1010 -26430 1020 -26420
rect 2500 -26430 2700 -26420
rect 3160 -26430 3360 -26420
rect 3820 -26430 4020 -26420
rect 4700 -26430 4900 -26420
rect 5360 -26430 5560 -26420
rect 6020 -26430 6220 -26420
rect 6900 -26430 7100 -26420
rect 7560 -26430 7760 -26420
rect 8220 -26430 8420 -26420
rect 9100 -26430 9300 -26420
rect 9760 -26430 9960 -26420
rect 10420 -26430 10620 -26420
rect 11300 -26430 11500 -26420
rect 11960 -26430 12160 -26420
rect 12620 -26430 12820 -26420
rect 13500 -26430 13700 -26420
rect 14160 -26430 14360 -26420
rect 14820 -26430 15020 -26420
rect 15700 -26430 15900 -26420
rect 16360 -26430 16560 -26420
rect 17020 -26430 17220 -26420
rect 17900 -26430 18100 -26420
rect 18560 -26430 18760 -26420
rect 19220 -26430 19420 -26420
rect 20500 -26430 20510 -26420
rect 20690 -26360 20700 -26350
rect 20690 -26420 22140 -26360
rect 20690 -26430 20700 -26420
rect 820 -26440 1020 -26430
rect 20500 -26440 20700 -26430
rect 1220 -26490 1420 -26480
rect 20900 -26490 21100 -26480
rect 1220 -26500 1230 -26490
rect -260 -26560 1230 -26500
rect 1220 -26570 1230 -26560
rect 1410 -26500 1420 -26490
rect 2500 -26500 2700 -26490
rect 3160 -26500 3360 -26490
rect 3820 -26500 4020 -26490
rect 4700 -26500 4900 -26490
rect 5360 -26500 5560 -26490
rect 6020 -26500 6220 -26490
rect 6900 -26500 7100 -26490
rect 7560 -26500 7760 -26490
rect 8220 -26500 8420 -26490
rect 9100 -26500 9300 -26490
rect 9760 -26500 9960 -26490
rect 10420 -26500 10620 -26490
rect 11300 -26500 11500 -26490
rect 11960 -26500 12160 -26490
rect 12620 -26500 12820 -26490
rect 13500 -26500 13700 -26490
rect 14160 -26500 14360 -26490
rect 14820 -26500 15020 -26490
rect 15700 -26500 15900 -26490
rect 16360 -26500 16560 -26490
rect 17020 -26500 17220 -26490
rect 17900 -26500 18100 -26490
rect 18560 -26500 18760 -26490
rect 19220 -26500 19420 -26490
rect 20900 -26500 20910 -26490
rect 1410 -26560 6910 -26500
rect 7090 -26560 7570 -26500
rect 7750 -26560 8230 -26500
rect 8410 -26560 9110 -26500
rect 9290 -26560 9770 -26500
rect 9950 -26560 10430 -26500
rect 10610 -26560 11310 -26500
rect 11490 -26560 11970 -26500
rect 12150 -26560 12630 -26500
rect 12810 -26560 13510 -26500
rect 13690 -26560 14170 -26500
rect 14350 -26560 14830 -26500
rect 15010 -26560 20910 -26500
rect 1410 -26570 1420 -26560
rect 2500 -26570 2700 -26560
rect 3160 -26570 3360 -26560
rect 3820 -26570 4020 -26560
rect 4700 -26570 4900 -26560
rect 5360 -26570 5560 -26560
rect 6020 -26570 6220 -26560
rect 6900 -26570 7100 -26560
rect 7560 -26570 7760 -26560
rect 8220 -26570 8420 -26560
rect 9100 -26570 9300 -26560
rect 9760 -26570 9960 -26560
rect 10420 -26570 10620 -26560
rect 11300 -26570 11500 -26560
rect 11960 -26570 12160 -26560
rect 12620 -26570 12820 -26560
rect 13500 -26570 13700 -26560
rect 14160 -26570 14360 -26560
rect 14820 -26570 15020 -26560
rect 15700 -26570 15900 -26560
rect 16360 -26570 16560 -26560
rect 17020 -26570 17220 -26560
rect 17900 -26570 18100 -26560
rect 18560 -26570 18760 -26560
rect 19220 -26570 19420 -26560
rect 20900 -26570 20910 -26560
rect 21090 -26500 21100 -26490
rect 21090 -26560 22140 -26500
rect 21090 -26570 21100 -26560
rect 1220 -26580 1420 -26570
rect 20900 -26580 21100 -26570
rect 420 -26630 620 -26620
rect 420 -26710 430 -26630
rect 610 -26710 620 -26630
rect 1620 -26630 1820 -26620
rect 1620 -26640 1630 -26630
rect 1600 -26700 1630 -26640
rect 420 -26720 620 -26710
rect 1620 -26710 1630 -26700
rect 1810 -26640 1820 -26630
rect 20100 -26630 20300 -26620
rect 20100 -26640 20110 -26630
rect 1810 -26670 20110 -26640
rect 1810 -26700 4710 -26670
rect 1810 -26710 1820 -26700
rect 1620 -26720 1820 -26710
rect 4700 -26730 4710 -26700
rect 6210 -26700 6910 -26670
rect 6210 -26730 6220 -26700
rect 4700 -26740 6220 -26730
rect 6900 -26730 6910 -26700
rect 8410 -26700 9110 -26670
rect 8410 -26730 8420 -26700
rect 6900 -26740 8420 -26730
rect 9100 -26730 9110 -26700
rect 10610 -26700 11310 -26670
rect 10610 -26730 10620 -26700
rect 9100 -26740 10620 -26730
rect 11300 -26730 11310 -26700
rect 12810 -26700 13510 -26670
rect 12810 -26730 12820 -26700
rect 11300 -26740 12820 -26730
rect 13500 -26730 13510 -26700
rect 15010 -26700 15710 -26670
rect 15010 -26730 15020 -26700
rect 13500 -26740 15020 -26730
rect 15700 -26730 15710 -26700
rect 17210 -26700 20110 -26670
rect 17210 -26730 17220 -26700
rect 20100 -26710 20110 -26700
rect 20290 -26640 20300 -26630
rect 21300 -26630 21500 -26620
rect 20290 -26700 20320 -26640
rect 20290 -26710 20300 -26700
rect 20100 -26720 20300 -26710
rect 21300 -26710 21310 -26630
rect 21490 -26710 21500 -26630
rect 21300 -26720 21500 -26710
rect 15700 -26740 17220 -26730
rect -110 -26810 30 -26780
rect -110 -27060 -80 -26810
rect 0 -27060 30 -26810
rect -110 -27080 30 -27060
rect 2090 -26810 2230 -26780
rect 2090 -27060 2120 -26810
rect 2200 -27060 2230 -26810
rect 2090 -27080 2230 -27060
rect 4290 -26810 4430 -26780
rect 4290 -27060 4320 -26810
rect 4400 -27060 4430 -26810
rect 4290 -27080 4430 -27060
rect 6490 -26810 6630 -26780
rect 6490 -27060 6520 -26810
rect 6600 -27060 6630 -26810
rect 6490 -27080 6630 -27060
rect 8690 -26810 8830 -26780
rect 8690 -27060 8720 -26810
rect 8800 -27060 8830 -26810
rect 8690 -27080 8830 -27060
rect 10890 -26810 11030 -26780
rect 10890 -27060 10920 -26810
rect 11000 -27060 11030 -26810
rect 10890 -27080 11030 -27060
rect 13090 -26810 13230 -26780
rect 13090 -27060 13120 -26810
rect 13200 -27060 13230 -26810
rect 13090 -27080 13230 -27060
rect 15290 -26810 15430 -26780
rect 15290 -27060 15320 -26810
rect 15400 -27060 15430 -26810
rect 15290 -27080 15430 -27060
rect 17490 -26810 17630 -26780
rect 17490 -27060 17520 -26810
rect 17600 -27060 17630 -26810
rect 17490 -27080 17630 -27060
rect 19690 -26810 19830 -26780
rect 19690 -27060 19720 -26810
rect 19800 -27060 19830 -26810
rect 19690 -27080 19830 -27060
rect 21890 -26810 22030 -26780
rect 21890 -27060 21920 -26810
rect 22000 -27060 22030 -26810
rect 21890 -27080 22030 -27060
rect 820 -27150 1020 -27140
rect 20500 -27150 20700 -27140
rect 820 -27160 830 -27150
rect -260 -27220 830 -27160
rect 820 -27230 830 -27220
rect 1010 -27160 1020 -27150
rect 2500 -27160 2700 -27150
rect 3160 -27160 3360 -27150
rect 3820 -27160 4020 -27150
rect 4700 -27160 4900 -27150
rect 5360 -27160 5560 -27150
rect 6020 -27160 6220 -27150
rect 6900 -27160 7100 -27150
rect 7560 -27160 7760 -27150
rect 8220 -27160 8420 -27150
rect 9100 -27160 9300 -27150
rect 9760 -27160 9960 -27150
rect 10420 -27160 10620 -27150
rect 11300 -27160 11500 -27150
rect 11960 -27160 12160 -27150
rect 12620 -27160 12820 -27150
rect 13500 -27160 13700 -27150
rect 14160 -27160 14360 -27150
rect 14820 -27160 15020 -27150
rect 15700 -27160 15900 -27150
rect 16360 -27160 16560 -27150
rect 17020 -27160 17220 -27150
rect 17900 -27160 18100 -27150
rect 18560 -27160 18760 -27150
rect 19220 -27160 19420 -27150
rect 20500 -27160 20510 -27150
rect 1010 -27220 6910 -27160
rect 7090 -27220 7570 -27160
rect 7750 -27220 8230 -27160
rect 8410 -27220 9110 -27160
rect 9290 -27220 9770 -27160
rect 9950 -27220 10430 -27160
rect 10610 -27220 11310 -27160
rect 11490 -27220 11970 -27160
rect 12150 -27220 12630 -27160
rect 12810 -27220 13510 -27160
rect 13690 -27220 14170 -27160
rect 14350 -27220 14830 -27160
rect 15010 -27220 20510 -27160
rect 1010 -27230 1020 -27220
rect 2500 -27230 2700 -27220
rect 3160 -27230 3360 -27220
rect 3820 -27230 4020 -27220
rect 4700 -27230 4900 -27220
rect 5360 -27230 5560 -27220
rect 6020 -27230 6220 -27220
rect 6900 -27230 7100 -27220
rect 7560 -27230 7760 -27220
rect 8220 -27230 8420 -27220
rect 9100 -27230 9300 -27220
rect 9760 -27230 9960 -27220
rect 10420 -27230 10620 -27220
rect 11300 -27230 11500 -27220
rect 11960 -27230 12160 -27220
rect 12620 -27230 12820 -27220
rect 13500 -27230 13700 -27220
rect 14160 -27230 14360 -27220
rect 14820 -27230 15020 -27220
rect 15700 -27230 15900 -27220
rect 16360 -27230 16560 -27220
rect 17020 -27230 17220 -27220
rect 17900 -27230 18100 -27220
rect 18560 -27230 18760 -27220
rect 19220 -27230 19420 -27220
rect 20500 -27230 20510 -27220
rect 20690 -27160 20700 -27150
rect 20690 -27220 22140 -27160
rect 20690 -27230 20700 -27220
rect 820 -27240 1020 -27230
rect 20500 -27240 20700 -27230
rect 1220 -27290 1420 -27280
rect 20900 -27290 21100 -27280
rect 1220 -27300 1230 -27290
rect -260 -27360 1230 -27300
rect 1220 -27370 1230 -27360
rect 1410 -27300 1420 -27290
rect 2500 -27300 2700 -27290
rect 3160 -27300 3360 -27290
rect 3820 -27300 4020 -27290
rect 4700 -27300 4900 -27290
rect 5360 -27300 5560 -27290
rect 6020 -27300 6220 -27290
rect 6900 -27300 7100 -27290
rect 7560 -27300 7760 -27290
rect 8220 -27300 8420 -27290
rect 9100 -27300 9300 -27290
rect 9760 -27300 9960 -27290
rect 10420 -27300 10620 -27290
rect 11300 -27300 11500 -27290
rect 11960 -27300 12160 -27290
rect 12620 -27300 12820 -27290
rect 13500 -27300 13700 -27290
rect 14160 -27300 14360 -27290
rect 14820 -27300 15020 -27290
rect 15700 -27300 15900 -27290
rect 16360 -27300 16560 -27290
rect 17020 -27300 17220 -27290
rect 17900 -27300 18100 -27290
rect 18560 -27300 18760 -27290
rect 19220 -27300 19420 -27290
rect 20900 -27300 20910 -27290
rect 1410 -27360 2510 -27300
rect 2690 -27360 3170 -27300
rect 3350 -27360 3830 -27300
rect 4010 -27360 4710 -27300
rect 4890 -27360 5370 -27300
rect 5550 -27360 6030 -27300
rect 6210 -27360 15710 -27300
rect 15890 -27360 16370 -27300
rect 16550 -27360 17030 -27300
rect 17210 -27360 17910 -27300
rect 18090 -27360 18570 -27300
rect 18750 -27360 19230 -27300
rect 19410 -27360 20910 -27300
rect 1410 -27370 1420 -27360
rect 2500 -27370 2700 -27360
rect 3160 -27370 3360 -27360
rect 3820 -27370 4020 -27360
rect 4700 -27370 4900 -27360
rect 5360 -27370 5560 -27360
rect 6020 -27370 6220 -27360
rect 6900 -27370 7100 -27360
rect 7560 -27370 7760 -27360
rect 8220 -27370 8420 -27360
rect 9100 -27370 9300 -27360
rect 9760 -27370 9960 -27360
rect 10420 -27370 10620 -27360
rect 11300 -27370 11500 -27360
rect 11960 -27370 12160 -27360
rect 12620 -27370 12820 -27360
rect 13500 -27370 13700 -27360
rect 14160 -27370 14360 -27360
rect 14820 -27370 15020 -27360
rect 15700 -27370 15900 -27360
rect 16360 -27370 16560 -27360
rect 17020 -27370 17220 -27360
rect 17900 -27370 18100 -27360
rect 18560 -27370 18760 -27360
rect 19220 -27370 19420 -27360
rect 20900 -27370 20910 -27360
rect 21090 -27300 21100 -27290
rect 21090 -27360 22140 -27300
rect 21090 -27370 21100 -27360
rect 1220 -27380 1420 -27370
rect 20900 -27380 21100 -27370
rect 420 -27430 620 -27420
rect 420 -27510 430 -27430
rect 610 -27510 620 -27430
rect 1620 -27430 1820 -27420
rect 1620 -27440 1630 -27430
rect 1600 -27500 1630 -27440
rect 420 -27520 620 -27510
rect 1620 -27510 1630 -27500
rect 1810 -27440 1820 -27430
rect 20100 -27430 20300 -27420
rect 20100 -27440 20110 -27430
rect 1810 -27470 20110 -27440
rect 1810 -27500 4710 -27470
rect 1810 -27510 1820 -27500
rect 1620 -27520 1820 -27510
rect 4700 -27530 4710 -27500
rect 6210 -27500 6910 -27470
rect 6210 -27530 6220 -27500
rect 4700 -27540 6220 -27530
rect 6900 -27530 6910 -27500
rect 8410 -27500 9110 -27470
rect 8410 -27530 8420 -27500
rect 6900 -27540 8420 -27530
rect 9100 -27530 9110 -27500
rect 10610 -27500 11310 -27470
rect 10610 -27530 10620 -27500
rect 9100 -27540 10620 -27530
rect 11300 -27530 11310 -27500
rect 12810 -27500 13510 -27470
rect 12810 -27530 12820 -27500
rect 11300 -27540 12820 -27530
rect 13500 -27530 13510 -27500
rect 15010 -27500 15710 -27470
rect 15010 -27530 15020 -27500
rect 13500 -27540 15020 -27530
rect 15700 -27530 15710 -27500
rect 17210 -27500 20110 -27470
rect 17210 -27530 17220 -27500
rect 20100 -27510 20110 -27500
rect 20290 -27440 20300 -27430
rect 21300 -27430 21500 -27420
rect 20290 -27500 20320 -27440
rect 20290 -27510 20300 -27500
rect 20100 -27520 20300 -27510
rect 21300 -27510 21310 -27430
rect 21490 -27510 21500 -27430
rect 21300 -27520 21500 -27510
rect 15700 -27540 17220 -27530
rect -110 -27610 30 -27580
rect -110 -27860 -80 -27610
rect 0 -27860 30 -27610
rect -110 -27880 30 -27860
rect 2090 -27610 2230 -27580
rect 2090 -27860 2120 -27610
rect 2200 -27860 2230 -27610
rect 2090 -27880 2230 -27860
rect 4290 -27610 4430 -27580
rect 4290 -27860 4320 -27610
rect 4400 -27860 4430 -27610
rect 4290 -27880 4430 -27860
rect 6490 -27610 6630 -27580
rect 6490 -27860 6520 -27610
rect 6600 -27860 6630 -27610
rect 6490 -27880 6630 -27860
rect 8690 -27610 8830 -27580
rect 8690 -27860 8720 -27610
rect 8800 -27860 8830 -27610
rect 8690 -27880 8830 -27860
rect 10890 -27610 11030 -27580
rect 10890 -27860 10920 -27610
rect 11000 -27860 11030 -27610
rect 10890 -27880 11030 -27860
rect 13090 -27610 13230 -27580
rect 13090 -27860 13120 -27610
rect 13200 -27860 13230 -27610
rect 13090 -27880 13230 -27860
rect 15290 -27610 15430 -27580
rect 15290 -27860 15320 -27610
rect 15400 -27860 15430 -27610
rect 15290 -27880 15430 -27860
rect 17490 -27610 17630 -27580
rect 17490 -27860 17520 -27610
rect 17600 -27860 17630 -27610
rect 17490 -27880 17630 -27860
rect 19690 -27610 19830 -27580
rect 19690 -27860 19720 -27610
rect 19800 -27860 19830 -27610
rect 19690 -27880 19830 -27860
rect 21890 -27610 22030 -27580
rect 21890 -27860 21920 -27610
rect 22000 -27860 22030 -27610
rect 21890 -27880 22030 -27860
rect 820 -27950 1020 -27940
rect 20500 -27950 20700 -27940
rect 820 -27960 830 -27950
rect -260 -28020 830 -27960
rect 820 -28030 830 -28020
rect 1010 -27960 1020 -27950
rect 2500 -27960 2700 -27950
rect 3160 -27960 3360 -27950
rect 3820 -27960 4020 -27950
rect 4700 -27960 4900 -27950
rect 5360 -27960 5560 -27950
rect 6020 -27960 6220 -27950
rect 6900 -27960 7100 -27950
rect 7560 -27960 7760 -27950
rect 8220 -27960 8420 -27950
rect 9100 -27960 9300 -27950
rect 9760 -27960 9960 -27950
rect 10420 -27960 10620 -27950
rect 11300 -27960 11500 -27950
rect 11960 -27960 12160 -27950
rect 12620 -27960 12820 -27950
rect 13500 -27960 13700 -27950
rect 14160 -27960 14360 -27950
rect 14820 -27960 15020 -27950
rect 15700 -27960 15900 -27950
rect 16360 -27960 16560 -27950
rect 17020 -27960 17220 -27950
rect 17900 -27960 18100 -27950
rect 18560 -27960 18760 -27950
rect 19220 -27960 19420 -27950
rect 20500 -27960 20510 -27950
rect 1010 -28020 2510 -27960
rect 2690 -28020 3170 -27960
rect 3350 -28020 3830 -27960
rect 4010 -28020 4710 -27960
rect 4890 -28020 5370 -27960
rect 5550 -28020 6030 -27960
rect 6210 -28020 15710 -27960
rect 15890 -28020 16370 -27960
rect 16550 -28020 17030 -27960
rect 17210 -28020 17910 -27960
rect 18090 -28020 18570 -27960
rect 18750 -28020 19230 -27960
rect 19410 -28020 20510 -27960
rect 1010 -28030 1020 -28020
rect 2500 -28030 2700 -28020
rect 3160 -28030 3360 -28020
rect 3820 -28030 4020 -28020
rect 4700 -28030 4900 -28020
rect 5360 -28030 5560 -28020
rect 6020 -28030 6220 -28020
rect 6900 -28030 7100 -28020
rect 7560 -28030 7760 -28020
rect 8220 -28030 8420 -28020
rect 9100 -28030 9300 -28020
rect 9760 -28030 9960 -28020
rect 10420 -28030 10620 -28020
rect 11300 -28030 11500 -28020
rect 11960 -28030 12160 -28020
rect 12620 -28030 12820 -28020
rect 13500 -28030 13700 -28020
rect 14160 -28030 14360 -28020
rect 14820 -28030 15020 -28020
rect 15700 -28030 15900 -28020
rect 16360 -28030 16560 -28020
rect 17020 -28030 17220 -28020
rect 17900 -28030 18100 -28020
rect 18560 -28030 18760 -28020
rect 19220 -28030 19420 -28020
rect 20500 -28030 20510 -28020
rect 20690 -27960 20700 -27950
rect 20690 -28020 22140 -27960
rect 20690 -28030 20700 -28020
rect 820 -28040 1020 -28030
rect 20500 -28040 20700 -28030
rect 1220 -28090 1420 -28080
rect 20900 -28090 21100 -28080
rect 1220 -28100 1230 -28090
rect -260 -28160 1230 -28100
rect 1220 -28170 1230 -28160
rect 1410 -28100 1420 -28090
rect 2500 -28100 2700 -28090
rect 3160 -28100 3360 -28090
rect 3820 -28100 4020 -28090
rect 4700 -28100 4900 -28090
rect 5360 -28100 5560 -28090
rect 6020 -28100 6220 -28090
rect 6900 -28100 7100 -28090
rect 7560 -28100 7760 -28090
rect 8220 -28100 8420 -28090
rect 9100 -28100 9300 -28090
rect 9760 -28100 9960 -28090
rect 10420 -28100 10620 -28090
rect 11300 -28100 11500 -28090
rect 11960 -28100 12160 -28090
rect 12620 -28100 12820 -28090
rect 13500 -28100 13700 -28090
rect 14160 -28100 14360 -28090
rect 14820 -28100 15020 -28090
rect 15700 -28100 15900 -28090
rect 16360 -28100 16560 -28090
rect 17020 -28100 17220 -28090
rect 17900 -28100 18100 -28090
rect 18560 -28100 18760 -28090
rect 19220 -28100 19420 -28090
rect 20900 -28100 20910 -28090
rect 1410 -28160 6910 -28100
rect 7090 -28160 7570 -28100
rect 7750 -28160 8230 -28100
rect 8410 -28160 9110 -28100
rect 9290 -28160 9770 -28100
rect 9950 -28160 10430 -28100
rect 10610 -28160 11310 -28100
rect 11490 -28160 11970 -28100
rect 12150 -28160 12630 -28100
rect 12810 -28160 13510 -28100
rect 13690 -28160 14170 -28100
rect 14350 -28160 14830 -28100
rect 15010 -28160 20910 -28100
rect 1410 -28170 1420 -28160
rect 2500 -28170 2700 -28160
rect 3160 -28170 3360 -28160
rect 3820 -28170 4020 -28160
rect 4700 -28170 4900 -28160
rect 5360 -28170 5560 -28160
rect 6020 -28170 6220 -28160
rect 6900 -28170 7100 -28160
rect 7560 -28170 7760 -28160
rect 8220 -28170 8420 -28160
rect 9100 -28170 9300 -28160
rect 9760 -28170 9960 -28160
rect 10420 -28170 10620 -28160
rect 11300 -28170 11500 -28160
rect 11960 -28170 12160 -28160
rect 12620 -28170 12820 -28160
rect 13500 -28170 13700 -28160
rect 14160 -28170 14360 -28160
rect 14820 -28170 15020 -28160
rect 15700 -28170 15900 -28160
rect 16360 -28170 16560 -28160
rect 17020 -28170 17220 -28160
rect 17900 -28170 18100 -28160
rect 18560 -28170 18760 -28160
rect 19220 -28170 19420 -28160
rect 20900 -28170 20910 -28160
rect 21090 -28100 21100 -28090
rect 21090 -28160 22140 -28100
rect 21090 -28170 21100 -28160
rect 1220 -28180 1420 -28170
rect 20900 -28180 21100 -28170
rect 420 -28230 620 -28220
rect 420 -28310 430 -28230
rect 610 -28310 620 -28230
rect 1620 -28230 1820 -28220
rect 1620 -28240 1630 -28230
rect 1600 -28300 1630 -28240
rect 420 -28320 620 -28310
rect 1620 -28310 1630 -28300
rect 1810 -28240 1820 -28230
rect 20100 -28230 20300 -28220
rect 20100 -28240 20110 -28230
rect 1810 -28270 20110 -28240
rect 1810 -28300 4710 -28270
rect 1810 -28310 1820 -28300
rect 1620 -28320 1820 -28310
rect 4700 -28330 4710 -28300
rect 6210 -28300 6910 -28270
rect 6210 -28330 6220 -28300
rect 4700 -28340 6220 -28330
rect 6900 -28330 6910 -28300
rect 8410 -28300 9110 -28270
rect 8410 -28330 8420 -28300
rect 6900 -28340 8420 -28330
rect 9100 -28330 9110 -28300
rect 10610 -28300 11310 -28270
rect 10610 -28330 10620 -28300
rect 9100 -28340 10620 -28330
rect 11300 -28330 11310 -28300
rect 12810 -28300 13510 -28270
rect 12810 -28330 12820 -28300
rect 11300 -28340 12820 -28330
rect 13500 -28330 13510 -28300
rect 15010 -28300 15710 -28270
rect 15010 -28330 15020 -28300
rect 13500 -28340 15020 -28330
rect 15700 -28330 15710 -28300
rect 17210 -28300 20110 -28270
rect 17210 -28330 17220 -28300
rect 20100 -28310 20110 -28300
rect 20290 -28240 20300 -28230
rect 21300 -28230 21500 -28220
rect 20290 -28300 20320 -28240
rect 20290 -28310 20300 -28300
rect 20100 -28320 20300 -28310
rect 21300 -28310 21310 -28230
rect 21490 -28310 21500 -28230
rect 21300 -28320 21500 -28310
rect 15700 -28340 17220 -28330
rect -110 -28410 30 -28380
rect -110 -28660 -80 -28410
rect 0 -28660 30 -28410
rect -110 -28680 30 -28660
rect 2090 -28410 2230 -28380
rect 2090 -28660 2120 -28410
rect 2200 -28660 2230 -28410
rect 2090 -28680 2230 -28660
rect 4290 -28410 4430 -28380
rect 4290 -28660 4320 -28410
rect 4400 -28660 4430 -28410
rect 4290 -28680 4430 -28660
rect 6490 -28410 6630 -28380
rect 6490 -28660 6520 -28410
rect 6600 -28660 6630 -28410
rect 6490 -28680 6630 -28660
rect 8690 -28410 8830 -28380
rect 8690 -28660 8720 -28410
rect 8800 -28660 8830 -28410
rect 8690 -28680 8830 -28660
rect 10890 -28410 11030 -28380
rect 10890 -28660 10920 -28410
rect 11000 -28660 11030 -28410
rect 10890 -28680 11030 -28660
rect 13090 -28410 13230 -28380
rect 13090 -28660 13120 -28410
rect 13200 -28660 13230 -28410
rect 13090 -28680 13230 -28660
rect 15290 -28410 15430 -28380
rect 15290 -28660 15320 -28410
rect 15400 -28660 15430 -28410
rect 15290 -28680 15430 -28660
rect 17490 -28410 17630 -28380
rect 17490 -28660 17520 -28410
rect 17600 -28660 17630 -28410
rect 17490 -28680 17630 -28660
rect 19690 -28410 19830 -28380
rect 19690 -28660 19720 -28410
rect 19800 -28660 19830 -28410
rect 19690 -28680 19830 -28660
rect 21890 -28410 22030 -28380
rect 21890 -28660 21920 -28410
rect 22000 -28660 22030 -28410
rect 21890 -28680 22030 -28660
rect 820 -28750 1020 -28740
rect 20500 -28750 20700 -28740
rect 820 -28760 830 -28750
rect -260 -28820 830 -28760
rect 820 -28830 830 -28820
rect 1010 -28760 1020 -28750
rect 2500 -28760 2700 -28750
rect 3160 -28760 3360 -28750
rect 3820 -28760 4020 -28750
rect 4700 -28760 4900 -28750
rect 5360 -28760 5560 -28750
rect 6020 -28760 6220 -28750
rect 6900 -28760 7100 -28750
rect 7560 -28760 7760 -28750
rect 8220 -28760 8420 -28750
rect 9100 -28760 9300 -28750
rect 9760 -28760 9960 -28750
rect 10420 -28760 10620 -28750
rect 11300 -28760 11500 -28750
rect 11960 -28760 12160 -28750
rect 12620 -28760 12820 -28750
rect 13500 -28760 13700 -28750
rect 14160 -28760 14360 -28750
rect 14820 -28760 15020 -28750
rect 15700 -28760 15900 -28750
rect 16360 -28760 16560 -28750
rect 17020 -28760 17220 -28750
rect 17900 -28760 18100 -28750
rect 18560 -28760 18760 -28750
rect 19220 -28760 19420 -28750
rect 20500 -28760 20510 -28750
rect 1010 -28820 2510 -28760
rect 2690 -28820 3170 -28760
rect 3350 -28820 3830 -28760
rect 4010 -28820 4710 -28760
rect 4890 -28820 5370 -28760
rect 5550 -28820 6030 -28760
rect 6210 -28820 15710 -28760
rect 15890 -28820 16370 -28760
rect 16550 -28820 17030 -28760
rect 17210 -28820 17910 -28760
rect 18090 -28820 18570 -28760
rect 18750 -28820 19230 -28760
rect 19410 -28820 20510 -28760
rect 1010 -28830 1020 -28820
rect 2500 -28830 2700 -28820
rect 3160 -28830 3360 -28820
rect 3820 -28830 4020 -28820
rect 4700 -28830 4900 -28820
rect 5360 -28830 5560 -28820
rect 6020 -28830 6220 -28820
rect 6900 -28830 7100 -28820
rect 7560 -28830 7760 -28820
rect 8220 -28830 8420 -28820
rect 9100 -28830 9300 -28820
rect 9760 -28830 9960 -28820
rect 10420 -28830 10620 -28820
rect 11300 -28830 11500 -28820
rect 11960 -28830 12160 -28820
rect 12620 -28830 12820 -28820
rect 13500 -28830 13700 -28820
rect 14160 -28830 14360 -28820
rect 14820 -28830 15020 -28820
rect 15700 -28830 15900 -28820
rect 16360 -28830 16560 -28820
rect 17020 -28830 17220 -28820
rect 17900 -28830 18100 -28820
rect 18560 -28830 18760 -28820
rect 19220 -28830 19420 -28820
rect 20500 -28830 20510 -28820
rect 20690 -28760 20700 -28750
rect 20690 -28820 22140 -28760
rect 20690 -28830 20700 -28820
rect 820 -28840 1020 -28830
rect 20500 -28840 20700 -28830
rect 1220 -28890 1420 -28880
rect 20900 -28890 21100 -28880
rect 1220 -28900 1230 -28890
rect -260 -28960 1230 -28900
rect 1220 -28970 1230 -28960
rect 1410 -28900 1420 -28890
rect 2500 -28900 2700 -28890
rect 3160 -28900 3360 -28890
rect 3820 -28900 4020 -28890
rect 4700 -28900 4900 -28890
rect 5360 -28900 5560 -28890
rect 6020 -28900 6220 -28890
rect 6900 -28900 7100 -28890
rect 7560 -28900 7760 -28890
rect 8220 -28900 8420 -28890
rect 9100 -28900 9300 -28890
rect 9760 -28900 9960 -28890
rect 10420 -28900 10620 -28890
rect 11300 -28900 11500 -28890
rect 11960 -28900 12160 -28890
rect 12620 -28900 12820 -28890
rect 13500 -28900 13700 -28890
rect 14160 -28900 14360 -28890
rect 14820 -28900 15020 -28890
rect 15700 -28900 15900 -28890
rect 16360 -28900 16560 -28890
rect 17020 -28900 17220 -28890
rect 17900 -28900 18100 -28890
rect 18560 -28900 18760 -28890
rect 19220 -28900 19420 -28890
rect 20900 -28900 20910 -28890
rect 1410 -28960 6910 -28900
rect 7090 -28960 7570 -28900
rect 7750 -28960 8230 -28900
rect 8410 -28960 9110 -28900
rect 9290 -28960 9770 -28900
rect 9950 -28960 10430 -28900
rect 10610 -28960 11310 -28900
rect 11490 -28960 11970 -28900
rect 12150 -28960 12630 -28900
rect 12810 -28960 13510 -28900
rect 13690 -28960 14170 -28900
rect 14350 -28960 14830 -28900
rect 15010 -28960 20910 -28900
rect 1410 -28970 1420 -28960
rect 2500 -28970 2700 -28960
rect 3160 -28970 3360 -28960
rect 3820 -28970 4020 -28960
rect 4700 -28970 4900 -28960
rect 5360 -28970 5560 -28960
rect 6020 -28970 6220 -28960
rect 6900 -28970 7100 -28960
rect 7560 -28970 7760 -28960
rect 8220 -28970 8420 -28960
rect 9100 -28970 9300 -28960
rect 9760 -28970 9960 -28960
rect 10420 -28970 10620 -28960
rect 11300 -28970 11500 -28960
rect 11960 -28970 12160 -28960
rect 12620 -28970 12820 -28960
rect 13500 -28970 13700 -28960
rect 14160 -28970 14360 -28960
rect 14820 -28970 15020 -28960
rect 15700 -28970 15900 -28960
rect 16360 -28970 16560 -28960
rect 17020 -28970 17220 -28960
rect 17900 -28970 18100 -28960
rect 18560 -28970 18760 -28960
rect 19220 -28970 19420 -28960
rect 20900 -28970 20910 -28960
rect 21090 -28900 21100 -28890
rect 21090 -28960 22140 -28900
rect 21090 -28970 21100 -28960
rect 1220 -28980 1420 -28970
rect 20900 -28980 21100 -28970
rect 420 -29030 620 -29020
rect 420 -29110 430 -29030
rect 610 -29110 620 -29030
rect 1620 -29030 1820 -29020
rect 1620 -29040 1630 -29030
rect 1600 -29100 1630 -29040
rect 420 -29120 620 -29110
rect 1620 -29110 1630 -29100
rect 1810 -29040 1820 -29030
rect 20100 -29030 20300 -29020
rect 20100 -29040 20110 -29030
rect 1810 -29070 20110 -29040
rect 1810 -29100 4710 -29070
rect 1810 -29110 1820 -29100
rect 1620 -29120 1820 -29110
rect 4700 -29130 4710 -29100
rect 6210 -29100 6910 -29070
rect 6210 -29130 6220 -29100
rect 4700 -29140 6220 -29130
rect 6900 -29130 6910 -29100
rect 8410 -29100 9110 -29070
rect 8410 -29130 8420 -29100
rect 6900 -29140 8420 -29130
rect 9100 -29130 9110 -29100
rect 10610 -29100 11310 -29070
rect 10610 -29130 10620 -29100
rect 9100 -29140 10620 -29130
rect 11300 -29130 11310 -29100
rect 12810 -29100 13510 -29070
rect 12810 -29130 12820 -29100
rect 11300 -29140 12820 -29130
rect 13500 -29130 13510 -29100
rect 15010 -29100 15710 -29070
rect 15010 -29130 15020 -29100
rect 13500 -29140 15020 -29130
rect 15700 -29130 15710 -29100
rect 17210 -29100 20110 -29070
rect 17210 -29130 17220 -29100
rect 20100 -29110 20110 -29100
rect 20290 -29040 20300 -29030
rect 21300 -29030 21500 -29020
rect 20290 -29100 20320 -29040
rect 20290 -29110 20300 -29100
rect 20100 -29120 20300 -29110
rect 21300 -29110 21310 -29030
rect 21490 -29110 21500 -29030
rect 21300 -29120 21500 -29110
rect 15700 -29140 17220 -29130
rect -110 -29210 30 -29180
rect -110 -29460 -80 -29210
rect 0 -29460 30 -29210
rect -110 -29480 30 -29460
rect 2090 -29210 2230 -29180
rect 2090 -29460 2120 -29210
rect 2200 -29460 2230 -29210
rect 2090 -29480 2230 -29460
rect 4290 -29210 4430 -29180
rect 4290 -29460 4320 -29210
rect 4400 -29460 4430 -29210
rect 4290 -29480 4430 -29460
rect 6490 -29210 6630 -29180
rect 6490 -29460 6520 -29210
rect 6600 -29460 6630 -29210
rect 6490 -29480 6630 -29460
rect 8690 -29210 8830 -29180
rect 8690 -29460 8720 -29210
rect 8800 -29460 8830 -29210
rect 8690 -29480 8830 -29460
rect 10890 -29210 11030 -29180
rect 10890 -29460 10920 -29210
rect 11000 -29460 11030 -29210
rect 10890 -29480 11030 -29460
rect 13090 -29210 13230 -29180
rect 13090 -29460 13120 -29210
rect 13200 -29460 13230 -29210
rect 13090 -29480 13230 -29460
rect 15290 -29210 15430 -29180
rect 15290 -29460 15320 -29210
rect 15400 -29460 15430 -29210
rect 15290 -29480 15430 -29460
rect 17490 -29210 17630 -29180
rect 17490 -29460 17520 -29210
rect 17600 -29460 17630 -29210
rect 17490 -29480 17630 -29460
rect 19690 -29210 19830 -29180
rect 19690 -29460 19720 -29210
rect 19800 -29460 19830 -29210
rect 19690 -29480 19830 -29460
rect 21890 -29210 22030 -29180
rect 21890 -29460 21920 -29210
rect 22000 -29460 22030 -29210
rect 21890 -29480 22030 -29460
rect 820 -29550 1020 -29540
rect 20500 -29550 20700 -29540
rect 820 -29560 830 -29550
rect -260 -29620 830 -29560
rect 820 -29630 830 -29620
rect 1010 -29560 1020 -29550
rect 2500 -29560 2700 -29550
rect 3160 -29560 3360 -29550
rect 3820 -29560 4020 -29550
rect 4700 -29560 4900 -29550
rect 5360 -29560 5560 -29550
rect 6020 -29560 6220 -29550
rect 6900 -29560 7100 -29550
rect 7560 -29560 7760 -29550
rect 8220 -29560 8420 -29550
rect 9100 -29560 9300 -29550
rect 9760 -29560 9960 -29550
rect 10420 -29560 10620 -29550
rect 11300 -29560 11500 -29550
rect 11960 -29560 12160 -29550
rect 12620 -29560 12820 -29550
rect 13500 -29560 13700 -29550
rect 14160 -29560 14360 -29550
rect 14820 -29560 15020 -29550
rect 15700 -29560 15900 -29550
rect 16360 -29560 16560 -29550
rect 17020 -29560 17220 -29550
rect 17900 -29560 18100 -29550
rect 18560 -29560 18760 -29550
rect 19220 -29560 19420 -29550
rect 20500 -29560 20510 -29550
rect 1010 -29620 6910 -29560
rect 7090 -29620 7570 -29560
rect 7750 -29620 8230 -29560
rect 8410 -29620 9110 -29560
rect 9290 -29620 9770 -29560
rect 9950 -29620 10430 -29560
rect 10610 -29620 11310 -29560
rect 11490 -29620 11970 -29560
rect 12150 -29620 12630 -29560
rect 12810 -29620 13510 -29560
rect 13690 -29620 14170 -29560
rect 14350 -29620 14830 -29560
rect 15010 -29620 20510 -29560
rect 1010 -29630 1020 -29620
rect 2500 -29630 2700 -29620
rect 3160 -29630 3360 -29620
rect 3820 -29630 4020 -29620
rect 4700 -29630 4900 -29620
rect 5360 -29630 5560 -29620
rect 6020 -29630 6220 -29620
rect 6900 -29630 7100 -29620
rect 7560 -29630 7760 -29620
rect 8220 -29630 8420 -29620
rect 9100 -29630 9300 -29620
rect 9760 -29630 9960 -29620
rect 10420 -29630 10620 -29620
rect 11300 -29630 11500 -29620
rect 11960 -29630 12160 -29620
rect 12620 -29630 12820 -29620
rect 13500 -29630 13700 -29620
rect 14160 -29630 14360 -29620
rect 14820 -29630 15020 -29620
rect 15700 -29630 15900 -29620
rect 16360 -29630 16560 -29620
rect 17020 -29630 17220 -29620
rect 17900 -29630 18100 -29620
rect 18560 -29630 18760 -29620
rect 19220 -29630 19420 -29620
rect 20500 -29630 20510 -29620
rect 20690 -29560 20700 -29550
rect 20690 -29620 22140 -29560
rect 20690 -29630 20700 -29620
rect 820 -29640 1020 -29630
rect 20500 -29640 20700 -29630
rect 1220 -29690 1420 -29680
rect 20900 -29690 21100 -29680
rect 1220 -29700 1230 -29690
rect -260 -29760 1230 -29700
rect 1220 -29770 1230 -29760
rect 1410 -29700 1420 -29690
rect 2500 -29700 2700 -29690
rect 3160 -29700 3360 -29690
rect 3820 -29700 4020 -29690
rect 4700 -29700 4900 -29690
rect 5360 -29700 5560 -29690
rect 6020 -29700 6220 -29690
rect 6900 -29700 7100 -29690
rect 7560 -29700 7760 -29690
rect 8220 -29700 8420 -29690
rect 9100 -29700 9300 -29690
rect 9760 -29700 9960 -29690
rect 10420 -29700 10620 -29690
rect 11300 -29700 11500 -29690
rect 11960 -29700 12160 -29690
rect 12620 -29700 12820 -29690
rect 13500 -29700 13700 -29690
rect 14160 -29700 14360 -29690
rect 14820 -29700 15020 -29690
rect 15700 -29700 15900 -29690
rect 16360 -29700 16560 -29690
rect 17020 -29700 17220 -29690
rect 17900 -29700 18100 -29690
rect 18560 -29700 18760 -29690
rect 19220 -29700 19420 -29690
rect 20900 -29700 20910 -29690
rect 1410 -29760 2510 -29700
rect 2690 -29760 3170 -29700
rect 3350 -29760 3830 -29700
rect 4010 -29760 4710 -29700
rect 4890 -29760 5370 -29700
rect 5550 -29760 6030 -29700
rect 6210 -29760 15710 -29700
rect 15890 -29760 16370 -29700
rect 16550 -29760 17030 -29700
rect 17210 -29760 17910 -29700
rect 18090 -29760 18570 -29700
rect 18750 -29760 19230 -29700
rect 19410 -29760 20910 -29700
rect 1410 -29770 1420 -29760
rect 2500 -29770 2700 -29760
rect 3160 -29770 3360 -29760
rect 3820 -29770 4020 -29760
rect 4700 -29770 4900 -29760
rect 5360 -29770 5560 -29760
rect 6020 -29770 6220 -29760
rect 6900 -29770 7100 -29760
rect 7560 -29770 7760 -29760
rect 8220 -29770 8420 -29760
rect 9100 -29770 9300 -29760
rect 9760 -29770 9960 -29760
rect 10420 -29770 10620 -29760
rect 11300 -29770 11500 -29760
rect 11960 -29770 12160 -29760
rect 12620 -29770 12820 -29760
rect 13500 -29770 13700 -29760
rect 14160 -29770 14360 -29760
rect 14820 -29770 15020 -29760
rect 15700 -29770 15900 -29760
rect 16360 -29770 16560 -29760
rect 17020 -29770 17220 -29760
rect 17900 -29770 18100 -29760
rect 18560 -29770 18760 -29760
rect 19220 -29770 19420 -29760
rect 20900 -29770 20910 -29760
rect 21090 -29700 21100 -29690
rect 21090 -29760 22140 -29700
rect 21090 -29770 21100 -29760
rect 1220 -29780 1420 -29770
rect 20900 -29780 21100 -29770
rect 1620 -29830 1820 -29820
rect 1620 -29840 1630 -29830
rect 1600 -29900 1630 -29840
rect 1620 -29910 1630 -29900
rect 1810 -29840 1820 -29830
rect 20100 -29830 20300 -29820
rect 20100 -29840 20110 -29830
rect 1810 -29870 20110 -29840
rect 1810 -29900 2510 -29870
rect 1810 -29910 1820 -29900
rect 1620 -29920 1820 -29910
rect 2500 -29930 2510 -29900
rect 4010 -29900 4710 -29870
rect 4010 -29930 4020 -29900
rect 2500 -29940 4020 -29930
rect 4700 -29930 4710 -29900
rect 6210 -29900 6910 -29870
rect 6210 -29930 6220 -29900
rect 4700 -29940 6220 -29930
rect 6900 -29930 6910 -29900
rect 8410 -29900 9110 -29870
rect 8410 -29930 8420 -29900
rect 6900 -29940 8420 -29930
rect 9100 -29930 9110 -29900
rect 10610 -29900 11310 -29870
rect 10610 -29930 10620 -29900
rect 9100 -29940 10620 -29930
rect 11300 -29930 11310 -29900
rect 12810 -29900 13510 -29870
rect 12810 -29930 12820 -29900
rect 11300 -29940 12820 -29930
rect 13500 -29930 13510 -29900
rect 15010 -29900 15710 -29870
rect 15010 -29930 15020 -29900
rect 13500 -29940 15020 -29930
rect 15700 -29930 15710 -29900
rect 17210 -29900 17910 -29870
rect 17210 -29930 17220 -29900
rect 15700 -29940 17220 -29930
rect 17900 -29930 17910 -29900
rect 19410 -29900 20110 -29870
rect 19410 -29930 19420 -29900
rect 20100 -29910 20110 -29900
rect 20290 -29840 20300 -29830
rect 20290 -29900 20320 -29840
rect 20290 -29910 20300 -29900
rect 20100 -29920 20300 -29910
rect 17900 -29940 19420 -29930
rect -110 -30010 30 -29980
rect -110 -30260 -80 -30010
rect 0 -30260 30 -30010
rect -110 -30280 30 -30260
rect 2090 -30010 2230 -29980
rect 2090 -30260 2120 -30010
rect 2200 -30260 2230 -30010
rect 2090 -30280 2230 -30260
rect 4290 -30010 4430 -29980
rect 4290 -30260 4320 -30010
rect 4400 -30260 4430 -30010
rect 4290 -30280 4430 -30260
rect 6490 -30010 6630 -29980
rect 6490 -30260 6520 -30010
rect 6600 -30260 6630 -30010
rect 6490 -30280 6630 -30260
rect 8690 -30010 8830 -29980
rect 8690 -30260 8720 -30010
rect 8800 -30260 8830 -30010
rect 8690 -30280 8830 -30260
rect 10890 -30010 11030 -29980
rect 10890 -30260 10920 -30010
rect 11000 -30260 11030 -30010
rect 10890 -30280 11030 -30260
rect 13090 -30010 13230 -29980
rect 13090 -30260 13120 -30010
rect 13200 -30260 13230 -30010
rect 13090 -30280 13230 -30260
rect 15290 -30010 15430 -29980
rect 15290 -30260 15320 -30010
rect 15400 -30260 15430 -30010
rect 15290 -30280 15430 -30260
rect 17490 -30010 17630 -29980
rect 17490 -30260 17520 -30010
rect 17600 -30260 17630 -30010
rect 17490 -30280 17630 -30260
rect 19690 -30010 19830 -29980
rect 19690 -30260 19720 -30010
rect 19800 -30260 19830 -30010
rect 19690 -30280 19830 -30260
rect 21890 -30010 22030 -29980
rect 21890 -30260 21920 -30010
rect 22000 -30260 22030 -30010
rect 21890 -30280 22030 -30260
rect 820 -30350 1020 -30340
rect 20500 -30350 20700 -30340
rect 820 -30360 830 -30350
rect -260 -30420 830 -30360
rect 820 -30430 830 -30420
rect 1010 -30360 1020 -30350
rect 2500 -30360 2700 -30350
rect 3160 -30360 3360 -30350
rect 3820 -30360 4020 -30350
rect 4700 -30360 4900 -30350
rect 5360 -30360 5560 -30350
rect 6020 -30360 6220 -30350
rect 6900 -30360 7100 -30350
rect 7560 -30360 7760 -30350
rect 8220 -30360 8420 -30350
rect 9100 -30360 9300 -30350
rect 9760 -30360 9960 -30350
rect 10420 -30360 10620 -30350
rect 11300 -30360 11500 -30350
rect 11960 -30360 12160 -30350
rect 12620 -30360 12820 -30350
rect 13500 -30360 13700 -30350
rect 14160 -30360 14360 -30350
rect 14820 -30360 15020 -30350
rect 15700 -30360 15900 -30350
rect 16360 -30360 16560 -30350
rect 17020 -30360 17220 -30350
rect 17900 -30360 18100 -30350
rect 18560 -30360 18760 -30350
rect 19220 -30360 19420 -30350
rect 20500 -30360 20510 -30350
rect 1010 -30420 2510 -30360
rect 2690 -30420 3170 -30360
rect 3350 -30420 3830 -30360
rect 4010 -30420 4710 -30360
rect 4890 -30420 5370 -30360
rect 5550 -30420 6030 -30360
rect 6210 -30420 15710 -30360
rect 15890 -30420 16370 -30360
rect 16550 -30420 17030 -30360
rect 17210 -30420 17910 -30360
rect 18090 -30420 18570 -30360
rect 18750 -30420 19230 -30360
rect 19410 -30420 20510 -30360
rect 1010 -30430 1020 -30420
rect 2500 -30430 2700 -30420
rect 3160 -30430 3360 -30420
rect 3820 -30430 4020 -30420
rect 4700 -30430 4900 -30420
rect 5360 -30430 5560 -30420
rect 6020 -30430 6220 -30420
rect 6900 -30430 7100 -30420
rect 7560 -30430 7760 -30420
rect 8220 -30430 8420 -30420
rect 9100 -30430 9300 -30420
rect 9760 -30430 9960 -30420
rect 10420 -30430 10620 -30420
rect 11300 -30430 11500 -30420
rect 11960 -30430 12160 -30420
rect 12620 -30430 12820 -30420
rect 13500 -30430 13700 -30420
rect 14160 -30430 14360 -30420
rect 14820 -30430 15020 -30420
rect 15700 -30430 15900 -30420
rect 16360 -30430 16560 -30420
rect 17020 -30430 17220 -30420
rect 17900 -30430 18100 -30420
rect 18560 -30430 18760 -30420
rect 19220 -30430 19420 -30420
rect 20500 -30430 20510 -30420
rect 20690 -30360 20700 -30350
rect 20690 -30420 22140 -30360
rect 20690 -30430 20700 -30420
rect 820 -30440 1020 -30430
rect 20500 -30440 20700 -30430
rect 1220 -30490 1420 -30480
rect 20900 -30490 21100 -30480
rect 1220 -30500 1230 -30490
rect -260 -30560 1230 -30500
rect 1220 -30570 1230 -30560
rect 1410 -30500 1420 -30490
rect 2500 -30500 2700 -30490
rect 3160 -30500 3360 -30490
rect 3820 -30500 4020 -30490
rect 4700 -30500 4900 -30490
rect 5360 -30500 5560 -30490
rect 6020 -30500 6220 -30490
rect 6900 -30500 7100 -30490
rect 7560 -30500 7760 -30490
rect 8220 -30500 8420 -30490
rect 9100 -30500 9300 -30490
rect 9760 -30500 9960 -30490
rect 10420 -30500 10620 -30490
rect 11300 -30500 11500 -30490
rect 11960 -30500 12160 -30490
rect 12620 -30500 12820 -30490
rect 13500 -30500 13700 -30490
rect 14160 -30500 14360 -30490
rect 14820 -30500 15020 -30490
rect 15700 -30500 15900 -30490
rect 16360 -30500 16560 -30490
rect 17020 -30500 17220 -30490
rect 17900 -30500 18100 -30490
rect 18560 -30500 18760 -30490
rect 19220 -30500 19420 -30490
rect 20900 -30500 20910 -30490
rect 1410 -30560 6910 -30500
rect 7090 -30560 7570 -30500
rect 7750 -30560 8230 -30500
rect 8410 -30560 9110 -30500
rect 9290 -30560 9770 -30500
rect 9950 -30560 10430 -30500
rect 10610 -30560 11310 -30500
rect 11490 -30560 11970 -30500
rect 12150 -30560 12630 -30500
rect 12810 -30560 13510 -30500
rect 13690 -30560 14170 -30500
rect 14350 -30560 14830 -30500
rect 15010 -30560 20910 -30500
rect 1410 -30570 1420 -30560
rect 2500 -30570 2700 -30560
rect 3160 -30570 3360 -30560
rect 3820 -30570 4020 -30560
rect 4700 -30570 4900 -30560
rect 5360 -30570 5560 -30560
rect 6020 -30570 6220 -30560
rect 6900 -30570 7100 -30560
rect 7560 -30570 7760 -30560
rect 8220 -30570 8420 -30560
rect 9100 -30570 9300 -30560
rect 9760 -30570 9960 -30560
rect 10420 -30570 10620 -30560
rect 11300 -30570 11500 -30560
rect 11960 -30570 12160 -30560
rect 12620 -30570 12820 -30560
rect 13500 -30570 13700 -30560
rect 14160 -30570 14360 -30560
rect 14820 -30570 15020 -30560
rect 15700 -30570 15900 -30560
rect 16360 -30570 16560 -30560
rect 17020 -30570 17220 -30560
rect 17900 -30570 18100 -30560
rect 18560 -30570 18760 -30560
rect 19220 -30570 19420 -30560
rect 20900 -30570 20910 -30560
rect 21090 -30500 21100 -30490
rect 21090 -30560 22140 -30500
rect 21090 -30570 21100 -30560
rect 1220 -30580 1420 -30570
rect 20900 -30580 21100 -30570
rect 1620 -30630 1820 -30620
rect 1620 -30640 1630 -30630
rect 1600 -30700 1630 -30640
rect 1620 -30710 1630 -30700
rect 1810 -30640 1820 -30630
rect 20100 -30630 20300 -30620
rect 20100 -30640 20110 -30630
rect 1810 -30670 20110 -30640
rect 1810 -30700 2510 -30670
rect 1810 -30710 1820 -30700
rect 1620 -30720 1820 -30710
rect 2500 -30730 2510 -30700
rect 4010 -30700 4710 -30670
rect 4010 -30730 4020 -30700
rect 2500 -30740 4020 -30730
rect 4700 -30730 4710 -30700
rect 6210 -30700 6910 -30670
rect 6210 -30730 6220 -30700
rect 4700 -30740 6220 -30730
rect 6900 -30730 6910 -30700
rect 8410 -30700 9110 -30670
rect 8410 -30730 8420 -30700
rect 6900 -30740 8420 -30730
rect 9100 -30730 9110 -30700
rect 10610 -30700 11310 -30670
rect 10610 -30730 10620 -30700
rect 9100 -30740 10620 -30730
rect 11300 -30730 11310 -30700
rect 12810 -30700 13510 -30670
rect 12810 -30730 12820 -30700
rect 11300 -30740 12820 -30730
rect 13500 -30730 13510 -30700
rect 15010 -30700 15710 -30670
rect 15010 -30730 15020 -30700
rect 13500 -30740 15020 -30730
rect 15700 -30730 15710 -30700
rect 17210 -30700 17910 -30670
rect 17210 -30730 17220 -30700
rect 15700 -30740 17220 -30730
rect 17900 -30730 17910 -30700
rect 19410 -30700 20110 -30670
rect 19410 -30730 19420 -30700
rect 20100 -30710 20110 -30700
rect 20290 -30640 20300 -30630
rect 20290 -30700 20320 -30640
rect 20290 -30710 20300 -30700
rect 20100 -30720 20300 -30710
rect 17900 -30740 19420 -30730
rect -110 -30810 30 -30780
rect -110 -31060 -80 -30810
rect 0 -31060 30 -30810
rect -110 -31080 30 -31060
rect 2090 -30810 2230 -30780
rect 2090 -31060 2120 -30810
rect 2200 -31060 2230 -30810
rect 2090 -31080 2230 -31060
rect 4290 -30810 4430 -30780
rect 4290 -31060 4320 -30810
rect 4400 -31060 4430 -30810
rect 4290 -31080 4430 -31060
rect 6490 -30810 6630 -30780
rect 6490 -31060 6520 -30810
rect 6600 -31060 6630 -30810
rect 6490 -31080 6630 -31060
rect 8690 -30810 8830 -30780
rect 8690 -31060 8720 -30810
rect 8800 -31060 8830 -30810
rect 8690 -31080 8830 -31060
rect 10890 -30810 11030 -30780
rect 10890 -31060 10920 -30810
rect 11000 -31060 11030 -30810
rect 10890 -31080 11030 -31060
rect 13090 -30810 13230 -30780
rect 13090 -31060 13120 -30810
rect 13200 -31060 13230 -30810
rect 13090 -31080 13230 -31060
rect 15290 -30810 15430 -30780
rect 15290 -31060 15320 -30810
rect 15400 -31060 15430 -30810
rect 15290 -31080 15430 -31060
rect 17490 -30810 17630 -30780
rect 17490 -31060 17520 -30810
rect 17600 -31060 17630 -30810
rect 17490 -31080 17630 -31060
rect 19690 -30810 19830 -30780
rect 19690 -31060 19720 -30810
rect 19800 -31060 19830 -30810
rect 19690 -31080 19830 -31060
rect 21890 -30810 22030 -30780
rect 21890 -31060 21920 -30810
rect 22000 -31060 22030 -30810
rect 21890 -31080 22030 -31060
rect 820 -31150 1020 -31140
rect 20500 -31150 20700 -31140
rect 820 -31160 830 -31150
rect -260 -31220 830 -31160
rect 820 -31230 830 -31220
rect 1010 -31160 1020 -31150
rect 2500 -31160 2700 -31150
rect 3160 -31160 3360 -31150
rect 3820 -31160 4020 -31150
rect 4700 -31160 4900 -31150
rect 5360 -31160 5560 -31150
rect 6020 -31160 6220 -31150
rect 6900 -31160 7100 -31150
rect 7560 -31160 7760 -31150
rect 8220 -31160 8420 -31150
rect 9100 -31160 9300 -31150
rect 9760 -31160 9960 -31150
rect 10420 -31160 10620 -31150
rect 11300 -31160 11500 -31150
rect 11960 -31160 12160 -31150
rect 12620 -31160 12820 -31150
rect 13500 -31160 13700 -31150
rect 14160 -31160 14360 -31150
rect 14820 -31160 15020 -31150
rect 15700 -31160 15900 -31150
rect 16360 -31160 16560 -31150
rect 17020 -31160 17220 -31150
rect 17900 -31160 18100 -31150
rect 18560 -31160 18760 -31150
rect 19220 -31160 19420 -31150
rect 20500 -31160 20510 -31150
rect 1010 -31220 6910 -31160
rect 7090 -31220 7570 -31160
rect 7750 -31220 8230 -31160
rect 8410 -31220 9110 -31160
rect 9290 -31220 9770 -31160
rect 9950 -31220 10430 -31160
rect 10610 -31220 11310 -31160
rect 11490 -31220 11970 -31160
rect 12150 -31220 12630 -31160
rect 12810 -31220 13510 -31160
rect 13690 -31220 14170 -31160
rect 14350 -31220 14830 -31160
rect 15010 -31220 20510 -31160
rect 1010 -31230 1020 -31220
rect 2500 -31230 2700 -31220
rect 3160 -31230 3360 -31220
rect 3820 -31230 4020 -31220
rect 4700 -31230 4900 -31220
rect 5360 -31230 5560 -31220
rect 6020 -31230 6220 -31220
rect 6900 -31230 7100 -31220
rect 7560 -31230 7760 -31220
rect 8220 -31230 8420 -31220
rect 9100 -31230 9300 -31220
rect 9760 -31230 9960 -31220
rect 10420 -31230 10620 -31220
rect 11300 -31230 11500 -31220
rect 11960 -31230 12160 -31220
rect 12620 -31230 12820 -31220
rect 13500 -31230 13700 -31220
rect 14160 -31230 14360 -31220
rect 14820 -31230 15020 -31220
rect 15700 -31230 15900 -31220
rect 16360 -31230 16560 -31220
rect 17020 -31230 17220 -31220
rect 17900 -31230 18100 -31220
rect 18560 -31230 18760 -31220
rect 19220 -31230 19420 -31220
rect 20500 -31230 20510 -31220
rect 20690 -31160 20700 -31150
rect 20690 -31220 22140 -31160
rect 20690 -31230 20700 -31220
rect 820 -31240 1020 -31230
rect 20500 -31240 20700 -31230
rect 1220 -31290 1420 -31280
rect 20900 -31290 21100 -31280
rect 1220 -31300 1230 -31290
rect -260 -31360 1230 -31300
rect 1220 -31370 1230 -31360
rect 1410 -31300 1420 -31290
rect 2500 -31300 2700 -31290
rect 3160 -31300 3360 -31290
rect 3820 -31300 4020 -31290
rect 4700 -31300 4900 -31290
rect 5360 -31300 5560 -31290
rect 6020 -31300 6220 -31290
rect 6900 -31300 7100 -31290
rect 7560 -31300 7760 -31290
rect 8220 -31300 8420 -31290
rect 9100 -31300 9300 -31290
rect 9760 -31300 9960 -31290
rect 10420 -31300 10620 -31290
rect 11300 -31300 11500 -31290
rect 11960 -31300 12160 -31290
rect 12620 -31300 12820 -31290
rect 13500 -31300 13700 -31290
rect 14160 -31300 14360 -31290
rect 14820 -31300 15020 -31290
rect 15700 -31300 15900 -31290
rect 16360 -31300 16560 -31290
rect 17020 -31300 17220 -31290
rect 17900 -31300 18100 -31290
rect 18560 -31300 18760 -31290
rect 19220 -31300 19420 -31290
rect 20900 -31300 20910 -31290
rect 1410 -31360 2510 -31300
rect 2690 -31360 3170 -31300
rect 3350 -31360 3830 -31300
rect 4010 -31360 4710 -31300
rect 4890 -31360 5370 -31300
rect 5550 -31360 6030 -31300
rect 6210 -31360 15710 -31300
rect 15890 -31360 16370 -31300
rect 16550 -31360 17030 -31300
rect 17210 -31360 17910 -31300
rect 18090 -31360 18570 -31300
rect 18750 -31360 19230 -31300
rect 19410 -31360 20910 -31300
rect 1410 -31370 1420 -31360
rect 2500 -31370 2700 -31360
rect 3160 -31370 3360 -31360
rect 3820 -31370 4020 -31360
rect 4700 -31370 4900 -31360
rect 5360 -31370 5560 -31360
rect 6020 -31370 6220 -31360
rect 6900 -31370 7100 -31360
rect 7560 -31370 7760 -31360
rect 8220 -31370 8420 -31360
rect 9100 -31370 9300 -31360
rect 9760 -31370 9960 -31360
rect 10420 -31370 10620 -31360
rect 11300 -31370 11500 -31360
rect 11960 -31370 12160 -31360
rect 12620 -31370 12820 -31360
rect 13500 -31370 13700 -31360
rect 14160 -31370 14360 -31360
rect 14820 -31370 15020 -31360
rect 15700 -31370 15900 -31360
rect 16360 -31370 16560 -31360
rect 17020 -31370 17220 -31360
rect 17900 -31370 18100 -31360
rect 18560 -31370 18760 -31360
rect 19220 -31370 19420 -31360
rect 20900 -31370 20910 -31360
rect 21090 -31300 21100 -31290
rect 21090 -31360 22140 -31300
rect 21090 -31370 21100 -31360
rect 1220 -31380 1420 -31370
rect 20900 -31380 21100 -31370
<< via3 >>
rect 830 11170 1010 11250
rect 20510 11170 20690 11250
rect 1230 11030 1410 11110
rect 20910 11030 21090 11110
rect -80 10930 0 10940
rect -80 10870 -70 10930
rect -70 10870 -10 10930
rect -10 10870 0 10930
rect -80 10690 0 10870
rect 2120 10930 2200 10940
rect 2120 10870 2130 10930
rect 2130 10870 2190 10930
rect 2190 10870 2200 10930
rect 2120 10690 2200 10870
rect 4320 10930 4400 10940
rect 4320 10870 4330 10930
rect 4330 10870 4390 10930
rect 4390 10870 4400 10930
rect 4320 10690 4400 10870
rect 6520 10930 6600 10940
rect 6520 10870 6530 10930
rect 6530 10870 6590 10930
rect 6590 10870 6600 10930
rect 6520 10690 6600 10870
rect 8720 10930 8800 10940
rect 8720 10870 8730 10930
rect 8730 10870 8790 10930
rect 8790 10870 8800 10930
rect 8720 10690 8800 10870
rect 10920 10930 11000 10940
rect 10920 10870 10930 10930
rect 10930 10870 10990 10930
rect 10990 10870 11000 10930
rect 10920 10690 11000 10870
rect 13120 10930 13200 10940
rect 13120 10870 13130 10930
rect 13130 10870 13190 10930
rect 13190 10870 13200 10930
rect 13120 10690 13200 10870
rect 15320 10930 15400 10940
rect 15320 10870 15330 10930
rect 15330 10870 15390 10930
rect 15390 10870 15400 10930
rect 15320 10690 15400 10870
rect 17520 10930 17600 10940
rect 17520 10870 17530 10930
rect 17530 10870 17590 10930
rect 17590 10870 17600 10930
rect 17520 10690 17600 10870
rect 19720 10930 19800 10940
rect 19720 10870 19730 10930
rect 19730 10870 19790 10930
rect 19790 10870 19800 10930
rect 19720 10690 19800 10870
rect 21920 10930 22000 10940
rect 21920 10870 21930 10930
rect 21930 10870 21990 10930
rect 21990 10870 22000 10930
rect 21920 10690 22000 10870
rect 1630 10510 1810 10590
rect 20110 10510 20290 10590
rect 830 10370 1010 10450
rect 20510 10370 20690 10450
rect 1230 10230 1410 10310
rect 20910 10230 21090 10310
rect -80 10130 0 10140
rect -80 10070 -70 10130
rect -70 10070 -10 10130
rect -10 10070 0 10130
rect -80 9890 0 10070
rect 2120 10130 2200 10140
rect 2120 10070 2130 10130
rect 2130 10070 2190 10130
rect 2190 10070 2200 10130
rect 2120 9890 2200 10070
rect 4320 10130 4400 10140
rect 4320 10070 4330 10130
rect 4330 10070 4390 10130
rect 4390 10070 4400 10130
rect 4320 9890 4400 10070
rect 6520 10130 6600 10140
rect 6520 10070 6530 10130
rect 6530 10070 6590 10130
rect 6590 10070 6600 10130
rect 6520 9890 6600 10070
rect 8720 10130 8800 10140
rect 8720 10070 8730 10130
rect 8730 10070 8790 10130
rect 8790 10070 8800 10130
rect 8720 9890 8800 10070
rect 10920 10130 11000 10140
rect 10920 10070 10930 10130
rect 10930 10070 10990 10130
rect 10990 10070 11000 10130
rect 10920 9890 11000 10070
rect 13120 10130 13200 10140
rect 13120 10070 13130 10130
rect 13130 10070 13190 10130
rect 13190 10070 13200 10130
rect 13120 9890 13200 10070
rect 15320 10130 15400 10140
rect 15320 10070 15330 10130
rect 15330 10070 15390 10130
rect 15390 10070 15400 10130
rect 15320 9890 15400 10070
rect 17520 10130 17600 10140
rect 17520 10070 17530 10130
rect 17530 10070 17590 10130
rect 17590 10070 17600 10130
rect 17520 9890 17600 10070
rect 19720 10130 19800 10140
rect 19720 10070 19730 10130
rect 19730 10070 19790 10130
rect 19790 10070 19800 10130
rect 19720 9890 19800 10070
rect 21920 10130 22000 10140
rect 21920 10070 21930 10130
rect 21930 10070 21990 10130
rect 21990 10070 22000 10130
rect 21920 9890 22000 10070
rect 1630 9710 1810 9790
rect 20110 9710 20290 9790
rect 830 9570 1010 9650
rect 20510 9570 20690 9650
rect 1230 9430 1410 9510
rect 20910 9430 21090 9510
rect -80 9330 0 9340
rect -80 9270 -70 9330
rect -70 9270 -10 9330
rect -10 9270 0 9330
rect -80 9090 0 9270
rect 2120 9330 2200 9340
rect 2120 9270 2130 9330
rect 2130 9270 2190 9330
rect 2190 9270 2200 9330
rect 2120 9090 2200 9270
rect 4320 9330 4400 9340
rect 4320 9270 4330 9330
rect 4330 9270 4390 9330
rect 4390 9270 4400 9330
rect 4320 9090 4400 9270
rect 6520 9330 6600 9340
rect 6520 9270 6530 9330
rect 6530 9270 6590 9330
rect 6590 9270 6600 9330
rect 6520 9090 6600 9270
rect 8720 9330 8800 9340
rect 8720 9270 8730 9330
rect 8730 9270 8790 9330
rect 8790 9270 8800 9330
rect 8720 9090 8800 9270
rect 10920 9330 11000 9340
rect 10920 9270 10930 9330
rect 10930 9270 10990 9330
rect 10990 9270 11000 9330
rect 10920 9090 11000 9270
rect 13120 9330 13200 9340
rect 13120 9270 13130 9330
rect 13130 9270 13190 9330
rect 13190 9270 13200 9330
rect 13120 9090 13200 9270
rect 15320 9330 15400 9340
rect 15320 9270 15330 9330
rect 15330 9270 15390 9330
rect 15390 9270 15400 9330
rect 15320 9090 15400 9270
rect 17520 9330 17600 9340
rect 17520 9270 17530 9330
rect 17530 9270 17590 9330
rect 17590 9270 17600 9330
rect 17520 9090 17600 9270
rect 19720 9330 19800 9340
rect 19720 9270 19730 9330
rect 19730 9270 19790 9330
rect 19790 9270 19800 9330
rect 19720 9090 19800 9270
rect 21920 9330 22000 9340
rect 21920 9270 21930 9330
rect 21930 9270 21990 9330
rect 21990 9270 22000 9330
rect 21920 9090 22000 9270
rect 430 8910 610 8990
rect 1630 8910 1810 8990
rect 20110 8910 20290 8990
rect 21310 8910 21490 8990
rect 830 8770 1010 8850
rect 20510 8770 20690 8850
rect 1230 8630 1410 8710
rect 20910 8630 21090 8710
rect -80 8530 0 8540
rect -80 8470 -70 8530
rect -70 8470 -10 8530
rect -10 8470 0 8530
rect -80 8290 0 8470
rect 2120 8530 2200 8540
rect 2120 8470 2130 8530
rect 2130 8470 2190 8530
rect 2190 8470 2200 8530
rect 2120 8290 2200 8470
rect 4320 8530 4400 8540
rect 4320 8470 4330 8530
rect 4330 8470 4390 8530
rect 4390 8470 4400 8530
rect 4320 8290 4400 8470
rect 6520 8530 6600 8540
rect 6520 8470 6530 8530
rect 6530 8470 6590 8530
rect 6590 8470 6600 8530
rect 6520 8290 6600 8470
rect 8720 8530 8800 8540
rect 8720 8470 8730 8530
rect 8730 8470 8790 8530
rect 8790 8470 8800 8530
rect 8720 8290 8800 8470
rect 10920 8530 11000 8540
rect 10920 8470 10930 8530
rect 10930 8470 10990 8530
rect 10990 8470 11000 8530
rect 10920 8290 11000 8470
rect 13120 8530 13200 8540
rect 13120 8470 13130 8530
rect 13130 8470 13190 8530
rect 13190 8470 13200 8530
rect 13120 8290 13200 8470
rect 15320 8530 15400 8540
rect 15320 8470 15330 8530
rect 15330 8470 15390 8530
rect 15390 8470 15400 8530
rect 15320 8290 15400 8470
rect 17520 8530 17600 8540
rect 17520 8470 17530 8530
rect 17530 8470 17590 8530
rect 17590 8470 17600 8530
rect 17520 8290 17600 8470
rect 19720 8530 19800 8540
rect 19720 8470 19730 8530
rect 19730 8470 19790 8530
rect 19790 8470 19800 8530
rect 19720 8290 19800 8470
rect 21920 8530 22000 8540
rect 21920 8470 21930 8530
rect 21930 8470 21990 8530
rect 21990 8470 22000 8530
rect 21920 8290 22000 8470
rect 430 8110 610 8190
rect 1630 8110 1810 8190
rect 20110 8110 20290 8190
rect 21310 8110 21490 8190
rect 830 7970 1010 8050
rect 20510 7970 20690 8050
rect 1230 7830 1410 7910
rect 20910 7830 21090 7910
rect -80 7730 0 7740
rect -80 7670 -70 7730
rect -70 7670 -10 7730
rect -10 7670 0 7730
rect -80 7490 0 7670
rect 2120 7730 2200 7740
rect 2120 7670 2130 7730
rect 2130 7670 2190 7730
rect 2190 7670 2200 7730
rect 2120 7490 2200 7670
rect 4320 7730 4400 7740
rect 4320 7670 4330 7730
rect 4330 7670 4390 7730
rect 4390 7670 4400 7730
rect 4320 7490 4400 7670
rect 6520 7730 6600 7740
rect 6520 7670 6530 7730
rect 6530 7670 6590 7730
rect 6590 7670 6600 7730
rect 6520 7490 6600 7670
rect 8720 7730 8800 7740
rect 8720 7670 8730 7730
rect 8730 7670 8790 7730
rect 8790 7670 8800 7730
rect 8720 7490 8800 7670
rect 10920 7730 11000 7740
rect 10920 7670 10930 7730
rect 10930 7670 10990 7730
rect 10990 7670 11000 7730
rect 10920 7490 11000 7670
rect 13120 7730 13200 7740
rect 13120 7670 13130 7730
rect 13130 7670 13190 7730
rect 13190 7670 13200 7730
rect 13120 7490 13200 7670
rect 15320 7730 15400 7740
rect 15320 7670 15330 7730
rect 15330 7670 15390 7730
rect 15390 7670 15400 7730
rect 15320 7490 15400 7670
rect 17520 7730 17600 7740
rect 17520 7670 17530 7730
rect 17530 7670 17590 7730
rect 17590 7670 17600 7730
rect 17520 7490 17600 7670
rect 19720 7730 19800 7740
rect 19720 7670 19730 7730
rect 19730 7670 19790 7730
rect 19790 7670 19800 7730
rect 19720 7490 19800 7670
rect 21920 7730 22000 7740
rect 21920 7670 21930 7730
rect 21930 7670 21990 7730
rect 21990 7670 22000 7730
rect 21920 7490 22000 7670
rect 430 7310 610 7390
rect 1630 7310 1810 7390
rect 20110 7310 20290 7390
rect 21310 7310 21490 7390
rect 830 7170 1010 7250
rect 20510 7170 20690 7250
rect 1230 7030 1410 7110
rect 20910 7030 21090 7110
rect -80 6930 0 6940
rect -80 6870 -70 6930
rect -70 6870 -10 6930
rect -10 6870 0 6930
rect -80 6690 0 6870
rect 2120 6930 2200 6940
rect 2120 6870 2130 6930
rect 2130 6870 2190 6930
rect 2190 6870 2200 6930
rect 2120 6690 2200 6870
rect 4320 6930 4400 6940
rect 4320 6870 4330 6930
rect 4330 6870 4390 6930
rect 4390 6870 4400 6930
rect 4320 6690 4400 6870
rect 6520 6930 6600 6940
rect 6520 6870 6530 6930
rect 6530 6870 6590 6930
rect 6590 6870 6600 6930
rect 6520 6690 6600 6870
rect 8720 6930 8800 6940
rect 8720 6870 8730 6930
rect 8730 6870 8790 6930
rect 8790 6870 8800 6930
rect 8720 6690 8800 6870
rect 10920 6930 11000 6940
rect 10920 6870 10930 6930
rect 10930 6870 10990 6930
rect 10990 6870 11000 6930
rect 10920 6690 11000 6870
rect 13120 6930 13200 6940
rect 13120 6870 13130 6930
rect 13130 6870 13190 6930
rect 13190 6870 13200 6930
rect 13120 6690 13200 6870
rect 15320 6930 15400 6940
rect 15320 6870 15330 6930
rect 15330 6870 15390 6930
rect 15390 6870 15400 6930
rect 15320 6690 15400 6870
rect 17520 6930 17600 6940
rect 17520 6870 17530 6930
rect 17530 6870 17590 6930
rect 17590 6870 17600 6930
rect 17520 6690 17600 6870
rect 19720 6930 19800 6940
rect 19720 6870 19730 6930
rect 19730 6870 19790 6930
rect 19790 6870 19800 6930
rect 19720 6690 19800 6870
rect 21920 6930 22000 6940
rect 21920 6870 21930 6930
rect 21930 6870 21990 6930
rect 21990 6870 22000 6930
rect 21920 6690 22000 6870
rect 430 6510 610 6590
rect 1630 6510 1810 6590
rect 20110 6510 20290 6590
rect 21310 6510 21490 6590
rect 830 6370 1010 6450
rect 20510 6370 20690 6450
rect 1230 6230 1410 6310
rect 20910 6230 21090 6310
rect -80 6130 0 6140
rect -80 6070 -70 6130
rect -70 6070 -10 6130
rect -10 6070 0 6130
rect -80 5890 0 6070
rect 2120 6130 2200 6140
rect 2120 6070 2130 6130
rect 2130 6070 2190 6130
rect 2190 6070 2200 6130
rect 2120 5890 2200 6070
rect 4320 6130 4400 6140
rect 4320 6070 4330 6130
rect 4330 6070 4390 6130
rect 4390 6070 4400 6130
rect 4320 5890 4400 6070
rect 6520 6130 6600 6140
rect 6520 6070 6530 6130
rect 6530 6070 6590 6130
rect 6590 6070 6600 6130
rect 6520 5890 6600 6070
rect 8720 6130 8800 6140
rect 8720 6070 8730 6130
rect 8730 6070 8790 6130
rect 8790 6070 8800 6130
rect 8720 5890 8800 6070
rect 10920 6130 11000 6140
rect 10920 6070 10930 6130
rect 10930 6070 10990 6130
rect 10990 6070 11000 6130
rect 10920 5890 11000 6070
rect 13120 6130 13200 6140
rect 13120 6070 13130 6130
rect 13130 6070 13190 6130
rect 13190 6070 13200 6130
rect 13120 5890 13200 6070
rect 15320 6130 15400 6140
rect 15320 6070 15330 6130
rect 15330 6070 15390 6130
rect 15390 6070 15400 6130
rect 15320 5890 15400 6070
rect 17520 6130 17600 6140
rect 17520 6070 17530 6130
rect 17530 6070 17590 6130
rect 17590 6070 17600 6130
rect 17520 5890 17600 6070
rect 19720 6130 19800 6140
rect 19720 6070 19730 6130
rect 19730 6070 19790 6130
rect 19790 6070 19800 6130
rect 19720 5890 19800 6070
rect 21920 6130 22000 6140
rect 21920 6070 21930 6130
rect 21930 6070 21990 6130
rect 21990 6070 22000 6130
rect 21920 5890 22000 6070
rect 1630 5710 1810 5790
rect 20110 5710 20290 5790
rect 830 5570 1010 5650
rect 20510 5570 20690 5650
rect 1230 5430 1410 5510
rect 20910 5430 21090 5510
rect -80 5330 0 5340
rect -80 5270 -70 5330
rect -70 5270 -10 5330
rect -10 5270 0 5330
rect -80 5090 0 5270
rect 2120 5330 2200 5340
rect 2120 5270 2130 5330
rect 2130 5270 2190 5330
rect 2190 5270 2200 5330
rect 2120 5090 2200 5270
rect 4320 5330 4400 5340
rect 4320 5270 4330 5330
rect 4330 5270 4390 5330
rect 4390 5270 4400 5330
rect 4320 5090 4400 5270
rect 6520 5330 6600 5340
rect 6520 5270 6530 5330
rect 6530 5270 6590 5330
rect 6590 5270 6600 5330
rect 6520 5090 6600 5270
rect 8720 5330 8800 5340
rect 8720 5270 8730 5330
rect 8730 5270 8790 5330
rect 8790 5270 8800 5330
rect 8720 5090 8800 5270
rect 10920 5330 11000 5340
rect 10920 5270 10930 5330
rect 10930 5270 10990 5330
rect 10990 5270 11000 5330
rect 10920 5090 11000 5270
rect 13120 5330 13200 5340
rect 13120 5270 13130 5330
rect 13130 5270 13190 5330
rect 13190 5270 13200 5330
rect 13120 5090 13200 5270
rect 15320 5330 15400 5340
rect 15320 5270 15330 5330
rect 15330 5270 15390 5330
rect 15390 5270 15400 5330
rect 15320 5090 15400 5270
rect 17520 5330 17600 5340
rect 17520 5270 17530 5330
rect 17530 5270 17590 5330
rect 17590 5270 17600 5330
rect 17520 5090 17600 5270
rect 19720 5330 19800 5340
rect 19720 5270 19730 5330
rect 19730 5270 19790 5330
rect 19790 5270 19800 5330
rect 19720 5090 19800 5270
rect 21920 5330 22000 5340
rect 21920 5270 21930 5330
rect 21930 5270 21990 5330
rect 21990 5270 22000 5330
rect 21920 5090 22000 5270
rect 1630 4910 1810 4990
rect 20110 4910 20290 4990
rect 430 3550 610 3730
rect 21310 3550 21490 3730
rect 1630 3150 1810 3330
rect 20110 3150 20290 3330
rect 14910 1300 15030 1960
rect 1630 -5350 1810 -5170
rect 20910 -5350 21090 -5170
rect 830 -5750 1010 -5570
rect 20510 -5750 20690 -5570
rect 14910 -6610 15030 -6490
rect 830 -7350 1010 -7170
rect 20510 -7350 20530 -7170
rect 20530 -7350 20690 -7170
rect 1230 -7750 1410 -7570
rect 22070 -7750 22250 -7570
rect 1630 -23450 1810 -23270
rect 20110 -23450 20290 -23270
rect 430 -23850 610 -23670
rect 21310 -23850 21490 -23670
rect 1630 -25110 1810 -25030
rect 20110 -25110 20290 -25030
rect -80 -25390 0 -25210
rect -80 -25450 -70 -25390
rect -70 -25450 -10 -25390
rect -10 -25450 0 -25390
rect -80 -25460 0 -25450
rect 2120 -25390 2200 -25210
rect 2120 -25450 2130 -25390
rect 2130 -25450 2190 -25390
rect 2190 -25450 2200 -25390
rect 2120 -25460 2200 -25450
rect 4320 -25390 4400 -25210
rect 4320 -25450 4330 -25390
rect 4330 -25450 4390 -25390
rect 4390 -25450 4400 -25390
rect 4320 -25460 4400 -25450
rect 6520 -25390 6600 -25210
rect 6520 -25450 6530 -25390
rect 6530 -25450 6590 -25390
rect 6590 -25450 6600 -25390
rect 6520 -25460 6600 -25450
rect 8720 -25390 8800 -25210
rect 8720 -25450 8730 -25390
rect 8730 -25450 8790 -25390
rect 8790 -25450 8800 -25390
rect 8720 -25460 8800 -25450
rect 10920 -25390 11000 -25210
rect 10920 -25450 10930 -25390
rect 10930 -25450 10990 -25390
rect 10990 -25450 11000 -25390
rect 10920 -25460 11000 -25450
rect 13120 -25390 13200 -25210
rect 13120 -25450 13130 -25390
rect 13130 -25450 13190 -25390
rect 13190 -25450 13200 -25390
rect 13120 -25460 13200 -25450
rect 15320 -25390 15400 -25210
rect 15320 -25450 15330 -25390
rect 15330 -25450 15390 -25390
rect 15390 -25450 15400 -25390
rect 15320 -25460 15400 -25450
rect 17520 -25390 17600 -25210
rect 17520 -25450 17530 -25390
rect 17530 -25450 17590 -25390
rect 17590 -25450 17600 -25390
rect 17520 -25460 17600 -25450
rect 19720 -25390 19800 -25210
rect 19720 -25450 19730 -25390
rect 19730 -25450 19790 -25390
rect 19790 -25450 19800 -25390
rect 19720 -25460 19800 -25450
rect 21920 -25390 22000 -25210
rect 21920 -25450 21930 -25390
rect 21930 -25450 21990 -25390
rect 21990 -25450 22000 -25390
rect 21920 -25460 22000 -25450
rect 830 -25630 1010 -25550
rect 20510 -25630 20690 -25550
rect 1230 -25770 1410 -25690
rect 20910 -25770 21090 -25690
rect 1630 -25910 1810 -25830
rect 20110 -25910 20290 -25830
rect -80 -26190 0 -26010
rect -80 -26250 -70 -26190
rect -70 -26250 -10 -26190
rect -10 -26250 0 -26190
rect -80 -26260 0 -26250
rect 2120 -26190 2200 -26010
rect 2120 -26250 2130 -26190
rect 2130 -26250 2190 -26190
rect 2190 -26250 2200 -26190
rect 2120 -26260 2200 -26250
rect 4320 -26190 4400 -26010
rect 4320 -26250 4330 -26190
rect 4330 -26250 4390 -26190
rect 4390 -26250 4400 -26190
rect 4320 -26260 4400 -26250
rect 6520 -26190 6600 -26010
rect 6520 -26250 6530 -26190
rect 6530 -26250 6590 -26190
rect 6590 -26250 6600 -26190
rect 6520 -26260 6600 -26250
rect 8720 -26190 8800 -26010
rect 8720 -26250 8730 -26190
rect 8730 -26250 8790 -26190
rect 8790 -26250 8800 -26190
rect 8720 -26260 8800 -26250
rect 10920 -26190 11000 -26010
rect 10920 -26250 10930 -26190
rect 10930 -26250 10990 -26190
rect 10990 -26250 11000 -26190
rect 10920 -26260 11000 -26250
rect 13120 -26190 13200 -26010
rect 13120 -26250 13130 -26190
rect 13130 -26250 13190 -26190
rect 13190 -26250 13200 -26190
rect 13120 -26260 13200 -26250
rect 15320 -26190 15400 -26010
rect 15320 -26250 15330 -26190
rect 15330 -26250 15390 -26190
rect 15390 -26250 15400 -26190
rect 15320 -26260 15400 -26250
rect 17520 -26190 17600 -26010
rect 17520 -26250 17530 -26190
rect 17530 -26250 17590 -26190
rect 17590 -26250 17600 -26190
rect 17520 -26260 17600 -26250
rect 19720 -26190 19800 -26010
rect 19720 -26250 19730 -26190
rect 19730 -26250 19790 -26190
rect 19790 -26250 19800 -26190
rect 19720 -26260 19800 -26250
rect 21920 -26190 22000 -26010
rect 21920 -26250 21930 -26190
rect 21930 -26250 21990 -26190
rect 21990 -26250 22000 -26190
rect 21920 -26260 22000 -26250
rect 830 -26430 1010 -26350
rect 20510 -26430 20690 -26350
rect 1230 -26570 1410 -26490
rect 20910 -26570 21090 -26490
rect 430 -26710 610 -26630
rect 1630 -26710 1810 -26630
rect 20110 -26710 20290 -26630
rect 21310 -26710 21490 -26630
rect -80 -26990 0 -26810
rect -80 -27050 -70 -26990
rect -70 -27050 -10 -26990
rect -10 -27050 0 -26990
rect -80 -27060 0 -27050
rect 2120 -26990 2200 -26810
rect 2120 -27050 2130 -26990
rect 2130 -27050 2190 -26990
rect 2190 -27050 2200 -26990
rect 2120 -27060 2200 -27050
rect 4320 -26990 4400 -26810
rect 4320 -27050 4330 -26990
rect 4330 -27050 4390 -26990
rect 4390 -27050 4400 -26990
rect 4320 -27060 4400 -27050
rect 6520 -26990 6600 -26810
rect 6520 -27050 6530 -26990
rect 6530 -27050 6590 -26990
rect 6590 -27050 6600 -26990
rect 6520 -27060 6600 -27050
rect 8720 -26990 8800 -26810
rect 8720 -27050 8730 -26990
rect 8730 -27050 8790 -26990
rect 8790 -27050 8800 -26990
rect 8720 -27060 8800 -27050
rect 10920 -26990 11000 -26810
rect 10920 -27050 10930 -26990
rect 10930 -27050 10990 -26990
rect 10990 -27050 11000 -26990
rect 10920 -27060 11000 -27050
rect 13120 -26990 13200 -26810
rect 13120 -27050 13130 -26990
rect 13130 -27050 13190 -26990
rect 13190 -27050 13200 -26990
rect 13120 -27060 13200 -27050
rect 15320 -26990 15400 -26810
rect 15320 -27050 15330 -26990
rect 15330 -27050 15390 -26990
rect 15390 -27050 15400 -26990
rect 15320 -27060 15400 -27050
rect 17520 -26990 17600 -26810
rect 17520 -27050 17530 -26990
rect 17530 -27050 17590 -26990
rect 17590 -27050 17600 -26990
rect 17520 -27060 17600 -27050
rect 19720 -26990 19800 -26810
rect 19720 -27050 19730 -26990
rect 19730 -27050 19790 -26990
rect 19790 -27050 19800 -26990
rect 19720 -27060 19800 -27050
rect 21920 -26990 22000 -26810
rect 21920 -27050 21930 -26990
rect 21930 -27050 21990 -26990
rect 21990 -27050 22000 -26990
rect 21920 -27060 22000 -27050
rect 830 -27230 1010 -27150
rect 20510 -27230 20690 -27150
rect 1230 -27370 1410 -27290
rect 20910 -27370 21090 -27290
rect 430 -27510 610 -27430
rect 1630 -27510 1810 -27430
rect 20110 -27510 20290 -27430
rect 21310 -27510 21490 -27430
rect -80 -27790 0 -27610
rect -80 -27850 -70 -27790
rect -70 -27850 -10 -27790
rect -10 -27850 0 -27790
rect -80 -27860 0 -27850
rect 2120 -27790 2200 -27610
rect 2120 -27850 2130 -27790
rect 2130 -27850 2190 -27790
rect 2190 -27850 2200 -27790
rect 2120 -27860 2200 -27850
rect 4320 -27790 4400 -27610
rect 4320 -27850 4330 -27790
rect 4330 -27850 4390 -27790
rect 4390 -27850 4400 -27790
rect 4320 -27860 4400 -27850
rect 6520 -27790 6600 -27610
rect 6520 -27850 6530 -27790
rect 6530 -27850 6590 -27790
rect 6590 -27850 6600 -27790
rect 6520 -27860 6600 -27850
rect 8720 -27790 8800 -27610
rect 8720 -27850 8730 -27790
rect 8730 -27850 8790 -27790
rect 8790 -27850 8800 -27790
rect 8720 -27860 8800 -27850
rect 10920 -27790 11000 -27610
rect 10920 -27850 10930 -27790
rect 10930 -27850 10990 -27790
rect 10990 -27850 11000 -27790
rect 10920 -27860 11000 -27850
rect 13120 -27790 13200 -27610
rect 13120 -27850 13130 -27790
rect 13130 -27850 13190 -27790
rect 13190 -27850 13200 -27790
rect 13120 -27860 13200 -27850
rect 15320 -27790 15400 -27610
rect 15320 -27850 15330 -27790
rect 15330 -27850 15390 -27790
rect 15390 -27850 15400 -27790
rect 15320 -27860 15400 -27850
rect 17520 -27790 17600 -27610
rect 17520 -27850 17530 -27790
rect 17530 -27850 17590 -27790
rect 17590 -27850 17600 -27790
rect 17520 -27860 17600 -27850
rect 19720 -27790 19800 -27610
rect 19720 -27850 19730 -27790
rect 19730 -27850 19790 -27790
rect 19790 -27850 19800 -27790
rect 19720 -27860 19800 -27850
rect 21920 -27790 22000 -27610
rect 21920 -27850 21930 -27790
rect 21930 -27850 21990 -27790
rect 21990 -27850 22000 -27790
rect 21920 -27860 22000 -27850
rect 830 -28030 1010 -27950
rect 20510 -28030 20690 -27950
rect 1230 -28170 1410 -28090
rect 20910 -28170 21090 -28090
rect 430 -28310 610 -28230
rect 1630 -28310 1810 -28230
rect 20110 -28310 20290 -28230
rect 21310 -28310 21490 -28230
rect -80 -28590 0 -28410
rect -80 -28650 -70 -28590
rect -70 -28650 -10 -28590
rect -10 -28650 0 -28590
rect -80 -28660 0 -28650
rect 2120 -28590 2200 -28410
rect 2120 -28650 2130 -28590
rect 2130 -28650 2190 -28590
rect 2190 -28650 2200 -28590
rect 2120 -28660 2200 -28650
rect 4320 -28590 4400 -28410
rect 4320 -28650 4330 -28590
rect 4330 -28650 4390 -28590
rect 4390 -28650 4400 -28590
rect 4320 -28660 4400 -28650
rect 6520 -28590 6600 -28410
rect 6520 -28650 6530 -28590
rect 6530 -28650 6590 -28590
rect 6590 -28650 6600 -28590
rect 6520 -28660 6600 -28650
rect 8720 -28590 8800 -28410
rect 8720 -28650 8730 -28590
rect 8730 -28650 8790 -28590
rect 8790 -28650 8800 -28590
rect 8720 -28660 8800 -28650
rect 10920 -28590 11000 -28410
rect 10920 -28650 10930 -28590
rect 10930 -28650 10990 -28590
rect 10990 -28650 11000 -28590
rect 10920 -28660 11000 -28650
rect 13120 -28590 13200 -28410
rect 13120 -28650 13130 -28590
rect 13130 -28650 13190 -28590
rect 13190 -28650 13200 -28590
rect 13120 -28660 13200 -28650
rect 15320 -28590 15400 -28410
rect 15320 -28650 15330 -28590
rect 15330 -28650 15390 -28590
rect 15390 -28650 15400 -28590
rect 15320 -28660 15400 -28650
rect 17520 -28590 17600 -28410
rect 17520 -28650 17530 -28590
rect 17530 -28650 17590 -28590
rect 17590 -28650 17600 -28590
rect 17520 -28660 17600 -28650
rect 19720 -28590 19800 -28410
rect 19720 -28650 19730 -28590
rect 19730 -28650 19790 -28590
rect 19790 -28650 19800 -28590
rect 19720 -28660 19800 -28650
rect 21920 -28590 22000 -28410
rect 21920 -28650 21930 -28590
rect 21930 -28650 21990 -28590
rect 21990 -28650 22000 -28590
rect 21920 -28660 22000 -28650
rect 830 -28830 1010 -28750
rect 20510 -28830 20690 -28750
rect 1230 -28970 1410 -28890
rect 20910 -28970 21090 -28890
rect 430 -29110 610 -29030
rect 1630 -29110 1810 -29030
rect 20110 -29110 20290 -29030
rect 21310 -29110 21490 -29030
rect -80 -29390 0 -29210
rect -80 -29450 -70 -29390
rect -70 -29450 -10 -29390
rect -10 -29450 0 -29390
rect -80 -29460 0 -29450
rect 2120 -29390 2200 -29210
rect 2120 -29450 2130 -29390
rect 2130 -29450 2190 -29390
rect 2190 -29450 2200 -29390
rect 2120 -29460 2200 -29450
rect 4320 -29390 4400 -29210
rect 4320 -29450 4330 -29390
rect 4330 -29450 4390 -29390
rect 4390 -29450 4400 -29390
rect 4320 -29460 4400 -29450
rect 6520 -29390 6600 -29210
rect 6520 -29450 6530 -29390
rect 6530 -29450 6590 -29390
rect 6590 -29450 6600 -29390
rect 6520 -29460 6600 -29450
rect 8720 -29390 8800 -29210
rect 8720 -29450 8730 -29390
rect 8730 -29450 8790 -29390
rect 8790 -29450 8800 -29390
rect 8720 -29460 8800 -29450
rect 10920 -29390 11000 -29210
rect 10920 -29450 10930 -29390
rect 10930 -29450 10990 -29390
rect 10990 -29450 11000 -29390
rect 10920 -29460 11000 -29450
rect 13120 -29390 13200 -29210
rect 13120 -29450 13130 -29390
rect 13130 -29450 13190 -29390
rect 13190 -29450 13200 -29390
rect 13120 -29460 13200 -29450
rect 15320 -29390 15400 -29210
rect 15320 -29450 15330 -29390
rect 15330 -29450 15390 -29390
rect 15390 -29450 15400 -29390
rect 15320 -29460 15400 -29450
rect 17520 -29390 17600 -29210
rect 17520 -29450 17530 -29390
rect 17530 -29450 17590 -29390
rect 17590 -29450 17600 -29390
rect 17520 -29460 17600 -29450
rect 19720 -29390 19800 -29210
rect 19720 -29450 19730 -29390
rect 19730 -29450 19790 -29390
rect 19790 -29450 19800 -29390
rect 19720 -29460 19800 -29450
rect 21920 -29390 22000 -29210
rect 21920 -29450 21930 -29390
rect 21930 -29450 21990 -29390
rect 21990 -29450 22000 -29390
rect 21920 -29460 22000 -29450
rect 830 -29630 1010 -29550
rect 20510 -29630 20690 -29550
rect 1230 -29770 1410 -29690
rect 20910 -29770 21090 -29690
rect 1630 -29910 1810 -29830
rect 20110 -29910 20290 -29830
rect -80 -30190 0 -30010
rect -80 -30250 -70 -30190
rect -70 -30250 -10 -30190
rect -10 -30250 0 -30190
rect -80 -30260 0 -30250
rect 2120 -30190 2200 -30010
rect 2120 -30250 2130 -30190
rect 2130 -30250 2190 -30190
rect 2190 -30250 2200 -30190
rect 2120 -30260 2200 -30250
rect 4320 -30190 4400 -30010
rect 4320 -30250 4330 -30190
rect 4330 -30250 4390 -30190
rect 4390 -30250 4400 -30190
rect 4320 -30260 4400 -30250
rect 6520 -30190 6600 -30010
rect 6520 -30250 6530 -30190
rect 6530 -30250 6590 -30190
rect 6590 -30250 6600 -30190
rect 6520 -30260 6600 -30250
rect 8720 -30190 8800 -30010
rect 8720 -30250 8730 -30190
rect 8730 -30250 8790 -30190
rect 8790 -30250 8800 -30190
rect 8720 -30260 8800 -30250
rect 10920 -30190 11000 -30010
rect 10920 -30250 10930 -30190
rect 10930 -30250 10990 -30190
rect 10990 -30250 11000 -30190
rect 10920 -30260 11000 -30250
rect 13120 -30190 13200 -30010
rect 13120 -30250 13130 -30190
rect 13130 -30250 13190 -30190
rect 13190 -30250 13200 -30190
rect 13120 -30260 13200 -30250
rect 15320 -30190 15400 -30010
rect 15320 -30250 15330 -30190
rect 15330 -30250 15390 -30190
rect 15390 -30250 15400 -30190
rect 15320 -30260 15400 -30250
rect 17520 -30190 17600 -30010
rect 17520 -30250 17530 -30190
rect 17530 -30250 17590 -30190
rect 17590 -30250 17600 -30190
rect 17520 -30260 17600 -30250
rect 19720 -30190 19800 -30010
rect 19720 -30250 19730 -30190
rect 19730 -30250 19790 -30190
rect 19790 -30250 19800 -30190
rect 19720 -30260 19800 -30250
rect 21920 -30190 22000 -30010
rect 21920 -30250 21930 -30190
rect 21930 -30250 21990 -30190
rect 21990 -30250 22000 -30190
rect 21920 -30260 22000 -30250
rect 830 -30430 1010 -30350
rect 20510 -30430 20690 -30350
rect 1230 -30570 1410 -30490
rect 20910 -30570 21090 -30490
rect 1630 -30710 1810 -30630
rect 20110 -30710 20290 -30630
rect -80 -30990 0 -30810
rect -80 -31050 -70 -30990
rect -70 -31050 -10 -30990
rect -10 -31050 0 -30990
rect -80 -31060 0 -31050
rect 2120 -30990 2200 -30810
rect 2120 -31050 2130 -30990
rect 2130 -31050 2190 -30990
rect 2190 -31050 2200 -30990
rect 2120 -31060 2200 -31050
rect 4320 -30990 4400 -30810
rect 4320 -31050 4330 -30990
rect 4330 -31050 4390 -30990
rect 4390 -31050 4400 -30990
rect 4320 -31060 4400 -31050
rect 6520 -30990 6600 -30810
rect 6520 -31050 6530 -30990
rect 6530 -31050 6590 -30990
rect 6590 -31050 6600 -30990
rect 6520 -31060 6600 -31050
rect 8720 -30990 8800 -30810
rect 8720 -31050 8730 -30990
rect 8730 -31050 8790 -30990
rect 8790 -31050 8800 -30990
rect 8720 -31060 8800 -31050
rect 10920 -30990 11000 -30810
rect 10920 -31050 10930 -30990
rect 10930 -31050 10990 -30990
rect 10990 -31050 11000 -30990
rect 10920 -31060 11000 -31050
rect 13120 -30990 13200 -30810
rect 13120 -31050 13130 -30990
rect 13130 -31050 13190 -30990
rect 13190 -31050 13200 -30990
rect 13120 -31060 13200 -31050
rect 15320 -30990 15400 -30810
rect 15320 -31050 15330 -30990
rect 15330 -31050 15390 -30990
rect 15390 -31050 15400 -30990
rect 15320 -31060 15400 -31050
rect 17520 -30990 17600 -30810
rect 17520 -31050 17530 -30990
rect 17530 -31050 17590 -30990
rect 17590 -31050 17600 -30990
rect 17520 -31060 17600 -31050
rect 19720 -30990 19800 -30810
rect 19720 -31050 19730 -30990
rect 19730 -31050 19790 -30990
rect 19790 -31050 19800 -30990
rect 19720 -31060 19800 -31050
rect 21920 -30990 22000 -30810
rect 21920 -31050 21930 -30990
rect 21930 -31050 21990 -30990
rect 21990 -31050 22000 -30990
rect 21920 -31060 22000 -31050
rect 830 -31230 1010 -31150
rect 20510 -31230 20690 -31150
rect 1230 -31370 1410 -31290
rect 20910 -31370 21090 -31290
<< metal4 >>
rect -180 10940 100 11900
rect -180 10690 -80 10940
rect 0 10690 100 10940
rect -180 10140 100 10690
rect -180 9890 -80 10140
rect 0 9890 100 10140
rect -180 9340 100 9890
rect -180 9090 -80 9340
rect 0 9090 100 9340
rect -180 8540 100 9090
rect -180 8290 -80 8540
rect 0 8290 100 8540
rect -180 7740 100 8290
rect -180 7490 -80 7740
rect 0 7490 100 7740
rect -180 6940 100 7490
rect -180 6690 -80 6940
rect 0 6690 100 6940
rect -180 6140 100 6690
rect -180 5890 -80 6140
rect 0 5890 100 6140
rect -180 5340 100 5890
rect -180 5090 -80 5340
rect 0 5090 100 5340
rect -180 2480 100 5090
rect 420 8990 620 11300
rect 420 8910 430 8990
rect 610 8910 620 8990
rect 420 8190 620 8910
rect 420 8110 430 8190
rect 610 8110 620 8190
rect 420 7390 620 8110
rect 420 7310 430 7390
rect 610 7310 620 7390
rect 420 6590 620 7310
rect 420 6510 430 6590
rect 610 6510 620 6590
rect 420 3730 620 6510
rect 420 3550 430 3730
rect 610 3550 620 3730
rect 420 3540 620 3550
rect 820 11250 1020 11300
rect 820 11170 830 11250
rect 1010 11170 1020 11250
rect 820 10450 1020 11170
rect 820 10370 830 10450
rect 1010 10370 1020 10450
rect 820 9650 1020 10370
rect 820 9570 830 9650
rect 1010 9570 1020 9650
rect 820 8850 1020 9570
rect 820 8770 830 8850
rect 1010 8770 1020 8850
rect 820 8050 1020 8770
rect 820 7970 830 8050
rect 1010 7970 1020 8050
rect 820 7250 1020 7970
rect 820 7170 830 7250
rect 1010 7170 1020 7250
rect 820 6450 1020 7170
rect 820 6370 830 6450
rect 1010 6370 1020 6450
rect 820 5650 1020 6370
rect 820 5570 830 5650
rect 1010 5570 1020 5650
rect 820 -5570 1020 5570
rect 820 -5750 830 -5570
rect 1010 -5750 1020 -5570
rect 820 -5760 1020 -5750
rect 1220 11110 1420 11300
rect 1220 11030 1230 11110
rect 1410 11030 1420 11110
rect 1220 10310 1420 11030
rect 1220 10230 1230 10310
rect 1410 10230 1420 10310
rect 1220 9510 1420 10230
rect 1220 9430 1230 9510
rect 1410 9430 1420 9510
rect 1220 8710 1420 9430
rect 1220 8630 1230 8710
rect 1410 8630 1420 8710
rect 1220 7910 1420 8630
rect 1220 7830 1230 7910
rect 1410 7830 1420 7910
rect 1220 7110 1420 7830
rect 1220 7030 1230 7110
rect 1410 7030 1420 7110
rect 1220 6310 1420 7030
rect 1220 6230 1230 6310
rect 1410 6230 1420 6310
rect 1220 5510 1420 6230
rect 1220 5430 1230 5510
rect 1410 5430 1420 5510
rect 820 -7170 1020 -7160
rect 820 -7350 830 -7170
rect 1010 -7350 1020 -7170
rect -180 -25210 100 -23180
rect -180 -25460 -80 -25210
rect 0 -25460 100 -25210
rect -180 -26010 100 -25460
rect -180 -26260 -80 -26010
rect 0 -26260 100 -26010
rect -180 -26810 100 -26260
rect -180 -27060 -80 -26810
rect 0 -27060 100 -26810
rect -180 -27610 100 -27060
rect -180 -27860 -80 -27610
rect 0 -27860 100 -27610
rect -180 -28410 100 -27860
rect -180 -28660 -80 -28410
rect 0 -28660 100 -28410
rect -180 -29210 100 -28660
rect -180 -29460 -80 -29210
rect 0 -29460 100 -29210
rect -180 -30010 100 -29460
rect -180 -30260 -80 -30010
rect 0 -30260 100 -30010
rect -180 -30810 100 -30260
rect -180 -31060 -80 -30810
rect 0 -31060 100 -30810
rect -180 -32020 100 -31060
rect 420 -23670 620 -23660
rect 420 -23850 430 -23670
rect 610 -23850 620 -23670
rect 420 -26630 620 -23850
rect 420 -26710 430 -26630
rect 610 -26710 620 -26630
rect 420 -27430 620 -26710
rect 420 -27510 430 -27430
rect 610 -27510 620 -27430
rect 420 -28230 620 -27510
rect 420 -28310 430 -28230
rect 610 -28310 620 -28230
rect 420 -29030 620 -28310
rect 420 -29110 430 -29030
rect 610 -29110 620 -29030
rect 420 -31420 620 -29110
rect 820 -25550 1020 -7350
rect 1220 -7570 1420 5430
rect 1620 10590 1820 11300
rect 1620 10510 1630 10590
rect 1810 10510 1820 10590
rect 1620 9790 1820 10510
rect 1620 9710 1630 9790
rect 1810 9710 1820 9790
rect 1620 8990 1820 9710
rect 1620 8910 1630 8990
rect 1810 8910 1820 8990
rect 1620 8190 1820 8910
rect 1620 8110 1630 8190
rect 1810 8110 1820 8190
rect 1620 7390 1820 8110
rect 1620 7310 1630 7390
rect 1810 7310 1820 7390
rect 1620 6590 1820 7310
rect 1620 6510 1630 6590
rect 1810 6510 1820 6590
rect 1620 5790 1820 6510
rect 1620 5710 1630 5790
rect 1810 5710 1820 5790
rect 1620 4990 1820 5710
rect 1620 4910 1630 4990
rect 1810 4910 1820 4990
rect 1620 3330 1820 4910
rect 2020 10940 2300 11900
rect 2020 10690 2120 10940
rect 2200 10690 2300 10940
rect 2020 10140 2300 10690
rect 2020 9890 2120 10140
rect 2200 9890 2300 10140
rect 2020 9340 2300 9890
rect 2020 9090 2120 9340
rect 2200 9090 2300 9340
rect 2020 8540 2300 9090
rect 2020 8290 2120 8540
rect 2200 8290 2300 8540
rect 2020 7740 2300 8290
rect 2020 7490 2120 7740
rect 2200 7490 2300 7740
rect 2020 6940 2300 7490
rect 2020 6690 2120 6940
rect 2200 6690 2300 6940
rect 2020 6140 2300 6690
rect 2020 5890 2120 6140
rect 2200 5890 2300 6140
rect 2020 5340 2300 5890
rect 2020 5090 2120 5340
rect 2200 5090 2300 5340
rect 2020 3660 2300 5090
rect 4220 10940 4500 11900
rect 4220 10690 4320 10940
rect 4400 10690 4500 10940
rect 4220 10140 4500 10690
rect 4220 9890 4320 10140
rect 4400 9890 4500 10140
rect 4220 9340 4500 9890
rect 4220 9090 4320 9340
rect 4400 9090 4500 9340
rect 4220 8540 4500 9090
rect 4220 8290 4320 8540
rect 4400 8290 4500 8540
rect 4220 7740 4500 8290
rect 4220 7490 4320 7740
rect 4400 7490 4500 7740
rect 4220 6940 4500 7490
rect 4220 6690 4320 6940
rect 4400 6690 4500 6940
rect 4220 6140 4500 6690
rect 4220 5890 4320 6140
rect 4400 5890 4500 6140
rect 4220 5340 4500 5890
rect 4220 5090 4320 5340
rect 4400 5090 4500 5340
rect 4220 3660 4500 5090
rect 6420 10940 6700 11900
rect 6420 10690 6520 10940
rect 6600 10690 6700 10940
rect 6420 10140 6700 10690
rect 6420 9890 6520 10140
rect 6600 9890 6700 10140
rect 6420 9340 6700 9890
rect 6420 9090 6520 9340
rect 6600 9090 6700 9340
rect 6420 8540 6700 9090
rect 6420 8290 6520 8540
rect 6600 8290 6700 8540
rect 6420 7740 6700 8290
rect 6420 7490 6520 7740
rect 6600 7490 6700 7740
rect 6420 6940 6700 7490
rect 6420 6690 6520 6940
rect 6600 6690 6700 6940
rect 6420 6140 6700 6690
rect 6420 5890 6520 6140
rect 6600 5890 6700 6140
rect 6420 5340 6700 5890
rect 6420 5090 6520 5340
rect 6600 5090 6700 5340
rect 6420 3660 6700 5090
rect 8620 10940 8900 11900
rect 8620 10690 8720 10940
rect 8800 10690 8900 10940
rect 8620 10140 8900 10690
rect 8620 9890 8720 10140
rect 8800 9890 8900 10140
rect 8620 9340 8900 9890
rect 8620 9090 8720 9340
rect 8800 9090 8900 9340
rect 8620 8540 8900 9090
rect 8620 8290 8720 8540
rect 8800 8290 8900 8540
rect 8620 7740 8900 8290
rect 8620 7490 8720 7740
rect 8800 7490 8900 7740
rect 8620 6940 8900 7490
rect 8620 6690 8720 6940
rect 8800 6690 8900 6940
rect 8620 6140 8900 6690
rect 8620 5890 8720 6140
rect 8800 5890 8900 6140
rect 8620 5340 8900 5890
rect 8620 5090 8720 5340
rect 8800 5090 8900 5340
rect 8620 3660 8900 5090
rect 10820 10940 11100 11900
rect 10820 10690 10920 10940
rect 11000 10690 11100 10940
rect 10820 10140 11100 10690
rect 10820 9890 10920 10140
rect 11000 9890 11100 10140
rect 10820 9340 11100 9890
rect 10820 9090 10920 9340
rect 11000 9090 11100 9340
rect 10820 8540 11100 9090
rect 10820 8290 10920 8540
rect 11000 8290 11100 8540
rect 10820 7740 11100 8290
rect 10820 7490 10920 7740
rect 11000 7490 11100 7740
rect 10820 6940 11100 7490
rect 10820 6690 10920 6940
rect 11000 6690 11100 6940
rect 10820 6140 11100 6690
rect 10820 5890 10920 6140
rect 11000 5890 11100 6140
rect 10820 5340 11100 5890
rect 10820 5090 10920 5340
rect 11000 5090 11100 5340
rect 10820 3660 11100 5090
rect 13020 10940 13300 11900
rect 13020 10690 13120 10940
rect 13200 10690 13300 10940
rect 13020 10140 13300 10690
rect 13020 9890 13120 10140
rect 13200 9890 13300 10140
rect 13020 9340 13300 9890
rect 13020 9090 13120 9340
rect 13200 9090 13300 9340
rect 13020 8540 13300 9090
rect 13020 8290 13120 8540
rect 13200 8290 13300 8540
rect 13020 7740 13300 8290
rect 13020 7490 13120 7740
rect 13200 7490 13300 7740
rect 13020 6940 13300 7490
rect 13020 6690 13120 6940
rect 13200 6690 13300 6940
rect 13020 6140 13300 6690
rect 13020 5890 13120 6140
rect 13200 5890 13300 6140
rect 13020 5340 13300 5890
rect 13020 5090 13120 5340
rect 13200 5090 13300 5340
rect 13020 3660 13300 5090
rect 15220 10940 15500 11900
rect 15220 10690 15320 10940
rect 15400 10690 15500 10940
rect 15220 10140 15500 10690
rect 15220 9890 15320 10140
rect 15400 9890 15500 10140
rect 15220 9340 15500 9890
rect 15220 9090 15320 9340
rect 15400 9090 15500 9340
rect 15220 8540 15500 9090
rect 15220 8290 15320 8540
rect 15400 8290 15500 8540
rect 15220 7740 15500 8290
rect 15220 7490 15320 7740
rect 15400 7490 15500 7740
rect 15220 6940 15500 7490
rect 15220 6690 15320 6940
rect 15400 6690 15500 6940
rect 15220 6140 15500 6690
rect 15220 5890 15320 6140
rect 15400 5890 15500 6140
rect 15220 5340 15500 5890
rect 15220 5090 15320 5340
rect 15400 5090 15500 5340
rect 15220 3660 15500 5090
rect 17420 10940 17700 11900
rect 17420 10690 17520 10940
rect 17600 10690 17700 10940
rect 17420 10140 17700 10690
rect 17420 9890 17520 10140
rect 17600 9890 17700 10140
rect 17420 9340 17700 9890
rect 17420 9090 17520 9340
rect 17600 9090 17700 9340
rect 17420 8540 17700 9090
rect 17420 8290 17520 8540
rect 17600 8290 17700 8540
rect 17420 7740 17700 8290
rect 17420 7490 17520 7740
rect 17600 7490 17700 7740
rect 17420 6940 17700 7490
rect 17420 6690 17520 6940
rect 17600 6690 17700 6940
rect 17420 6140 17700 6690
rect 17420 5890 17520 6140
rect 17600 5890 17700 6140
rect 17420 5340 17700 5890
rect 17420 5090 17520 5340
rect 17600 5090 17700 5340
rect 17420 3660 17700 5090
rect 19620 10940 19900 11900
rect 19620 10690 19720 10940
rect 19800 10690 19900 10940
rect 19620 10140 19900 10690
rect 19620 9890 19720 10140
rect 19800 9890 19900 10140
rect 19620 9340 19900 9890
rect 19620 9090 19720 9340
rect 19800 9090 19900 9340
rect 19620 8540 19900 9090
rect 19620 8290 19720 8540
rect 19800 8290 19900 8540
rect 19620 7740 19900 8290
rect 19620 7490 19720 7740
rect 19800 7490 19900 7740
rect 19620 6940 19900 7490
rect 19620 6690 19720 6940
rect 19800 6690 19900 6940
rect 19620 6140 19900 6690
rect 19620 5890 19720 6140
rect 19800 5890 19900 6140
rect 19620 5340 19900 5890
rect 19620 5090 19720 5340
rect 19800 5090 19900 5340
rect 19620 3660 19900 5090
rect 20100 10590 20300 11300
rect 20100 10510 20110 10590
rect 20290 10510 20300 10590
rect 20100 9790 20300 10510
rect 20100 9710 20110 9790
rect 20290 9710 20300 9790
rect 20100 8990 20300 9710
rect 20100 8910 20110 8990
rect 20290 8910 20300 8990
rect 20100 8190 20300 8910
rect 20100 8110 20110 8190
rect 20290 8110 20300 8190
rect 20100 7390 20300 8110
rect 20100 7310 20110 7390
rect 20290 7310 20300 7390
rect 20100 6590 20300 7310
rect 20100 6510 20110 6590
rect 20290 6510 20300 6590
rect 20100 5790 20300 6510
rect 20100 5710 20110 5790
rect 20290 5710 20300 5790
rect 20100 4990 20300 5710
rect 20100 4910 20110 4990
rect 20290 4910 20300 4990
rect 1620 3150 1630 3330
rect 1810 3150 1820 3330
rect 1620 3140 1820 3150
rect 20100 3330 20300 4910
rect 20100 3150 20110 3330
rect 20290 3150 20300 3330
rect 20100 3140 20300 3150
rect 20500 11250 20700 11300
rect 20500 11170 20510 11250
rect 20690 11170 20700 11250
rect 20500 10450 20700 11170
rect 20500 10370 20510 10450
rect 20690 10370 20700 10450
rect 20500 9650 20700 10370
rect 20500 9570 20510 9650
rect 20690 9570 20700 9650
rect 20500 8850 20700 9570
rect 20500 8770 20510 8850
rect 20690 8770 20700 8850
rect 20500 8050 20700 8770
rect 20500 7970 20510 8050
rect 20690 7970 20700 8050
rect 20500 7250 20700 7970
rect 20500 7170 20510 7250
rect 20690 7170 20700 7250
rect 20500 6450 20700 7170
rect 20500 6370 20510 6450
rect 20690 6370 20700 6450
rect 20500 5650 20700 6370
rect 20500 5570 20510 5650
rect 20690 5570 20700 5650
rect 14900 1960 15040 1990
rect 14900 1300 14910 1960
rect 15030 1300 15040 1960
rect 1220 -7750 1230 -7570
rect 1410 -7750 1420 -7570
rect 1220 -7760 1420 -7750
rect 1620 -5170 1820 -5160
rect 1620 -5350 1630 -5170
rect 1810 -5350 1820 -5170
rect 1620 -8040 1820 -5350
rect 14900 -6490 15040 1300
rect 20500 -5570 20700 5570
rect 20900 11110 21100 11300
rect 20900 11030 20910 11110
rect 21090 11030 21100 11110
rect 20900 10310 21100 11030
rect 20900 10230 20910 10310
rect 21090 10230 21100 10310
rect 20900 9510 21100 10230
rect 20900 9430 20910 9510
rect 21090 9430 21100 9510
rect 20900 8710 21100 9430
rect 20900 8630 20910 8710
rect 21090 8630 21100 8710
rect 20900 7910 21100 8630
rect 20900 7830 20910 7910
rect 21090 7830 21100 7910
rect 20900 7110 21100 7830
rect 20900 7030 20910 7110
rect 21090 7030 21100 7110
rect 20900 6310 21100 7030
rect 20900 6230 20910 6310
rect 21090 6230 21100 6310
rect 20900 5510 21100 6230
rect 20900 5430 20910 5510
rect 21090 5430 21100 5510
rect 20900 3340 21100 5430
rect 21300 8990 21500 11300
rect 21300 8910 21310 8990
rect 21490 8910 21500 8990
rect 21300 8190 21500 8910
rect 21300 8110 21310 8190
rect 21490 8110 21500 8190
rect 21300 7390 21500 8110
rect 21300 7310 21310 7390
rect 21490 7310 21500 7390
rect 21300 6590 21500 7310
rect 21300 6510 21310 6590
rect 21490 6510 21500 6590
rect 21300 3730 21500 6510
rect 21300 3550 21310 3730
rect 21490 3550 21500 3730
rect 21820 10940 22100 11900
rect 21820 10690 21920 10940
rect 22000 10690 22100 10940
rect 21820 10140 22100 10690
rect 21820 9890 21920 10140
rect 22000 9890 22100 10140
rect 21820 9340 22100 9890
rect 21820 9090 21920 9340
rect 22000 9090 22100 9340
rect 21820 8540 22100 9090
rect 21820 8290 21920 8540
rect 22000 8290 22100 8540
rect 21820 7740 22100 8290
rect 21820 7490 21920 7740
rect 22000 7490 22100 7740
rect 21820 6940 22100 7490
rect 21820 6690 21920 6940
rect 22000 6690 22100 6940
rect 21820 6140 22100 6690
rect 21820 5890 21920 6140
rect 22000 5890 22100 6140
rect 21820 5340 22100 5890
rect 21820 5090 21920 5340
rect 22000 5090 22100 5340
rect 21820 3660 22100 5090
rect 21300 3540 21500 3550
rect 20900 3140 22260 3340
rect 20500 -5750 20510 -5570
rect 20690 -5750 20700 -5570
rect 20500 -5760 20700 -5750
rect 20900 -5170 21100 -5160
rect 20900 -5350 20910 -5170
rect 21090 -5350 21100 -5170
rect 14900 -6610 14910 -6490
rect 15030 -6610 15040 -6490
rect 14900 -6620 15040 -6610
rect 820 -25630 830 -25550
rect 1010 -25630 1020 -25550
rect 820 -26350 1020 -25630
rect 820 -26430 830 -26350
rect 1010 -26430 1020 -26350
rect 820 -27150 1020 -26430
rect 820 -27230 830 -27150
rect 1010 -27230 1020 -27150
rect 820 -27950 1020 -27230
rect 820 -28030 830 -27950
rect 1010 -28030 1020 -27950
rect 820 -28750 1020 -28030
rect 820 -28830 830 -28750
rect 1010 -28830 1020 -28750
rect 820 -29550 1020 -28830
rect 820 -29630 830 -29550
rect 1010 -29630 1020 -29550
rect 820 -30350 1020 -29630
rect 820 -30430 830 -30350
rect 1010 -30430 1020 -30350
rect 820 -31150 1020 -30430
rect 820 -31230 830 -31150
rect 1010 -31230 1020 -31150
rect 820 -31420 1020 -31230
rect 1220 -8240 1820 -8040
rect 20500 -7170 20700 -7160
rect 20500 -7350 20510 -7170
rect 20690 -7350 20700 -7170
rect 1220 -25690 1420 -8240
rect 1220 -25770 1230 -25690
rect 1410 -25770 1420 -25690
rect 1220 -26490 1420 -25770
rect 1220 -26570 1230 -26490
rect 1410 -26570 1420 -26490
rect 1220 -27290 1420 -26570
rect 1220 -27370 1230 -27290
rect 1410 -27370 1420 -27290
rect 1220 -28090 1420 -27370
rect 1220 -28170 1230 -28090
rect 1410 -28170 1420 -28090
rect 1220 -28890 1420 -28170
rect 1220 -28970 1230 -28890
rect 1410 -28970 1420 -28890
rect 1220 -29690 1420 -28970
rect 1220 -29770 1230 -29690
rect 1410 -29770 1420 -29690
rect 1220 -30490 1420 -29770
rect 1220 -30570 1230 -30490
rect 1410 -30570 1420 -30490
rect 1220 -31290 1420 -30570
rect 1220 -31370 1230 -31290
rect 1410 -31370 1420 -31290
rect 1220 -31420 1420 -31370
rect 1620 -23270 1820 -23260
rect 1620 -23450 1630 -23270
rect 1810 -23450 1820 -23270
rect 1620 -25030 1820 -23450
rect 20100 -23270 20300 -23260
rect 20100 -23450 20110 -23270
rect 20290 -23450 20300 -23270
rect 1620 -25110 1630 -25030
rect 1810 -25110 1820 -25030
rect 1620 -25830 1820 -25110
rect 1620 -25910 1630 -25830
rect 1810 -25910 1820 -25830
rect 1620 -26630 1820 -25910
rect 1620 -26710 1630 -26630
rect 1810 -26710 1820 -26630
rect 1620 -27430 1820 -26710
rect 1620 -27510 1630 -27430
rect 1810 -27510 1820 -27430
rect 1620 -28230 1820 -27510
rect 1620 -28310 1630 -28230
rect 1810 -28310 1820 -28230
rect 1620 -29030 1820 -28310
rect 1620 -29110 1630 -29030
rect 1810 -29110 1820 -29030
rect 1620 -29830 1820 -29110
rect 1620 -29910 1630 -29830
rect 1810 -29910 1820 -29830
rect 1620 -30630 1820 -29910
rect 1620 -30710 1630 -30630
rect 1810 -30710 1820 -30630
rect 1620 -31420 1820 -30710
rect 2020 -25210 2300 -23780
rect 2020 -25460 2120 -25210
rect 2200 -25460 2300 -25210
rect 2020 -26010 2300 -25460
rect 2020 -26260 2120 -26010
rect 2200 -26260 2300 -26010
rect 2020 -26810 2300 -26260
rect 2020 -27060 2120 -26810
rect 2200 -27060 2300 -26810
rect 2020 -27610 2300 -27060
rect 2020 -27860 2120 -27610
rect 2200 -27860 2300 -27610
rect 2020 -28410 2300 -27860
rect 2020 -28660 2120 -28410
rect 2200 -28660 2300 -28410
rect 2020 -29210 2300 -28660
rect 2020 -29460 2120 -29210
rect 2200 -29460 2300 -29210
rect 2020 -30010 2300 -29460
rect 2020 -30260 2120 -30010
rect 2200 -30260 2300 -30010
rect 2020 -30810 2300 -30260
rect 2020 -31060 2120 -30810
rect 2200 -31060 2300 -30810
rect 2020 -32020 2300 -31060
rect 4220 -25210 4500 -23780
rect 4220 -25460 4320 -25210
rect 4400 -25460 4500 -25210
rect 4220 -26010 4500 -25460
rect 4220 -26260 4320 -26010
rect 4400 -26260 4500 -26010
rect 4220 -26810 4500 -26260
rect 4220 -27060 4320 -26810
rect 4400 -27060 4500 -26810
rect 4220 -27610 4500 -27060
rect 4220 -27860 4320 -27610
rect 4400 -27860 4500 -27610
rect 4220 -28410 4500 -27860
rect 4220 -28660 4320 -28410
rect 4400 -28660 4500 -28410
rect 4220 -29210 4500 -28660
rect 4220 -29460 4320 -29210
rect 4400 -29460 4500 -29210
rect 4220 -30010 4500 -29460
rect 4220 -30260 4320 -30010
rect 4400 -30260 4500 -30010
rect 4220 -30810 4500 -30260
rect 4220 -31060 4320 -30810
rect 4400 -31060 4500 -30810
rect 4220 -32020 4500 -31060
rect 6420 -25210 6700 -23780
rect 6420 -25460 6520 -25210
rect 6600 -25460 6700 -25210
rect 6420 -26010 6700 -25460
rect 6420 -26260 6520 -26010
rect 6600 -26260 6700 -26010
rect 6420 -26810 6700 -26260
rect 6420 -27060 6520 -26810
rect 6600 -27060 6700 -26810
rect 6420 -27610 6700 -27060
rect 6420 -27860 6520 -27610
rect 6600 -27860 6700 -27610
rect 6420 -28410 6700 -27860
rect 6420 -28660 6520 -28410
rect 6600 -28660 6700 -28410
rect 6420 -29210 6700 -28660
rect 6420 -29460 6520 -29210
rect 6600 -29460 6700 -29210
rect 6420 -30010 6700 -29460
rect 6420 -30260 6520 -30010
rect 6600 -30260 6700 -30010
rect 6420 -30810 6700 -30260
rect 6420 -31060 6520 -30810
rect 6600 -31060 6700 -30810
rect 6420 -32020 6700 -31060
rect 8620 -25210 8900 -23780
rect 8620 -25460 8720 -25210
rect 8800 -25460 8900 -25210
rect 8620 -26010 8900 -25460
rect 8620 -26260 8720 -26010
rect 8800 -26260 8900 -26010
rect 8620 -26810 8900 -26260
rect 8620 -27060 8720 -26810
rect 8800 -27060 8900 -26810
rect 8620 -27610 8900 -27060
rect 8620 -27860 8720 -27610
rect 8800 -27860 8900 -27610
rect 8620 -28410 8900 -27860
rect 8620 -28660 8720 -28410
rect 8800 -28660 8900 -28410
rect 8620 -29210 8900 -28660
rect 8620 -29460 8720 -29210
rect 8800 -29460 8900 -29210
rect 8620 -30010 8900 -29460
rect 8620 -30260 8720 -30010
rect 8800 -30260 8900 -30010
rect 8620 -30810 8900 -30260
rect 8620 -31060 8720 -30810
rect 8800 -31060 8900 -30810
rect 8620 -32020 8900 -31060
rect 10820 -25210 11100 -23780
rect 10820 -25460 10920 -25210
rect 11000 -25460 11100 -25210
rect 10820 -26010 11100 -25460
rect 10820 -26260 10920 -26010
rect 11000 -26260 11100 -26010
rect 10820 -26810 11100 -26260
rect 10820 -27060 10920 -26810
rect 11000 -27060 11100 -26810
rect 10820 -27610 11100 -27060
rect 10820 -27860 10920 -27610
rect 11000 -27860 11100 -27610
rect 10820 -28410 11100 -27860
rect 10820 -28660 10920 -28410
rect 11000 -28660 11100 -28410
rect 10820 -29210 11100 -28660
rect 10820 -29460 10920 -29210
rect 11000 -29460 11100 -29210
rect 10820 -30010 11100 -29460
rect 10820 -30260 10920 -30010
rect 11000 -30260 11100 -30010
rect 10820 -30810 11100 -30260
rect 10820 -31060 10920 -30810
rect 11000 -31060 11100 -30810
rect 10820 -32020 11100 -31060
rect 13020 -25210 13300 -23780
rect 13020 -25460 13120 -25210
rect 13200 -25460 13300 -25210
rect 13020 -26010 13300 -25460
rect 13020 -26260 13120 -26010
rect 13200 -26260 13300 -26010
rect 13020 -26810 13300 -26260
rect 13020 -27060 13120 -26810
rect 13200 -27060 13300 -26810
rect 13020 -27610 13300 -27060
rect 13020 -27860 13120 -27610
rect 13200 -27860 13300 -27610
rect 13020 -28410 13300 -27860
rect 13020 -28660 13120 -28410
rect 13200 -28660 13300 -28410
rect 13020 -29210 13300 -28660
rect 13020 -29460 13120 -29210
rect 13200 -29460 13300 -29210
rect 13020 -30010 13300 -29460
rect 13020 -30260 13120 -30010
rect 13200 -30260 13300 -30010
rect 13020 -30810 13300 -30260
rect 13020 -31060 13120 -30810
rect 13200 -31060 13300 -30810
rect 13020 -32020 13300 -31060
rect 15220 -25210 15500 -23780
rect 15220 -25460 15320 -25210
rect 15400 -25460 15500 -25210
rect 15220 -26010 15500 -25460
rect 15220 -26260 15320 -26010
rect 15400 -26260 15500 -26010
rect 15220 -26810 15500 -26260
rect 15220 -27060 15320 -26810
rect 15400 -27060 15500 -26810
rect 15220 -27610 15500 -27060
rect 15220 -27860 15320 -27610
rect 15400 -27860 15500 -27610
rect 15220 -28410 15500 -27860
rect 15220 -28660 15320 -28410
rect 15400 -28660 15500 -28410
rect 15220 -29210 15500 -28660
rect 15220 -29460 15320 -29210
rect 15400 -29460 15500 -29210
rect 15220 -30010 15500 -29460
rect 15220 -30260 15320 -30010
rect 15400 -30260 15500 -30010
rect 15220 -30810 15500 -30260
rect 15220 -31060 15320 -30810
rect 15400 -31060 15500 -30810
rect 15220 -32020 15500 -31060
rect 17420 -25210 17700 -23780
rect 17420 -25460 17520 -25210
rect 17600 -25460 17700 -25210
rect 17420 -26010 17700 -25460
rect 17420 -26260 17520 -26010
rect 17600 -26260 17700 -26010
rect 17420 -26810 17700 -26260
rect 17420 -27060 17520 -26810
rect 17600 -27060 17700 -26810
rect 17420 -27610 17700 -27060
rect 17420 -27860 17520 -27610
rect 17600 -27860 17700 -27610
rect 17420 -28410 17700 -27860
rect 17420 -28660 17520 -28410
rect 17600 -28660 17700 -28410
rect 17420 -29210 17700 -28660
rect 17420 -29460 17520 -29210
rect 17600 -29460 17700 -29210
rect 17420 -30010 17700 -29460
rect 17420 -30260 17520 -30010
rect 17600 -30260 17700 -30010
rect 17420 -30810 17700 -30260
rect 17420 -31060 17520 -30810
rect 17600 -31060 17700 -30810
rect 17420 -32020 17700 -31060
rect 19620 -25210 19900 -23780
rect 19620 -25460 19720 -25210
rect 19800 -25460 19900 -25210
rect 19620 -26010 19900 -25460
rect 19620 -26260 19720 -26010
rect 19800 -26260 19900 -26010
rect 19620 -26810 19900 -26260
rect 19620 -27060 19720 -26810
rect 19800 -27060 19900 -26810
rect 19620 -27610 19900 -27060
rect 19620 -27860 19720 -27610
rect 19800 -27860 19900 -27610
rect 19620 -28410 19900 -27860
rect 19620 -28660 19720 -28410
rect 19800 -28660 19900 -28410
rect 19620 -29210 19900 -28660
rect 19620 -29460 19720 -29210
rect 19800 -29460 19900 -29210
rect 19620 -30010 19900 -29460
rect 19620 -30260 19720 -30010
rect 19800 -30260 19900 -30010
rect 19620 -30810 19900 -30260
rect 19620 -31060 19720 -30810
rect 19800 -31060 19900 -30810
rect 19620 -32020 19900 -31060
rect 20100 -25030 20300 -23450
rect 20100 -25110 20110 -25030
rect 20290 -25110 20300 -25030
rect 20100 -25830 20300 -25110
rect 20100 -25910 20110 -25830
rect 20290 -25910 20300 -25830
rect 20100 -26630 20300 -25910
rect 20100 -26710 20110 -26630
rect 20290 -26710 20300 -26630
rect 20100 -27430 20300 -26710
rect 20100 -27510 20110 -27430
rect 20290 -27510 20300 -27430
rect 20100 -28230 20300 -27510
rect 20100 -28310 20110 -28230
rect 20290 -28310 20300 -28230
rect 20100 -29030 20300 -28310
rect 20100 -29110 20110 -29030
rect 20290 -29110 20300 -29030
rect 20100 -29830 20300 -29110
rect 20100 -29910 20110 -29830
rect 20290 -29910 20300 -29830
rect 20100 -30630 20300 -29910
rect 20100 -30710 20110 -30630
rect 20290 -30710 20300 -30630
rect 20100 -31420 20300 -30710
rect 20500 -25550 20700 -7350
rect 20500 -25630 20510 -25550
rect 20690 -25630 20700 -25550
rect 20500 -26350 20700 -25630
rect 20500 -26430 20510 -26350
rect 20690 -26430 20700 -26350
rect 20500 -27150 20700 -26430
rect 20500 -27230 20510 -27150
rect 20690 -27230 20700 -27150
rect 20500 -27950 20700 -27230
rect 20500 -28030 20510 -27950
rect 20690 -28030 20700 -27950
rect 20500 -28750 20700 -28030
rect 20500 -28830 20510 -28750
rect 20690 -28830 20700 -28750
rect 20500 -29550 20700 -28830
rect 20500 -29630 20510 -29550
rect 20690 -29630 20700 -29550
rect 20500 -30350 20700 -29630
rect 20500 -30430 20510 -30350
rect 20690 -30430 20700 -30350
rect 20500 -31150 20700 -30430
rect 20500 -31230 20510 -31150
rect 20690 -31230 20700 -31150
rect 20500 -31420 20700 -31230
rect 20900 -25690 21100 -5350
rect 22060 -7570 22260 3140
rect 22060 -7750 22070 -7570
rect 22250 -7750 22260 -7570
rect 22060 -7760 22260 -7750
rect 20900 -25770 20910 -25690
rect 21090 -25770 21100 -25690
rect 20900 -26490 21100 -25770
rect 20900 -26570 20910 -26490
rect 21090 -26570 21100 -26490
rect 20900 -27290 21100 -26570
rect 20900 -27370 20910 -27290
rect 21090 -27370 21100 -27290
rect 20900 -28090 21100 -27370
rect 20900 -28170 20910 -28090
rect 21090 -28170 21100 -28090
rect 20900 -28890 21100 -28170
rect 20900 -28970 20910 -28890
rect 21090 -28970 21100 -28890
rect 20900 -29690 21100 -28970
rect 20900 -29770 20910 -29690
rect 21090 -29770 21100 -29690
rect 20900 -30490 21100 -29770
rect 20900 -30570 20910 -30490
rect 21090 -30570 21100 -30490
rect 20900 -31290 21100 -30570
rect 20900 -31370 20910 -31290
rect 21090 -31370 21100 -31290
rect 20900 -31420 21100 -31370
rect 21300 -23670 21500 -23660
rect 21300 -23850 21310 -23670
rect 21490 -23850 21500 -23670
rect 21300 -26630 21500 -23850
rect 21300 -26710 21310 -26630
rect 21490 -26710 21500 -26630
rect 21300 -27430 21500 -26710
rect 21300 -27510 21310 -27430
rect 21490 -27510 21500 -27430
rect 21300 -28230 21500 -27510
rect 21300 -28310 21310 -28230
rect 21490 -28310 21500 -28230
rect 21300 -29030 21500 -28310
rect 21300 -29110 21310 -29030
rect 21490 -29110 21500 -29030
rect 21300 -31420 21500 -29110
rect 21820 -25210 22100 -23780
rect 21820 -25460 21920 -25210
rect 22000 -25460 22100 -25210
rect 21820 -26010 22100 -25460
rect 21820 -26260 21920 -26010
rect 22000 -26260 22100 -26010
rect 21820 -26810 22100 -26260
rect 21820 -27060 21920 -26810
rect 22000 -27060 22100 -26810
rect 21820 -27610 22100 -27060
rect 21820 -27860 21920 -27610
rect 22000 -27860 22100 -27610
rect 21820 -28410 22100 -27860
rect 21820 -28660 21920 -28410
rect 22000 -28660 22100 -28410
rect 21820 -29210 22100 -28660
rect 21820 -29460 21920 -29210
rect 22000 -29460 22100 -29210
rect 21820 -30010 22100 -29460
rect 21820 -30260 21920 -30010
rect 22000 -30260 22100 -30010
rect 21820 -30810 22100 -30260
rect 21820 -31060 21920 -30810
rect 22000 -31060 22100 -30810
rect 21820 -32020 22100 -31060
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_9
timestamp 1713067540
transform 0 1 5458 -1 0 5178
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_10
timestamp 1713067540
transform 0 1 5458 -1 0 5978
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_11
timestamp 1713067540
transform 0 1 5458 -1 0 6778
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_12
timestamp 1713067540
transform 0 1 5458 -1 0 7578
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_13
timestamp 1713067540
transform 0 1 5458 -1 0 8378
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_14
timestamp 1713067540
transform 0 1 5458 -1 0 9178
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_15
timestamp 1713067540
transform 0 1 5458 -1 0 9978
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_17
timestamp 1713067540
transform 0 1 3258 -1 0 5178
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_18
timestamp 1713067540
transform 0 1 3258 -1 0 5978
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_19
timestamp 1713067540
transform 0 1 3258 -1 0 6778
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_20
timestamp 1713067540
transform 0 1 3258 -1 0 7578
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_21
timestamp 1713067540
transform 0 1 3258 -1 0 8378
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_22
timestamp 1713067540
transform 0 1 3258 -1 0 9178
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_23
timestamp 1713067540
transform 0 1 3258 -1 0 9978
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_25
timestamp 1713067540
transform 0 1 7658 -1 0 5178
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_26
timestamp 1713067540
transform 0 1 7658 -1 0 5978
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_27
timestamp 1713067540
transform 0 1 7658 -1 0 6778
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_28
timestamp 1713067540
transform 0 1 7658 -1 0 7578
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_29
timestamp 1713067540
transform 0 1 7658 -1 0 8378
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_30
timestamp 1713067540
transform 0 1 7658 -1 0 9178
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_31
timestamp 1713067540
transform 0 1 7658 -1 0 9978
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_32
timestamp 1713067540
transform 0 1 12058 -1 0 9978
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_33
timestamp 1713067540
transform 0 1 12058 -1 0 9178
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_34
timestamp 1713067540
transform 0 1 12058 -1 0 8378
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_35
timestamp 1713067540
transform 0 1 12058 -1 0 7578
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_36
timestamp 1713067540
transform 0 1 12058 -1 0 6778
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_37
timestamp 1713067540
transform 0 1 12058 -1 0 5978
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_38
timestamp 1713067540
transform 0 1 12058 -1 0 5178
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_40
timestamp 1713067540
transform 0 1 9858 -1 0 9978
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_41
timestamp 1713067540
transform 0 1 9858 -1 0 9178
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_42
timestamp 1713067540
transform 0 1 9858 -1 0 8378
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_43
timestamp 1713067540
transform 0 1 9858 -1 0 7578
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_44
timestamp 1713067540
transform 0 1 9858 -1 0 6778
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_45
timestamp 1713067540
transform 0 1 9858 -1 0 5978
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_46
timestamp 1713067540
transform 0 1 9858 -1 0 5178
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_49
timestamp 1713067540
transform 0 1 14258 -1 0 7578
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_50
timestamp 1713067540
transform 0 1 14258 -1 0 6778
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_51
timestamp 1713067540
transform 0 1 14258 -1 0 5978
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_52
timestamp 1713067540
transform 0 1 14258 -1 0 5178
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_53
timestamp 1713067540
transform 0 1 14258 -1 0 9978
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_54
timestamp 1713067540
transform 0 1 14258 -1 0 9178
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_55
timestamp 1713067540
transform 0 1 14258 -1 0 8378
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_57
timestamp 1713067540
transform 0 1 16458 -1 0 7578
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_58
timestamp 1713067540
transform 0 1 16458 -1 0 6778
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_59
timestamp 1713067540
transform 0 1 16458 -1 0 5978
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_60
timestamp 1713067540
transform 0 1 16458 -1 0 5178
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_61
timestamp 1713067540
transform 0 1 16458 -1 0 9978
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_62
timestamp 1713067540
transform 0 1 16458 -1 0 9178
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_63
timestamp 1713067540
transform 0 1 16458 -1 0 8378
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_73
timestamp 1713067540
transform 0 1 3258 -1 0 10778
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_74
timestamp 1713067540
transform 0 1 5458 -1 0 10778
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_75
timestamp 1713067540
transform 0 1 7658 -1 0 10778
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_76
timestamp 1713067540
transform 0 1 9858 -1 0 10778
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_77
timestamp 1713067540
transform 0 1 12058 -1 0 10778
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_78
timestamp 1713067540
transform 0 1 14258 -1 0 10778
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_79
timestamp 1713067540
transform 0 1 16458 -1 0 10778
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_81
timestamp 1713067540
transform 0 1 18658 -1 0 10778
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_82
timestamp 1713067540
transform 0 1 18658 -1 0 9978
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_83
timestamp 1713067540
transform 0 1 18658 -1 0 9178
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_84
timestamp 1713067540
transform 0 1 18658 -1 0 8378
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_85
timestamp 1713067540
transform 0 1 18658 -1 0 7578
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_86
timestamp 1713067540
transform 0 1 18658 -1 0 6778
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_87
timestamp 1713067540
transform 0 1 18658 -1 0 5978
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_88
timestamp 1713067540
transform 0 1 18658 -1 0 5178
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_T8W2FW  sky130_fd_pr__nfet_g5v0d10v5_T8W2FW_0
timestamp 1713067540
transform 0 1 1059 -1 0 9179
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_T8W2FW  sky130_fd_pr__nfet_g5v0d10v5_T8W2FW_1
timestamp 1713067540
transform 0 1 1059 -1 0 9979
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_T8W2FW  sky130_fd_pr__nfet_g5v0d10v5_T8W2FW_2
timestamp 1713067540
transform 0 1 1059 -1 0 10779
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_T8W2FW  sky130_fd_pr__nfet_g5v0d10v5_T8W2FW_3
timestamp 1713067540
transform 0 1 1059 -1 0 11579
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_T8W2FW  sky130_fd_pr__nfet_g5v0d10v5_T8W2FW_4
timestamp 1713067540
transform 0 1 1059 -1 0 8379
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_T8W2FW  sky130_fd_pr__nfet_g5v0d10v5_T8W2FW_5
timestamp 1713067540
transform 0 1 1059 -1 0 7579
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_T8W2FW  sky130_fd_pr__nfet_g5v0d10v5_T8W2FW_6
timestamp 1713067540
transform 0 1 1059 -1 0 4379
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_T8W2FW  sky130_fd_pr__nfet_g5v0d10v5_T8W2FW_7
timestamp 1713067540
transform 0 1 1059 -1 0 6779
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_T8W2FW  sky130_fd_pr__nfet_g5v0d10v5_T8W2FW_8
timestamp 1713067540
transform 0 1 1059 -1 0 5979
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_T8W2FW  sky130_fd_pr__nfet_g5v0d10v5_T8W2FW_9
timestamp 1713067540
transform 0 1 1059 -1 0 5179
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_T8W2FW  sky130_fd_pr__nfet_g5v0d10v5_T8W2FW_10
timestamp 1713067540
transform 0 1 3259 -1 0 4379
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_T8W2FW  sky130_fd_pr__nfet_g5v0d10v5_T8W2FW_11
timestamp 1713067540
transform 0 1 5459 -1 0 4379
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_T8W2FW  sky130_fd_pr__nfet_g5v0d10v5_T8W2FW_12
timestamp 1713067540
transform 0 1 7659 -1 0 4379
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_T8W2FW  sky130_fd_pr__nfet_g5v0d10v5_T8W2FW_13
timestamp 1713067540
transform 0 1 9859 -1 0 4379
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_T8W2FW  sky130_fd_pr__nfet_g5v0d10v5_T8W2FW_14
timestamp 1713067540
transform 0 1 12059 -1 0 4379
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_T8W2FW  sky130_fd_pr__nfet_g5v0d10v5_T8W2FW_15
timestamp 1713067540
transform 0 1 14259 -1 0 4379
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_T8W2FW  sky130_fd_pr__nfet_g5v0d10v5_T8W2FW_16
timestamp 1713067540
transform 0 1 16459 -1 0 4379
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_T8W2FW  sky130_fd_pr__nfet_g5v0d10v5_T8W2FW_17
timestamp 1713067540
transform 0 1 18659 -1 0 4379
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_T8W2FW  sky130_fd_pr__nfet_g5v0d10v5_T8W2FW_18
timestamp 1713067540
transform 0 1 3259 -1 0 11579
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_T8W2FW  sky130_fd_pr__nfet_g5v0d10v5_T8W2FW_19
timestamp 1713067540
transform 0 1 20859 -1 0 4379
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_T8W2FW  sky130_fd_pr__nfet_g5v0d10v5_T8W2FW_20
timestamp 1713067540
transform 0 1 20859 -1 0 5179
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_T8W2FW  sky130_fd_pr__nfet_g5v0d10v5_T8W2FW_21
timestamp 1713067540
transform 0 1 20859 -1 0 5979
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_T8W2FW  sky130_fd_pr__nfet_g5v0d10v5_T8W2FW_22
timestamp 1713067540
transform 0 1 20859 -1 0 6779
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_T8W2FW  sky130_fd_pr__nfet_g5v0d10v5_T8W2FW_23
timestamp 1713067540
transform 0 1 20859 -1 0 7579
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_T8W2FW  sky130_fd_pr__nfet_g5v0d10v5_T8W2FW_24
timestamp 1713067540
transform 0 1 20859 -1 0 8379
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_T8W2FW  sky130_fd_pr__nfet_g5v0d10v5_T8W2FW_25
timestamp 1713067540
transform 0 1 20859 -1 0 9179
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_T8W2FW  sky130_fd_pr__nfet_g5v0d10v5_T8W2FW_26
timestamp 1713067540
transform 0 1 20859 -1 0 9979
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_T8W2FW  sky130_fd_pr__nfet_g5v0d10v5_T8W2FW_27
timestamp 1713067540
transform 0 1 20859 -1 0 10779
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_T8W2FW  sky130_fd_pr__nfet_g5v0d10v5_T8W2FW_28
timestamp 1713067540
transform 0 1 20859 -1 0 11579
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_T8W2FW  sky130_fd_pr__nfet_g5v0d10v5_T8W2FW_29
timestamp 1713067540
transform 0 1 18659 -1 0 11579
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_T8W2FW  sky130_fd_pr__nfet_g5v0d10v5_T8W2FW_30
timestamp 1713067540
transform 0 1 16459 -1 0 11579
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_T8W2FW  sky130_fd_pr__nfet_g5v0d10v5_T8W2FW_31
timestamp 1713067540
transform 0 1 14259 -1 0 11579
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_T8W2FW  sky130_fd_pr__nfet_g5v0d10v5_T8W2FW_32
timestamp 1713067540
transform 0 1 12059 -1 0 11579
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_T8W2FW  sky130_fd_pr__nfet_g5v0d10v5_T8W2FW_33
timestamp 1713067540
transform 0 1 9859 -1 0 11579
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_T8W2FW  sky130_fd_pr__nfet_g5v0d10v5_T8W2FW_34
timestamp 1713067540
transform 0 1 7659 -1 0 11579
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_T8W2FW  sky130_fd_pr__nfet_g5v0d10v5_T8W2FW_35
timestamp 1713067540
transform 0 1 5459 -1 0 11579
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_V7WNNP  sky130_fd_pr__nfet_g5v0d10v5_V7WNNP_0
array 0 3 -1800 0 23 1600
timestamp 1713067540
transform 0 1 568 -1 0 -4597
box -328 -767 328 767
use sky130_fd_pr__nfet_g5v0d10v5_WGHV7X  sky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0
array 0 3 -1800 0 23 1600
timestamp 1713067540
transform 0 1 568 -1 0 -3771
box -628 -767 628 767
use sky130_fd_pr__pfet_g5v0d10v5_CRL9SD  sky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0
array 0 7 -800 0 7 2200
timestamp 1713067540
transform 0 1 3267 -1 0 -30902
box -408 -1097 408 1097
use sky130_fd_pr__pfet_g5v0d10v5_CS979Q  sky130_fd_pr__pfet_g5v0d10v5_CS979Q_0
array 0 7 -1800 0 23 1600
timestamp 1713067540
transform 0 1 575 -1 0 -21742
box -658 -815 658 815
use sky130_fd_pr__pfet_g5v0d10v5_GHE6GF  sky130_fd_pr__pfet_g5v0d10v5_GHE6GF_0
array 0 7 -1800 0 23 1600
timestamp 1713067540
transform 0 1 575 -1 0 -20916
box -358 -815 358 815
use sky130_fd_pr__pfet_g5v0d10v5_PJ2Z6Q  sky130_fd_pr__pfet_g5v0d10v5_PJ2Z6Q_0
timestamp 1713076297
transform 1 0 31625 0 1 10462
box -545 -662 545 662
use sky130_fd_pr__pfet_g5v0d10v5_PJ2Z6Q  sky130_fd_pr__pfet_g5v0d10v5_PJ2Z6Q_1
timestamp 1713076297
transform 1 0 29545 0 1 10462
box -545 -662 545 662
use sky130_fd_pr__pfet_g5v0d10v5_PJ2Z6Q  sky130_fd_pr__pfet_g5v0d10v5_PJ2Z6Q_2
timestamp 1713076297
transform 1 0 30585 0 1 10462
box -545 -662 545 662
use sky130_fd_pr__pfet_g5v0d10v5_PJ2ZJN  sky130_fd_pr__pfet_g5v0d10v5_PJ2ZJN_0
timestamp 1713076297
transform 1 0 29545 0 1 9162
box -545 -662 545 662
use sky130_fd_pr__pfet_g5v0d10v5_PJ2ZJN  sky130_fd_pr__pfet_g5v0d10v5_PJ2ZJN_1
timestamp 1713076297
transform 1 0 30585 0 1 9162
box -545 -662 545 662
use sky130_fd_pr__pfet_g5v0d10v5_PJ2ZJN  sky130_fd_pr__pfet_g5v0d10v5_PJ2ZJN_2
timestamp 1713076297
transform 1 0 31625 0 1 9162
box -545 -662 545 662
use sky130_fd_pr__pfet_g5v0d10v5_PNRDLC  sky130_fd_pr__pfet_g5v0d10v5_PNRDLC_0
timestamp 1713074216
transform 0 1 20867 -1 0 -25302
box -408 -1097 408 1097
use sky130_fd_pr__pfet_g5v0d10v5_PNRDLC  sky130_fd_pr__pfet_g5v0d10v5_PNRDLC_1
timestamp 1713074216
transform 0 1 3267 -1 0 -31702
box -408 -1097 408 1097
use sky130_fd_pr__pfet_g5v0d10v5_PNRDLC  sky130_fd_pr__pfet_g5v0d10v5_PNRDLC_2
timestamp 1713074216
transform 0 1 5467 -1 0 -31702
box -408 -1097 408 1097
use sky130_fd_pr__pfet_g5v0d10v5_PNRDLC  sky130_fd_pr__pfet_g5v0d10v5_PNRDLC_3
timestamp 1713074216
transform 0 1 7667 -1 0 -31702
box -408 -1097 408 1097
use sky130_fd_pr__pfet_g5v0d10v5_PNRDLC  sky130_fd_pr__pfet_g5v0d10v5_PNRDLC_4
timestamp 1713074216
transform 0 1 9867 -1 0 -31702
box -408 -1097 408 1097
use sky130_fd_pr__pfet_g5v0d10v5_PNRDLC  sky130_fd_pr__pfet_g5v0d10v5_PNRDLC_5
timestamp 1713074216
transform 0 1 12067 -1 0 -31702
box -408 -1097 408 1097
use sky130_fd_pr__pfet_g5v0d10v5_PNRDLC  sky130_fd_pr__pfet_g5v0d10v5_PNRDLC_6
timestamp 1713074216
transform 0 1 14267 -1 0 -31702
box -408 -1097 408 1097
use sky130_fd_pr__pfet_g5v0d10v5_PNRDLC  sky130_fd_pr__pfet_g5v0d10v5_PNRDLC_7
timestamp 1713074216
transform 0 1 16467 -1 0 -31702
box -408 -1097 408 1097
use sky130_fd_pr__pfet_g5v0d10v5_PNRDLC  sky130_fd_pr__pfet_g5v0d10v5_PNRDLC_8
timestamp 1713074216
transform 0 1 18667 -1 0 -31702
box -408 -1097 408 1097
use sky130_fd_pr__pfet_g5v0d10v5_PNRDLC  sky130_fd_pr__pfet_g5v0d10v5_PNRDLC_9
timestamp 1713074216
transform 0 1 20867 -1 0 -31702
box -408 -1097 408 1097
use sky130_fd_pr__pfet_g5v0d10v5_PNRDLC  sky130_fd_pr__pfet_g5v0d10v5_PNRDLC_10
timestamp 1713074216
transform 0 1 20867 -1 0 -30902
box -408 -1097 408 1097
use sky130_fd_pr__pfet_g5v0d10v5_PNRDLC  sky130_fd_pr__pfet_g5v0d10v5_PNRDLC_11
timestamp 1713074216
transform 0 1 20867 -1 0 -30102
box -408 -1097 408 1097
use sky130_fd_pr__pfet_g5v0d10v5_PNRDLC  sky130_fd_pr__pfet_g5v0d10v5_PNRDLC_12
timestamp 1713074216
transform 0 1 20867 -1 0 -29302
box -408 -1097 408 1097
use sky130_fd_pr__pfet_g5v0d10v5_PNRDLC  sky130_fd_pr__pfet_g5v0d10v5_PNRDLC_13
timestamp 1713074216
transform 0 1 20867 -1 0 -28502
box -408 -1097 408 1097
use sky130_fd_pr__pfet_g5v0d10v5_PNRDLC  sky130_fd_pr__pfet_g5v0d10v5_PNRDLC_14
timestamp 1713074216
transform 0 1 20867 -1 0 -27702
box -408 -1097 408 1097
use sky130_fd_pr__pfet_g5v0d10v5_PNRDLC  sky130_fd_pr__pfet_g5v0d10v5_PNRDLC_15
timestamp 1713074216
transform 0 1 20867 -1 0 -26902
box -408 -1097 408 1097
use sky130_fd_pr__pfet_g5v0d10v5_PNRDLC  sky130_fd_pr__pfet_g5v0d10v5_PNRDLC_16
timestamp 1713074216
transform 0 1 20867 -1 0 -26102
box -408 -1097 408 1097
use sky130_fd_pr__pfet_g5v0d10v5_PNRDLC  sky130_fd_pr__pfet_g5v0d10v5_PNRDLC_17
timestamp 1713074216
transform 0 1 1067 -1 0 -31702
box -408 -1097 408 1097
use sky130_fd_pr__pfet_g5v0d10v5_PNRDLC  sky130_fd_pr__pfet_g5v0d10v5_PNRDLC_18
timestamp 1713074216
transform 0 1 20867 -1 0 -24502
box -408 -1097 408 1097
use sky130_fd_pr__pfet_g5v0d10v5_PNRDLC  sky130_fd_pr__pfet_g5v0d10v5_PNRDLC_19
timestamp 1713074216
transform 0 1 18667 -1 0 -24502
box -408 -1097 408 1097
use sky130_fd_pr__pfet_g5v0d10v5_PNRDLC  sky130_fd_pr__pfet_g5v0d10v5_PNRDLC_20
timestamp 1713074216
transform 0 1 16467 -1 0 -24502
box -408 -1097 408 1097
use sky130_fd_pr__pfet_g5v0d10v5_PNRDLC  sky130_fd_pr__pfet_g5v0d10v5_PNRDLC_21
timestamp 1713074216
transform 0 1 14267 -1 0 -24502
box -408 -1097 408 1097
use sky130_fd_pr__pfet_g5v0d10v5_PNRDLC  sky130_fd_pr__pfet_g5v0d10v5_PNRDLC_22
timestamp 1713074216
transform 0 1 12067 -1 0 -24502
box -408 -1097 408 1097
use sky130_fd_pr__pfet_g5v0d10v5_PNRDLC  sky130_fd_pr__pfet_g5v0d10v5_PNRDLC_23
timestamp 1713074216
transform 0 1 9867 -1 0 -24502
box -408 -1097 408 1097
use sky130_fd_pr__pfet_g5v0d10v5_PNRDLC  sky130_fd_pr__pfet_g5v0d10v5_PNRDLC_24
timestamp 1713074216
transform 0 1 7667 -1 0 -24502
box -408 -1097 408 1097
use sky130_fd_pr__pfet_g5v0d10v5_PNRDLC  sky130_fd_pr__pfet_g5v0d10v5_PNRDLC_25
timestamp 1713074216
transform 0 1 5467 -1 0 -24502
box -408 -1097 408 1097
use sky130_fd_pr__pfet_g5v0d10v5_PNRDLC  sky130_fd_pr__pfet_g5v0d10v5_PNRDLC_26
timestamp 1713074216
transform 0 1 3267 -1 0 -24502
box -408 -1097 408 1097
use sky130_fd_pr__pfet_g5v0d10v5_PNRDLC  sky130_fd_pr__pfet_g5v0d10v5_PNRDLC_27
timestamp 1713074216
transform 0 1 1067 -1 0 -24502
box -408 -1097 408 1097
use sky130_fd_pr__pfet_g5v0d10v5_PNRDLC  sky130_fd_pr__pfet_g5v0d10v5_PNRDLC_28
timestamp 1713074216
transform 0 1 1067 -1 0 -25302
box -408 -1097 408 1097
use sky130_fd_pr__pfet_g5v0d10v5_PNRDLC  sky130_fd_pr__pfet_g5v0d10v5_PNRDLC_29
timestamp 1713074216
transform 0 1 1067 -1 0 -26102
box -408 -1097 408 1097
use sky130_fd_pr__pfet_g5v0d10v5_PNRDLC  sky130_fd_pr__pfet_g5v0d10v5_PNRDLC_30
timestamp 1713074216
transform 0 1 1067 -1 0 -26902
box -408 -1097 408 1097
use sky130_fd_pr__pfet_g5v0d10v5_PNRDLC  sky130_fd_pr__pfet_g5v0d10v5_PNRDLC_31
timestamp 1713074216
transform 0 1 1067 -1 0 -27702
box -408 -1097 408 1097
use sky130_fd_pr__pfet_g5v0d10v5_PNRDLC  sky130_fd_pr__pfet_g5v0d10v5_PNRDLC_32
timestamp 1713074216
transform 0 1 1067 -1 0 -28502
box -408 -1097 408 1097
use sky130_fd_pr__pfet_g5v0d10v5_PNRDLC  sky130_fd_pr__pfet_g5v0d10v5_PNRDLC_33
timestamp 1713074216
transform 0 1 1067 -1 0 -29302
box -408 -1097 408 1097
use sky130_fd_pr__pfet_g5v0d10v5_PNRDLC  sky130_fd_pr__pfet_g5v0d10v5_PNRDLC_34
timestamp 1713074216
transform 0 1 1067 -1 0 -30102
box -408 -1097 408 1097
use sky130_fd_pr__pfet_g5v0d10v5_PNRDLC  sky130_fd_pr__pfet_g5v0d10v5_PNRDLC_35
timestamp 1713074216
transform 0 1 1067 -1 0 -30902
box -408 -1097 408 1097
use sky130_fd_pr__res_high_po_2p85_XPXHHN  sky130_fd_pr__res_high_po_2p85_XPXHHN_0
timestamp 1713072694
transform 1 0 25715 0 1 8278
box -3115 -2878 3115 2878
<< end >>
