magic
tech sky130A
magscale 1 2
timestamp 1713067540
<< nwell >>
rect -358 -815 358 815
<< mvpmos >>
rect -100 118 100 518
rect -100 -518 100 -118
<< mvpdiff >>
rect -158 506 -100 518
rect -158 130 -146 506
rect -112 130 -100 506
rect -158 118 -100 130
rect 100 506 158 518
rect 100 130 112 506
rect 146 130 158 506
rect 100 118 158 130
rect -158 -130 -100 -118
rect -158 -506 -146 -130
rect -112 -506 -100 -130
rect -158 -518 -100 -506
rect 100 -130 158 -118
rect 100 -506 112 -130
rect 146 -506 158 -130
rect 100 -518 158 -506
<< mvpdiffc >>
rect -146 130 -112 506
rect 112 130 146 506
rect -146 -506 -112 -130
rect 112 -506 146 -130
<< mvnsubdiff >>
rect -292 737 292 749
rect -292 703 -184 737
rect 184 703 292 737
rect -292 691 292 703
rect -292 641 -234 691
rect -292 -641 -280 641
rect -246 -641 -234 641
rect 234 641 292 691
rect -292 -691 -234 -641
rect 234 -641 246 641
rect 280 -641 292 641
rect 234 -691 292 -641
rect -292 -703 292 -691
rect -292 -737 -184 -703
rect 184 -737 292 -703
rect -292 -749 292 -737
<< mvnsubdiffcont >>
rect -184 703 184 737
rect -280 -641 -246 641
rect 246 -641 280 641
rect -184 -737 184 -703
<< poly >>
rect -100 599 100 615
rect -100 565 -84 599
rect 84 565 100 599
rect -100 518 100 565
rect -100 71 100 118
rect -100 37 -84 71
rect 84 37 100 71
rect -100 21 100 37
rect -100 -37 100 -21
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -100 -118 100 -71
rect -100 -565 100 -518
rect -100 -599 -84 -565
rect 84 -599 100 -565
rect -100 -615 100 -599
<< polycont >>
rect -84 565 84 599
rect -84 37 84 71
rect -84 -71 84 -37
rect -84 -599 84 -565
<< locali >>
rect -280 703 -184 737
rect 184 703 280 737
rect -280 641 -246 703
rect 246 641 280 703
rect -100 565 -84 599
rect 84 565 100 599
rect -146 506 -112 522
rect -146 114 -112 130
rect 112 506 146 522
rect 112 114 146 130
rect -100 37 -84 71
rect 84 37 100 71
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -146 -130 -112 -114
rect -146 -522 -112 -506
rect 112 -130 146 -114
rect 112 -522 146 -506
rect -100 -599 -84 -565
rect 84 -599 100 -565
rect -280 -703 -246 -641
rect 246 -703 280 -641
rect -280 -737 -184 -703
rect 184 -737 280 -703
<< viali >>
rect -67 565 67 599
rect -146 130 -112 506
rect 112 130 146 506
rect -67 37 67 71
rect -67 -71 67 -37
rect -146 -506 -112 -130
rect 112 -506 146 -130
rect -67 -599 67 -565
<< metal1 >>
rect -79 599 79 605
rect -79 565 -67 599
rect 67 565 79 599
rect -79 559 79 565
rect -152 506 -106 518
rect -152 130 -146 506
rect -112 130 -106 506
rect -152 118 -106 130
rect 106 506 152 518
rect 106 130 112 506
rect 146 130 152 506
rect 106 118 152 130
rect -79 71 79 77
rect -79 37 -67 71
rect 67 37 79 71
rect -79 31 79 37
rect -79 -37 79 -31
rect -79 -71 -67 -37
rect 67 -71 79 -37
rect -79 -77 79 -71
rect -152 -130 -106 -118
rect -152 -506 -146 -130
rect -112 -506 -106 -130
rect -152 -518 -106 -506
rect 106 -130 152 -118
rect 106 -506 112 -130
rect 146 -506 152 -130
rect 106 -518 152 -506
rect -79 -565 79 -559
rect -79 -599 -67 -565
rect 67 -599 79 -565
rect -79 -605 79 -599
<< properties >>
string FIXED_BBOX -263 -720 263 720
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 2 l 1 m 2 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 80 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
