magic
tech sky130A
magscale 1 2
timestamp 1713594760
<< error_p >>
rect -111 131 -47 137
rect 47 131 111 137
rect -111 97 -99 131
rect 47 97 59 131
rect -111 91 -47 97
rect 47 91 111 97
rect -111 -97 -47 -91
rect 47 -97 111 -91
rect -111 -131 -99 -97
rect 47 -131 59 -97
rect -111 -137 -47 -131
rect 47 -137 111 -131
<< nwell >>
rect -387 -347 387 347
<< mvpmos >>
rect -129 -50 -29 50
rect 29 -50 129 50
<< mvpdiff >>
rect -187 38 -129 50
rect -187 -38 -175 38
rect -141 -38 -129 38
rect -187 -50 -129 -38
rect -29 38 29 50
rect -29 -38 -17 38
rect 17 -38 29 38
rect -29 -50 29 -38
rect 129 38 187 50
rect 129 -38 141 38
rect 175 -38 187 38
rect 129 -50 187 -38
<< mvpdiffc >>
rect -175 -38 -141 38
rect -17 -38 17 38
rect 141 -38 175 38
<< mvnsubdiff >>
rect -321 269 321 281
rect -321 235 -213 269
rect 213 235 321 269
rect -321 223 321 235
rect -321 173 -263 223
rect -321 -173 -309 173
rect -275 -173 -263 173
rect 263 173 321 223
rect -321 -223 -263 -173
rect 263 -173 275 173
rect 309 -173 321 173
rect 263 -223 321 -173
rect -321 -235 321 -223
rect -321 -269 -213 -235
rect 213 -269 321 -235
rect -321 -281 321 -269
<< mvnsubdiffcont >>
rect -213 235 213 269
rect -309 -173 -275 173
rect 275 -173 309 173
rect -213 -269 213 -235
<< poly >>
rect -129 131 -29 147
rect -129 97 -113 131
rect -45 97 -29 131
rect -129 50 -29 97
rect 29 131 129 147
rect 29 97 45 131
rect 113 97 129 131
rect 29 50 129 97
rect -129 -97 -29 -50
rect -129 -131 -113 -97
rect -45 -131 -29 -97
rect -129 -147 -29 -131
rect 29 -97 129 -50
rect 29 -131 45 -97
rect 113 -131 129 -97
rect 29 -147 129 -131
<< polycont >>
rect -113 97 -45 131
rect 45 97 113 131
rect -113 -131 -45 -97
rect 45 -131 113 -97
<< locali >>
rect -309 235 -220 269
rect 220 235 309 269
rect -309 188 -275 235
rect 275 188 309 235
rect -129 97 -113 131
rect -45 97 -29 131
rect 29 97 45 131
rect 113 97 129 131
rect -175 38 -141 54
rect -175 -54 -141 -38
rect -17 38 17 54
rect -17 -54 17 -38
rect 141 38 175 54
rect 141 -54 175 -38
rect -129 -131 -113 -97
rect -45 -131 -29 -97
rect 29 -131 45 -97
rect 113 -131 129 -97
rect -309 -235 -275 -188
rect 275 -235 309 -188
rect -309 -269 -213 -235
rect 213 -269 309 -235
<< viali >>
rect -220 235 -213 269
rect -213 235 213 269
rect 213 235 220 269
rect -309 173 -275 188
rect -309 -173 -275 173
rect 275 173 309 188
rect -99 97 -59 131
rect 59 97 99 131
rect -175 -38 -141 38
rect -17 -38 17 38
rect 141 -38 175 38
rect -99 -131 -59 -97
rect 59 -131 99 -97
rect -309 -188 -275 -173
rect 275 -173 309 173
rect 275 -188 309 -173
<< metal1 >>
rect -232 269 232 275
rect -232 235 -220 269
rect 220 235 232 269
rect -232 229 232 235
rect -315 188 -269 200
rect -315 -188 -309 188
rect -275 -188 -269 188
rect 269 188 315 200
rect -111 131 -47 137
rect -111 97 -99 131
rect -59 97 -47 131
rect -111 91 -47 97
rect 47 131 111 137
rect 47 97 59 131
rect 99 97 111 131
rect 47 91 111 97
rect -181 38 -135 50
rect -181 -38 -175 38
rect -141 -38 -135 38
rect -181 -50 -135 -38
rect -23 38 23 50
rect -23 -38 -17 38
rect 17 -38 23 38
rect -23 -50 23 -38
rect 135 38 181 50
rect 135 -38 141 38
rect 175 -38 181 38
rect 135 -50 181 -38
rect -111 -97 -47 -91
rect -111 -131 -99 -97
rect -59 -131 -47 -97
rect -111 -137 -47 -131
rect 47 -97 111 -91
rect 47 -131 59 -97
rect 99 -131 111 -97
rect 47 -137 111 -131
rect -315 -200 -269 -188
rect 269 -188 275 188
rect 309 -188 315 188
rect 269 -200 315 -188
<< properties >>
string FIXED_BBOX -292 -252 292 252
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 0.5 l 0.50 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 60 viagb 0 viagr 80 viagl 80 viagt 80
<< end >>
