magic
tech sky130A
magscale 1 2
timestamp 1713575337
<< nwell >>
rect -1087 -815 1087 815
<< mvpmos >>
rect -829 118 -29 518
rect 29 118 829 518
rect -829 -518 -29 -118
rect 29 -518 829 -118
<< mvpdiff >>
rect -887 506 -829 518
rect -887 130 -875 506
rect -841 130 -829 506
rect -887 118 -829 130
rect -29 506 29 518
rect -29 130 -17 506
rect 17 130 29 506
rect -29 118 29 130
rect 829 506 887 518
rect 829 130 841 506
rect 875 130 887 506
rect 829 118 887 130
rect -887 -130 -829 -118
rect -887 -506 -875 -130
rect -841 -506 -829 -130
rect -887 -518 -829 -506
rect -29 -130 29 -118
rect -29 -506 -17 -130
rect 17 -506 29 -130
rect -29 -518 29 -506
rect 829 -130 887 -118
rect 829 -506 841 -130
rect 875 -506 887 -130
rect 829 -518 887 -506
<< mvpdiffc >>
rect -875 130 -841 506
rect -17 130 17 506
rect 841 130 875 506
rect -875 -506 -841 -130
rect -17 -506 17 -130
rect 841 -506 875 -130
<< mvnsubdiff >>
rect -1021 737 1021 749
rect -1021 703 -913 737
rect 913 703 1021 737
rect -1021 691 1021 703
rect -1021 641 -963 691
rect -1021 -641 -1009 641
rect -975 -641 -963 641
rect 963 641 1021 691
rect -1021 -691 -963 -641
rect 963 -641 975 641
rect 1009 -641 1021 641
rect 963 -691 1021 -641
rect -1021 -703 1021 -691
rect -1021 -737 -913 -703
rect 913 -737 1021 -703
rect -1021 -749 1021 -737
<< mvnsubdiffcont >>
rect -913 703 913 737
rect -1009 -641 -975 641
rect 975 -641 1009 641
rect -913 -737 913 -703
<< poly >>
rect -829 599 -29 615
rect -829 565 -813 599
rect -45 565 -29 599
rect -829 518 -29 565
rect 29 599 829 615
rect 29 565 45 599
rect 813 565 829 599
rect 29 518 829 565
rect -829 71 -29 118
rect -829 37 -813 71
rect -45 37 -29 71
rect -829 21 -29 37
rect 29 71 829 118
rect 29 37 45 71
rect 813 37 829 71
rect 29 21 829 37
rect -829 -37 -29 -21
rect -829 -71 -813 -37
rect -45 -71 -29 -37
rect -829 -118 -29 -71
rect 29 -37 829 -21
rect 29 -71 45 -37
rect 813 -71 829 -37
rect 29 -118 829 -71
rect -829 -565 -29 -518
rect -829 -599 -813 -565
rect -45 -599 -29 -565
rect -829 -615 -29 -599
rect 29 -565 829 -518
rect 29 -599 45 -565
rect 813 -599 829 -565
rect 29 -615 829 -599
<< polycont >>
rect -813 565 -45 599
rect 45 565 813 599
rect -813 37 -45 71
rect 45 37 813 71
rect -813 -71 -45 -37
rect 45 -71 813 -37
rect -813 -599 -45 -565
rect 45 -599 813 -565
<< locali >>
rect -1009 703 -913 737
rect 913 703 1009 737
rect -1009 641 -975 703
rect 975 641 1009 703
rect -829 565 -813 599
rect -45 565 -29 599
rect 29 565 45 599
rect 813 565 829 599
rect -875 506 -841 522
rect -875 114 -841 130
rect -17 506 17 522
rect -17 114 17 130
rect 841 506 875 522
rect 841 114 875 130
rect -829 37 -813 71
rect -45 37 -29 71
rect 29 37 45 71
rect 813 37 829 71
rect -829 -71 -813 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 813 -71 829 -37
rect -875 -130 -841 -114
rect -875 -522 -841 -506
rect -17 -130 17 -114
rect -17 -522 17 -506
rect 841 -130 875 -114
rect 841 -522 875 -506
rect -829 -599 -813 -565
rect -45 -599 -29 -565
rect 29 -599 45 -565
rect 813 -599 829 -565
rect -1009 -703 -975 -641
rect 975 -703 1009 -641
rect -1009 -737 -913 -703
rect 913 -737 1009 -703
<< viali >>
rect -780 703 780 737
rect -813 565 -45 599
rect 45 565 813 599
rect -875 130 -841 506
rect -17 130 17 506
rect 841 130 875 506
rect -813 37 -45 71
rect 45 37 813 71
rect -813 -71 -45 -37
rect 45 -71 813 -37
rect -875 -506 -841 -130
rect -17 -506 17 -130
rect 841 -506 875 -130
rect 975 -562 1009 562
rect -813 -599 -45 -565
rect 45 -599 813 -565
<< metal1 >>
rect -792 737 792 743
rect -792 703 -780 737
rect 780 703 792 737
rect -792 697 792 703
rect -825 599 -33 605
rect -825 565 -813 599
rect -45 565 -33 599
rect -825 559 -33 565
rect 33 599 825 605
rect 33 565 45 599
rect 813 565 825 599
rect 33 559 825 565
rect 969 562 1015 574
rect -881 506 -835 518
rect -881 130 -875 506
rect -841 130 -835 506
rect -881 118 -835 130
rect -23 506 23 518
rect -23 130 -17 506
rect 17 130 23 506
rect -23 118 23 130
rect 835 506 881 518
rect 835 130 841 506
rect 875 130 881 506
rect 835 118 881 130
rect -825 71 -33 77
rect -825 37 -813 71
rect -45 37 -33 71
rect -825 31 -33 37
rect 33 71 825 77
rect 33 37 45 71
rect 813 37 825 71
rect 33 31 825 37
rect -825 -37 -33 -31
rect -825 -71 -813 -37
rect -45 -71 -33 -37
rect -825 -77 -33 -71
rect 33 -37 825 -31
rect 33 -71 45 -37
rect 813 -71 825 -37
rect 33 -77 825 -71
rect -881 -130 -835 -118
rect -881 -506 -875 -130
rect -841 -506 -835 -130
rect -881 -518 -835 -506
rect -23 -130 23 -118
rect -23 -506 -17 -130
rect 17 -506 23 -130
rect -23 -518 23 -506
rect 835 -130 881 -118
rect 835 -506 841 -130
rect 875 -506 881 -130
rect 835 -518 881 -506
rect -825 -565 -33 -559
rect -825 -599 -813 -565
rect -45 -599 -33 -565
rect -825 -605 -33 -599
rect 33 -565 825 -559
rect 33 -599 45 -565
rect 813 -599 825 -565
rect 969 -562 975 562
rect 1009 -562 1015 562
rect 969 -574 1015 -562
rect 33 -605 825 -599
<< properties >>
string FIXED_BBOX -992 -720 992 720
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 2 l 4 m 2 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 80 viagl 0 viagt 80
<< end >>
