magic
tech sky130A
magscale 1 2
timestamp 1713382499
<< nwell >>
rect 27700 10800 29024 11670
rect 29932 10800 36542 11204
rect 27700 10210 36542 10800
rect 27700 6600 32200 10210
rect 32760 8858 34450 9078
rect 32760 8020 35702 8858
rect 32760 7840 34450 8020
rect 27700 5380 29024 6600
rect 29460 6560 32194 6600
rect 27700 4060 29016 5380
rect -200 -7958 38400 -7600
rect -240 -22400 38400 -7958
rect -200 -23800 38400 -22400
rect -200 -32200 27370 -23800
rect 30200 -29200 38400 -23800
rect 31600 -29218 38210 -29200
rect 31612 -31800 38222 -30806
<< pwell >>
rect -200 3600 27400 12200
rect 29986 11985 30178 11986
rect 31670 11985 31780 11986
rect 31912 11985 31956 11986
rect 32186 11985 32378 11986
rect 33870 11985 33980 11986
rect 34112 11985 34156 11986
rect 34386 11985 34578 11986
rect 36070 11985 36180 11986
rect 36312 11985 36356 11986
rect 29920 11269 32111 11985
rect 32120 11269 34311 11985
rect 34320 11269 36511 11985
rect 31710 11264 31754 11269
rect 33910 11264 33954 11269
rect 36110 11264 36154 11269
rect 29500 6400 30816 6416
rect 30840 6400 32156 6416
rect 32600 6400 35800 7800
rect 29500 5760 35800 6400
rect 36200 6182 38200 6200
rect 29600 5156 35800 5760
rect 29500 4600 35800 5156
rect 29500 4500 30816 4600
rect 30840 4500 32156 4600
rect 32540 3600 34202 4216
rect 34730 3600 35602 4216
rect 36190 3720 38200 6182
rect 36200 3600 38200 3720
rect -200 -5000 38200 3600
rect 27740 -25370 28996 -24454
rect 27740 -26390 28994 -25370
rect 27740 -27430 28994 -26400
rect 27740 -28470 28994 -27440
rect 27740 -29510 28994 -28480
rect 31988 -29283 32032 -29278
rect 34188 -29283 34232 -29278
rect 36388 -29283 36432 -29278
rect 27740 -30550 28994 -29520
rect 31631 -29999 33822 -29283
rect 33831 -29999 36022 -29283
rect 36031 -29999 38222 -29283
rect 31786 -30000 31830 -29999
rect 31962 -30000 32072 -29999
rect 33564 -30000 33756 -29999
rect 33986 -30000 34030 -29999
rect 34162 -30000 34272 -29999
rect 35764 -30000 35956 -29999
rect 36186 -30000 36230 -29999
rect 36362 -30000 36472 -29999
rect 37964 -30000 38156 -29999
rect 31666 -30025 31858 -30024
rect 33350 -30025 33460 -30024
rect 33592 -30025 33636 -30024
rect 33866 -30025 34058 -30024
rect 35550 -30025 35660 -30024
rect 35792 -30025 35836 -30024
rect 36066 -30025 36258 -30024
rect 37750 -30025 37860 -30024
rect 37992 -30025 38036 -30024
rect 27740 -31590 28994 -30560
rect 31600 -30741 33791 -30025
rect 33800 -30741 35991 -30025
rect 36000 -30741 38191 -30025
rect 33390 -30746 33434 -30741
rect 35590 -30746 35634 -30741
rect 37790 -30746 37834 -30741
<< nmos >>
rect 34636 7130 34666 7330
rect 35056 7130 35086 7330
rect 35476 7130 35506 7330
<< pmos >>
rect 32956 8059 33156 8859
rect 33214 8059 33414 8859
rect 33796 8059 33996 8859
rect 34054 8059 34254 8859
rect 34636 8239 34666 8639
rect 35056 8239 35086 8639
rect 35476 8239 35506 8639
<< mvnmos >>
rect 259 11429 1859 11729
rect 2459 11429 4059 11729
rect 4659 11429 6259 11729
rect 6859 11429 8459 11729
rect 9059 11429 10659 11729
rect 11259 11429 12859 11729
rect 13459 11429 15059 11729
rect 15659 11429 17259 11729
rect 17859 11429 19459 11729
rect 20059 11429 21659 11729
rect 259 10629 1859 10929
rect 2458 10628 4058 10928
rect 4658 10628 6258 10928
rect 6858 10628 8458 10928
rect 9058 10628 10658 10928
rect 11258 10628 12858 10928
rect 13458 10628 15058 10928
rect 15658 10628 17258 10928
rect 17858 10628 19458 10928
rect 20059 10629 21659 10929
rect 259 9829 1859 10129
rect 2458 9828 4058 10128
rect 4658 9828 6258 10128
rect 6858 9828 8458 10128
rect 9058 9828 10658 10128
rect 11258 9828 12858 10128
rect 13458 9828 15058 10128
rect 15658 9828 17258 10128
rect 17858 9828 19458 10128
rect 20059 9829 21659 10129
rect 259 9029 1859 9329
rect 2458 9028 4058 9328
rect 4658 9028 6258 9328
rect 6858 9028 8458 9328
rect 9058 9028 10658 9328
rect 11258 9028 12858 9328
rect 13458 9028 15058 9328
rect 15658 9028 17258 9328
rect 17858 9028 19458 9328
rect 20059 9029 21659 9329
rect 259 8229 1859 8529
rect 2458 8228 4058 8528
rect 4658 8228 6258 8528
rect 6858 8228 8458 8528
rect 9058 8228 10658 8528
rect 11258 8228 12858 8528
rect 13458 8228 15058 8528
rect 15658 8228 17258 8528
rect 17858 8228 19458 8528
rect 20059 8229 21659 8529
rect 259 7429 1859 7729
rect 2458 7428 4058 7728
rect 4658 7428 6258 7728
rect 6858 7428 8458 7728
rect 9058 7428 10658 7728
rect 11258 7428 12858 7728
rect 13458 7428 15058 7728
rect 15658 7428 17258 7728
rect 17858 7428 19458 7728
rect 20059 7429 21659 7729
rect 259 6629 1859 6929
rect 2458 6628 4058 6928
rect 4658 6628 6258 6928
rect 6858 6628 8458 6928
rect 9058 6628 10658 6928
rect 11258 6628 12858 6928
rect 13458 6628 15058 6928
rect 15658 6628 17258 6928
rect 17858 6628 19458 6928
rect 20059 6629 21659 6929
rect 259 5829 1859 6129
rect 2458 5828 4058 6128
rect 4658 5828 6258 6128
rect 6858 5828 8458 6128
rect 9058 5828 10658 6128
rect 11258 5828 12858 6128
rect 13458 5828 15058 6128
rect 15658 5828 17258 6128
rect 17858 5828 19458 6128
rect 20059 5829 21659 6129
rect 259 5029 1859 5329
rect 2458 5028 4058 5328
rect 4658 5028 6258 5328
rect 6858 5028 8458 5328
rect 9058 5028 10658 5328
rect 11258 5028 12858 5328
rect 13458 5028 15058 5328
rect 15658 5028 17258 5328
rect 17858 5028 19458 5328
rect 20059 5029 21659 5329
rect 259 4229 1859 4529
rect 2459 4229 4059 4529
rect 4659 4229 6259 4529
rect 6859 4229 8459 4529
rect 9060 4230 10660 4530
rect 11260 4230 12860 4530
rect 13459 4229 15059 4529
rect 15659 4229 17259 4529
rect 17859 4229 19459 4529
rect 20059 4229 21659 4529
rect 30148 11527 30248 11727
rect 30306 11527 30406 11727
rect 30464 11527 30564 11727
rect 30903 11527 31003 11727
rect 31343 11527 31443 11727
rect 31783 11527 31883 11727
rect 32348 11527 32448 11727
rect 32506 11527 32606 11727
rect 32664 11527 32764 11727
rect 33103 11527 33203 11727
rect 33543 11527 33643 11727
rect 33983 11527 34083 11727
rect 34548 11527 34648 11727
rect 34706 11527 34806 11727
rect 34864 11527 34964 11727
rect 35303 11527 35403 11727
rect 35743 11527 35843 11727
rect 36183 11527 36283 11727
rect 33518 7038 33618 7438
rect 33676 7038 33776 7438
rect 33834 7038 33934 7438
rect 33992 7038 34092 7438
rect 29758 5988 30558 6188
rect 31098 5988 31898 6188
rect 29968 5408 30368 5508
rect 31278 5408 31678 5508
rect 29758 4728 30558 4928
rect 31098 4728 31898 4928
rect 17148 2516 17248 3316
rect 17306 2516 17406 3316
rect 17464 2516 17564 3316
rect 17622 2516 17722 3316
rect 32768 3558 32868 3958
rect 32926 3558 33026 3958
rect 33084 3558 33184 3958
rect 33242 3558 33342 3958
rect 33400 3558 33500 3958
rect 33558 3558 33658 3958
rect 33716 3558 33816 3958
rect 33874 3558 33974 3958
rect 34958 3558 35058 3958
rect 35116 3558 35216 3958
rect 35274 3558 35374 3958
rect 36448 5754 36848 5954
rect 36448 5496 36848 5696
rect 36448 5238 36848 5438
rect 36448 4980 36848 5180
rect 36448 4722 36848 4922
rect 36448 4464 36848 4664
rect 36448 4206 36848 4406
rect 36448 3948 36848 4148
rect 37234 5754 37634 5954
rect 37234 5496 37634 5696
rect 37234 5238 37634 5438
rect 37234 4980 37634 5180
rect 37234 4722 37634 4922
rect 37234 4464 37634 4664
rect 37234 4206 37634 4406
rect 37234 3948 37634 4148
rect 32438 2628 32538 3028
rect 32596 2628 32696 3028
rect 34038 2628 34138 3028
rect 34196 2628 34296 3028
rect 35638 2628 35738 3028
rect 35796 2628 35896 3028
rect 59 1249 459 2049
rect 677 1249 1077 2049
rect 59 703 459 903
rect 677 703 1077 903
rect 1659 1249 2059 2049
rect 2277 1249 2677 2049
rect 1659 703 2059 903
rect 2277 703 2677 903
rect 3259 1249 3659 2049
rect 3877 1249 4277 2049
rect 3259 703 3659 903
rect 3877 703 4277 903
rect 4859 1249 5259 2049
rect 5477 1249 5877 2049
rect 4859 703 5259 903
rect 5477 703 5877 903
rect 6459 1249 6859 2049
rect 7077 1249 7477 2049
rect 6459 703 6859 903
rect 7077 703 7477 903
rect 8059 1249 8459 2049
rect 8677 1249 9077 2049
rect 8059 703 8459 903
rect 8677 703 9077 903
rect 9659 1249 10059 2049
rect 10277 1249 10677 2049
rect 9659 703 10059 903
rect 10277 703 10677 903
rect 11259 1249 11659 2049
rect 11877 1249 12277 2049
rect 11259 703 11659 903
rect 11877 703 12277 903
rect 12859 1249 13259 2049
rect 13477 1249 13877 2049
rect 12859 703 13259 903
rect 13477 703 13877 903
rect 14459 1249 14859 2049
rect 15077 1249 15477 2049
rect 14459 703 14859 903
rect 15077 703 15477 903
rect 16059 1249 16459 2049
rect 16677 1249 17077 2049
rect 16059 703 16459 903
rect 16677 703 17077 903
rect 17659 1249 18059 2049
rect 18277 1249 18677 2049
rect 17659 703 18059 903
rect 18277 703 18677 903
rect 19259 1249 19659 2049
rect 19877 1249 20277 2049
rect 19259 703 19659 903
rect 19877 703 20277 903
rect 20859 1249 21259 2049
rect 21477 1249 21877 2049
rect 20859 703 21259 903
rect 21477 703 21877 903
rect 22459 1249 22859 2049
rect 23077 1249 23477 2049
rect 22459 703 22859 903
rect 23077 703 23477 903
rect 24059 1249 24459 2049
rect 24677 1249 25077 2049
rect 24059 703 24459 903
rect 24677 703 25077 903
rect 25659 1249 26059 2049
rect 26277 1249 26677 2049
rect 25659 703 26059 903
rect 26277 703 26677 903
rect 27259 1249 27659 2049
rect 27877 1249 28277 2049
rect 27259 703 27659 903
rect 27877 703 28277 903
rect 28859 1249 29259 2049
rect 29477 1249 29877 2049
rect 28859 703 29259 903
rect 29477 703 29877 903
rect 30459 1249 30859 2049
rect 31077 1249 31477 2049
rect 30459 703 30859 903
rect 31077 703 31477 903
rect 32059 1249 32459 2049
rect 32677 1249 33077 2049
rect 32059 703 32459 903
rect 32677 703 33077 903
rect 33659 1249 34059 2049
rect 34277 1249 34677 2049
rect 33659 703 34059 903
rect 34277 703 34677 903
rect 35259 1249 35659 2049
rect 35877 1249 36277 2049
rect 35259 703 35659 903
rect 35877 703 36277 903
rect 36859 1249 37259 2049
rect 37477 1249 37877 2049
rect 36859 703 37259 903
rect 37477 703 37877 903
rect 59 -551 459 249
rect 677 -551 1077 249
rect 59 -1097 459 -897
rect 677 -1097 1077 -897
rect 1659 -551 2059 249
rect 2277 -551 2677 249
rect 1659 -1097 2059 -897
rect 2277 -1097 2677 -897
rect 3259 -551 3659 249
rect 3877 -551 4277 249
rect 3259 -1097 3659 -897
rect 3877 -1097 4277 -897
rect 4859 -551 5259 249
rect 5477 -551 5877 249
rect 4859 -1097 5259 -897
rect 5477 -1097 5877 -897
rect 6459 -551 6859 249
rect 7077 -551 7477 249
rect 6459 -1097 6859 -897
rect 7077 -1097 7477 -897
rect 8059 -551 8459 249
rect 8677 -551 9077 249
rect 8059 -1097 8459 -897
rect 8677 -1097 9077 -897
rect 9659 -551 10059 249
rect 10277 -551 10677 249
rect 9659 -1097 10059 -897
rect 10277 -1097 10677 -897
rect 11259 -551 11659 249
rect 11877 -551 12277 249
rect 11259 -1097 11659 -897
rect 11877 -1097 12277 -897
rect 12859 -551 13259 249
rect 13477 -551 13877 249
rect 12859 -1097 13259 -897
rect 13477 -1097 13877 -897
rect 14459 -551 14859 249
rect 15077 -551 15477 249
rect 14459 -1097 14859 -897
rect 15077 -1097 15477 -897
rect 16059 -551 16459 249
rect 16677 -551 17077 249
rect 16059 -1097 16459 -897
rect 16677 -1097 17077 -897
rect 17659 -551 18059 249
rect 18277 -551 18677 249
rect 17659 -1097 18059 -897
rect 18277 -1097 18677 -897
rect 19259 -551 19659 249
rect 19877 -551 20277 249
rect 19259 -1097 19659 -897
rect 19877 -1097 20277 -897
rect 20859 -551 21259 249
rect 21477 -551 21877 249
rect 20859 -1097 21259 -897
rect 21477 -1097 21877 -897
rect 22459 -551 22859 249
rect 23077 -551 23477 249
rect 22459 -1097 22859 -897
rect 23077 -1097 23477 -897
rect 24059 -551 24459 249
rect 24677 -551 25077 249
rect 24059 -1097 24459 -897
rect 24677 -1097 25077 -897
rect 25659 -551 26059 249
rect 26277 -551 26677 249
rect 25659 -1097 26059 -897
rect 26277 -1097 26677 -897
rect 27259 -551 27659 249
rect 27877 -551 28277 249
rect 27259 -1097 27659 -897
rect 27877 -1097 28277 -897
rect 28859 -551 29259 249
rect 29477 -551 29877 249
rect 28859 -1097 29259 -897
rect 29477 -1097 29877 -897
rect 30459 -551 30859 249
rect 31077 -551 31477 249
rect 30459 -1097 30859 -897
rect 31077 -1097 31477 -897
rect 32059 -551 32459 249
rect 32677 -551 33077 249
rect 32059 -1097 32459 -897
rect 32677 -1097 33077 -897
rect 33659 -551 34059 249
rect 34277 -551 34677 249
rect 33659 -1097 34059 -897
rect 34277 -1097 34677 -897
rect 35259 -551 35659 249
rect 35877 -551 36277 249
rect 35259 -1097 35659 -897
rect 35877 -1097 36277 -897
rect 36859 -551 37259 249
rect 37477 -551 37877 249
rect 36859 -1097 37259 -897
rect 37477 -1097 37877 -897
rect 59 -2351 459 -1551
rect 677 -2351 1077 -1551
rect 59 -2897 459 -2697
rect 677 -2897 1077 -2697
rect 1659 -2351 2059 -1551
rect 2277 -2351 2677 -1551
rect 1659 -2897 2059 -2697
rect 2277 -2897 2677 -2697
rect 3259 -2351 3659 -1551
rect 3877 -2351 4277 -1551
rect 3259 -2897 3659 -2697
rect 3877 -2897 4277 -2697
rect 4859 -2351 5259 -1551
rect 5477 -2351 5877 -1551
rect 4859 -2897 5259 -2697
rect 5477 -2897 5877 -2697
rect 6459 -2351 6859 -1551
rect 7077 -2351 7477 -1551
rect 6459 -2897 6859 -2697
rect 7077 -2897 7477 -2697
rect 8059 -2351 8459 -1551
rect 8677 -2351 9077 -1551
rect 8059 -2897 8459 -2697
rect 8677 -2897 9077 -2697
rect 9659 -2351 10059 -1551
rect 10277 -2351 10677 -1551
rect 9659 -2897 10059 -2697
rect 10277 -2897 10677 -2697
rect 11259 -2351 11659 -1551
rect 11877 -2351 12277 -1551
rect 11259 -2897 11659 -2697
rect 11877 -2897 12277 -2697
rect 12859 -2351 13259 -1551
rect 13477 -2351 13877 -1551
rect 12859 -2897 13259 -2697
rect 13477 -2897 13877 -2697
rect 14459 -2351 14859 -1551
rect 15077 -2351 15477 -1551
rect 14459 -2897 14859 -2697
rect 15077 -2897 15477 -2697
rect 16059 -2351 16459 -1551
rect 16677 -2351 17077 -1551
rect 16059 -2897 16459 -2697
rect 16677 -2897 17077 -2697
rect 17659 -2351 18059 -1551
rect 18277 -2351 18677 -1551
rect 17659 -2897 18059 -2697
rect 18277 -2897 18677 -2697
rect 19259 -2351 19659 -1551
rect 19877 -2351 20277 -1551
rect 19259 -2897 19659 -2697
rect 19877 -2897 20277 -2697
rect 20859 -2351 21259 -1551
rect 21477 -2351 21877 -1551
rect 20859 -2897 21259 -2697
rect 21477 -2897 21877 -2697
rect 22459 -2351 22859 -1551
rect 23077 -2351 23477 -1551
rect 22459 -2897 22859 -2697
rect 23077 -2897 23477 -2697
rect 24059 -2351 24459 -1551
rect 24677 -2351 25077 -1551
rect 24059 -2897 24459 -2697
rect 24677 -2897 25077 -2697
rect 25659 -2351 26059 -1551
rect 26277 -2351 26677 -1551
rect 25659 -2897 26059 -2697
rect 26277 -2897 26677 -2697
rect 27259 -2351 27659 -1551
rect 27877 -2351 28277 -1551
rect 27259 -2897 27659 -2697
rect 27877 -2897 28277 -2697
rect 28859 -2351 29259 -1551
rect 29477 -2351 29877 -1551
rect 28859 -2897 29259 -2697
rect 29477 -2897 29877 -2697
rect 30459 -2351 30859 -1551
rect 31077 -2351 31477 -1551
rect 30459 -2897 30859 -2697
rect 31077 -2897 31477 -2697
rect 32059 -2351 32459 -1551
rect 32677 -2351 33077 -1551
rect 32059 -2897 32459 -2697
rect 32677 -2897 33077 -2697
rect 33659 -2351 34059 -1551
rect 34277 -2351 34677 -1551
rect 33659 -2897 34059 -2697
rect 34277 -2897 34677 -2697
rect 35259 -2351 35659 -1551
rect 35877 -2351 36277 -1551
rect 35259 -2897 35659 -2697
rect 35877 -2897 36277 -2697
rect 36859 -2351 37259 -1551
rect 37477 -2351 37877 -1551
rect 36859 -2897 37259 -2697
rect 37477 -2897 37877 -2697
rect 59 -4151 459 -3351
rect 677 -4151 1077 -3351
rect 59 -4697 459 -4497
rect 677 -4697 1077 -4497
rect 1659 -4151 2059 -3351
rect 2277 -4151 2677 -3351
rect 1659 -4697 2059 -4497
rect 2277 -4697 2677 -4497
rect 3259 -4151 3659 -3351
rect 3877 -4151 4277 -3351
rect 3259 -4697 3659 -4497
rect 3877 -4697 4277 -4497
rect 4859 -4151 5259 -3351
rect 5477 -4151 5877 -3351
rect 4859 -4697 5259 -4497
rect 5477 -4697 5877 -4497
rect 6459 -4151 6859 -3351
rect 7077 -4151 7477 -3351
rect 6459 -4697 6859 -4497
rect 7077 -4697 7477 -4497
rect 8059 -4151 8459 -3351
rect 8677 -4151 9077 -3351
rect 8059 -4697 8459 -4497
rect 8677 -4697 9077 -4497
rect 9659 -4151 10059 -3351
rect 10277 -4151 10677 -3351
rect 9659 -4697 10059 -4497
rect 10277 -4697 10677 -4497
rect 11259 -4151 11659 -3351
rect 11877 -4151 12277 -3351
rect 11259 -4697 11659 -4497
rect 11877 -4697 12277 -4497
rect 12859 -4151 13259 -3351
rect 13477 -4151 13877 -3351
rect 12859 -4697 13259 -4497
rect 13477 -4697 13877 -4497
rect 14459 -4151 14859 -3351
rect 15077 -4151 15477 -3351
rect 14459 -4697 14859 -4497
rect 15077 -4697 15477 -4497
rect 16059 -4151 16459 -3351
rect 16677 -4151 17077 -3351
rect 16059 -4697 16459 -4497
rect 16677 -4697 17077 -4497
rect 17659 -4151 18059 -3351
rect 18277 -4151 18677 -3351
rect 17659 -4697 18059 -4497
rect 18277 -4697 18677 -4497
rect 19259 -4151 19659 -3351
rect 19877 -4151 20277 -3351
rect 19259 -4697 19659 -4497
rect 19877 -4697 20277 -4497
rect 20859 -4151 21259 -3351
rect 21477 -4151 21877 -3351
rect 20859 -4697 21259 -4497
rect 21477 -4697 21877 -4497
rect 22459 -4151 22859 -3351
rect 23077 -4151 23477 -3351
rect 22459 -4697 22859 -4497
rect 23077 -4697 23477 -4497
rect 24059 -4151 24459 -3351
rect 24677 -4151 25077 -3351
rect 24059 -4697 24459 -4497
rect 24677 -4697 25077 -4497
rect 25659 -4151 26059 -3351
rect 26277 -4151 26677 -3351
rect 25659 -4697 26059 -4497
rect 26277 -4697 26677 -4497
rect 27259 -4151 27659 -3351
rect 27877 -4151 28277 -3351
rect 27259 -4697 27659 -4497
rect 27877 -4697 28277 -4497
rect 28859 -4151 29259 -3351
rect 29477 -4151 29877 -3351
rect 28859 -4697 29259 -4497
rect 29477 -4697 29877 -4497
rect 30459 -4151 30859 -3351
rect 31077 -4151 31477 -3351
rect 30459 -4697 30859 -4497
rect 31077 -4697 31477 -4497
rect 32059 -4151 32459 -3351
rect 32677 -4151 33077 -3351
rect 32059 -4697 32459 -4497
rect 32677 -4697 33077 -4497
rect 33659 -4151 34059 -3351
rect 34277 -4151 34677 -3351
rect 33659 -4697 34059 -4497
rect 34277 -4697 34677 -4497
rect 35259 -4151 35659 -3351
rect 35877 -4151 36277 -3351
rect 35259 -4697 35659 -4497
rect 35877 -4697 36277 -4497
rect 36859 -4151 37259 -3351
rect 37477 -4151 37877 -3351
rect 36859 -4697 37259 -4497
rect 37477 -4697 37877 -4497
rect 27968 -25112 28768 -24712
rect 27936 -25688 28736 -25588
rect 27936 -25846 28736 -25746
rect 27936 -26004 28736 -25904
rect 27936 -26162 28736 -26062
rect 27936 -26728 28736 -26628
rect 27936 -26886 28736 -26786
rect 27936 -27044 28736 -26944
rect 27936 -27202 28736 -27102
rect 27936 -27768 28736 -27668
rect 27936 -27926 28736 -27826
rect 27936 -28084 28736 -27984
rect 27936 -28242 28736 -28142
rect 27936 -28808 28736 -28708
rect 27936 -28966 28736 -28866
rect 27936 -29124 28736 -29024
rect 27936 -29282 28736 -29182
rect 27936 -29848 28736 -29748
rect 27936 -30006 28736 -29906
rect 27936 -30164 28736 -30064
rect 27936 -30322 28736 -30222
rect 31859 -29741 31959 -29541
rect 32299 -29741 32399 -29541
rect 32739 -29741 32839 -29541
rect 33178 -29741 33278 -29541
rect 33336 -29741 33436 -29541
rect 33494 -29741 33594 -29541
rect 34059 -29741 34159 -29541
rect 34499 -29741 34599 -29541
rect 34939 -29741 35039 -29541
rect 35378 -29741 35478 -29541
rect 35536 -29741 35636 -29541
rect 35694 -29741 35794 -29541
rect 36259 -29741 36359 -29541
rect 36699 -29741 36799 -29541
rect 37139 -29741 37239 -29541
rect 37578 -29741 37678 -29541
rect 37736 -29741 37836 -29541
rect 37894 -29741 37994 -29541
rect 27936 -30888 28736 -30788
rect 27936 -31046 28736 -30946
rect 27936 -31204 28736 -31104
rect 27936 -31362 28736 -31262
rect 31828 -30483 31928 -30283
rect 31986 -30483 32086 -30283
rect 32144 -30483 32244 -30283
rect 32583 -30483 32683 -30283
rect 33023 -30483 33123 -30283
rect 33463 -30483 33563 -30283
rect 34028 -30483 34128 -30283
rect 34186 -30483 34286 -30283
rect 34344 -30483 34444 -30283
rect 34783 -30483 34883 -30283
rect 35223 -30483 35323 -30283
rect 35663 -30483 35763 -30283
rect 36228 -30483 36328 -30283
rect 36386 -30483 36486 -30283
rect 36544 -30483 36644 -30283
rect 36983 -30483 37083 -30283
rect 37423 -30483 37523 -30283
rect 37863 -30483 37963 -30283
<< mvpmos >>
rect 27926 11312 28726 11412
rect 27926 11154 28726 11254
rect 27926 10996 28726 11096
rect 27926 10838 28726 10938
rect 30190 10807 30590 10907
rect 27926 10272 28726 10372
rect 27926 10114 28726 10214
rect 27926 9956 28726 10056
rect 27926 9798 28726 9898
rect 30904 10507 31004 10907
rect 31344 10507 31444 10907
rect 31784 10507 31884 10907
rect 32390 10807 32790 10907
rect 33104 10507 33204 10907
rect 33544 10507 33644 10907
rect 33984 10507 34084 10907
rect 34590 10807 34990 10907
rect 35304 10507 35404 10907
rect 35744 10507 35844 10907
rect 36184 10507 36284 10907
rect 27926 9232 28726 9332
rect 27926 9074 28726 9174
rect 27926 8916 28726 9016
rect 27926 8758 28726 8858
rect 29778 9197 30578 9597
rect 30636 9197 31436 9597
rect 27926 8192 28726 8292
rect 27926 8034 28726 8134
rect 27926 7876 28726 7976
rect 27926 7718 28726 7818
rect 27926 7152 28726 7252
rect 27926 6994 28726 7094
rect 27926 6836 28726 6936
rect 27926 6678 28726 6778
rect 29778 8193 30578 8593
rect 30636 8193 31436 8593
rect 29778 7557 30578 7957
rect 30636 7557 31436 7957
rect 29757 6818 30557 7018
rect 31097 6818 31897 7018
rect 27926 6112 28726 6212
rect 27926 5954 28726 6054
rect 27926 5796 28726 5896
rect 27926 5638 28726 5738
rect 27958 4357 28758 5157
rect 57 -8416 457 -8216
rect 693 -8416 1093 -8216
rect 57 -9542 457 -8742
rect 693 -9542 1093 -8742
rect 1657 -8416 2057 -8216
rect 2293 -8416 2693 -8216
rect 1657 -9542 2057 -8742
rect 2293 -9542 2693 -8742
rect 3257 -8416 3657 -8216
rect 3893 -8416 4293 -8216
rect 3257 -9542 3657 -8742
rect 3893 -9542 4293 -8742
rect 4857 -8416 5257 -8216
rect 5493 -8416 5893 -8216
rect 4857 -9542 5257 -8742
rect 5493 -9542 5893 -8742
rect 6457 -8416 6857 -8216
rect 7093 -8416 7493 -8216
rect 6457 -9542 6857 -8742
rect 7093 -9542 7493 -8742
rect 8057 -8416 8457 -8216
rect 8693 -8416 9093 -8216
rect 8057 -9542 8457 -8742
rect 8693 -9542 9093 -8742
rect 9657 -8416 10057 -8216
rect 10293 -8416 10693 -8216
rect 9657 -9542 10057 -8742
rect 10293 -9542 10693 -8742
rect 11257 -8416 11657 -8216
rect 11893 -8416 12293 -8216
rect 11257 -9542 11657 -8742
rect 11893 -9542 12293 -8742
rect 12857 -8416 13257 -8216
rect 13493 -8416 13893 -8216
rect 12857 -9542 13257 -8742
rect 13493 -9542 13893 -8742
rect 14457 -8416 14857 -8216
rect 15093 -8416 15493 -8216
rect 14457 -9542 14857 -8742
rect 15093 -9542 15493 -8742
rect 16057 -8416 16457 -8216
rect 16693 -8416 17093 -8216
rect 16057 -9542 16457 -8742
rect 16693 -9542 17093 -8742
rect 17657 -8416 18057 -8216
rect 18293 -8416 18693 -8216
rect 17657 -9542 18057 -8742
rect 18293 -9542 18693 -8742
rect 19257 -8416 19657 -8216
rect 19893 -8416 20293 -8216
rect 19257 -9542 19657 -8742
rect 19893 -9542 20293 -8742
rect 20857 -8416 21257 -8216
rect 21493 -8416 21893 -8216
rect 20857 -9542 21257 -8742
rect 21493 -9542 21893 -8742
rect 22457 -8416 22857 -8216
rect 23093 -8416 23493 -8216
rect 22457 -9542 22857 -8742
rect 23093 -9542 23493 -8742
rect 24057 -8416 24457 -8216
rect 24693 -8416 25093 -8216
rect 24057 -9542 24457 -8742
rect 24693 -9542 25093 -8742
rect 25657 -8416 26057 -8216
rect 26293 -8416 26693 -8216
rect 25657 -9542 26057 -8742
rect 26293 -9542 26693 -8742
rect 27257 -8416 27657 -8216
rect 27893 -8416 28293 -8216
rect 27257 -9542 27657 -8742
rect 27893 -9542 28293 -8742
rect 28857 -8416 29257 -8216
rect 29493 -8416 29893 -8216
rect 28857 -9542 29257 -8742
rect 29493 -9542 29893 -8742
rect 30457 -8416 30857 -8216
rect 31093 -8416 31493 -8216
rect 30457 -9542 30857 -8742
rect 31093 -9542 31493 -8742
rect 32057 -8416 32457 -8216
rect 32693 -8416 33093 -8216
rect 32057 -9542 32457 -8742
rect 32693 -9542 33093 -8742
rect 33657 -8416 34057 -8216
rect 34293 -8416 34693 -8216
rect 33657 -9542 34057 -8742
rect 34293 -9542 34693 -8742
rect 35257 -8416 35657 -8216
rect 35893 -8416 36293 -8216
rect 35257 -9542 35657 -8742
rect 35893 -9542 36293 -8742
rect 36857 -8416 37257 -8216
rect 37493 -8416 37893 -8216
rect 36857 -9542 37257 -8742
rect 37493 -9542 37893 -8742
rect 57 -10216 457 -10016
rect 693 -10216 1093 -10016
rect 57 -11342 457 -10542
rect 693 -11342 1093 -10542
rect 1657 -10216 2057 -10016
rect 2293 -10216 2693 -10016
rect 1657 -11342 2057 -10542
rect 2293 -11342 2693 -10542
rect 3257 -10216 3657 -10016
rect 3893 -10216 4293 -10016
rect 3257 -11342 3657 -10542
rect 3893 -11342 4293 -10542
rect 4857 -10216 5257 -10016
rect 5493 -10216 5893 -10016
rect 4857 -11342 5257 -10542
rect 5493 -11342 5893 -10542
rect 6457 -10216 6857 -10016
rect 7093 -10216 7493 -10016
rect 6457 -11342 6857 -10542
rect 7093 -11342 7493 -10542
rect 8057 -10216 8457 -10016
rect 8693 -10216 9093 -10016
rect 8057 -11342 8457 -10542
rect 8693 -11342 9093 -10542
rect 9657 -10216 10057 -10016
rect 10293 -10216 10693 -10016
rect 9657 -11342 10057 -10542
rect 10293 -11342 10693 -10542
rect 11257 -10216 11657 -10016
rect 11893 -10216 12293 -10016
rect 11257 -11342 11657 -10542
rect 11893 -11342 12293 -10542
rect 12857 -10216 13257 -10016
rect 13493 -10216 13893 -10016
rect 12857 -11342 13257 -10542
rect 13493 -11342 13893 -10542
rect 14457 -10216 14857 -10016
rect 15093 -10216 15493 -10016
rect 14457 -11342 14857 -10542
rect 15093 -11342 15493 -10542
rect 16057 -10216 16457 -10016
rect 16693 -10216 17093 -10016
rect 16057 -11342 16457 -10542
rect 16693 -11342 17093 -10542
rect 17657 -10216 18057 -10016
rect 18293 -10216 18693 -10016
rect 17657 -11342 18057 -10542
rect 18293 -11342 18693 -10542
rect 19257 -10216 19657 -10016
rect 19893 -10216 20293 -10016
rect 19257 -11342 19657 -10542
rect 19893 -11342 20293 -10542
rect 20857 -10216 21257 -10016
rect 21493 -10216 21893 -10016
rect 20857 -11342 21257 -10542
rect 21493 -11342 21893 -10542
rect 22457 -10216 22857 -10016
rect 23093 -10216 23493 -10016
rect 22457 -11342 22857 -10542
rect 23093 -11342 23493 -10542
rect 24057 -10216 24457 -10016
rect 24693 -10216 25093 -10016
rect 24057 -11342 24457 -10542
rect 24693 -11342 25093 -10542
rect 25657 -10216 26057 -10016
rect 26293 -10216 26693 -10016
rect 25657 -11342 26057 -10542
rect 26293 -11342 26693 -10542
rect 27257 -10216 27657 -10016
rect 27893 -10216 28293 -10016
rect 27257 -11342 27657 -10542
rect 27893 -11342 28293 -10542
rect 28857 -10216 29257 -10016
rect 29493 -10216 29893 -10016
rect 28857 -11342 29257 -10542
rect 29493 -11342 29893 -10542
rect 30457 -10216 30857 -10016
rect 31093 -10216 31493 -10016
rect 30457 -11342 30857 -10542
rect 31093 -11342 31493 -10542
rect 32057 -10216 32457 -10016
rect 32693 -10216 33093 -10016
rect 32057 -11342 32457 -10542
rect 32693 -11342 33093 -10542
rect 33657 -10216 34057 -10016
rect 34293 -10216 34693 -10016
rect 33657 -11342 34057 -10542
rect 34293 -11342 34693 -10542
rect 35257 -10216 35657 -10016
rect 35893 -10216 36293 -10016
rect 35257 -11342 35657 -10542
rect 35893 -11342 36293 -10542
rect 36857 -10216 37257 -10016
rect 37493 -10216 37893 -10016
rect 36857 -11342 37257 -10542
rect 37493 -11342 37893 -10542
rect 57 -12016 457 -11816
rect 693 -12016 1093 -11816
rect 57 -13142 457 -12342
rect 693 -13142 1093 -12342
rect 1657 -12016 2057 -11816
rect 2293 -12016 2693 -11816
rect 1657 -13142 2057 -12342
rect 2293 -13142 2693 -12342
rect 3257 -12016 3657 -11816
rect 3893 -12016 4293 -11816
rect 3257 -13142 3657 -12342
rect 3893 -13142 4293 -12342
rect 4857 -12016 5257 -11816
rect 5493 -12016 5893 -11816
rect 4857 -13142 5257 -12342
rect 5493 -13142 5893 -12342
rect 6457 -12016 6857 -11816
rect 7093 -12016 7493 -11816
rect 6457 -13142 6857 -12342
rect 7093 -13142 7493 -12342
rect 8057 -12016 8457 -11816
rect 8693 -12016 9093 -11816
rect 8057 -13142 8457 -12342
rect 8693 -13142 9093 -12342
rect 9657 -12016 10057 -11816
rect 10293 -12016 10693 -11816
rect 9657 -13142 10057 -12342
rect 10293 -13142 10693 -12342
rect 11257 -12016 11657 -11816
rect 11893 -12016 12293 -11816
rect 11257 -13142 11657 -12342
rect 11893 -13142 12293 -12342
rect 12857 -12016 13257 -11816
rect 13493 -12016 13893 -11816
rect 12857 -13142 13257 -12342
rect 13493 -13142 13893 -12342
rect 14457 -12016 14857 -11816
rect 15093 -12016 15493 -11816
rect 14457 -13142 14857 -12342
rect 15093 -13142 15493 -12342
rect 16057 -12016 16457 -11816
rect 16693 -12016 17093 -11816
rect 16057 -13142 16457 -12342
rect 16693 -13142 17093 -12342
rect 17657 -12016 18057 -11816
rect 18293 -12016 18693 -11816
rect 17657 -13142 18057 -12342
rect 18293 -13142 18693 -12342
rect 19257 -12016 19657 -11816
rect 19893 -12016 20293 -11816
rect 19257 -13142 19657 -12342
rect 19893 -13142 20293 -12342
rect 20857 -12016 21257 -11816
rect 21493 -12016 21893 -11816
rect 20857 -13142 21257 -12342
rect 21493 -13142 21893 -12342
rect 22457 -12016 22857 -11816
rect 23093 -12016 23493 -11816
rect 22457 -13142 22857 -12342
rect 23093 -13142 23493 -12342
rect 24057 -12016 24457 -11816
rect 24693 -12016 25093 -11816
rect 24057 -13142 24457 -12342
rect 24693 -13142 25093 -12342
rect 25657 -12016 26057 -11816
rect 26293 -12016 26693 -11816
rect 25657 -13142 26057 -12342
rect 26293 -13142 26693 -12342
rect 27257 -12016 27657 -11816
rect 27893 -12016 28293 -11816
rect 27257 -13142 27657 -12342
rect 27893 -13142 28293 -12342
rect 28857 -12016 29257 -11816
rect 29493 -12016 29893 -11816
rect 28857 -13142 29257 -12342
rect 29493 -13142 29893 -12342
rect 30457 -12016 30857 -11816
rect 31093 -12016 31493 -11816
rect 30457 -13142 30857 -12342
rect 31093 -13142 31493 -12342
rect 32057 -12016 32457 -11816
rect 32693 -12016 33093 -11816
rect 32057 -13142 32457 -12342
rect 32693 -13142 33093 -12342
rect 33657 -12016 34057 -11816
rect 34293 -12016 34693 -11816
rect 33657 -13142 34057 -12342
rect 34293 -13142 34693 -12342
rect 35257 -12016 35657 -11816
rect 35893 -12016 36293 -11816
rect 35257 -13142 35657 -12342
rect 35893 -13142 36293 -12342
rect 36857 -12016 37257 -11816
rect 37493 -12016 37893 -11816
rect 36857 -13142 37257 -12342
rect 37493 -13142 37893 -12342
rect 57 -13816 457 -13616
rect 693 -13816 1093 -13616
rect 57 -14942 457 -14142
rect 693 -14942 1093 -14142
rect 1657 -13816 2057 -13616
rect 2293 -13816 2693 -13616
rect 1657 -14942 2057 -14142
rect 2293 -14942 2693 -14142
rect 3257 -13816 3657 -13616
rect 3893 -13816 4293 -13616
rect 3257 -14942 3657 -14142
rect 3893 -14942 4293 -14142
rect 4857 -13816 5257 -13616
rect 5493 -13816 5893 -13616
rect 4857 -14942 5257 -14142
rect 5493 -14942 5893 -14142
rect 6457 -13816 6857 -13616
rect 7093 -13816 7493 -13616
rect 6457 -14942 6857 -14142
rect 7093 -14942 7493 -14142
rect 8057 -13816 8457 -13616
rect 8693 -13816 9093 -13616
rect 8057 -14942 8457 -14142
rect 8693 -14942 9093 -14142
rect 9657 -13816 10057 -13616
rect 10293 -13816 10693 -13616
rect 9657 -14942 10057 -14142
rect 10293 -14942 10693 -14142
rect 11257 -13816 11657 -13616
rect 11893 -13816 12293 -13616
rect 11257 -14942 11657 -14142
rect 11893 -14942 12293 -14142
rect 12857 -13816 13257 -13616
rect 13493 -13816 13893 -13616
rect 12857 -14942 13257 -14142
rect 13493 -14942 13893 -14142
rect 14457 -13816 14857 -13616
rect 15093 -13816 15493 -13616
rect 14457 -14942 14857 -14142
rect 15093 -14942 15493 -14142
rect 16057 -13816 16457 -13616
rect 16693 -13816 17093 -13616
rect 16057 -14942 16457 -14142
rect 16693 -14942 17093 -14142
rect 17657 -13816 18057 -13616
rect 18293 -13816 18693 -13616
rect 17657 -14942 18057 -14142
rect 18293 -14942 18693 -14142
rect 19257 -13816 19657 -13616
rect 19893 -13816 20293 -13616
rect 19257 -14942 19657 -14142
rect 19893 -14942 20293 -14142
rect 20857 -13816 21257 -13616
rect 21493 -13816 21893 -13616
rect 20857 -14942 21257 -14142
rect 21493 -14942 21893 -14142
rect 22457 -13816 22857 -13616
rect 23093 -13816 23493 -13616
rect 22457 -14942 22857 -14142
rect 23093 -14942 23493 -14142
rect 24057 -13816 24457 -13616
rect 24693 -13816 25093 -13616
rect 24057 -14942 24457 -14142
rect 24693 -14942 25093 -14142
rect 25657 -13816 26057 -13616
rect 26293 -13816 26693 -13616
rect 25657 -14942 26057 -14142
rect 26293 -14942 26693 -14142
rect 27257 -13816 27657 -13616
rect 27893 -13816 28293 -13616
rect 27257 -14942 27657 -14142
rect 27893 -14942 28293 -14142
rect 28857 -13816 29257 -13616
rect 29493 -13816 29893 -13616
rect 28857 -14942 29257 -14142
rect 29493 -14942 29893 -14142
rect 30457 -13816 30857 -13616
rect 31093 -13816 31493 -13616
rect 30457 -14942 30857 -14142
rect 31093 -14942 31493 -14142
rect 32057 -13816 32457 -13616
rect 32693 -13816 33093 -13616
rect 32057 -14942 32457 -14142
rect 32693 -14942 33093 -14142
rect 33657 -13816 34057 -13616
rect 34293 -13816 34693 -13616
rect 33657 -14942 34057 -14142
rect 34293 -14942 34693 -14142
rect 35257 -13816 35657 -13616
rect 35893 -13816 36293 -13616
rect 35257 -14942 35657 -14142
rect 35893 -14942 36293 -14142
rect 36857 -13816 37257 -13616
rect 37493 -13816 37893 -13616
rect 36857 -14942 37257 -14142
rect 37493 -14942 37893 -14142
rect 57 -15616 457 -15416
rect 693 -15616 1093 -15416
rect 57 -16742 457 -15942
rect 693 -16742 1093 -15942
rect 1657 -15616 2057 -15416
rect 2293 -15616 2693 -15416
rect 1657 -16742 2057 -15942
rect 2293 -16742 2693 -15942
rect 3257 -15616 3657 -15416
rect 3893 -15616 4293 -15416
rect 3257 -16742 3657 -15942
rect 3893 -16742 4293 -15942
rect 4857 -15616 5257 -15416
rect 5493 -15616 5893 -15416
rect 4857 -16742 5257 -15942
rect 5493 -16742 5893 -15942
rect 6457 -15616 6857 -15416
rect 7093 -15616 7493 -15416
rect 6457 -16742 6857 -15942
rect 7093 -16742 7493 -15942
rect 8057 -15616 8457 -15416
rect 8693 -15616 9093 -15416
rect 8057 -16742 8457 -15942
rect 8693 -16742 9093 -15942
rect 9657 -15616 10057 -15416
rect 10293 -15616 10693 -15416
rect 9657 -16742 10057 -15942
rect 10293 -16742 10693 -15942
rect 11257 -15616 11657 -15416
rect 11893 -15616 12293 -15416
rect 11257 -16742 11657 -15942
rect 11893 -16742 12293 -15942
rect 12857 -15616 13257 -15416
rect 13493 -15616 13893 -15416
rect 12857 -16742 13257 -15942
rect 13493 -16742 13893 -15942
rect 14457 -15616 14857 -15416
rect 15093 -15616 15493 -15416
rect 14457 -16742 14857 -15942
rect 15093 -16742 15493 -15942
rect 16057 -15616 16457 -15416
rect 16693 -15616 17093 -15416
rect 16057 -16742 16457 -15942
rect 16693 -16742 17093 -15942
rect 17657 -15616 18057 -15416
rect 18293 -15616 18693 -15416
rect 17657 -16742 18057 -15942
rect 18293 -16742 18693 -15942
rect 19257 -15616 19657 -15416
rect 19893 -15616 20293 -15416
rect 19257 -16742 19657 -15942
rect 19893 -16742 20293 -15942
rect 20857 -15616 21257 -15416
rect 21493 -15616 21893 -15416
rect 20857 -16742 21257 -15942
rect 21493 -16742 21893 -15942
rect 22457 -15616 22857 -15416
rect 23093 -15616 23493 -15416
rect 22457 -16742 22857 -15942
rect 23093 -16742 23493 -15942
rect 24057 -15616 24457 -15416
rect 24693 -15616 25093 -15416
rect 24057 -16742 24457 -15942
rect 24693 -16742 25093 -15942
rect 25657 -15616 26057 -15416
rect 26293 -15616 26693 -15416
rect 25657 -16742 26057 -15942
rect 26293 -16742 26693 -15942
rect 27257 -15616 27657 -15416
rect 27893 -15616 28293 -15416
rect 27257 -16742 27657 -15942
rect 27893 -16742 28293 -15942
rect 28857 -15616 29257 -15416
rect 29493 -15616 29893 -15416
rect 28857 -16742 29257 -15942
rect 29493 -16742 29893 -15942
rect 30457 -15616 30857 -15416
rect 31093 -15616 31493 -15416
rect 30457 -16742 30857 -15942
rect 31093 -16742 31493 -15942
rect 32057 -15616 32457 -15416
rect 32693 -15616 33093 -15416
rect 32057 -16742 32457 -15942
rect 32693 -16742 33093 -15942
rect 33657 -15616 34057 -15416
rect 34293 -15616 34693 -15416
rect 33657 -16742 34057 -15942
rect 34293 -16742 34693 -15942
rect 35257 -15616 35657 -15416
rect 35893 -15616 36293 -15416
rect 35257 -16742 35657 -15942
rect 35893 -16742 36293 -15942
rect 36857 -15616 37257 -15416
rect 37493 -15616 37893 -15416
rect 36857 -16742 37257 -15942
rect 37493 -16742 37893 -15942
rect 57 -17416 457 -17216
rect 693 -17416 1093 -17216
rect 57 -18542 457 -17742
rect 693 -18542 1093 -17742
rect 1657 -17416 2057 -17216
rect 2293 -17416 2693 -17216
rect 1657 -18542 2057 -17742
rect 2293 -18542 2693 -17742
rect 3257 -17416 3657 -17216
rect 3893 -17416 4293 -17216
rect 3257 -18542 3657 -17742
rect 3893 -18542 4293 -17742
rect 4857 -17416 5257 -17216
rect 5493 -17416 5893 -17216
rect 4857 -18542 5257 -17742
rect 5493 -18542 5893 -17742
rect 6457 -17416 6857 -17216
rect 7093 -17416 7493 -17216
rect 6457 -18542 6857 -17742
rect 7093 -18542 7493 -17742
rect 8057 -17416 8457 -17216
rect 8693 -17416 9093 -17216
rect 8057 -18542 8457 -17742
rect 8693 -18542 9093 -17742
rect 9657 -17416 10057 -17216
rect 10293 -17416 10693 -17216
rect 9657 -18542 10057 -17742
rect 10293 -18542 10693 -17742
rect 11257 -17416 11657 -17216
rect 11893 -17416 12293 -17216
rect 11257 -18542 11657 -17742
rect 11893 -18542 12293 -17742
rect 12857 -17416 13257 -17216
rect 13493 -17416 13893 -17216
rect 12857 -18542 13257 -17742
rect 13493 -18542 13893 -17742
rect 14457 -17416 14857 -17216
rect 15093 -17416 15493 -17216
rect 14457 -18542 14857 -17742
rect 15093 -18542 15493 -17742
rect 16057 -17416 16457 -17216
rect 16693 -17416 17093 -17216
rect 16057 -18542 16457 -17742
rect 16693 -18542 17093 -17742
rect 17657 -17416 18057 -17216
rect 18293 -17416 18693 -17216
rect 17657 -18542 18057 -17742
rect 18293 -18542 18693 -17742
rect 19257 -17416 19657 -17216
rect 19893 -17416 20293 -17216
rect 19257 -18542 19657 -17742
rect 19893 -18542 20293 -17742
rect 20857 -17416 21257 -17216
rect 21493 -17416 21893 -17216
rect 20857 -18542 21257 -17742
rect 21493 -18542 21893 -17742
rect 22457 -17416 22857 -17216
rect 23093 -17416 23493 -17216
rect 22457 -18542 22857 -17742
rect 23093 -18542 23493 -17742
rect 24057 -17416 24457 -17216
rect 24693 -17416 25093 -17216
rect 24057 -18542 24457 -17742
rect 24693 -18542 25093 -17742
rect 25657 -17416 26057 -17216
rect 26293 -17416 26693 -17216
rect 25657 -18542 26057 -17742
rect 26293 -18542 26693 -17742
rect 27257 -17416 27657 -17216
rect 27893 -17416 28293 -17216
rect 27257 -18542 27657 -17742
rect 27893 -18542 28293 -17742
rect 28857 -17416 29257 -17216
rect 29493 -17416 29893 -17216
rect 28857 -18542 29257 -17742
rect 29493 -18542 29893 -17742
rect 30457 -17416 30857 -17216
rect 31093 -17416 31493 -17216
rect 30457 -18542 30857 -17742
rect 31093 -18542 31493 -17742
rect 32057 -17416 32457 -17216
rect 32693 -17416 33093 -17216
rect 32057 -18542 32457 -17742
rect 32693 -18542 33093 -17742
rect 33657 -17416 34057 -17216
rect 34293 -17416 34693 -17216
rect 33657 -18542 34057 -17742
rect 34293 -18542 34693 -17742
rect 35257 -17416 35657 -17216
rect 35893 -17416 36293 -17216
rect 35257 -18542 35657 -17742
rect 35893 -18542 36293 -17742
rect 36857 -17416 37257 -17216
rect 37493 -17416 37893 -17216
rect 36857 -18542 37257 -17742
rect 37493 -18542 37893 -17742
rect 57 -19216 457 -19016
rect 693 -19216 1093 -19016
rect 57 -20342 457 -19542
rect 693 -20342 1093 -19542
rect 1657 -19216 2057 -19016
rect 2293 -19216 2693 -19016
rect 1657 -20342 2057 -19542
rect 2293 -20342 2693 -19542
rect 3257 -19216 3657 -19016
rect 3893 -19216 4293 -19016
rect 3257 -20342 3657 -19542
rect 3893 -20342 4293 -19542
rect 4857 -19216 5257 -19016
rect 5493 -19216 5893 -19016
rect 4857 -20342 5257 -19542
rect 5493 -20342 5893 -19542
rect 6457 -19216 6857 -19016
rect 7093 -19216 7493 -19016
rect 6457 -20342 6857 -19542
rect 7093 -20342 7493 -19542
rect 8057 -19216 8457 -19016
rect 8693 -19216 9093 -19016
rect 8057 -20342 8457 -19542
rect 8693 -20342 9093 -19542
rect 9657 -19216 10057 -19016
rect 10293 -19216 10693 -19016
rect 9657 -20342 10057 -19542
rect 10293 -20342 10693 -19542
rect 11257 -19216 11657 -19016
rect 11893 -19216 12293 -19016
rect 11257 -20342 11657 -19542
rect 11893 -20342 12293 -19542
rect 12857 -19216 13257 -19016
rect 13493 -19216 13893 -19016
rect 12857 -20342 13257 -19542
rect 13493 -20342 13893 -19542
rect 14457 -19216 14857 -19016
rect 15093 -19216 15493 -19016
rect 14457 -20342 14857 -19542
rect 15093 -20342 15493 -19542
rect 16057 -19216 16457 -19016
rect 16693 -19216 17093 -19016
rect 16057 -20342 16457 -19542
rect 16693 -20342 17093 -19542
rect 17657 -19216 18057 -19016
rect 18293 -19216 18693 -19016
rect 17657 -20342 18057 -19542
rect 18293 -20342 18693 -19542
rect 19257 -19216 19657 -19016
rect 19893 -19216 20293 -19016
rect 19257 -20342 19657 -19542
rect 19893 -20342 20293 -19542
rect 20857 -19216 21257 -19016
rect 21493 -19216 21893 -19016
rect 20857 -20342 21257 -19542
rect 21493 -20342 21893 -19542
rect 22457 -19216 22857 -19016
rect 23093 -19216 23493 -19016
rect 22457 -20342 22857 -19542
rect 23093 -20342 23493 -19542
rect 24057 -19216 24457 -19016
rect 24693 -19216 25093 -19016
rect 24057 -20342 24457 -19542
rect 24693 -20342 25093 -19542
rect 25657 -19216 26057 -19016
rect 26293 -19216 26693 -19016
rect 25657 -20342 26057 -19542
rect 26293 -20342 26693 -19542
rect 27257 -19216 27657 -19016
rect 27893 -19216 28293 -19016
rect 27257 -20342 27657 -19542
rect 27893 -20342 28293 -19542
rect 28857 -19216 29257 -19016
rect 29493 -19216 29893 -19016
rect 28857 -20342 29257 -19542
rect 29493 -20342 29893 -19542
rect 30457 -19216 30857 -19016
rect 31093 -19216 31493 -19016
rect 30457 -20342 30857 -19542
rect 31093 -20342 31493 -19542
rect 32057 -19216 32457 -19016
rect 32693 -19216 33093 -19016
rect 32057 -20342 32457 -19542
rect 32693 -20342 33093 -19542
rect 33657 -19216 34057 -19016
rect 34293 -19216 34693 -19016
rect 33657 -20342 34057 -19542
rect 34293 -20342 34693 -19542
rect 35257 -19216 35657 -19016
rect 35893 -19216 36293 -19016
rect 35257 -20342 35657 -19542
rect 35893 -20342 36293 -19542
rect 36857 -19216 37257 -19016
rect 37493 -19216 37893 -19016
rect 36857 -20342 37257 -19542
rect 37493 -20342 37893 -19542
rect 57 -21016 457 -20816
rect 693 -21016 1093 -20816
rect 57 -22142 457 -21342
rect 693 -22142 1093 -21342
rect 1657 -21016 2057 -20816
rect 2293 -21016 2693 -20816
rect 1657 -22142 2057 -21342
rect 2293 -22142 2693 -21342
rect 3257 -21016 3657 -20816
rect 3893 -21016 4293 -20816
rect 3257 -22142 3657 -21342
rect 3893 -22142 4293 -21342
rect 4857 -21016 5257 -20816
rect 5493 -21016 5893 -20816
rect 4857 -22142 5257 -21342
rect 5493 -22142 5893 -21342
rect 6457 -21016 6857 -20816
rect 7093 -21016 7493 -20816
rect 6457 -22142 6857 -21342
rect 7093 -22142 7493 -21342
rect 8057 -21016 8457 -20816
rect 8693 -21016 9093 -20816
rect 8057 -22142 8457 -21342
rect 8693 -22142 9093 -21342
rect 9657 -21016 10057 -20816
rect 10293 -21016 10693 -20816
rect 9657 -22142 10057 -21342
rect 10293 -22142 10693 -21342
rect 11257 -21016 11657 -20816
rect 11893 -21016 12293 -20816
rect 11257 -22142 11657 -21342
rect 11893 -22142 12293 -21342
rect 12857 -21016 13257 -20816
rect 13493 -21016 13893 -20816
rect 12857 -22142 13257 -21342
rect 13493 -22142 13893 -21342
rect 14457 -21016 14857 -20816
rect 15093 -21016 15493 -20816
rect 14457 -22142 14857 -21342
rect 15093 -22142 15493 -21342
rect 16057 -21016 16457 -20816
rect 16693 -21016 17093 -20816
rect 16057 -22142 16457 -21342
rect 16693 -22142 17093 -21342
rect 17657 -21016 18057 -20816
rect 18293 -21016 18693 -20816
rect 17657 -22142 18057 -21342
rect 18293 -22142 18693 -21342
rect 19257 -21016 19657 -20816
rect 19893 -21016 20293 -20816
rect 19257 -22142 19657 -21342
rect 19893 -22142 20293 -21342
rect 20857 -21016 21257 -20816
rect 21493 -21016 21893 -20816
rect 20857 -22142 21257 -21342
rect 21493 -22142 21893 -21342
rect 22457 -21016 22857 -20816
rect 23093 -21016 23493 -20816
rect 22457 -22142 22857 -21342
rect 23093 -22142 23493 -21342
rect 24057 -21016 24457 -20816
rect 24693 -21016 25093 -20816
rect 24057 -22142 24457 -21342
rect 24693 -22142 25093 -21342
rect 25657 -21016 26057 -20816
rect 26293 -21016 26693 -20816
rect 25657 -22142 26057 -21342
rect 26293 -22142 26693 -21342
rect 27257 -21016 27657 -20816
rect 27893 -21016 28293 -20816
rect 27257 -22142 27657 -21342
rect 27893 -22142 28293 -21342
rect 28857 -21016 29257 -20816
rect 29493 -21016 29893 -20816
rect 28857 -22142 29257 -21342
rect 29493 -22142 29893 -21342
rect 30457 -21016 30857 -20816
rect 31093 -21016 31493 -20816
rect 30457 -22142 30857 -21342
rect 31093 -22142 31493 -21342
rect 32057 -21016 32457 -20816
rect 32693 -21016 33093 -20816
rect 32057 -22142 32457 -21342
rect 32693 -22142 33093 -21342
rect 33657 -21016 34057 -20816
rect 34293 -21016 34693 -20816
rect 33657 -22142 34057 -21342
rect 34293 -22142 34693 -21342
rect 35257 -21016 35657 -20816
rect 35893 -21016 36293 -20816
rect 35257 -22142 35657 -21342
rect 35893 -22142 36293 -21342
rect 36857 -21016 37257 -20816
rect 37493 -21016 37893 -20816
rect 36857 -22142 37257 -21342
rect 37493 -22142 37893 -21342
rect 28398 -23472 28498 -22672
rect 28556 -23472 28656 -22672
rect 28714 -23472 28814 -22672
rect 28872 -23472 28972 -22672
rect 32678 -23023 32778 -22623
rect 32836 -23023 32936 -22623
rect 32994 -23023 33094 -22623
rect 33152 -23023 33252 -22623
rect 34048 -23043 34148 -22643
rect 34206 -23043 34306 -22643
rect 267 -24652 1867 -24352
rect 2467 -24652 4067 -24352
rect 4667 -24652 6267 -24352
rect 6867 -24652 8467 -24352
rect 9067 -24652 10667 -24352
rect 11267 -24652 12867 -24352
rect 13467 -24652 15067 -24352
rect 15667 -24652 17267 -24352
rect 17867 -24652 19467 -24352
rect 20067 -24652 21667 -24352
rect 33216 -24165 33316 -23765
rect 33374 -24165 33474 -23765
rect 33532 -24165 33632 -23765
rect 33690 -24165 33790 -23765
rect 33848 -24165 33948 -23765
rect 34006 -24165 34106 -23765
rect 34588 -24163 34688 -23763
rect 34746 -24163 34846 -23763
rect 34904 -24163 35004 -23763
rect 35062 -24163 35162 -23763
rect 35220 -24163 35320 -23763
rect 35378 -24163 35478 -23763
rect 35536 -24163 35636 -23763
rect 35694 -24163 35794 -23763
rect 35852 -24163 35952 -23763
rect 36010 -24163 36110 -23763
rect 36168 -24163 36268 -23763
rect 36326 -24163 36426 -23763
rect 36484 -24163 36584 -23763
rect 36642 -24163 36742 -23763
rect 36800 -24163 36900 -23763
rect 36958 -24163 37058 -23763
rect 267 -25452 1867 -25152
rect 2467 -25452 4067 -25152
rect 4667 -25452 6267 -25152
rect 6867 -25452 8467 -25152
rect 9067 -25452 10667 -25152
rect 11267 -25452 12867 -25152
rect 13467 -25452 15067 -25152
rect 15667 -25452 17267 -25152
rect 17867 -25452 19467 -25152
rect 20067 -25452 21667 -25152
rect 267 -26252 1867 -25952
rect 2467 -26252 4067 -25952
rect 4667 -26252 6267 -25952
rect 6867 -26252 8467 -25952
rect 9067 -26252 10667 -25952
rect 11267 -26252 12867 -25952
rect 13467 -26252 15067 -25952
rect 15667 -26252 17267 -25952
rect 17867 -26252 19467 -25952
rect 20067 -26252 21667 -25952
rect 267 -27052 1867 -26752
rect 2467 -27052 4067 -26752
rect 4667 -27052 6267 -26752
rect 6867 -27052 8467 -26752
rect 9067 -27052 10667 -26752
rect 11267 -27052 12867 -26752
rect 13467 -27052 15067 -26752
rect 15667 -27052 17267 -26752
rect 17867 -27052 19467 -26752
rect 20067 -27052 21667 -26752
rect 267 -27852 1867 -27552
rect 2467 -27852 4067 -27552
rect 4667 -27852 6267 -27552
rect 6867 -27852 8467 -27552
rect 9067 -27852 10667 -27552
rect 11267 -27852 12867 -27552
rect 13467 -27852 15067 -27552
rect 15667 -27852 17267 -27552
rect 17867 -27852 19467 -27552
rect 20067 -27852 21667 -27552
rect 267 -28652 1867 -28352
rect 2467 -28652 4067 -28352
rect 4667 -28652 6267 -28352
rect 6867 -28652 8467 -28352
rect 9067 -28652 10667 -28352
rect 11267 -28652 12867 -28352
rect 13467 -28652 15067 -28352
rect 15667 -28652 17267 -28352
rect 17867 -28652 19467 -28352
rect 20067 -28652 21667 -28352
rect 267 -29452 1867 -29152
rect 2467 -29452 4067 -29152
rect 4667 -29452 6267 -29152
rect 6867 -29452 8467 -29152
rect 9067 -29452 10667 -29152
rect 11267 -29452 12867 -29152
rect 13467 -29452 15067 -29152
rect 15667 -29452 17267 -29152
rect 17867 -29452 19467 -29152
rect 20067 -29452 21667 -29152
rect 267 -30252 1867 -29952
rect 2467 -30252 4067 -29952
rect 4667 -30252 6267 -29952
rect 6867 -30252 8467 -29952
rect 9067 -30252 10667 -29952
rect 11267 -30252 12867 -29952
rect 13467 -30252 15067 -29952
rect 15667 -30252 17267 -29952
rect 17867 -30252 19467 -29952
rect 20067 -30252 21667 -29952
rect 267 -31052 1867 -30752
rect 2467 -31052 4067 -30752
rect 4667 -31052 6267 -30752
rect 6867 -31052 8467 -30752
rect 9067 -31052 10667 -30752
rect 11267 -31052 12867 -30752
rect 13467 -31052 15067 -30752
rect 15667 -31052 17267 -30752
rect 17867 -31052 19467 -30752
rect 20067 -31052 21667 -30752
rect 267 -31852 1867 -31552
rect 2467 -31852 4067 -31552
rect 4667 -31852 6267 -31552
rect 6867 -31852 8467 -31552
rect 9067 -31852 10667 -31552
rect 11267 -31852 12867 -31552
rect 13467 -31852 15067 -31552
rect 15667 -31852 17267 -31552
rect 17867 -31852 19467 -31552
rect 20067 -31852 21667 -31552
rect 34977 -25076 35777 -24876
rect 34977 -25334 35777 -25134
rect 34977 -25592 35777 -25392
rect 34977 -25850 35777 -25650
rect 34977 -26108 35777 -25908
rect 34977 -26366 35777 -26166
rect 34977 -26624 35777 -26424
rect 34977 -26882 35777 -26682
rect 36317 -25076 37117 -24876
rect 36317 -25334 37117 -25134
rect 36317 -25592 37117 -25392
rect 36317 -25850 37117 -25650
rect 36317 -26108 37117 -25908
rect 36317 -26366 37117 -26166
rect 36317 -26624 37117 -26424
rect 36317 -26882 37117 -26682
rect 31858 -28921 31958 -28521
rect 32298 -28921 32398 -28521
rect 32738 -28921 32838 -28521
rect 33152 -28921 33552 -28821
rect 34058 -28921 34158 -28521
rect 34498 -28921 34598 -28521
rect 34938 -28921 35038 -28521
rect 35352 -28921 35752 -28821
rect 36258 -28921 36358 -28521
rect 36698 -28921 36798 -28521
rect 37138 -28921 37238 -28521
rect 37552 -28921 37952 -28821
rect 31870 -31203 32270 -31103
rect 32584 -31503 32684 -31103
rect 33024 -31503 33124 -31103
rect 33464 -31503 33564 -31103
rect 34070 -31203 34470 -31103
rect 34784 -31503 34884 -31103
rect 35224 -31503 35324 -31103
rect 35664 -31503 35764 -31103
rect 36270 -31203 36670 -31103
rect 36984 -31503 37084 -31103
rect 37424 -31503 37524 -31103
rect 37864 -31503 37964 -31103
<< ndiff >>
rect 34578 7318 34636 7330
rect 34578 7142 34590 7318
rect 34624 7142 34636 7318
rect 34578 7130 34636 7142
rect 34666 7318 34724 7330
rect 34666 7142 34678 7318
rect 34712 7142 34724 7318
rect 34666 7130 34724 7142
rect 34998 7318 35056 7330
rect 34998 7142 35010 7318
rect 35044 7142 35056 7318
rect 34998 7130 35056 7142
rect 35086 7318 35144 7330
rect 35086 7142 35098 7318
rect 35132 7142 35144 7318
rect 35086 7130 35144 7142
rect 35418 7318 35476 7330
rect 35418 7142 35430 7318
rect 35464 7142 35476 7318
rect 35418 7130 35476 7142
rect 35506 7318 35564 7330
rect 35506 7142 35518 7318
rect 35552 7142 35564 7318
rect 35506 7130 35564 7142
<< pdiff >>
rect 32898 8847 32956 8859
rect 32898 8071 32910 8847
rect 32944 8071 32956 8847
rect 32898 8059 32956 8071
rect 33156 8847 33214 8859
rect 33156 8071 33168 8847
rect 33202 8071 33214 8847
rect 33156 8059 33214 8071
rect 33414 8847 33472 8859
rect 33414 8071 33426 8847
rect 33460 8071 33472 8847
rect 33414 8059 33472 8071
rect 33738 8847 33796 8859
rect 33738 8071 33750 8847
rect 33784 8071 33796 8847
rect 33738 8059 33796 8071
rect 33996 8847 34054 8859
rect 33996 8071 34008 8847
rect 34042 8071 34054 8847
rect 33996 8059 34054 8071
rect 34254 8847 34312 8859
rect 34254 8071 34266 8847
rect 34300 8071 34312 8847
rect 34254 8059 34312 8071
rect 34578 8627 34636 8639
rect 34578 8251 34590 8627
rect 34624 8251 34636 8627
rect 34578 8239 34636 8251
rect 34666 8627 34724 8639
rect 34666 8251 34678 8627
rect 34712 8251 34724 8627
rect 34666 8239 34724 8251
rect 34998 8627 35056 8639
rect 34998 8251 35010 8627
rect 35044 8251 35056 8627
rect 34998 8239 35056 8251
rect 35086 8627 35144 8639
rect 35086 8251 35098 8627
rect 35132 8251 35144 8627
rect 35086 8239 35144 8251
rect 35418 8627 35476 8639
rect 35418 8251 35430 8627
rect 35464 8251 35476 8627
rect 35418 8239 35476 8251
rect 35506 8627 35564 8639
rect 35506 8251 35518 8627
rect 35552 8251 35564 8627
rect 35506 8239 35564 8251
<< mvndiff >>
rect 259 11775 1859 11787
rect 259 11741 271 11775
rect 1847 11741 1859 11775
rect 259 11729 1859 11741
rect 259 11417 1859 11429
rect 259 11383 271 11417
rect 1847 11383 1859 11417
rect 259 11371 1859 11383
rect 2459 11775 4059 11787
rect 2459 11741 2471 11775
rect 4047 11741 4059 11775
rect 2459 11729 4059 11741
rect 2459 11417 4059 11429
rect 2459 11383 2471 11417
rect 4047 11383 4059 11417
rect 2459 11371 4059 11383
rect 4659 11775 6259 11787
rect 4659 11741 4671 11775
rect 6247 11741 6259 11775
rect 4659 11729 6259 11741
rect 4659 11417 6259 11429
rect 4659 11383 4671 11417
rect 6247 11383 6259 11417
rect 4659 11371 6259 11383
rect 6859 11775 8459 11787
rect 6859 11741 6871 11775
rect 8447 11741 8459 11775
rect 6859 11729 8459 11741
rect 6859 11417 8459 11429
rect 6859 11383 6871 11417
rect 8447 11383 8459 11417
rect 6859 11371 8459 11383
rect 9059 11775 10659 11787
rect 9059 11741 9071 11775
rect 10647 11741 10659 11775
rect 9059 11729 10659 11741
rect 9059 11417 10659 11429
rect 9059 11383 9071 11417
rect 10647 11383 10659 11417
rect 9059 11371 10659 11383
rect 11259 11775 12859 11787
rect 11259 11741 11271 11775
rect 12847 11741 12859 11775
rect 11259 11729 12859 11741
rect 11259 11417 12859 11429
rect 11259 11383 11271 11417
rect 12847 11383 12859 11417
rect 11259 11371 12859 11383
rect 13459 11775 15059 11787
rect 13459 11741 13471 11775
rect 15047 11741 15059 11775
rect 13459 11729 15059 11741
rect 13459 11417 15059 11429
rect 13459 11383 13471 11417
rect 15047 11383 15059 11417
rect 13459 11371 15059 11383
rect 15659 11775 17259 11787
rect 15659 11741 15671 11775
rect 17247 11741 17259 11775
rect 15659 11729 17259 11741
rect 15659 11417 17259 11429
rect 15659 11383 15671 11417
rect 17247 11383 17259 11417
rect 15659 11371 17259 11383
rect 17859 11775 19459 11787
rect 17859 11741 17871 11775
rect 19447 11741 19459 11775
rect 17859 11729 19459 11741
rect 17859 11417 19459 11429
rect 17859 11383 17871 11417
rect 19447 11383 19459 11417
rect 17859 11371 19459 11383
rect 20059 11775 21659 11787
rect 20059 11741 20071 11775
rect 21647 11741 21659 11775
rect 20059 11729 21659 11741
rect 20059 11417 21659 11429
rect 20059 11383 20071 11417
rect 21647 11383 21659 11417
rect 20059 11371 21659 11383
rect 259 10975 1859 10987
rect 259 10941 271 10975
rect 1847 10941 1859 10975
rect 259 10929 1859 10941
rect 259 10617 1859 10629
rect 259 10583 271 10617
rect 1847 10583 1859 10617
rect 259 10571 1859 10583
rect 2458 10974 4058 10986
rect 2458 10940 2470 10974
rect 4046 10940 4058 10974
rect 2458 10928 4058 10940
rect 2458 10616 4058 10628
rect 2458 10582 2470 10616
rect 4046 10582 4058 10616
rect 2458 10570 4058 10582
rect 4658 10974 6258 10986
rect 4658 10940 4670 10974
rect 6246 10940 6258 10974
rect 4658 10928 6258 10940
rect 4658 10616 6258 10628
rect 4658 10582 4670 10616
rect 6246 10582 6258 10616
rect 4658 10570 6258 10582
rect 6858 10974 8458 10986
rect 6858 10940 6870 10974
rect 8446 10940 8458 10974
rect 6858 10928 8458 10940
rect 6858 10616 8458 10628
rect 6858 10582 6870 10616
rect 8446 10582 8458 10616
rect 6858 10570 8458 10582
rect 9058 10974 10658 10986
rect 9058 10940 9070 10974
rect 10646 10940 10658 10974
rect 9058 10928 10658 10940
rect 9058 10616 10658 10628
rect 9058 10582 9070 10616
rect 10646 10582 10658 10616
rect 9058 10570 10658 10582
rect 11258 10974 12858 10986
rect 11258 10940 11270 10974
rect 12846 10940 12858 10974
rect 11258 10928 12858 10940
rect 11258 10616 12858 10628
rect 11258 10582 11270 10616
rect 12846 10582 12858 10616
rect 11258 10570 12858 10582
rect 13458 10974 15058 10986
rect 13458 10940 13470 10974
rect 15046 10940 15058 10974
rect 13458 10928 15058 10940
rect 13458 10616 15058 10628
rect 13458 10582 13470 10616
rect 15046 10582 15058 10616
rect 13458 10570 15058 10582
rect 15658 10974 17258 10986
rect 15658 10940 15670 10974
rect 17246 10940 17258 10974
rect 15658 10928 17258 10940
rect 15658 10616 17258 10628
rect 15658 10582 15670 10616
rect 17246 10582 17258 10616
rect 15658 10570 17258 10582
rect 17858 10974 19458 10986
rect 17858 10940 17870 10974
rect 19446 10940 19458 10974
rect 17858 10928 19458 10940
rect 17858 10616 19458 10628
rect 17858 10582 17870 10616
rect 19446 10582 19458 10616
rect 17858 10570 19458 10582
rect 20059 10975 21659 10987
rect 20059 10941 20071 10975
rect 21647 10941 21659 10975
rect 20059 10929 21659 10941
rect 20059 10617 21659 10629
rect 20059 10583 20071 10617
rect 21647 10583 21659 10617
rect 20059 10571 21659 10583
rect 259 10175 1859 10187
rect 259 10141 271 10175
rect 1847 10141 1859 10175
rect 259 10129 1859 10141
rect 259 9817 1859 9829
rect 259 9783 271 9817
rect 1847 9783 1859 9817
rect 259 9771 1859 9783
rect 2458 10174 4058 10186
rect 2458 10140 2470 10174
rect 4046 10140 4058 10174
rect 2458 10128 4058 10140
rect 2458 9816 4058 9828
rect 2458 9782 2470 9816
rect 4046 9782 4058 9816
rect 2458 9770 4058 9782
rect 4658 10174 6258 10186
rect 4658 10140 4670 10174
rect 6246 10140 6258 10174
rect 4658 10128 6258 10140
rect 4658 9816 6258 9828
rect 4658 9782 4670 9816
rect 6246 9782 6258 9816
rect 4658 9770 6258 9782
rect 6858 10174 8458 10186
rect 6858 10140 6870 10174
rect 8446 10140 8458 10174
rect 6858 10128 8458 10140
rect 6858 9816 8458 9828
rect 6858 9782 6870 9816
rect 8446 9782 8458 9816
rect 6858 9770 8458 9782
rect 9058 10174 10658 10186
rect 9058 10140 9070 10174
rect 10646 10140 10658 10174
rect 9058 10128 10658 10140
rect 9058 9816 10658 9828
rect 9058 9782 9070 9816
rect 10646 9782 10658 9816
rect 9058 9770 10658 9782
rect 11258 10174 12858 10186
rect 11258 10140 11270 10174
rect 12846 10140 12858 10174
rect 11258 10128 12858 10140
rect 11258 9816 12858 9828
rect 11258 9782 11270 9816
rect 12846 9782 12858 9816
rect 11258 9770 12858 9782
rect 13458 10174 15058 10186
rect 13458 10140 13470 10174
rect 15046 10140 15058 10174
rect 13458 10128 15058 10140
rect 13458 9816 15058 9828
rect 13458 9782 13470 9816
rect 15046 9782 15058 9816
rect 13458 9770 15058 9782
rect 15658 10174 17258 10186
rect 15658 10140 15670 10174
rect 17246 10140 17258 10174
rect 15658 10128 17258 10140
rect 15658 9816 17258 9828
rect 15658 9782 15670 9816
rect 17246 9782 17258 9816
rect 15658 9770 17258 9782
rect 17858 10174 19458 10186
rect 17858 10140 17870 10174
rect 19446 10140 19458 10174
rect 17858 10128 19458 10140
rect 17858 9816 19458 9828
rect 17858 9782 17870 9816
rect 19446 9782 19458 9816
rect 17858 9770 19458 9782
rect 20059 10175 21659 10187
rect 20059 10141 20071 10175
rect 21647 10141 21659 10175
rect 20059 10129 21659 10141
rect 20059 9817 21659 9829
rect 20059 9783 20071 9817
rect 21647 9783 21659 9817
rect 20059 9771 21659 9783
rect 259 9375 1859 9387
rect 259 9341 271 9375
rect 1847 9341 1859 9375
rect 259 9329 1859 9341
rect 259 9017 1859 9029
rect 259 8983 271 9017
rect 1847 8983 1859 9017
rect 259 8971 1859 8983
rect 2458 9374 4058 9386
rect 2458 9340 2470 9374
rect 4046 9340 4058 9374
rect 2458 9328 4058 9340
rect 2458 9016 4058 9028
rect 2458 8982 2470 9016
rect 4046 8982 4058 9016
rect 2458 8970 4058 8982
rect 4658 9374 6258 9386
rect 4658 9340 4670 9374
rect 6246 9340 6258 9374
rect 4658 9328 6258 9340
rect 4658 9016 6258 9028
rect 4658 8982 4670 9016
rect 6246 8982 6258 9016
rect 4658 8970 6258 8982
rect 6858 9374 8458 9386
rect 6858 9340 6870 9374
rect 8446 9340 8458 9374
rect 6858 9328 8458 9340
rect 6858 9016 8458 9028
rect 6858 8982 6870 9016
rect 8446 8982 8458 9016
rect 6858 8970 8458 8982
rect 9058 9374 10658 9386
rect 9058 9340 9070 9374
rect 10646 9340 10658 9374
rect 9058 9328 10658 9340
rect 9058 9016 10658 9028
rect 9058 8982 9070 9016
rect 10646 8982 10658 9016
rect 9058 8970 10658 8982
rect 11258 9374 12858 9386
rect 11258 9340 11270 9374
rect 12846 9340 12858 9374
rect 11258 9328 12858 9340
rect 11258 9016 12858 9028
rect 11258 8982 11270 9016
rect 12846 8982 12858 9016
rect 11258 8970 12858 8982
rect 13458 9374 15058 9386
rect 13458 9340 13470 9374
rect 15046 9340 15058 9374
rect 13458 9328 15058 9340
rect 13458 9016 15058 9028
rect 13458 8982 13470 9016
rect 15046 8982 15058 9016
rect 13458 8970 15058 8982
rect 15658 9374 17258 9386
rect 15658 9340 15670 9374
rect 17246 9340 17258 9374
rect 15658 9328 17258 9340
rect 15658 9016 17258 9028
rect 15658 8982 15670 9016
rect 17246 8982 17258 9016
rect 15658 8970 17258 8982
rect 17858 9374 19458 9386
rect 17858 9340 17870 9374
rect 19446 9340 19458 9374
rect 17858 9328 19458 9340
rect 17858 9016 19458 9028
rect 17858 8982 17870 9016
rect 19446 8982 19458 9016
rect 17858 8970 19458 8982
rect 20059 9375 21659 9387
rect 20059 9341 20071 9375
rect 21647 9341 21659 9375
rect 20059 9329 21659 9341
rect 20059 9017 21659 9029
rect 20059 8983 20071 9017
rect 21647 8983 21659 9017
rect 20059 8971 21659 8983
rect 259 8575 1859 8587
rect 259 8541 271 8575
rect 1847 8541 1859 8575
rect 259 8529 1859 8541
rect 259 8217 1859 8229
rect 259 8183 271 8217
rect 1847 8183 1859 8217
rect 259 8171 1859 8183
rect 2458 8574 4058 8586
rect 2458 8540 2470 8574
rect 4046 8540 4058 8574
rect 2458 8528 4058 8540
rect 2458 8216 4058 8228
rect 2458 8182 2470 8216
rect 4046 8182 4058 8216
rect 2458 8170 4058 8182
rect 4658 8574 6258 8586
rect 4658 8540 4670 8574
rect 6246 8540 6258 8574
rect 4658 8528 6258 8540
rect 4658 8216 6258 8228
rect 4658 8182 4670 8216
rect 6246 8182 6258 8216
rect 4658 8170 6258 8182
rect 6858 8574 8458 8586
rect 6858 8540 6870 8574
rect 8446 8540 8458 8574
rect 6858 8528 8458 8540
rect 6858 8216 8458 8228
rect 6858 8182 6870 8216
rect 8446 8182 8458 8216
rect 6858 8170 8458 8182
rect 9058 8574 10658 8586
rect 9058 8540 9070 8574
rect 10646 8540 10658 8574
rect 9058 8528 10658 8540
rect 9058 8216 10658 8228
rect 9058 8182 9070 8216
rect 10646 8182 10658 8216
rect 9058 8170 10658 8182
rect 11258 8574 12858 8586
rect 11258 8540 11270 8574
rect 12846 8540 12858 8574
rect 11258 8528 12858 8540
rect 11258 8216 12858 8228
rect 11258 8182 11270 8216
rect 12846 8182 12858 8216
rect 11258 8170 12858 8182
rect 13458 8574 15058 8586
rect 13458 8540 13470 8574
rect 15046 8540 15058 8574
rect 13458 8528 15058 8540
rect 13458 8216 15058 8228
rect 13458 8182 13470 8216
rect 15046 8182 15058 8216
rect 13458 8170 15058 8182
rect 15658 8574 17258 8586
rect 15658 8540 15670 8574
rect 17246 8540 17258 8574
rect 15658 8528 17258 8540
rect 15658 8216 17258 8228
rect 15658 8182 15670 8216
rect 17246 8182 17258 8216
rect 15658 8170 17258 8182
rect 17858 8574 19458 8586
rect 17858 8540 17870 8574
rect 19446 8540 19458 8574
rect 17858 8528 19458 8540
rect 17858 8216 19458 8228
rect 17858 8182 17870 8216
rect 19446 8182 19458 8216
rect 17858 8170 19458 8182
rect 20059 8575 21659 8587
rect 20059 8541 20071 8575
rect 21647 8541 21659 8575
rect 20059 8529 21659 8541
rect 20059 8217 21659 8229
rect 20059 8183 20071 8217
rect 21647 8183 21659 8217
rect 20059 8171 21659 8183
rect 259 7775 1859 7787
rect 259 7741 271 7775
rect 1847 7741 1859 7775
rect 259 7729 1859 7741
rect 259 7417 1859 7429
rect 259 7383 271 7417
rect 1847 7383 1859 7417
rect 259 7371 1859 7383
rect 2458 7774 4058 7786
rect 2458 7740 2470 7774
rect 4046 7740 4058 7774
rect 2458 7728 4058 7740
rect 2458 7416 4058 7428
rect 2458 7382 2470 7416
rect 4046 7382 4058 7416
rect 2458 7370 4058 7382
rect 4658 7774 6258 7786
rect 4658 7740 4670 7774
rect 6246 7740 6258 7774
rect 4658 7728 6258 7740
rect 4658 7416 6258 7428
rect 4658 7382 4670 7416
rect 6246 7382 6258 7416
rect 4658 7370 6258 7382
rect 6858 7774 8458 7786
rect 6858 7740 6870 7774
rect 8446 7740 8458 7774
rect 6858 7728 8458 7740
rect 6858 7416 8458 7428
rect 6858 7382 6870 7416
rect 8446 7382 8458 7416
rect 6858 7370 8458 7382
rect 9058 7774 10658 7786
rect 9058 7740 9070 7774
rect 10646 7740 10658 7774
rect 9058 7728 10658 7740
rect 9058 7416 10658 7428
rect 9058 7382 9070 7416
rect 10646 7382 10658 7416
rect 9058 7370 10658 7382
rect 11258 7774 12858 7786
rect 11258 7740 11270 7774
rect 12846 7740 12858 7774
rect 11258 7728 12858 7740
rect 11258 7416 12858 7428
rect 11258 7382 11270 7416
rect 12846 7382 12858 7416
rect 11258 7370 12858 7382
rect 13458 7774 15058 7786
rect 13458 7740 13470 7774
rect 15046 7740 15058 7774
rect 13458 7728 15058 7740
rect 13458 7416 15058 7428
rect 13458 7382 13470 7416
rect 15046 7382 15058 7416
rect 13458 7370 15058 7382
rect 15658 7774 17258 7786
rect 15658 7740 15670 7774
rect 17246 7740 17258 7774
rect 15658 7728 17258 7740
rect 15658 7416 17258 7428
rect 15658 7382 15670 7416
rect 17246 7382 17258 7416
rect 15658 7370 17258 7382
rect 17858 7774 19458 7786
rect 17858 7740 17870 7774
rect 19446 7740 19458 7774
rect 17858 7728 19458 7740
rect 17858 7416 19458 7428
rect 17858 7382 17870 7416
rect 19446 7382 19458 7416
rect 17858 7370 19458 7382
rect 20059 7775 21659 7787
rect 20059 7741 20071 7775
rect 21647 7741 21659 7775
rect 20059 7729 21659 7741
rect 20059 7417 21659 7429
rect 20059 7383 20071 7417
rect 21647 7383 21659 7417
rect 20059 7371 21659 7383
rect 259 6975 1859 6987
rect 259 6941 271 6975
rect 1847 6941 1859 6975
rect 259 6929 1859 6941
rect 259 6617 1859 6629
rect 259 6583 271 6617
rect 1847 6583 1859 6617
rect 259 6571 1859 6583
rect 2458 6974 4058 6986
rect 2458 6940 2470 6974
rect 4046 6940 4058 6974
rect 2458 6928 4058 6940
rect 2458 6616 4058 6628
rect 2458 6582 2470 6616
rect 4046 6582 4058 6616
rect 2458 6570 4058 6582
rect 4658 6974 6258 6986
rect 4658 6940 4670 6974
rect 6246 6940 6258 6974
rect 4658 6928 6258 6940
rect 4658 6616 6258 6628
rect 4658 6582 4670 6616
rect 6246 6582 6258 6616
rect 4658 6570 6258 6582
rect 6858 6974 8458 6986
rect 6858 6940 6870 6974
rect 8446 6940 8458 6974
rect 6858 6928 8458 6940
rect 6858 6616 8458 6628
rect 6858 6582 6870 6616
rect 8446 6582 8458 6616
rect 6858 6570 8458 6582
rect 9058 6974 10658 6986
rect 9058 6940 9070 6974
rect 10646 6940 10658 6974
rect 9058 6928 10658 6940
rect 9058 6616 10658 6628
rect 9058 6582 9070 6616
rect 10646 6582 10658 6616
rect 9058 6570 10658 6582
rect 11258 6974 12858 6986
rect 11258 6940 11270 6974
rect 12846 6940 12858 6974
rect 11258 6928 12858 6940
rect 11258 6616 12858 6628
rect 11258 6582 11270 6616
rect 12846 6582 12858 6616
rect 11258 6570 12858 6582
rect 13458 6974 15058 6986
rect 13458 6940 13470 6974
rect 15046 6940 15058 6974
rect 13458 6928 15058 6940
rect 13458 6616 15058 6628
rect 13458 6582 13470 6616
rect 15046 6582 15058 6616
rect 13458 6570 15058 6582
rect 15658 6974 17258 6986
rect 15658 6940 15670 6974
rect 17246 6940 17258 6974
rect 15658 6928 17258 6940
rect 15658 6616 17258 6628
rect 15658 6582 15670 6616
rect 17246 6582 17258 6616
rect 15658 6570 17258 6582
rect 17858 6974 19458 6986
rect 17858 6940 17870 6974
rect 19446 6940 19458 6974
rect 17858 6928 19458 6940
rect 17858 6616 19458 6628
rect 17858 6582 17870 6616
rect 19446 6582 19458 6616
rect 17858 6570 19458 6582
rect 20059 6975 21659 6987
rect 20059 6941 20071 6975
rect 21647 6941 21659 6975
rect 20059 6929 21659 6941
rect 20059 6617 21659 6629
rect 20059 6583 20071 6617
rect 21647 6583 21659 6617
rect 20059 6571 21659 6583
rect 259 6175 1859 6187
rect 259 6141 271 6175
rect 1847 6141 1859 6175
rect 259 6129 1859 6141
rect 259 5817 1859 5829
rect 259 5783 271 5817
rect 1847 5783 1859 5817
rect 259 5771 1859 5783
rect 2458 6174 4058 6186
rect 2458 6140 2470 6174
rect 4046 6140 4058 6174
rect 2458 6128 4058 6140
rect 2458 5816 4058 5828
rect 2458 5782 2470 5816
rect 4046 5782 4058 5816
rect 2458 5770 4058 5782
rect 4658 6174 6258 6186
rect 4658 6140 4670 6174
rect 6246 6140 6258 6174
rect 4658 6128 6258 6140
rect 4658 5816 6258 5828
rect 4658 5782 4670 5816
rect 6246 5782 6258 5816
rect 4658 5770 6258 5782
rect 6858 6174 8458 6186
rect 6858 6140 6870 6174
rect 8446 6140 8458 6174
rect 6858 6128 8458 6140
rect 6858 5816 8458 5828
rect 6858 5782 6870 5816
rect 8446 5782 8458 5816
rect 6858 5770 8458 5782
rect 9058 6174 10658 6186
rect 9058 6140 9070 6174
rect 10646 6140 10658 6174
rect 9058 6128 10658 6140
rect 9058 5816 10658 5828
rect 9058 5782 9070 5816
rect 10646 5782 10658 5816
rect 9058 5770 10658 5782
rect 11258 6174 12858 6186
rect 11258 6140 11270 6174
rect 12846 6140 12858 6174
rect 11258 6128 12858 6140
rect 11258 5816 12858 5828
rect 11258 5782 11270 5816
rect 12846 5782 12858 5816
rect 11258 5770 12858 5782
rect 13458 6174 15058 6186
rect 13458 6140 13470 6174
rect 15046 6140 15058 6174
rect 13458 6128 15058 6140
rect 13458 5816 15058 5828
rect 13458 5782 13470 5816
rect 15046 5782 15058 5816
rect 13458 5770 15058 5782
rect 15658 6174 17258 6186
rect 15658 6140 15670 6174
rect 17246 6140 17258 6174
rect 15658 6128 17258 6140
rect 15658 5816 17258 5828
rect 15658 5782 15670 5816
rect 17246 5782 17258 5816
rect 15658 5770 17258 5782
rect 17858 6174 19458 6186
rect 17858 6140 17870 6174
rect 19446 6140 19458 6174
rect 17858 6128 19458 6140
rect 17858 5816 19458 5828
rect 17858 5782 17870 5816
rect 19446 5782 19458 5816
rect 17858 5770 19458 5782
rect 20059 6175 21659 6187
rect 20059 6141 20071 6175
rect 21647 6141 21659 6175
rect 20059 6129 21659 6141
rect 20059 5817 21659 5829
rect 20059 5783 20071 5817
rect 21647 5783 21659 5817
rect 20059 5771 21659 5783
rect 259 5375 1859 5387
rect 259 5341 271 5375
rect 1847 5341 1859 5375
rect 259 5329 1859 5341
rect 259 5017 1859 5029
rect 259 4983 271 5017
rect 1847 4983 1859 5017
rect 259 4971 1859 4983
rect 2458 5374 4058 5386
rect 2458 5340 2470 5374
rect 4046 5340 4058 5374
rect 2458 5328 4058 5340
rect 2458 5016 4058 5028
rect 2458 4982 2470 5016
rect 4046 4982 4058 5016
rect 2458 4970 4058 4982
rect 4658 5374 6258 5386
rect 4658 5340 4670 5374
rect 6246 5340 6258 5374
rect 4658 5328 6258 5340
rect 4658 5016 6258 5028
rect 4658 4982 4670 5016
rect 6246 4982 6258 5016
rect 4658 4970 6258 4982
rect 6858 5374 8458 5386
rect 6858 5340 6870 5374
rect 8446 5340 8458 5374
rect 6858 5328 8458 5340
rect 6858 5016 8458 5028
rect 6858 4982 6870 5016
rect 8446 4982 8458 5016
rect 6858 4970 8458 4982
rect 9058 5374 10658 5386
rect 9058 5340 9070 5374
rect 10646 5340 10658 5374
rect 9058 5328 10658 5340
rect 9058 5016 10658 5028
rect 9058 4982 9070 5016
rect 10646 4982 10658 5016
rect 9058 4970 10658 4982
rect 11258 5374 12858 5386
rect 11258 5340 11270 5374
rect 12846 5340 12858 5374
rect 11258 5328 12858 5340
rect 11258 5016 12858 5028
rect 11258 4982 11270 5016
rect 12846 4982 12858 5016
rect 11258 4970 12858 4982
rect 13458 5374 15058 5386
rect 13458 5340 13470 5374
rect 15046 5340 15058 5374
rect 13458 5328 15058 5340
rect 13458 5016 15058 5028
rect 13458 4982 13470 5016
rect 15046 4982 15058 5016
rect 13458 4970 15058 4982
rect 15658 5374 17258 5386
rect 15658 5340 15670 5374
rect 17246 5340 17258 5374
rect 15658 5328 17258 5340
rect 15658 5016 17258 5028
rect 15658 4982 15670 5016
rect 17246 4982 17258 5016
rect 15658 4970 17258 4982
rect 17858 5374 19458 5386
rect 17858 5340 17870 5374
rect 19446 5340 19458 5374
rect 17858 5328 19458 5340
rect 17858 5016 19458 5028
rect 17858 4982 17870 5016
rect 19446 4982 19458 5016
rect 17858 4970 19458 4982
rect 20059 5375 21659 5387
rect 20059 5341 20071 5375
rect 21647 5341 21659 5375
rect 20059 5329 21659 5341
rect 20059 5017 21659 5029
rect 20059 4983 20071 5017
rect 21647 4983 21659 5017
rect 20059 4971 21659 4983
rect 259 4575 1859 4587
rect 259 4541 271 4575
rect 1847 4541 1859 4575
rect 259 4529 1859 4541
rect 259 4217 1859 4229
rect 259 4183 271 4217
rect 1847 4183 1859 4217
rect 259 4171 1859 4183
rect 2459 4575 4059 4587
rect 2459 4541 2471 4575
rect 4047 4541 4059 4575
rect 2459 4529 4059 4541
rect 2459 4217 4059 4229
rect 2459 4183 2471 4217
rect 4047 4183 4059 4217
rect 2459 4171 4059 4183
rect 4659 4575 6259 4587
rect 4659 4541 4671 4575
rect 6247 4541 6259 4575
rect 4659 4529 6259 4541
rect 4659 4217 6259 4229
rect 4659 4183 4671 4217
rect 6247 4183 6259 4217
rect 4659 4171 6259 4183
rect 6859 4575 8459 4587
rect 6859 4541 6871 4575
rect 8447 4541 8459 4575
rect 6859 4529 8459 4541
rect 6859 4217 8459 4229
rect 6859 4183 6871 4217
rect 8447 4183 8459 4217
rect 6859 4171 8459 4183
rect 9060 4576 10660 4588
rect 9060 4542 9072 4576
rect 10648 4542 10660 4576
rect 9060 4530 10660 4542
rect 9060 4218 10660 4230
rect 9060 4184 9072 4218
rect 10648 4184 10660 4218
rect 9060 4172 10660 4184
rect 11260 4576 12860 4588
rect 11260 4542 11272 4576
rect 12848 4542 12860 4576
rect 11260 4530 12860 4542
rect 11260 4218 12860 4230
rect 11260 4184 11272 4218
rect 12848 4184 12860 4218
rect 11260 4172 12860 4184
rect 13459 4575 15059 4587
rect 13459 4541 13471 4575
rect 15047 4541 15059 4575
rect 13459 4529 15059 4541
rect 13459 4217 15059 4229
rect 13459 4183 13471 4217
rect 15047 4183 15059 4217
rect 13459 4171 15059 4183
rect 15659 4575 17259 4587
rect 15659 4541 15671 4575
rect 17247 4541 17259 4575
rect 15659 4529 17259 4541
rect 15659 4217 17259 4229
rect 15659 4183 15671 4217
rect 17247 4183 17259 4217
rect 15659 4171 17259 4183
rect 17859 4575 19459 4587
rect 17859 4541 17871 4575
rect 19447 4541 19459 4575
rect 17859 4529 19459 4541
rect 17859 4217 19459 4229
rect 17859 4183 17871 4217
rect 19447 4183 19459 4217
rect 17859 4171 19459 4183
rect 20059 4575 21659 4587
rect 20059 4541 20071 4575
rect 21647 4541 21659 4575
rect 20059 4529 21659 4541
rect 20059 4217 21659 4229
rect 20059 4183 20071 4217
rect 21647 4183 21659 4217
rect 20059 4171 21659 4183
rect 30090 11715 30148 11727
rect 30090 11539 30102 11715
rect 30136 11539 30148 11715
rect 30090 11527 30148 11539
rect 30248 11715 30306 11727
rect 30248 11539 30260 11715
rect 30294 11539 30306 11715
rect 30248 11527 30306 11539
rect 30406 11715 30464 11727
rect 30406 11539 30418 11715
rect 30452 11539 30464 11715
rect 30406 11527 30464 11539
rect 30564 11715 30622 11727
rect 30564 11539 30576 11715
rect 30610 11539 30622 11715
rect 30564 11527 30622 11539
rect 30845 11715 30903 11727
rect 30845 11539 30857 11715
rect 30891 11539 30903 11715
rect 30845 11527 30903 11539
rect 31003 11715 31061 11727
rect 31003 11539 31015 11715
rect 31049 11539 31061 11715
rect 31003 11527 31061 11539
rect 31285 11715 31343 11727
rect 31285 11539 31297 11715
rect 31331 11539 31343 11715
rect 31285 11527 31343 11539
rect 31443 11715 31501 11727
rect 31443 11539 31455 11715
rect 31489 11539 31501 11715
rect 31443 11527 31501 11539
rect 31725 11715 31783 11727
rect 31725 11539 31737 11715
rect 31771 11539 31783 11715
rect 31725 11527 31783 11539
rect 31883 11715 31941 11727
rect 31883 11539 31895 11715
rect 31929 11539 31941 11715
rect 31883 11527 31941 11539
rect 32290 11715 32348 11727
rect 32290 11539 32302 11715
rect 32336 11539 32348 11715
rect 32290 11527 32348 11539
rect 32448 11715 32506 11727
rect 32448 11539 32460 11715
rect 32494 11539 32506 11715
rect 32448 11527 32506 11539
rect 32606 11715 32664 11727
rect 32606 11539 32618 11715
rect 32652 11539 32664 11715
rect 32606 11527 32664 11539
rect 32764 11715 32822 11727
rect 32764 11539 32776 11715
rect 32810 11539 32822 11715
rect 32764 11527 32822 11539
rect 33045 11715 33103 11727
rect 33045 11539 33057 11715
rect 33091 11539 33103 11715
rect 33045 11527 33103 11539
rect 33203 11715 33261 11727
rect 33203 11539 33215 11715
rect 33249 11539 33261 11715
rect 33203 11527 33261 11539
rect 33485 11715 33543 11727
rect 33485 11539 33497 11715
rect 33531 11539 33543 11715
rect 33485 11527 33543 11539
rect 33643 11715 33701 11727
rect 33643 11539 33655 11715
rect 33689 11539 33701 11715
rect 33643 11527 33701 11539
rect 33925 11715 33983 11727
rect 33925 11539 33937 11715
rect 33971 11539 33983 11715
rect 33925 11527 33983 11539
rect 34083 11715 34141 11727
rect 34083 11539 34095 11715
rect 34129 11539 34141 11715
rect 34083 11527 34141 11539
rect 34490 11715 34548 11727
rect 34490 11539 34502 11715
rect 34536 11539 34548 11715
rect 34490 11527 34548 11539
rect 34648 11715 34706 11727
rect 34648 11539 34660 11715
rect 34694 11539 34706 11715
rect 34648 11527 34706 11539
rect 34806 11715 34864 11727
rect 34806 11539 34818 11715
rect 34852 11539 34864 11715
rect 34806 11527 34864 11539
rect 34964 11715 35022 11727
rect 34964 11539 34976 11715
rect 35010 11539 35022 11715
rect 34964 11527 35022 11539
rect 35245 11715 35303 11727
rect 35245 11539 35257 11715
rect 35291 11539 35303 11715
rect 35245 11527 35303 11539
rect 35403 11715 35461 11727
rect 35403 11539 35415 11715
rect 35449 11539 35461 11715
rect 35403 11527 35461 11539
rect 35685 11715 35743 11727
rect 35685 11539 35697 11715
rect 35731 11539 35743 11715
rect 35685 11527 35743 11539
rect 35843 11715 35901 11727
rect 35843 11539 35855 11715
rect 35889 11539 35901 11715
rect 35843 11527 35901 11539
rect 36125 11715 36183 11727
rect 36125 11539 36137 11715
rect 36171 11539 36183 11715
rect 36125 11527 36183 11539
rect 36283 11715 36341 11727
rect 36283 11539 36295 11715
rect 36329 11539 36341 11715
rect 36283 11527 36341 11539
rect 33460 7426 33518 7438
rect 33460 7050 33472 7426
rect 33506 7050 33518 7426
rect 33460 7038 33518 7050
rect 33618 7426 33676 7438
rect 33618 7050 33630 7426
rect 33664 7050 33676 7426
rect 33618 7038 33676 7050
rect 33776 7426 33834 7438
rect 33776 7050 33788 7426
rect 33822 7050 33834 7426
rect 33776 7038 33834 7050
rect 33934 7426 33992 7438
rect 33934 7050 33946 7426
rect 33980 7050 33992 7426
rect 33934 7038 33992 7050
rect 34092 7426 34150 7438
rect 34092 7050 34104 7426
rect 34138 7050 34150 7426
rect 34092 7038 34150 7050
rect 29758 6234 30558 6246
rect 29758 6200 29770 6234
rect 30546 6200 30558 6234
rect 29758 6188 30558 6200
rect 29758 5976 30558 5988
rect 29758 5942 29770 5976
rect 30546 5942 30558 5976
rect 29758 5930 30558 5942
rect 31098 6234 31898 6246
rect 31098 6200 31110 6234
rect 31886 6200 31898 6234
rect 31098 6188 31898 6200
rect 31098 5976 31898 5988
rect 31098 5942 31110 5976
rect 31886 5942 31898 5976
rect 31098 5930 31898 5942
rect 29910 5496 29968 5508
rect 29910 5420 29922 5496
rect 29956 5420 29968 5496
rect 29910 5408 29968 5420
rect 30368 5496 30426 5508
rect 30368 5420 30380 5496
rect 30414 5420 30426 5496
rect 30368 5408 30426 5420
rect 31220 5496 31278 5508
rect 31220 5420 31232 5496
rect 31266 5420 31278 5496
rect 31220 5408 31278 5420
rect 31678 5496 31736 5508
rect 31678 5420 31690 5496
rect 31724 5420 31736 5496
rect 31678 5408 31736 5420
rect 29758 4974 30558 4986
rect 29758 4940 29770 4974
rect 30546 4940 30558 4974
rect 29758 4928 30558 4940
rect 29758 4716 30558 4728
rect 29758 4682 29770 4716
rect 30546 4682 30558 4716
rect 29758 4670 30558 4682
rect 31098 4974 31898 4986
rect 31098 4940 31110 4974
rect 31886 4940 31898 4974
rect 31098 4928 31898 4940
rect 31098 4716 31898 4728
rect 31098 4682 31110 4716
rect 31886 4682 31898 4716
rect 31098 4670 31898 4682
rect 17090 3304 17148 3316
rect 17090 2528 17102 3304
rect 17136 2528 17148 3304
rect 17090 2516 17148 2528
rect 17248 3304 17306 3316
rect 17248 2528 17260 3304
rect 17294 2528 17306 3304
rect 17248 2516 17306 2528
rect 17406 3304 17464 3316
rect 17406 2528 17418 3304
rect 17452 2528 17464 3304
rect 17406 2516 17464 2528
rect 17564 3304 17622 3316
rect 17564 2528 17576 3304
rect 17610 2528 17622 3304
rect 17564 2516 17622 2528
rect 17722 3304 17780 3316
rect 17722 2528 17734 3304
rect 17768 2528 17780 3304
rect 17722 2516 17780 2528
rect 32710 3946 32768 3958
rect 32710 3570 32722 3946
rect 32756 3570 32768 3946
rect 32710 3558 32768 3570
rect 32868 3946 32926 3958
rect 32868 3570 32880 3946
rect 32914 3570 32926 3946
rect 32868 3558 32926 3570
rect 33026 3946 33084 3958
rect 33026 3570 33038 3946
rect 33072 3570 33084 3946
rect 33026 3558 33084 3570
rect 33184 3946 33242 3958
rect 33184 3570 33196 3946
rect 33230 3570 33242 3946
rect 33184 3558 33242 3570
rect 33342 3946 33400 3958
rect 33342 3570 33354 3946
rect 33388 3570 33400 3946
rect 33342 3558 33400 3570
rect 33500 3946 33558 3958
rect 33500 3570 33512 3946
rect 33546 3570 33558 3946
rect 33500 3558 33558 3570
rect 33658 3946 33716 3958
rect 33658 3570 33670 3946
rect 33704 3570 33716 3946
rect 33658 3558 33716 3570
rect 33816 3946 33874 3958
rect 33816 3570 33828 3946
rect 33862 3570 33874 3946
rect 33816 3558 33874 3570
rect 33974 3946 34032 3958
rect 33974 3570 33986 3946
rect 34020 3570 34032 3946
rect 33974 3558 34032 3570
rect 34900 3946 34958 3958
rect 34900 3570 34912 3946
rect 34946 3570 34958 3946
rect 34900 3558 34958 3570
rect 35058 3946 35116 3958
rect 35058 3570 35070 3946
rect 35104 3570 35116 3946
rect 35058 3558 35116 3570
rect 35216 3946 35274 3958
rect 35216 3570 35228 3946
rect 35262 3570 35274 3946
rect 35216 3558 35274 3570
rect 35374 3946 35432 3958
rect 35374 3570 35386 3946
rect 35420 3570 35432 3946
rect 35374 3558 35432 3570
rect 36448 6000 36848 6012
rect 36448 5966 36460 6000
rect 36836 5966 36848 6000
rect 36448 5954 36848 5966
rect 36448 5742 36848 5754
rect 36448 5708 36460 5742
rect 36836 5708 36848 5742
rect 36448 5696 36848 5708
rect 36448 5484 36848 5496
rect 36448 5450 36460 5484
rect 36836 5450 36848 5484
rect 36448 5438 36848 5450
rect 36448 5226 36848 5238
rect 36448 5192 36460 5226
rect 36836 5192 36848 5226
rect 36448 5180 36848 5192
rect 36448 4968 36848 4980
rect 36448 4934 36460 4968
rect 36836 4934 36848 4968
rect 36448 4922 36848 4934
rect 36448 4710 36848 4722
rect 36448 4676 36460 4710
rect 36836 4676 36848 4710
rect 36448 4664 36848 4676
rect 36448 4452 36848 4464
rect 36448 4418 36460 4452
rect 36836 4418 36848 4452
rect 36448 4406 36848 4418
rect 36448 4194 36848 4206
rect 36448 4160 36460 4194
rect 36836 4160 36848 4194
rect 36448 4148 36848 4160
rect 36448 3936 36848 3948
rect 36448 3902 36460 3936
rect 36836 3902 36848 3936
rect 36448 3890 36848 3902
rect 37234 6000 37634 6012
rect 37234 5966 37246 6000
rect 37622 5966 37634 6000
rect 37234 5954 37634 5966
rect 37234 5742 37634 5754
rect 37234 5708 37246 5742
rect 37622 5708 37634 5742
rect 37234 5696 37634 5708
rect 37234 5484 37634 5496
rect 37234 5450 37246 5484
rect 37622 5450 37634 5484
rect 37234 5438 37634 5450
rect 37234 5226 37634 5238
rect 37234 5192 37246 5226
rect 37622 5192 37634 5226
rect 37234 5180 37634 5192
rect 37234 4968 37634 4980
rect 37234 4934 37246 4968
rect 37622 4934 37634 4968
rect 37234 4922 37634 4934
rect 37234 4710 37634 4722
rect 37234 4676 37246 4710
rect 37622 4676 37634 4710
rect 37234 4664 37634 4676
rect 37234 4452 37634 4464
rect 37234 4418 37246 4452
rect 37622 4418 37634 4452
rect 37234 4406 37634 4418
rect 37234 4194 37634 4206
rect 37234 4160 37246 4194
rect 37622 4160 37634 4194
rect 37234 4148 37634 4160
rect 37234 3936 37634 3948
rect 37234 3902 37246 3936
rect 37622 3902 37634 3936
rect 37234 3890 37634 3902
rect 32380 3016 32438 3028
rect 32380 2640 32392 3016
rect 32426 2640 32438 3016
rect 32380 2628 32438 2640
rect 32538 3016 32596 3028
rect 32538 2640 32550 3016
rect 32584 2640 32596 3016
rect 32538 2628 32596 2640
rect 32696 3016 32754 3028
rect 32696 2640 32708 3016
rect 32742 2640 32754 3016
rect 32696 2628 32754 2640
rect 33980 3016 34038 3028
rect 33980 2640 33992 3016
rect 34026 2640 34038 3016
rect 33980 2628 34038 2640
rect 34138 3016 34196 3028
rect 34138 2640 34150 3016
rect 34184 2640 34196 3016
rect 34138 2628 34196 2640
rect 34296 3016 34354 3028
rect 34296 2640 34308 3016
rect 34342 2640 34354 3016
rect 34296 2628 34354 2640
rect 35580 3016 35638 3028
rect 35580 2640 35592 3016
rect 35626 2640 35638 3016
rect 35580 2628 35638 2640
rect 35738 3016 35796 3028
rect 35738 2640 35750 3016
rect 35784 2640 35796 3016
rect 35738 2628 35796 2640
rect 35896 3016 35954 3028
rect 35896 2640 35908 3016
rect 35942 2640 35954 3016
rect 35896 2628 35954 2640
rect 59 2095 459 2107
rect 59 2061 71 2095
rect 447 2061 459 2095
rect 59 2049 459 2061
rect 677 2095 1077 2107
rect 677 2061 689 2095
rect 1065 2061 1077 2095
rect 677 2049 1077 2061
rect 59 1237 459 1249
rect 59 1203 71 1237
rect 447 1203 459 1237
rect 59 1191 459 1203
rect 677 1237 1077 1249
rect 677 1203 689 1237
rect 1065 1203 1077 1237
rect 677 1191 1077 1203
rect 59 949 459 961
rect 59 915 71 949
rect 447 915 459 949
rect 59 903 459 915
rect 677 949 1077 961
rect 677 915 689 949
rect 1065 915 1077 949
rect 677 903 1077 915
rect 59 691 459 703
rect 59 657 71 691
rect 447 657 459 691
rect 59 645 459 657
rect 677 691 1077 703
rect 677 657 689 691
rect 1065 657 1077 691
rect 677 645 1077 657
rect 1659 2095 2059 2107
rect 1659 2061 1671 2095
rect 2047 2061 2059 2095
rect 1659 2049 2059 2061
rect 2277 2095 2677 2107
rect 2277 2061 2289 2095
rect 2665 2061 2677 2095
rect 2277 2049 2677 2061
rect 1659 1237 2059 1249
rect 1659 1203 1671 1237
rect 2047 1203 2059 1237
rect 1659 1191 2059 1203
rect 2277 1237 2677 1249
rect 2277 1203 2289 1237
rect 2665 1203 2677 1237
rect 2277 1191 2677 1203
rect 1659 949 2059 961
rect 1659 915 1671 949
rect 2047 915 2059 949
rect 1659 903 2059 915
rect 2277 949 2677 961
rect 2277 915 2289 949
rect 2665 915 2677 949
rect 2277 903 2677 915
rect 1659 691 2059 703
rect 1659 657 1671 691
rect 2047 657 2059 691
rect 1659 645 2059 657
rect 2277 691 2677 703
rect 2277 657 2289 691
rect 2665 657 2677 691
rect 2277 645 2677 657
rect 3259 2095 3659 2107
rect 3259 2061 3271 2095
rect 3647 2061 3659 2095
rect 3259 2049 3659 2061
rect 3877 2095 4277 2107
rect 3877 2061 3889 2095
rect 4265 2061 4277 2095
rect 3877 2049 4277 2061
rect 3259 1237 3659 1249
rect 3259 1203 3271 1237
rect 3647 1203 3659 1237
rect 3259 1191 3659 1203
rect 3877 1237 4277 1249
rect 3877 1203 3889 1237
rect 4265 1203 4277 1237
rect 3877 1191 4277 1203
rect 3259 949 3659 961
rect 3259 915 3271 949
rect 3647 915 3659 949
rect 3259 903 3659 915
rect 3877 949 4277 961
rect 3877 915 3889 949
rect 4265 915 4277 949
rect 3877 903 4277 915
rect 3259 691 3659 703
rect 3259 657 3271 691
rect 3647 657 3659 691
rect 3259 645 3659 657
rect 3877 691 4277 703
rect 3877 657 3889 691
rect 4265 657 4277 691
rect 3877 645 4277 657
rect 4859 2095 5259 2107
rect 4859 2061 4871 2095
rect 5247 2061 5259 2095
rect 4859 2049 5259 2061
rect 5477 2095 5877 2107
rect 5477 2061 5489 2095
rect 5865 2061 5877 2095
rect 5477 2049 5877 2061
rect 4859 1237 5259 1249
rect 4859 1203 4871 1237
rect 5247 1203 5259 1237
rect 4859 1191 5259 1203
rect 5477 1237 5877 1249
rect 5477 1203 5489 1237
rect 5865 1203 5877 1237
rect 5477 1191 5877 1203
rect 4859 949 5259 961
rect 4859 915 4871 949
rect 5247 915 5259 949
rect 4859 903 5259 915
rect 5477 949 5877 961
rect 5477 915 5489 949
rect 5865 915 5877 949
rect 5477 903 5877 915
rect 4859 691 5259 703
rect 4859 657 4871 691
rect 5247 657 5259 691
rect 4859 645 5259 657
rect 5477 691 5877 703
rect 5477 657 5489 691
rect 5865 657 5877 691
rect 5477 645 5877 657
rect 6459 2095 6859 2107
rect 6459 2061 6471 2095
rect 6847 2061 6859 2095
rect 6459 2049 6859 2061
rect 7077 2095 7477 2107
rect 7077 2061 7089 2095
rect 7465 2061 7477 2095
rect 7077 2049 7477 2061
rect 6459 1237 6859 1249
rect 6459 1203 6471 1237
rect 6847 1203 6859 1237
rect 6459 1191 6859 1203
rect 7077 1237 7477 1249
rect 7077 1203 7089 1237
rect 7465 1203 7477 1237
rect 7077 1191 7477 1203
rect 6459 949 6859 961
rect 6459 915 6471 949
rect 6847 915 6859 949
rect 6459 903 6859 915
rect 7077 949 7477 961
rect 7077 915 7089 949
rect 7465 915 7477 949
rect 7077 903 7477 915
rect 6459 691 6859 703
rect 6459 657 6471 691
rect 6847 657 6859 691
rect 6459 645 6859 657
rect 7077 691 7477 703
rect 7077 657 7089 691
rect 7465 657 7477 691
rect 7077 645 7477 657
rect 8059 2095 8459 2107
rect 8059 2061 8071 2095
rect 8447 2061 8459 2095
rect 8059 2049 8459 2061
rect 8677 2095 9077 2107
rect 8677 2061 8689 2095
rect 9065 2061 9077 2095
rect 8677 2049 9077 2061
rect 8059 1237 8459 1249
rect 8059 1203 8071 1237
rect 8447 1203 8459 1237
rect 8059 1191 8459 1203
rect 8677 1237 9077 1249
rect 8677 1203 8689 1237
rect 9065 1203 9077 1237
rect 8677 1191 9077 1203
rect 8059 949 8459 961
rect 8059 915 8071 949
rect 8447 915 8459 949
rect 8059 903 8459 915
rect 8677 949 9077 961
rect 8677 915 8689 949
rect 9065 915 9077 949
rect 8677 903 9077 915
rect 8059 691 8459 703
rect 8059 657 8071 691
rect 8447 657 8459 691
rect 8059 645 8459 657
rect 8677 691 9077 703
rect 8677 657 8689 691
rect 9065 657 9077 691
rect 8677 645 9077 657
rect 9659 2095 10059 2107
rect 9659 2061 9671 2095
rect 10047 2061 10059 2095
rect 9659 2049 10059 2061
rect 10277 2095 10677 2107
rect 10277 2061 10289 2095
rect 10665 2061 10677 2095
rect 10277 2049 10677 2061
rect 9659 1237 10059 1249
rect 9659 1203 9671 1237
rect 10047 1203 10059 1237
rect 9659 1191 10059 1203
rect 10277 1237 10677 1249
rect 10277 1203 10289 1237
rect 10665 1203 10677 1237
rect 10277 1191 10677 1203
rect 9659 949 10059 961
rect 9659 915 9671 949
rect 10047 915 10059 949
rect 9659 903 10059 915
rect 10277 949 10677 961
rect 10277 915 10289 949
rect 10665 915 10677 949
rect 10277 903 10677 915
rect 9659 691 10059 703
rect 9659 657 9671 691
rect 10047 657 10059 691
rect 9659 645 10059 657
rect 10277 691 10677 703
rect 10277 657 10289 691
rect 10665 657 10677 691
rect 10277 645 10677 657
rect 11259 2095 11659 2107
rect 11259 2061 11271 2095
rect 11647 2061 11659 2095
rect 11259 2049 11659 2061
rect 11877 2095 12277 2107
rect 11877 2061 11889 2095
rect 12265 2061 12277 2095
rect 11877 2049 12277 2061
rect 11259 1237 11659 1249
rect 11259 1203 11271 1237
rect 11647 1203 11659 1237
rect 11259 1191 11659 1203
rect 11877 1237 12277 1249
rect 11877 1203 11889 1237
rect 12265 1203 12277 1237
rect 11877 1191 12277 1203
rect 11259 949 11659 961
rect 11259 915 11271 949
rect 11647 915 11659 949
rect 11259 903 11659 915
rect 11877 949 12277 961
rect 11877 915 11889 949
rect 12265 915 12277 949
rect 11877 903 12277 915
rect 11259 691 11659 703
rect 11259 657 11271 691
rect 11647 657 11659 691
rect 11259 645 11659 657
rect 11877 691 12277 703
rect 11877 657 11889 691
rect 12265 657 12277 691
rect 11877 645 12277 657
rect 12859 2095 13259 2107
rect 12859 2061 12871 2095
rect 13247 2061 13259 2095
rect 12859 2049 13259 2061
rect 13477 2095 13877 2107
rect 13477 2061 13489 2095
rect 13865 2061 13877 2095
rect 13477 2049 13877 2061
rect 12859 1237 13259 1249
rect 12859 1203 12871 1237
rect 13247 1203 13259 1237
rect 12859 1191 13259 1203
rect 13477 1237 13877 1249
rect 13477 1203 13489 1237
rect 13865 1203 13877 1237
rect 13477 1191 13877 1203
rect 12859 949 13259 961
rect 12859 915 12871 949
rect 13247 915 13259 949
rect 12859 903 13259 915
rect 13477 949 13877 961
rect 13477 915 13489 949
rect 13865 915 13877 949
rect 13477 903 13877 915
rect 12859 691 13259 703
rect 12859 657 12871 691
rect 13247 657 13259 691
rect 12859 645 13259 657
rect 13477 691 13877 703
rect 13477 657 13489 691
rect 13865 657 13877 691
rect 13477 645 13877 657
rect 14459 2095 14859 2107
rect 14459 2061 14471 2095
rect 14847 2061 14859 2095
rect 14459 2049 14859 2061
rect 15077 2095 15477 2107
rect 15077 2061 15089 2095
rect 15465 2061 15477 2095
rect 15077 2049 15477 2061
rect 14459 1237 14859 1249
rect 14459 1203 14471 1237
rect 14847 1203 14859 1237
rect 14459 1191 14859 1203
rect 15077 1237 15477 1249
rect 15077 1203 15089 1237
rect 15465 1203 15477 1237
rect 15077 1191 15477 1203
rect 14459 949 14859 961
rect 14459 915 14471 949
rect 14847 915 14859 949
rect 14459 903 14859 915
rect 15077 949 15477 961
rect 15077 915 15089 949
rect 15465 915 15477 949
rect 15077 903 15477 915
rect 14459 691 14859 703
rect 14459 657 14471 691
rect 14847 657 14859 691
rect 14459 645 14859 657
rect 15077 691 15477 703
rect 15077 657 15089 691
rect 15465 657 15477 691
rect 15077 645 15477 657
rect 16059 2095 16459 2107
rect 16059 2061 16071 2095
rect 16447 2061 16459 2095
rect 16059 2049 16459 2061
rect 16677 2095 17077 2107
rect 16677 2061 16689 2095
rect 17065 2061 17077 2095
rect 16677 2049 17077 2061
rect 16059 1237 16459 1249
rect 16059 1203 16071 1237
rect 16447 1203 16459 1237
rect 16059 1191 16459 1203
rect 16677 1237 17077 1249
rect 16677 1203 16689 1237
rect 17065 1203 17077 1237
rect 16677 1191 17077 1203
rect 16059 949 16459 961
rect 16059 915 16071 949
rect 16447 915 16459 949
rect 16059 903 16459 915
rect 16677 949 17077 961
rect 16677 915 16689 949
rect 17065 915 17077 949
rect 16677 903 17077 915
rect 16059 691 16459 703
rect 16059 657 16071 691
rect 16447 657 16459 691
rect 16059 645 16459 657
rect 16677 691 17077 703
rect 16677 657 16689 691
rect 17065 657 17077 691
rect 16677 645 17077 657
rect 17659 2095 18059 2107
rect 17659 2061 17671 2095
rect 18047 2061 18059 2095
rect 17659 2049 18059 2061
rect 18277 2095 18677 2107
rect 18277 2061 18289 2095
rect 18665 2061 18677 2095
rect 18277 2049 18677 2061
rect 17659 1237 18059 1249
rect 17659 1203 17671 1237
rect 18047 1203 18059 1237
rect 17659 1191 18059 1203
rect 18277 1237 18677 1249
rect 18277 1203 18289 1237
rect 18665 1203 18677 1237
rect 18277 1191 18677 1203
rect 17659 949 18059 961
rect 17659 915 17671 949
rect 18047 915 18059 949
rect 17659 903 18059 915
rect 18277 949 18677 961
rect 18277 915 18289 949
rect 18665 915 18677 949
rect 18277 903 18677 915
rect 17659 691 18059 703
rect 17659 657 17671 691
rect 18047 657 18059 691
rect 17659 645 18059 657
rect 18277 691 18677 703
rect 18277 657 18289 691
rect 18665 657 18677 691
rect 18277 645 18677 657
rect 19259 2095 19659 2107
rect 19259 2061 19271 2095
rect 19647 2061 19659 2095
rect 19259 2049 19659 2061
rect 19877 2095 20277 2107
rect 19877 2061 19889 2095
rect 20265 2061 20277 2095
rect 19877 2049 20277 2061
rect 19259 1237 19659 1249
rect 19259 1203 19271 1237
rect 19647 1203 19659 1237
rect 19259 1191 19659 1203
rect 19877 1237 20277 1249
rect 19877 1203 19889 1237
rect 20265 1203 20277 1237
rect 19877 1191 20277 1203
rect 19259 949 19659 961
rect 19259 915 19271 949
rect 19647 915 19659 949
rect 19259 903 19659 915
rect 19877 949 20277 961
rect 19877 915 19889 949
rect 20265 915 20277 949
rect 19877 903 20277 915
rect 19259 691 19659 703
rect 19259 657 19271 691
rect 19647 657 19659 691
rect 19259 645 19659 657
rect 19877 691 20277 703
rect 19877 657 19889 691
rect 20265 657 20277 691
rect 19877 645 20277 657
rect 20859 2095 21259 2107
rect 20859 2061 20871 2095
rect 21247 2061 21259 2095
rect 20859 2049 21259 2061
rect 21477 2095 21877 2107
rect 21477 2061 21489 2095
rect 21865 2061 21877 2095
rect 21477 2049 21877 2061
rect 20859 1237 21259 1249
rect 20859 1203 20871 1237
rect 21247 1203 21259 1237
rect 20859 1191 21259 1203
rect 21477 1237 21877 1249
rect 21477 1203 21489 1237
rect 21865 1203 21877 1237
rect 21477 1191 21877 1203
rect 20859 949 21259 961
rect 20859 915 20871 949
rect 21247 915 21259 949
rect 20859 903 21259 915
rect 21477 949 21877 961
rect 21477 915 21489 949
rect 21865 915 21877 949
rect 21477 903 21877 915
rect 20859 691 21259 703
rect 20859 657 20871 691
rect 21247 657 21259 691
rect 20859 645 21259 657
rect 21477 691 21877 703
rect 21477 657 21489 691
rect 21865 657 21877 691
rect 21477 645 21877 657
rect 22459 2095 22859 2107
rect 22459 2061 22471 2095
rect 22847 2061 22859 2095
rect 22459 2049 22859 2061
rect 23077 2095 23477 2107
rect 23077 2061 23089 2095
rect 23465 2061 23477 2095
rect 23077 2049 23477 2061
rect 22459 1237 22859 1249
rect 22459 1203 22471 1237
rect 22847 1203 22859 1237
rect 22459 1191 22859 1203
rect 23077 1237 23477 1249
rect 23077 1203 23089 1237
rect 23465 1203 23477 1237
rect 23077 1191 23477 1203
rect 22459 949 22859 961
rect 22459 915 22471 949
rect 22847 915 22859 949
rect 22459 903 22859 915
rect 23077 949 23477 961
rect 23077 915 23089 949
rect 23465 915 23477 949
rect 23077 903 23477 915
rect 22459 691 22859 703
rect 22459 657 22471 691
rect 22847 657 22859 691
rect 22459 645 22859 657
rect 23077 691 23477 703
rect 23077 657 23089 691
rect 23465 657 23477 691
rect 23077 645 23477 657
rect 24059 2095 24459 2107
rect 24059 2061 24071 2095
rect 24447 2061 24459 2095
rect 24059 2049 24459 2061
rect 24677 2095 25077 2107
rect 24677 2061 24689 2095
rect 25065 2061 25077 2095
rect 24677 2049 25077 2061
rect 24059 1237 24459 1249
rect 24059 1203 24071 1237
rect 24447 1203 24459 1237
rect 24059 1191 24459 1203
rect 24677 1237 25077 1249
rect 24677 1203 24689 1237
rect 25065 1203 25077 1237
rect 24677 1191 25077 1203
rect 24059 949 24459 961
rect 24059 915 24071 949
rect 24447 915 24459 949
rect 24059 903 24459 915
rect 24677 949 25077 961
rect 24677 915 24689 949
rect 25065 915 25077 949
rect 24677 903 25077 915
rect 24059 691 24459 703
rect 24059 657 24071 691
rect 24447 657 24459 691
rect 24059 645 24459 657
rect 24677 691 25077 703
rect 24677 657 24689 691
rect 25065 657 25077 691
rect 24677 645 25077 657
rect 25659 2095 26059 2107
rect 25659 2061 25671 2095
rect 26047 2061 26059 2095
rect 25659 2049 26059 2061
rect 26277 2095 26677 2107
rect 26277 2061 26289 2095
rect 26665 2061 26677 2095
rect 26277 2049 26677 2061
rect 25659 1237 26059 1249
rect 25659 1203 25671 1237
rect 26047 1203 26059 1237
rect 25659 1191 26059 1203
rect 26277 1237 26677 1249
rect 26277 1203 26289 1237
rect 26665 1203 26677 1237
rect 26277 1191 26677 1203
rect 25659 949 26059 961
rect 25659 915 25671 949
rect 26047 915 26059 949
rect 25659 903 26059 915
rect 26277 949 26677 961
rect 26277 915 26289 949
rect 26665 915 26677 949
rect 26277 903 26677 915
rect 25659 691 26059 703
rect 25659 657 25671 691
rect 26047 657 26059 691
rect 25659 645 26059 657
rect 26277 691 26677 703
rect 26277 657 26289 691
rect 26665 657 26677 691
rect 26277 645 26677 657
rect 27259 2095 27659 2107
rect 27259 2061 27271 2095
rect 27647 2061 27659 2095
rect 27259 2049 27659 2061
rect 27877 2095 28277 2107
rect 27877 2061 27889 2095
rect 28265 2061 28277 2095
rect 27877 2049 28277 2061
rect 27259 1237 27659 1249
rect 27259 1203 27271 1237
rect 27647 1203 27659 1237
rect 27259 1191 27659 1203
rect 27877 1237 28277 1249
rect 27877 1203 27889 1237
rect 28265 1203 28277 1237
rect 27877 1191 28277 1203
rect 27259 949 27659 961
rect 27259 915 27271 949
rect 27647 915 27659 949
rect 27259 903 27659 915
rect 27877 949 28277 961
rect 27877 915 27889 949
rect 28265 915 28277 949
rect 27877 903 28277 915
rect 27259 691 27659 703
rect 27259 657 27271 691
rect 27647 657 27659 691
rect 27259 645 27659 657
rect 27877 691 28277 703
rect 27877 657 27889 691
rect 28265 657 28277 691
rect 27877 645 28277 657
rect 28859 2095 29259 2107
rect 28859 2061 28871 2095
rect 29247 2061 29259 2095
rect 28859 2049 29259 2061
rect 29477 2095 29877 2107
rect 29477 2061 29489 2095
rect 29865 2061 29877 2095
rect 29477 2049 29877 2061
rect 28859 1237 29259 1249
rect 28859 1203 28871 1237
rect 29247 1203 29259 1237
rect 28859 1191 29259 1203
rect 29477 1237 29877 1249
rect 29477 1203 29489 1237
rect 29865 1203 29877 1237
rect 29477 1191 29877 1203
rect 28859 949 29259 961
rect 28859 915 28871 949
rect 29247 915 29259 949
rect 28859 903 29259 915
rect 29477 949 29877 961
rect 29477 915 29489 949
rect 29865 915 29877 949
rect 29477 903 29877 915
rect 28859 691 29259 703
rect 28859 657 28871 691
rect 29247 657 29259 691
rect 28859 645 29259 657
rect 29477 691 29877 703
rect 29477 657 29489 691
rect 29865 657 29877 691
rect 29477 645 29877 657
rect 30459 2095 30859 2107
rect 30459 2061 30471 2095
rect 30847 2061 30859 2095
rect 30459 2049 30859 2061
rect 31077 2095 31477 2107
rect 31077 2061 31089 2095
rect 31465 2061 31477 2095
rect 31077 2049 31477 2061
rect 30459 1237 30859 1249
rect 30459 1203 30471 1237
rect 30847 1203 30859 1237
rect 30459 1191 30859 1203
rect 31077 1237 31477 1249
rect 31077 1203 31089 1237
rect 31465 1203 31477 1237
rect 31077 1191 31477 1203
rect 30459 949 30859 961
rect 30459 915 30471 949
rect 30847 915 30859 949
rect 30459 903 30859 915
rect 31077 949 31477 961
rect 31077 915 31089 949
rect 31465 915 31477 949
rect 31077 903 31477 915
rect 30459 691 30859 703
rect 30459 657 30471 691
rect 30847 657 30859 691
rect 30459 645 30859 657
rect 31077 691 31477 703
rect 31077 657 31089 691
rect 31465 657 31477 691
rect 31077 645 31477 657
rect 32059 2095 32459 2107
rect 32059 2061 32071 2095
rect 32447 2061 32459 2095
rect 32059 2049 32459 2061
rect 32677 2095 33077 2107
rect 32677 2061 32689 2095
rect 33065 2061 33077 2095
rect 32677 2049 33077 2061
rect 32059 1237 32459 1249
rect 32059 1203 32071 1237
rect 32447 1203 32459 1237
rect 32059 1191 32459 1203
rect 32677 1237 33077 1249
rect 32677 1203 32689 1237
rect 33065 1203 33077 1237
rect 32677 1191 33077 1203
rect 32059 949 32459 961
rect 32059 915 32071 949
rect 32447 915 32459 949
rect 32059 903 32459 915
rect 32677 949 33077 961
rect 32677 915 32689 949
rect 33065 915 33077 949
rect 32677 903 33077 915
rect 32059 691 32459 703
rect 32059 657 32071 691
rect 32447 657 32459 691
rect 32059 645 32459 657
rect 32677 691 33077 703
rect 32677 657 32689 691
rect 33065 657 33077 691
rect 32677 645 33077 657
rect 33659 2095 34059 2107
rect 33659 2061 33671 2095
rect 34047 2061 34059 2095
rect 33659 2049 34059 2061
rect 34277 2095 34677 2107
rect 34277 2061 34289 2095
rect 34665 2061 34677 2095
rect 34277 2049 34677 2061
rect 33659 1237 34059 1249
rect 33659 1203 33671 1237
rect 34047 1203 34059 1237
rect 33659 1191 34059 1203
rect 34277 1237 34677 1249
rect 34277 1203 34289 1237
rect 34665 1203 34677 1237
rect 34277 1191 34677 1203
rect 33659 949 34059 961
rect 33659 915 33671 949
rect 34047 915 34059 949
rect 33659 903 34059 915
rect 34277 949 34677 961
rect 34277 915 34289 949
rect 34665 915 34677 949
rect 34277 903 34677 915
rect 33659 691 34059 703
rect 33659 657 33671 691
rect 34047 657 34059 691
rect 33659 645 34059 657
rect 34277 691 34677 703
rect 34277 657 34289 691
rect 34665 657 34677 691
rect 34277 645 34677 657
rect 35259 2095 35659 2107
rect 35259 2061 35271 2095
rect 35647 2061 35659 2095
rect 35259 2049 35659 2061
rect 35877 2095 36277 2107
rect 35877 2061 35889 2095
rect 36265 2061 36277 2095
rect 35877 2049 36277 2061
rect 35259 1237 35659 1249
rect 35259 1203 35271 1237
rect 35647 1203 35659 1237
rect 35259 1191 35659 1203
rect 35877 1237 36277 1249
rect 35877 1203 35889 1237
rect 36265 1203 36277 1237
rect 35877 1191 36277 1203
rect 35259 949 35659 961
rect 35259 915 35271 949
rect 35647 915 35659 949
rect 35259 903 35659 915
rect 35877 949 36277 961
rect 35877 915 35889 949
rect 36265 915 36277 949
rect 35877 903 36277 915
rect 35259 691 35659 703
rect 35259 657 35271 691
rect 35647 657 35659 691
rect 35259 645 35659 657
rect 35877 691 36277 703
rect 35877 657 35889 691
rect 36265 657 36277 691
rect 35877 645 36277 657
rect 36859 2095 37259 2107
rect 36859 2061 36871 2095
rect 37247 2061 37259 2095
rect 36859 2049 37259 2061
rect 37477 2095 37877 2107
rect 37477 2061 37489 2095
rect 37865 2061 37877 2095
rect 37477 2049 37877 2061
rect 36859 1237 37259 1249
rect 36859 1203 36871 1237
rect 37247 1203 37259 1237
rect 36859 1191 37259 1203
rect 37477 1237 37877 1249
rect 37477 1203 37489 1237
rect 37865 1203 37877 1237
rect 37477 1191 37877 1203
rect 36859 949 37259 961
rect 36859 915 36871 949
rect 37247 915 37259 949
rect 36859 903 37259 915
rect 37477 949 37877 961
rect 37477 915 37489 949
rect 37865 915 37877 949
rect 37477 903 37877 915
rect 36859 691 37259 703
rect 36859 657 36871 691
rect 37247 657 37259 691
rect 36859 645 37259 657
rect 37477 691 37877 703
rect 37477 657 37489 691
rect 37865 657 37877 691
rect 37477 645 37877 657
rect 59 295 459 307
rect 59 261 71 295
rect 447 261 459 295
rect 59 249 459 261
rect 677 295 1077 307
rect 677 261 689 295
rect 1065 261 1077 295
rect 677 249 1077 261
rect 59 -563 459 -551
rect 59 -597 71 -563
rect 447 -597 459 -563
rect 59 -609 459 -597
rect 677 -563 1077 -551
rect 677 -597 689 -563
rect 1065 -597 1077 -563
rect 677 -609 1077 -597
rect 59 -851 459 -839
rect 59 -885 71 -851
rect 447 -885 459 -851
rect 59 -897 459 -885
rect 677 -851 1077 -839
rect 677 -885 689 -851
rect 1065 -885 1077 -851
rect 677 -897 1077 -885
rect 59 -1109 459 -1097
rect 59 -1143 71 -1109
rect 447 -1143 459 -1109
rect 59 -1155 459 -1143
rect 677 -1109 1077 -1097
rect 677 -1143 689 -1109
rect 1065 -1143 1077 -1109
rect 677 -1155 1077 -1143
rect 1659 295 2059 307
rect 1659 261 1671 295
rect 2047 261 2059 295
rect 1659 249 2059 261
rect 2277 295 2677 307
rect 2277 261 2289 295
rect 2665 261 2677 295
rect 2277 249 2677 261
rect 1659 -563 2059 -551
rect 1659 -597 1671 -563
rect 2047 -597 2059 -563
rect 1659 -609 2059 -597
rect 2277 -563 2677 -551
rect 2277 -597 2289 -563
rect 2665 -597 2677 -563
rect 2277 -609 2677 -597
rect 1659 -851 2059 -839
rect 1659 -885 1671 -851
rect 2047 -885 2059 -851
rect 1659 -897 2059 -885
rect 2277 -851 2677 -839
rect 2277 -885 2289 -851
rect 2665 -885 2677 -851
rect 2277 -897 2677 -885
rect 1659 -1109 2059 -1097
rect 1659 -1143 1671 -1109
rect 2047 -1143 2059 -1109
rect 1659 -1155 2059 -1143
rect 2277 -1109 2677 -1097
rect 2277 -1143 2289 -1109
rect 2665 -1143 2677 -1109
rect 2277 -1155 2677 -1143
rect 3259 295 3659 307
rect 3259 261 3271 295
rect 3647 261 3659 295
rect 3259 249 3659 261
rect 3877 295 4277 307
rect 3877 261 3889 295
rect 4265 261 4277 295
rect 3877 249 4277 261
rect 3259 -563 3659 -551
rect 3259 -597 3271 -563
rect 3647 -597 3659 -563
rect 3259 -609 3659 -597
rect 3877 -563 4277 -551
rect 3877 -597 3889 -563
rect 4265 -597 4277 -563
rect 3877 -609 4277 -597
rect 3259 -851 3659 -839
rect 3259 -885 3271 -851
rect 3647 -885 3659 -851
rect 3259 -897 3659 -885
rect 3877 -851 4277 -839
rect 3877 -885 3889 -851
rect 4265 -885 4277 -851
rect 3877 -897 4277 -885
rect 3259 -1109 3659 -1097
rect 3259 -1143 3271 -1109
rect 3647 -1143 3659 -1109
rect 3259 -1155 3659 -1143
rect 3877 -1109 4277 -1097
rect 3877 -1143 3889 -1109
rect 4265 -1143 4277 -1109
rect 3877 -1155 4277 -1143
rect 4859 295 5259 307
rect 4859 261 4871 295
rect 5247 261 5259 295
rect 4859 249 5259 261
rect 5477 295 5877 307
rect 5477 261 5489 295
rect 5865 261 5877 295
rect 5477 249 5877 261
rect 4859 -563 5259 -551
rect 4859 -597 4871 -563
rect 5247 -597 5259 -563
rect 4859 -609 5259 -597
rect 5477 -563 5877 -551
rect 5477 -597 5489 -563
rect 5865 -597 5877 -563
rect 5477 -609 5877 -597
rect 4859 -851 5259 -839
rect 4859 -885 4871 -851
rect 5247 -885 5259 -851
rect 4859 -897 5259 -885
rect 5477 -851 5877 -839
rect 5477 -885 5489 -851
rect 5865 -885 5877 -851
rect 5477 -897 5877 -885
rect 4859 -1109 5259 -1097
rect 4859 -1143 4871 -1109
rect 5247 -1143 5259 -1109
rect 4859 -1155 5259 -1143
rect 5477 -1109 5877 -1097
rect 5477 -1143 5489 -1109
rect 5865 -1143 5877 -1109
rect 5477 -1155 5877 -1143
rect 6459 295 6859 307
rect 6459 261 6471 295
rect 6847 261 6859 295
rect 6459 249 6859 261
rect 7077 295 7477 307
rect 7077 261 7089 295
rect 7465 261 7477 295
rect 7077 249 7477 261
rect 6459 -563 6859 -551
rect 6459 -597 6471 -563
rect 6847 -597 6859 -563
rect 6459 -609 6859 -597
rect 7077 -563 7477 -551
rect 7077 -597 7089 -563
rect 7465 -597 7477 -563
rect 7077 -609 7477 -597
rect 6459 -851 6859 -839
rect 6459 -885 6471 -851
rect 6847 -885 6859 -851
rect 6459 -897 6859 -885
rect 7077 -851 7477 -839
rect 7077 -885 7089 -851
rect 7465 -885 7477 -851
rect 7077 -897 7477 -885
rect 6459 -1109 6859 -1097
rect 6459 -1143 6471 -1109
rect 6847 -1143 6859 -1109
rect 6459 -1155 6859 -1143
rect 7077 -1109 7477 -1097
rect 7077 -1143 7089 -1109
rect 7465 -1143 7477 -1109
rect 7077 -1155 7477 -1143
rect 8059 295 8459 307
rect 8059 261 8071 295
rect 8447 261 8459 295
rect 8059 249 8459 261
rect 8677 295 9077 307
rect 8677 261 8689 295
rect 9065 261 9077 295
rect 8677 249 9077 261
rect 8059 -563 8459 -551
rect 8059 -597 8071 -563
rect 8447 -597 8459 -563
rect 8059 -609 8459 -597
rect 8677 -563 9077 -551
rect 8677 -597 8689 -563
rect 9065 -597 9077 -563
rect 8677 -609 9077 -597
rect 8059 -851 8459 -839
rect 8059 -885 8071 -851
rect 8447 -885 8459 -851
rect 8059 -897 8459 -885
rect 8677 -851 9077 -839
rect 8677 -885 8689 -851
rect 9065 -885 9077 -851
rect 8677 -897 9077 -885
rect 8059 -1109 8459 -1097
rect 8059 -1143 8071 -1109
rect 8447 -1143 8459 -1109
rect 8059 -1155 8459 -1143
rect 8677 -1109 9077 -1097
rect 8677 -1143 8689 -1109
rect 9065 -1143 9077 -1109
rect 8677 -1155 9077 -1143
rect 9659 295 10059 307
rect 9659 261 9671 295
rect 10047 261 10059 295
rect 9659 249 10059 261
rect 10277 295 10677 307
rect 10277 261 10289 295
rect 10665 261 10677 295
rect 10277 249 10677 261
rect 9659 -563 10059 -551
rect 9659 -597 9671 -563
rect 10047 -597 10059 -563
rect 9659 -609 10059 -597
rect 10277 -563 10677 -551
rect 10277 -597 10289 -563
rect 10665 -597 10677 -563
rect 10277 -609 10677 -597
rect 9659 -851 10059 -839
rect 9659 -885 9671 -851
rect 10047 -885 10059 -851
rect 9659 -897 10059 -885
rect 10277 -851 10677 -839
rect 10277 -885 10289 -851
rect 10665 -885 10677 -851
rect 10277 -897 10677 -885
rect 9659 -1109 10059 -1097
rect 9659 -1143 9671 -1109
rect 10047 -1143 10059 -1109
rect 9659 -1155 10059 -1143
rect 10277 -1109 10677 -1097
rect 10277 -1143 10289 -1109
rect 10665 -1143 10677 -1109
rect 10277 -1155 10677 -1143
rect 11259 295 11659 307
rect 11259 261 11271 295
rect 11647 261 11659 295
rect 11259 249 11659 261
rect 11877 295 12277 307
rect 11877 261 11889 295
rect 12265 261 12277 295
rect 11877 249 12277 261
rect 11259 -563 11659 -551
rect 11259 -597 11271 -563
rect 11647 -597 11659 -563
rect 11259 -609 11659 -597
rect 11877 -563 12277 -551
rect 11877 -597 11889 -563
rect 12265 -597 12277 -563
rect 11877 -609 12277 -597
rect 11259 -851 11659 -839
rect 11259 -885 11271 -851
rect 11647 -885 11659 -851
rect 11259 -897 11659 -885
rect 11877 -851 12277 -839
rect 11877 -885 11889 -851
rect 12265 -885 12277 -851
rect 11877 -897 12277 -885
rect 11259 -1109 11659 -1097
rect 11259 -1143 11271 -1109
rect 11647 -1143 11659 -1109
rect 11259 -1155 11659 -1143
rect 11877 -1109 12277 -1097
rect 11877 -1143 11889 -1109
rect 12265 -1143 12277 -1109
rect 11877 -1155 12277 -1143
rect 12859 295 13259 307
rect 12859 261 12871 295
rect 13247 261 13259 295
rect 12859 249 13259 261
rect 13477 295 13877 307
rect 13477 261 13489 295
rect 13865 261 13877 295
rect 13477 249 13877 261
rect 12859 -563 13259 -551
rect 12859 -597 12871 -563
rect 13247 -597 13259 -563
rect 12859 -609 13259 -597
rect 13477 -563 13877 -551
rect 13477 -597 13489 -563
rect 13865 -597 13877 -563
rect 13477 -609 13877 -597
rect 12859 -851 13259 -839
rect 12859 -885 12871 -851
rect 13247 -885 13259 -851
rect 12859 -897 13259 -885
rect 13477 -851 13877 -839
rect 13477 -885 13489 -851
rect 13865 -885 13877 -851
rect 13477 -897 13877 -885
rect 12859 -1109 13259 -1097
rect 12859 -1143 12871 -1109
rect 13247 -1143 13259 -1109
rect 12859 -1155 13259 -1143
rect 13477 -1109 13877 -1097
rect 13477 -1143 13489 -1109
rect 13865 -1143 13877 -1109
rect 13477 -1155 13877 -1143
rect 14459 295 14859 307
rect 14459 261 14471 295
rect 14847 261 14859 295
rect 14459 249 14859 261
rect 15077 295 15477 307
rect 15077 261 15089 295
rect 15465 261 15477 295
rect 15077 249 15477 261
rect 14459 -563 14859 -551
rect 14459 -597 14471 -563
rect 14847 -597 14859 -563
rect 14459 -609 14859 -597
rect 15077 -563 15477 -551
rect 15077 -597 15089 -563
rect 15465 -597 15477 -563
rect 15077 -609 15477 -597
rect 14459 -851 14859 -839
rect 14459 -885 14471 -851
rect 14847 -885 14859 -851
rect 14459 -897 14859 -885
rect 15077 -851 15477 -839
rect 15077 -885 15089 -851
rect 15465 -885 15477 -851
rect 15077 -897 15477 -885
rect 14459 -1109 14859 -1097
rect 14459 -1143 14471 -1109
rect 14847 -1143 14859 -1109
rect 14459 -1155 14859 -1143
rect 15077 -1109 15477 -1097
rect 15077 -1143 15089 -1109
rect 15465 -1143 15477 -1109
rect 15077 -1155 15477 -1143
rect 16059 295 16459 307
rect 16059 261 16071 295
rect 16447 261 16459 295
rect 16059 249 16459 261
rect 16677 295 17077 307
rect 16677 261 16689 295
rect 17065 261 17077 295
rect 16677 249 17077 261
rect 16059 -563 16459 -551
rect 16059 -597 16071 -563
rect 16447 -597 16459 -563
rect 16059 -609 16459 -597
rect 16677 -563 17077 -551
rect 16677 -597 16689 -563
rect 17065 -597 17077 -563
rect 16677 -609 17077 -597
rect 16059 -851 16459 -839
rect 16059 -885 16071 -851
rect 16447 -885 16459 -851
rect 16059 -897 16459 -885
rect 16677 -851 17077 -839
rect 16677 -885 16689 -851
rect 17065 -885 17077 -851
rect 16677 -897 17077 -885
rect 16059 -1109 16459 -1097
rect 16059 -1143 16071 -1109
rect 16447 -1143 16459 -1109
rect 16059 -1155 16459 -1143
rect 16677 -1109 17077 -1097
rect 16677 -1143 16689 -1109
rect 17065 -1143 17077 -1109
rect 16677 -1155 17077 -1143
rect 17659 295 18059 307
rect 17659 261 17671 295
rect 18047 261 18059 295
rect 17659 249 18059 261
rect 18277 295 18677 307
rect 18277 261 18289 295
rect 18665 261 18677 295
rect 18277 249 18677 261
rect 17659 -563 18059 -551
rect 17659 -597 17671 -563
rect 18047 -597 18059 -563
rect 17659 -609 18059 -597
rect 18277 -563 18677 -551
rect 18277 -597 18289 -563
rect 18665 -597 18677 -563
rect 18277 -609 18677 -597
rect 17659 -851 18059 -839
rect 17659 -885 17671 -851
rect 18047 -885 18059 -851
rect 17659 -897 18059 -885
rect 18277 -851 18677 -839
rect 18277 -885 18289 -851
rect 18665 -885 18677 -851
rect 18277 -897 18677 -885
rect 17659 -1109 18059 -1097
rect 17659 -1143 17671 -1109
rect 18047 -1143 18059 -1109
rect 17659 -1155 18059 -1143
rect 18277 -1109 18677 -1097
rect 18277 -1143 18289 -1109
rect 18665 -1143 18677 -1109
rect 18277 -1155 18677 -1143
rect 19259 295 19659 307
rect 19259 261 19271 295
rect 19647 261 19659 295
rect 19259 249 19659 261
rect 19877 295 20277 307
rect 19877 261 19889 295
rect 20265 261 20277 295
rect 19877 249 20277 261
rect 19259 -563 19659 -551
rect 19259 -597 19271 -563
rect 19647 -597 19659 -563
rect 19259 -609 19659 -597
rect 19877 -563 20277 -551
rect 19877 -597 19889 -563
rect 20265 -597 20277 -563
rect 19877 -609 20277 -597
rect 19259 -851 19659 -839
rect 19259 -885 19271 -851
rect 19647 -885 19659 -851
rect 19259 -897 19659 -885
rect 19877 -851 20277 -839
rect 19877 -885 19889 -851
rect 20265 -885 20277 -851
rect 19877 -897 20277 -885
rect 19259 -1109 19659 -1097
rect 19259 -1143 19271 -1109
rect 19647 -1143 19659 -1109
rect 19259 -1155 19659 -1143
rect 19877 -1109 20277 -1097
rect 19877 -1143 19889 -1109
rect 20265 -1143 20277 -1109
rect 19877 -1155 20277 -1143
rect 20859 295 21259 307
rect 20859 261 20871 295
rect 21247 261 21259 295
rect 20859 249 21259 261
rect 21477 295 21877 307
rect 21477 261 21489 295
rect 21865 261 21877 295
rect 21477 249 21877 261
rect 20859 -563 21259 -551
rect 20859 -597 20871 -563
rect 21247 -597 21259 -563
rect 20859 -609 21259 -597
rect 21477 -563 21877 -551
rect 21477 -597 21489 -563
rect 21865 -597 21877 -563
rect 21477 -609 21877 -597
rect 20859 -851 21259 -839
rect 20859 -885 20871 -851
rect 21247 -885 21259 -851
rect 20859 -897 21259 -885
rect 21477 -851 21877 -839
rect 21477 -885 21489 -851
rect 21865 -885 21877 -851
rect 21477 -897 21877 -885
rect 20859 -1109 21259 -1097
rect 20859 -1143 20871 -1109
rect 21247 -1143 21259 -1109
rect 20859 -1155 21259 -1143
rect 21477 -1109 21877 -1097
rect 21477 -1143 21489 -1109
rect 21865 -1143 21877 -1109
rect 21477 -1155 21877 -1143
rect 22459 295 22859 307
rect 22459 261 22471 295
rect 22847 261 22859 295
rect 22459 249 22859 261
rect 23077 295 23477 307
rect 23077 261 23089 295
rect 23465 261 23477 295
rect 23077 249 23477 261
rect 22459 -563 22859 -551
rect 22459 -597 22471 -563
rect 22847 -597 22859 -563
rect 22459 -609 22859 -597
rect 23077 -563 23477 -551
rect 23077 -597 23089 -563
rect 23465 -597 23477 -563
rect 23077 -609 23477 -597
rect 22459 -851 22859 -839
rect 22459 -885 22471 -851
rect 22847 -885 22859 -851
rect 22459 -897 22859 -885
rect 23077 -851 23477 -839
rect 23077 -885 23089 -851
rect 23465 -885 23477 -851
rect 23077 -897 23477 -885
rect 22459 -1109 22859 -1097
rect 22459 -1143 22471 -1109
rect 22847 -1143 22859 -1109
rect 22459 -1155 22859 -1143
rect 23077 -1109 23477 -1097
rect 23077 -1143 23089 -1109
rect 23465 -1143 23477 -1109
rect 23077 -1155 23477 -1143
rect 24059 295 24459 307
rect 24059 261 24071 295
rect 24447 261 24459 295
rect 24059 249 24459 261
rect 24677 295 25077 307
rect 24677 261 24689 295
rect 25065 261 25077 295
rect 24677 249 25077 261
rect 24059 -563 24459 -551
rect 24059 -597 24071 -563
rect 24447 -597 24459 -563
rect 24059 -609 24459 -597
rect 24677 -563 25077 -551
rect 24677 -597 24689 -563
rect 25065 -597 25077 -563
rect 24677 -609 25077 -597
rect 24059 -851 24459 -839
rect 24059 -885 24071 -851
rect 24447 -885 24459 -851
rect 24059 -897 24459 -885
rect 24677 -851 25077 -839
rect 24677 -885 24689 -851
rect 25065 -885 25077 -851
rect 24677 -897 25077 -885
rect 24059 -1109 24459 -1097
rect 24059 -1143 24071 -1109
rect 24447 -1143 24459 -1109
rect 24059 -1155 24459 -1143
rect 24677 -1109 25077 -1097
rect 24677 -1143 24689 -1109
rect 25065 -1143 25077 -1109
rect 24677 -1155 25077 -1143
rect 25659 295 26059 307
rect 25659 261 25671 295
rect 26047 261 26059 295
rect 25659 249 26059 261
rect 26277 295 26677 307
rect 26277 261 26289 295
rect 26665 261 26677 295
rect 26277 249 26677 261
rect 25659 -563 26059 -551
rect 25659 -597 25671 -563
rect 26047 -597 26059 -563
rect 25659 -609 26059 -597
rect 26277 -563 26677 -551
rect 26277 -597 26289 -563
rect 26665 -597 26677 -563
rect 26277 -609 26677 -597
rect 25659 -851 26059 -839
rect 25659 -885 25671 -851
rect 26047 -885 26059 -851
rect 25659 -897 26059 -885
rect 26277 -851 26677 -839
rect 26277 -885 26289 -851
rect 26665 -885 26677 -851
rect 26277 -897 26677 -885
rect 25659 -1109 26059 -1097
rect 25659 -1143 25671 -1109
rect 26047 -1143 26059 -1109
rect 25659 -1155 26059 -1143
rect 26277 -1109 26677 -1097
rect 26277 -1143 26289 -1109
rect 26665 -1143 26677 -1109
rect 26277 -1155 26677 -1143
rect 27259 295 27659 307
rect 27259 261 27271 295
rect 27647 261 27659 295
rect 27259 249 27659 261
rect 27877 295 28277 307
rect 27877 261 27889 295
rect 28265 261 28277 295
rect 27877 249 28277 261
rect 27259 -563 27659 -551
rect 27259 -597 27271 -563
rect 27647 -597 27659 -563
rect 27259 -609 27659 -597
rect 27877 -563 28277 -551
rect 27877 -597 27889 -563
rect 28265 -597 28277 -563
rect 27877 -609 28277 -597
rect 27259 -851 27659 -839
rect 27259 -885 27271 -851
rect 27647 -885 27659 -851
rect 27259 -897 27659 -885
rect 27877 -851 28277 -839
rect 27877 -885 27889 -851
rect 28265 -885 28277 -851
rect 27877 -897 28277 -885
rect 27259 -1109 27659 -1097
rect 27259 -1143 27271 -1109
rect 27647 -1143 27659 -1109
rect 27259 -1155 27659 -1143
rect 27877 -1109 28277 -1097
rect 27877 -1143 27889 -1109
rect 28265 -1143 28277 -1109
rect 27877 -1155 28277 -1143
rect 28859 295 29259 307
rect 28859 261 28871 295
rect 29247 261 29259 295
rect 28859 249 29259 261
rect 29477 295 29877 307
rect 29477 261 29489 295
rect 29865 261 29877 295
rect 29477 249 29877 261
rect 28859 -563 29259 -551
rect 28859 -597 28871 -563
rect 29247 -597 29259 -563
rect 28859 -609 29259 -597
rect 29477 -563 29877 -551
rect 29477 -597 29489 -563
rect 29865 -597 29877 -563
rect 29477 -609 29877 -597
rect 28859 -851 29259 -839
rect 28859 -885 28871 -851
rect 29247 -885 29259 -851
rect 28859 -897 29259 -885
rect 29477 -851 29877 -839
rect 29477 -885 29489 -851
rect 29865 -885 29877 -851
rect 29477 -897 29877 -885
rect 28859 -1109 29259 -1097
rect 28859 -1143 28871 -1109
rect 29247 -1143 29259 -1109
rect 28859 -1155 29259 -1143
rect 29477 -1109 29877 -1097
rect 29477 -1143 29489 -1109
rect 29865 -1143 29877 -1109
rect 29477 -1155 29877 -1143
rect 30459 295 30859 307
rect 30459 261 30471 295
rect 30847 261 30859 295
rect 30459 249 30859 261
rect 31077 295 31477 307
rect 31077 261 31089 295
rect 31465 261 31477 295
rect 31077 249 31477 261
rect 30459 -563 30859 -551
rect 30459 -597 30471 -563
rect 30847 -597 30859 -563
rect 30459 -609 30859 -597
rect 31077 -563 31477 -551
rect 31077 -597 31089 -563
rect 31465 -597 31477 -563
rect 31077 -609 31477 -597
rect 30459 -851 30859 -839
rect 30459 -885 30471 -851
rect 30847 -885 30859 -851
rect 30459 -897 30859 -885
rect 31077 -851 31477 -839
rect 31077 -885 31089 -851
rect 31465 -885 31477 -851
rect 31077 -897 31477 -885
rect 30459 -1109 30859 -1097
rect 30459 -1143 30471 -1109
rect 30847 -1143 30859 -1109
rect 30459 -1155 30859 -1143
rect 31077 -1109 31477 -1097
rect 31077 -1143 31089 -1109
rect 31465 -1143 31477 -1109
rect 31077 -1155 31477 -1143
rect 32059 295 32459 307
rect 32059 261 32071 295
rect 32447 261 32459 295
rect 32059 249 32459 261
rect 32677 295 33077 307
rect 32677 261 32689 295
rect 33065 261 33077 295
rect 32677 249 33077 261
rect 32059 -563 32459 -551
rect 32059 -597 32071 -563
rect 32447 -597 32459 -563
rect 32059 -609 32459 -597
rect 32677 -563 33077 -551
rect 32677 -597 32689 -563
rect 33065 -597 33077 -563
rect 32677 -609 33077 -597
rect 32059 -851 32459 -839
rect 32059 -885 32071 -851
rect 32447 -885 32459 -851
rect 32059 -897 32459 -885
rect 32677 -851 33077 -839
rect 32677 -885 32689 -851
rect 33065 -885 33077 -851
rect 32677 -897 33077 -885
rect 32059 -1109 32459 -1097
rect 32059 -1143 32071 -1109
rect 32447 -1143 32459 -1109
rect 32059 -1155 32459 -1143
rect 32677 -1109 33077 -1097
rect 32677 -1143 32689 -1109
rect 33065 -1143 33077 -1109
rect 32677 -1155 33077 -1143
rect 33659 295 34059 307
rect 33659 261 33671 295
rect 34047 261 34059 295
rect 33659 249 34059 261
rect 34277 295 34677 307
rect 34277 261 34289 295
rect 34665 261 34677 295
rect 34277 249 34677 261
rect 33659 -563 34059 -551
rect 33659 -597 33671 -563
rect 34047 -597 34059 -563
rect 33659 -609 34059 -597
rect 34277 -563 34677 -551
rect 34277 -597 34289 -563
rect 34665 -597 34677 -563
rect 34277 -609 34677 -597
rect 33659 -851 34059 -839
rect 33659 -885 33671 -851
rect 34047 -885 34059 -851
rect 33659 -897 34059 -885
rect 34277 -851 34677 -839
rect 34277 -885 34289 -851
rect 34665 -885 34677 -851
rect 34277 -897 34677 -885
rect 33659 -1109 34059 -1097
rect 33659 -1143 33671 -1109
rect 34047 -1143 34059 -1109
rect 33659 -1155 34059 -1143
rect 34277 -1109 34677 -1097
rect 34277 -1143 34289 -1109
rect 34665 -1143 34677 -1109
rect 34277 -1155 34677 -1143
rect 35259 295 35659 307
rect 35259 261 35271 295
rect 35647 261 35659 295
rect 35259 249 35659 261
rect 35877 295 36277 307
rect 35877 261 35889 295
rect 36265 261 36277 295
rect 35877 249 36277 261
rect 35259 -563 35659 -551
rect 35259 -597 35271 -563
rect 35647 -597 35659 -563
rect 35259 -609 35659 -597
rect 35877 -563 36277 -551
rect 35877 -597 35889 -563
rect 36265 -597 36277 -563
rect 35877 -609 36277 -597
rect 35259 -851 35659 -839
rect 35259 -885 35271 -851
rect 35647 -885 35659 -851
rect 35259 -897 35659 -885
rect 35877 -851 36277 -839
rect 35877 -885 35889 -851
rect 36265 -885 36277 -851
rect 35877 -897 36277 -885
rect 35259 -1109 35659 -1097
rect 35259 -1143 35271 -1109
rect 35647 -1143 35659 -1109
rect 35259 -1155 35659 -1143
rect 35877 -1109 36277 -1097
rect 35877 -1143 35889 -1109
rect 36265 -1143 36277 -1109
rect 35877 -1155 36277 -1143
rect 36859 295 37259 307
rect 36859 261 36871 295
rect 37247 261 37259 295
rect 36859 249 37259 261
rect 37477 295 37877 307
rect 37477 261 37489 295
rect 37865 261 37877 295
rect 37477 249 37877 261
rect 36859 -563 37259 -551
rect 36859 -597 36871 -563
rect 37247 -597 37259 -563
rect 36859 -609 37259 -597
rect 37477 -563 37877 -551
rect 37477 -597 37489 -563
rect 37865 -597 37877 -563
rect 37477 -609 37877 -597
rect 36859 -851 37259 -839
rect 36859 -885 36871 -851
rect 37247 -885 37259 -851
rect 36859 -897 37259 -885
rect 37477 -851 37877 -839
rect 37477 -885 37489 -851
rect 37865 -885 37877 -851
rect 37477 -897 37877 -885
rect 36859 -1109 37259 -1097
rect 36859 -1143 36871 -1109
rect 37247 -1143 37259 -1109
rect 36859 -1155 37259 -1143
rect 37477 -1109 37877 -1097
rect 37477 -1143 37489 -1109
rect 37865 -1143 37877 -1109
rect 37477 -1155 37877 -1143
rect 59 -1505 459 -1493
rect 59 -1539 71 -1505
rect 447 -1539 459 -1505
rect 59 -1551 459 -1539
rect 677 -1505 1077 -1493
rect 677 -1539 689 -1505
rect 1065 -1539 1077 -1505
rect 677 -1551 1077 -1539
rect 59 -2363 459 -2351
rect 59 -2397 71 -2363
rect 447 -2397 459 -2363
rect 59 -2409 459 -2397
rect 677 -2363 1077 -2351
rect 677 -2397 689 -2363
rect 1065 -2397 1077 -2363
rect 677 -2409 1077 -2397
rect 59 -2651 459 -2639
rect 59 -2685 71 -2651
rect 447 -2685 459 -2651
rect 59 -2697 459 -2685
rect 677 -2651 1077 -2639
rect 677 -2685 689 -2651
rect 1065 -2685 1077 -2651
rect 677 -2697 1077 -2685
rect 59 -2909 459 -2897
rect 59 -2943 71 -2909
rect 447 -2943 459 -2909
rect 59 -2955 459 -2943
rect 677 -2909 1077 -2897
rect 677 -2943 689 -2909
rect 1065 -2943 1077 -2909
rect 677 -2955 1077 -2943
rect 1659 -1505 2059 -1493
rect 1659 -1539 1671 -1505
rect 2047 -1539 2059 -1505
rect 1659 -1551 2059 -1539
rect 2277 -1505 2677 -1493
rect 2277 -1539 2289 -1505
rect 2665 -1539 2677 -1505
rect 2277 -1551 2677 -1539
rect 1659 -2363 2059 -2351
rect 1659 -2397 1671 -2363
rect 2047 -2397 2059 -2363
rect 1659 -2409 2059 -2397
rect 2277 -2363 2677 -2351
rect 2277 -2397 2289 -2363
rect 2665 -2397 2677 -2363
rect 2277 -2409 2677 -2397
rect 1659 -2651 2059 -2639
rect 1659 -2685 1671 -2651
rect 2047 -2685 2059 -2651
rect 1659 -2697 2059 -2685
rect 2277 -2651 2677 -2639
rect 2277 -2685 2289 -2651
rect 2665 -2685 2677 -2651
rect 2277 -2697 2677 -2685
rect 1659 -2909 2059 -2897
rect 1659 -2943 1671 -2909
rect 2047 -2943 2059 -2909
rect 1659 -2955 2059 -2943
rect 2277 -2909 2677 -2897
rect 2277 -2943 2289 -2909
rect 2665 -2943 2677 -2909
rect 2277 -2955 2677 -2943
rect 3259 -1505 3659 -1493
rect 3259 -1539 3271 -1505
rect 3647 -1539 3659 -1505
rect 3259 -1551 3659 -1539
rect 3877 -1505 4277 -1493
rect 3877 -1539 3889 -1505
rect 4265 -1539 4277 -1505
rect 3877 -1551 4277 -1539
rect 3259 -2363 3659 -2351
rect 3259 -2397 3271 -2363
rect 3647 -2397 3659 -2363
rect 3259 -2409 3659 -2397
rect 3877 -2363 4277 -2351
rect 3877 -2397 3889 -2363
rect 4265 -2397 4277 -2363
rect 3877 -2409 4277 -2397
rect 3259 -2651 3659 -2639
rect 3259 -2685 3271 -2651
rect 3647 -2685 3659 -2651
rect 3259 -2697 3659 -2685
rect 3877 -2651 4277 -2639
rect 3877 -2685 3889 -2651
rect 4265 -2685 4277 -2651
rect 3877 -2697 4277 -2685
rect 3259 -2909 3659 -2897
rect 3259 -2943 3271 -2909
rect 3647 -2943 3659 -2909
rect 3259 -2955 3659 -2943
rect 3877 -2909 4277 -2897
rect 3877 -2943 3889 -2909
rect 4265 -2943 4277 -2909
rect 3877 -2955 4277 -2943
rect 4859 -1505 5259 -1493
rect 4859 -1539 4871 -1505
rect 5247 -1539 5259 -1505
rect 4859 -1551 5259 -1539
rect 5477 -1505 5877 -1493
rect 5477 -1539 5489 -1505
rect 5865 -1539 5877 -1505
rect 5477 -1551 5877 -1539
rect 4859 -2363 5259 -2351
rect 4859 -2397 4871 -2363
rect 5247 -2397 5259 -2363
rect 4859 -2409 5259 -2397
rect 5477 -2363 5877 -2351
rect 5477 -2397 5489 -2363
rect 5865 -2397 5877 -2363
rect 5477 -2409 5877 -2397
rect 4859 -2651 5259 -2639
rect 4859 -2685 4871 -2651
rect 5247 -2685 5259 -2651
rect 4859 -2697 5259 -2685
rect 5477 -2651 5877 -2639
rect 5477 -2685 5489 -2651
rect 5865 -2685 5877 -2651
rect 5477 -2697 5877 -2685
rect 4859 -2909 5259 -2897
rect 4859 -2943 4871 -2909
rect 5247 -2943 5259 -2909
rect 4859 -2955 5259 -2943
rect 5477 -2909 5877 -2897
rect 5477 -2943 5489 -2909
rect 5865 -2943 5877 -2909
rect 5477 -2955 5877 -2943
rect 6459 -1505 6859 -1493
rect 6459 -1539 6471 -1505
rect 6847 -1539 6859 -1505
rect 6459 -1551 6859 -1539
rect 7077 -1505 7477 -1493
rect 7077 -1539 7089 -1505
rect 7465 -1539 7477 -1505
rect 7077 -1551 7477 -1539
rect 6459 -2363 6859 -2351
rect 6459 -2397 6471 -2363
rect 6847 -2397 6859 -2363
rect 6459 -2409 6859 -2397
rect 7077 -2363 7477 -2351
rect 7077 -2397 7089 -2363
rect 7465 -2397 7477 -2363
rect 7077 -2409 7477 -2397
rect 6459 -2651 6859 -2639
rect 6459 -2685 6471 -2651
rect 6847 -2685 6859 -2651
rect 6459 -2697 6859 -2685
rect 7077 -2651 7477 -2639
rect 7077 -2685 7089 -2651
rect 7465 -2685 7477 -2651
rect 7077 -2697 7477 -2685
rect 6459 -2909 6859 -2897
rect 6459 -2943 6471 -2909
rect 6847 -2943 6859 -2909
rect 6459 -2955 6859 -2943
rect 7077 -2909 7477 -2897
rect 7077 -2943 7089 -2909
rect 7465 -2943 7477 -2909
rect 7077 -2955 7477 -2943
rect 8059 -1505 8459 -1493
rect 8059 -1539 8071 -1505
rect 8447 -1539 8459 -1505
rect 8059 -1551 8459 -1539
rect 8677 -1505 9077 -1493
rect 8677 -1539 8689 -1505
rect 9065 -1539 9077 -1505
rect 8677 -1551 9077 -1539
rect 8059 -2363 8459 -2351
rect 8059 -2397 8071 -2363
rect 8447 -2397 8459 -2363
rect 8059 -2409 8459 -2397
rect 8677 -2363 9077 -2351
rect 8677 -2397 8689 -2363
rect 9065 -2397 9077 -2363
rect 8677 -2409 9077 -2397
rect 8059 -2651 8459 -2639
rect 8059 -2685 8071 -2651
rect 8447 -2685 8459 -2651
rect 8059 -2697 8459 -2685
rect 8677 -2651 9077 -2639
rect 8677 -2685 8689 -2651
rect 9065 -2685 9077 -2651
rect 8677 -2697 9077 -2685
rect 8059 -2909 8459 -2897
rect 8059 -2943 8071 -2909
rect 8447 -2943 8459 -2909
rect 8059 -2955 8459 -2943
rect 8677 -2909 9077 -2897
rect 8677 -2943 8689 -2909
rect 9065 -2943 9077 -2909
rect 8677 -2955 9077 -2943
rect 9659 -1505 10059 -1493
rect 9659 -1539 9671 -1505
rect 10047 -1539 10059 -1505
rect 9659 -1551 10059 -1539
rect 10277 -1505 10677 -1493
rect 10277 -1539 10289 -1505
rect 10665 -1539 10677 -1505
rect 10277 -1551 10677 -1539
rect 9659 -2363 10059 -2351
rect 9659 -2397 9671 -2363
rect 10047 -2397 10059 -2363
rect 9659 -2409 10059 -2397
rect 10277 -2363 10677 -2351
rect 10277 -2397 10289 -2363
rect 10665 -2397 10677 -2363
rect 10277 -2409 10677 -2397
rect 9659 -2651 10059 -2639
rect 9659 -2685 9671 -2651
rect 10047 -2685 10059 -2651
rect 9659 -2697 10059 -2685
rect 10277 -2651 10677 -2639
rect 10277 -2685 10289 -2651
rect 10665 -2685 10677 -2651
rect 10277 -2697 10677 -2685
rect 9659 -2909 10059 -2897
rect 9659 -2943 9671 -2909
rect 10047 -2943 10059 -2909
rect 9659 -2955 10059 -2943
rect 10277 -2909 10677 -2897
rect 10277 -2943 10289 -2909
rect 10665 -2943 10677 -2909
rect 10277 -2955 10677 -2943
rect 11259 -1505 11659 -1493
rect 11259 -1539 11271 -1505
rect 11647 -1539 11659 -1505
rect 11259 -1551 11659 -1539
rect 11877 -1505 12277 -1493
rect 11877 -1539 11889 -1505
rect 12265 -1539 12277 -1505
rect 11877 -1551 12277 -1539
rect 11259 -2363 11659 -2351
rect 11259 -2397 11271 -2363
rect 11647 -2397 11659 -2363
rect 11259 -2409 11659 -2397
rect 11877 -2363 12277 -2351
rect 11877 -2397 11889 -2363
rect 12265 -2397 12277 -2363
rect 11877 -2409 12277 -2397
rect 11259 -2651 11659 -2639
rect 11259 -2685 11271 -2651
rect 11647 -2685 11659 -2651
rect 11259 -2697 11659 -2685
rect 11877 -2651 12277 -2639
rect 11877 -2685 11889 -2651
rect 12265 -2685 12277 -2651
rect 11877 -2697 12277 -2685
rect 11259 -2909 11659 -2897
rect 11259 -2943 11271 -2909
rect 11647 -2943 11659 -2909
rect 11259 -2955 11659 -2943
rect 11877 -2909 12277 -2897
rect 11877 -2943 11889 -2909
rect 12265 -2943 12277 -2909
rect 11877 -2955 12277 -2943
rect 12859 -1505 13259 -1493
rect 12859 -1539 12871 -1505
rect 13247 -1539 13259 -1505
rect 12859 -1551 13259 -1539
rect 13477 -1505 13877 -1493
rect 13477 -1539 13489 -1505
rect 13865 -1539 13877 -1505
rect 13477 -1551 13877 -1539
rect 12859 -2363 13259 -2351
rect 12859 -2397 12871 -2363
rect 13247 -2397 13259 -2363
rect 12859 -2409 13259 -2397
rect 13477 -2363 13877 -2351
rect 13477 -2397 13489 -2363
rect 13865 -2397 13877 -2363
rect 13477 -2409 13877 -2397
rect 12859 -2651 13259 -2639
rect 12859 -2685 12871 -2651
rect 13247 -2685 13259 -2651
rect 12859 -2697 13259 -2685
rect 13477 -2651 13877 -2639
rect 13477 -2685 13489 -2651
rect 13865 -2685 13877 -2651
rect 13477 -2697 13877 -2685
rect 12859 -2909 13259 -2897
rect 12859 -2943 12871 -2909
rect 13247 -2943 13259 -2909
rect 12859 -2955 13259 -2943
rect 13477 -2909 13877 -2897
rect 13477 -2943 13489 -2909
rect 13865 -2943 13877 -2909
rect 13477 -2955 13877 -2943
rect 14459 -1505 14859 -1493
rect 14459 -1539 14471 -1505
rect 14847 -1539 14859 -1505
rect 14459 -1551 14859 -1539
rect 15077 -1505 15477 -1493
rect 15077 -1539 15089 -1505
rect 15465 -1539 15477 -1505
rect 15077 -1551 15477 -1539
rect 14459 -2363 14859 -2351
rect 14459 -2397 14471 -2363
rect 14847 -2397 14859 -2363
rect 14459 -2409 14859 -2397
rect 15077 -2363 15477 -2351
rect 15077 -2397 15089 -2363
rect 15465 -2397 15477 -2363
rect 15077 -2409 15477 -2397
rect 14459 -2651 14859 -2639
rect 14459 -2685 14471 -2651
rect 14847 -2685 14859 -2651
rect 14459 -2697 14859 -2685
rect 15077 -2651 15477 -2639
rect 15077 -2685 15089 -2651
rect 15465 -2685 15477 -2651
rect 15077 -2697 15477 -2685
rect 14459 -2909 14859 -2897
rect 14459 -2943 14471 -2909
rect 14847 -2943 14859 -2909
rect 14459 -2955 14859 -2943
rect 15077 -2909 15477 -2897
rect 15077 -2943 15089 -2909
rect 15465 -2943 15477 -2909
rect 15077 -2955 15477 -2943
rect 16059 -1505 16459 -1493
rect 16059 -1539 16071 -1505
rect 16447 -1539 16459 -1505
rect 16059 -1551 16459 -1539
rect 16677 -1505 17077 -1493
rect 16677 -1539 16689 -1505
rect 17065 -1539 17077 -1505
rect 16677 -1551 17077 -1539
rect 16059 -2363 16459 -2351
rect 16059 -2397 16071 -2363
rect 16447 -2397 16459 -2363
rect 16059 -2409 16459 -2397
rect 16677 -2363 17077 -2351
rect 16677 -2397 16689 -2363
rect 17065 -2397 17077 -2363
rect 16677 -2409 17077 -2397
rect 16059 -2651 16459 -2639
rect 16059 -2685 16071 -2651
rect 16447 -2685 16459 -2651
rect 16059 -2697 16459 -2685
rect 16677 -2651 17077 -2639
rect 16677 -2685 16689 -2651
rect 17065 -2685 17077 -2651
rect 16677 -2697 17077 -2685
rect 16059 -2909 16459 -2897
rect 16059 -2943 16071 -2909
rect 16447 -2943 16459 -2909
rect 16059 -2955 16459 -2943
rect 16677 -2909 17077 -2897
rect 16677 -2943 16689 -2909
rect 17065 -2943 17077 -2909
rect 16677 -2955 17077 -2943
rect 17659 -1505 18059 -1493
rect 17659 -1539 17671 -1505
rect 18047 -1539 18059 -1505
rect 17659 -1551 18059 -1539
rect 18277 -1505 18677 -1493
rect 18277 -1539 18289 -1505
rect 18665 -1539 18677 -1505
rect 18277 -1551 18677 -1539
rect 17659 -2363 18059 -2351
rect 17659 -2397 17671 -2363
rect 18047 -2397 18059 -2363
rect 17659 -2409 18059 -2397
rect 18277 -2363 18677 -2351
rect 18277 -2397 18289 -2363
rect 18665 -2397 18677 -2363
rect 18277 -2409 18677 -2397
rect 17659 -2651 18059 -2639
rect 17659 -2685 17671 -2651
rect 18047 -2685 18059 -2651
rect 17659 -2697 18059 -2685
rect 18277 -2651 18677 -2639
rect 18277 -2685 18289 -2651
rect 18665 -2685 18677 -2651
rect 18277 -2697 18677 -2685
rect 17659 -2909 18059 -2897
rect 17659 -2943 17671 -2909
rect 18047 -2943 18059 -2909
rect 17659 -2955 18059 -2943
rect 18277 -2909 18677 -2897
rect 18277 -2943 18289 -2909
rect 18665 -2943 18677 -2909
rect 18277 -2955 18677 -2943
rect 19259 -1505 19659 -1493
rect 19259 -1539 19271 -1505
rect 19647 -1539 19659 -1505
rect 19259 -1551 19659 -1539
rect 19877 -1505 20277 -1493
rect 19877 -1539 19889 -1505
rect 20265 -1539 20277 -1505
rect 19877 -1551 20277 -1539
rect 19259 -2363 19659 -2351
rect 19259 -2397 19271 -2363
rect 19647 -2397 19659 -2363
rect 19259 -2409 19659 -2397
rect 19877 -2363 20277 -2351
rect 19877 -2397 19889 -2363
rect 20265 -2397 20277 -2363
rect 19877 -2409 20277 -2397
rect 19259 -2651 19659 -2639
rect 19259 -2685 19271 -2651
rect 19647 -2685 19659 -2651
rect 19259 -2697 19659 -2685
rect 19877 -2651 20277 -2639
rect 19877 -2685 19889 -2651
rect 20265 -2685 20277 -2651
rect 19877 -2697 20277 -2685
rect 19259 -2909 19659 -2897
rect 19259 -2943 19271 -2909
rect 19647 -2943 19659 -2909
rect 19259 -2955 19659 -2943
rect 19877 -2909 20277 -2897
rect 19877 -2943 19889 -2909
rect 20265 -2943 20277 -2909
rect 19877 -2955 20277 -2943
rect 20859 -1505 21259 -1493
rect 20859 -1539 20871 -1505
rect 21247 -1539 21259 -1505
rect 20859 -1551 21259 -1539
rect 21477 -1505 21877 -1493
rect 21477 -1539 21489 -1505
rect 21865 -1539 21877 -1505
rect 21477 -1551 21877 -1539
rect 20859 -2363 21259 -2351
rect 20859 -2397 20871 -2363
rect 21247 -2397 21259 -2363
rect 20859 -2409 21259 -2397
rect 21477 -2363 21877 -2351
rect 21477 -2397 21489 -2363
rect 21865 -2397 21877 -2363
rect 21477 -2409 21877 -2397
rect 20859 -2651 21259 -2639
rect 20859 -2685 20871 -2651
rect 21247 -2685 21259 -2651
rect 20859 -2697 21259 -2685
rect 21477 -2651 21877 -2639
rect 21477 -2685 21489 -2651
rect 21865 -2685 21877 -2651
rect 21477 -2697 21877 -2685
rect 20859 -2909 21259 -2897
rect 20859 -2943 20871 -2909
rect 21247 -2943 21259 -2909
rect 20859 -2955 21259 -2943
rect 21477 -2909 21877 -2897
rect 21477 -2943 21489 -2909
rect 21865 -2943 21877 -2909
rect 21477 -2955 21877 -2943
rect 22459 -1505 22859 -1493
rect 22459 -1539 22471 -1505
rect 22847 -1539 22859 -1505
rect 22459 -1551 22859 -1539
rect 23077 -1505 23477 -1493
rect 23077 -1539 23089 -1505
rect 23465 -1539 23477 -1505
rect 23077 -1551 23477 -1539
rect 22459 -2363 22859 -2351
rect 22459 -2397 22471 -2363
rect 22847 -2397 22859 -2363
rect 22459 -2409 22859 -2397
rect 23077 -2363 23477 -2351
rect 23077 -2397 23089 -2363
rect 23465 -2397 23477 -2363
rect 23077 -2409 23477 -2397
rect 22459 -2651 22859 -2639
rect 22459 -2685 22471 -2651
rect 22847 -2685 22859 -2651
rect 22459 -2697 22859 -2685
rect 23077 -2651 23477 -2639
rect 23077 -2685 23089 -2651
rect 23465 -2685 23477 -2651
rect 23077 -2697 23477 -2685
rect 22459 -2909 22859 -2897
rect 22459 -2943 22471 -2909
rect 22847 -2943 22859 -2909
rect 22459 -2955 22859 -2943
rect 23077 -2909 23477 -2897
rect 23077 -2943 23089 -2909
rect 23465 -2943 23477 -2909
rect 23077 -2955 23477 -2943
rect 24059 -1505 24459 -1493
rect 24059 -1539 24071 -1505
rect 24447 -1539 24459 -1505
rect 24059 -1551 24459 -1539
rect 24677 -1505 25077 -1493
rect 24677 -1539 24689 -1505
rect 25065 -1539 25077 -1505
rect 24677 -1551 25077 -1539
rect 24059 -2363 24459 -2351
rect 24059 -2397 24071 -2363
rect 24447 -2397 24459 -2363
rect 24059 -2409 24459 -2397
rect 24677 -2363 25077 -2351
rect 24677 -2397 24689 -2363
rect 25065 -2397 25077 -2363
rect 24677 -2409 25077 -2397
rect 24059 -2651 24459 -2639
rect 24059 -2685 24071 -2651
rect 24447 -2685 24459 -2651
rect 24059 -2697 24459 -2685
rect 24677 -2651 25077 -2639
rect 24677 -2685 24689 -2651
rect 25065 -2685 25077 -2651
rect 24677 -2697 25077 -2685
rect 24059 -2909 24459 -2897
rect 24059 -2943 24071 -2909
rect 24447 -2943 24459 -2909
rect 24059 -2955 24459 -2943
rect 24677 -2909 25077 -2897
rect 24677 -2943 24689 -2909
rect 25065 -2943 25077 -2909
rect 24677 -2955 25077 -2943
rect 25659 -1505 26059 -1493
rect 25659 -1539 25671 -1505
rect 26047 -1539 26059 -1505
rect 25659 -1551 26059 -1539
rect 26277 -1505 26677 -1493
rect 26277 -1539 26289 -1505
rect 26665 -1539 26677 -1505
rect 26277 -1551 26677 -1539
rect 25659 -2363 26059 -2351
rect 25659 -2397 25671 -2363
rect 26047 -2397 26059 -2363
rect 25659 -2409 26059 -2397
rect 26277 -2363 26677 -2351
rect 26277 -2397 26289 -2363
rect 26665 -2397 26677 -2363
rect 26277 -2409 26677 -2397
rect 25659 -2651 26059 -2639
rect 25659 -2685 25671 -2651
rect 26047 -2685 26059 -2651
rect 25659 -2697 26059 -2685
rect 26277 -2651 26677 -2639
rect 26277 -2685 26289 -2651
rect 26665 -2685 26677 -2651
rect 26277 -2697 26677 -2685
rect 25659 -2909 26059 -2897
rect 25659 -2943 25671 -2909
rect 26047 -2943 26059 -2909
rect 25659 -2955 26059 -2943
rect 26277 -2909 26677 -2897
rect 26277 -2943 26289 -2909
rect 26665 -2943 26677 -2909
rect 26277 -2955 26677 -2943
rect 27259 -1505 27659 -1493
rect 27259 -1539 27271 -1505
rect 27647 -1539 27659 -1505
rect 27259 -1551 27659 -1539
rect 27877 -1505 28277 -1493
rect 27877 -1539 27889 -1505
rect 28265 -1539 28277 -1505
rect 27877 -1551 28277 -1539
rect 27259 -2363 27659 -2351
rect 27259 -2397 27271 -2363
rect 27647 -2397 27659 -2363
rect 27259 -2409 27659 -2397
rect 27877 -2363 28277 -2351
rect 27877 -2397 27889 -2363
rect 28265 -2397 28277 -2363
rect 27877 -2409 28277 -2397
rect 27259 -2651 27659 -2639
rect 27259 -2685 27271 -2651
rect 27647 -2685 27659 -2651
rect 27259 -2697 27659 -2685
rect 27877 -2651 28277 -2639
rect 27877 -2685 27889 -2651
rect 28265 -2685 28277 -2651
rect 27877 -2697 28277 -2685
rect 27259 -2909 27659 -2897
rect 27259 -2943 27271 -2909
rect 27647 -2943 27659 -2909
rect 27259 -2955 27659 -2943
rect 27877 -2909 28277 -2897
rect 27877 -2943 27889 -2909
rect 28265 -2943 28277 -2909
rect 27877 -2955 28277 -2943
rect 28859 -1505 29259 -1493
rect 28859 -1539 28871 -1505
rect 29247 -1539 29259 -1505
rect 28859 -1551 29259 -1539
rect 29477 -1505 29877 -1493
rect 29477 -1539 29489 -1505
rect 29865 -1539 29877 -1505
rect 29477 -1551 29877 -1539
rect 28859 -2363 29259 -2351
rect 28859 -2397 28871 -2363
rect 29247 -2397 29259 -2363
rect 28859 -2409 29259 -2397
rect 29477 -2363 29877 -2351
rect 29477 -2397 29489 -2363
rect 29865 -2397 29877 -2363
rect 29477 -2409 29877 -2397
rect 28859 -2651 29259 -2639
rect 28859 -2685 28871 -2651
rect 29247 -2685 29259 -2651
rect 28859 -2697 29259 -2685
rect 29477 -2651 29877 -2639
rect 29477 -2685 29489 -2651
rect 29865 -2685 29877 -2651
rect 29477 -2697 29877 -2685
rect 28859 -2909 29259 -2897
rect 28859 -2943 28871 -2909
rect 29247 -2943 29259 -2909
rect 28859 -2955 29259 -2943
rect 29477 -2909 29877 -2897
rect 29477 -2943 29489 -2909
rect 29865 -2943 29877 -2909
rect 29477 -2955 29877 -2943
rect 30459 -1505 30859 -1493
rect 30459 -1539 30471 -1505
rect 30847 -1539 30859 -1505
rect 30459 -1551 30859 -1539
rect 31077 -1505 31477 -1493
rect 31077 -1539 31089 -1505
rect 31465 -1539 31477 -1505
rect 31077 -1551 31477 -1539
rect 30459 -2363 30859 -2351
rect 30459 -2397 30471 -2363
rect 30847 -2397 30859 -2363
rect 30459 -2409 30859 -2397
rect 31077 -2363 31477 -2351
rect 31077 -2397 31089 -2363
rect 31465 -2397 31477 -2363
rect 31077 -2409 31477 -2397
rect 30459 -2651 30859 -2639
rect 30459 -2685 30471 -2651
rect 30847 -2685 30859 -2651
rect 30459 -2697 30859 -2685
rect 31077 -2651 31477 -2639
rect 31077 -2685 31089 -2651
rect 31465 -2685 31477 -2651
rect 31077 -2697 31477 -2685
rect 30459 -2909 30859 -2897
rect 30459 -2943 30471 -2909
rect 30847 -2943 30859 -2909
rect 30459 -2955 30859 -2943
rect 31077 -2909 31477 -2897
rect 31077 -2943 31089 -2909
rect 31465 -2943 31477 -2909
rect 31077 -2955 31477 -2943
rect 32059 -1505 32459 -1493
rect 32059 -1539 32071 -1505
rect 32447 -1539 32459 -1505
rect 32059 -1551 32459 -1539
rect 32677 -1505 33077 -1493
rect 32677 -1539 32689 -1505
rect 33065 -1539 33077 -1505
rect 32677 -1551 33077 -1539
rect 32059 -2363 32459 -2351
rect 32059 -2397 32071 -2363
rect 32447 -2397 32459 -2363
rect 32059 -2409 32459 -2397
rect 32677 -2363 33077 -2351
rect 32677 -2397 32689 -2363
rect 33065 -2397 33077 -2363
rect 32677 -2409 33077 -2397
rect 32059 -2651 32459 -2639
rect 32059 -2685 32071 -2651
rect 32447 -2685 32459 -2651
rect 32059 -2697 32459 -2685
rect 32677 -2651 33077 -2639
rect 32677 -2685 32689 -2651
rect 33065 -2685 33077 -2651
rect 32677 -2697 33077 -2685
rect 32059 -2909 32459 -2897
rect 32059 -2943 32071 -2909
rect 32447 -2943 32459 -2909
rect 32059 -2955 32459 -2943
rect 32677 -2909 33077 -2897
rect 32677 -2943 32689 -2909
rect 33065 -2943 33077 -2909
rect 32677 -2955 33077 -2943
rect 33659 -1505 34059 -1493
rect 33659 -1539 33671 -1505
rect 34047 -1539 34059 -1505
rect 33659 -1551 34059 -1539
rect 34277 -1505 34677 -1493
rect 34277 -1539 34289 -1505
rect 34665 -1539 34677 -1505
rect 34277 -1551 34677 -1539
rect 33659 -2363 34059 -2351
rect 33659 -2397 33671 -2363
rect 34047 -2397 34059 -2363
rect 33659 -2409 34059 -2397
rect 34277 -2363 34677 -2351
rect 34277 -2397 34289 -2363
rect 34665 -2397 34677 -2363
rect 34277 -2409 34677 -2397
rect 33659 -2651 34059 -2639
rect 33659 -2685 33671 -2651
rect 34047 -2685 34059 -2651
rect 33659 -2697 34059 -2685
rect 34277 -2651 34677 -2639
rect 34277 -2685 34289 -2651
rect 34665 -2685 34677 -2651
rect 34277 -2697 34677 -2685
rect 33659 -2909 34059 -2897
rect 33659 -2943 33671 -2909
rect 34047 -2943 34059 -2909
rect 33659 -2955 34059 -2943
rect 34277 -2909 34677 -2897
rect 34277 -2943 34289 -2909
rect 34665 -2943 34677 -2909
rect 34277 -2955 34677 -2943
rect 35259 -1505 35659 -1493
rect 35259 -1539 35271 -1505
rect 35647 -1539 35659 -1505
rect 35259 -1551 35659 -1539
rect 35877 -1505 36277 -1493
rect 35877 -1539 35889 -1505
rect 36265 -1539 36277 -1505
rect 35877 -1551 36277 -1539
rect 35259 -2363 35659 -2351
rect 35259 -2397 35271 -2363
rect 35647 -2397 35659 -2363
rect 35259 -2409 35659 -2397
rect 35877 -2363 36277 -2351
rect 35877 -2397 35889 -2363
rect 36265 -2397 36277 -2363
rect 35877 -2409 36277 -2397
rect 35259 -2651 35659 -2639
rect 35259 -2685 35271 -2651
rect 35647 -2685 35659 -2651
rect 35259 -2697 35659 -2685
rect 35877 -2651 36277 -2639
rect 35877 -2685 35889 -2651
rect 36265 -2685 36277 -2651
rect 35877 -2697 36277 -2685
rect 35259 -2909 35659 -2897
rect 35259 -2943 35271 -2909
rect 35647 -2943 35659 -2909
rect 35259 -2955 35659 -2943
rect 35877 -2909 36277 -2897
rect 35877 -2943 35889 -2909
rect 36265 -2943 36277 -2909
rect 35877 -2955 36277 -2943
rect 36859 -1505 37259 -1493
rect 36859 -1539 36871 -1505
rect 37247 -1539 37259 -1505
rect 36859 -1551 37259 -1539
rect 37477 -1505 37877 -1493
rect 37477 -1539 37489 -1505
rect 37865 -1539 37877 -1505
rect 37477 -1551 37877 -1539
rect 36859 -2363 37259 -2351
rect 36859 -2397 36871 -2363
rect 37247 -2397 37259 -2363
rect 36859 -2409 37259 -2397
rect 37477 -2363 37877 -2351
rect 37477 -2397 37489 -2363
rect 37865 -2397 37877 -2363
rect 37477 -2409 37877 -2397
rect 36859 -2651 37259 -2639
rect 36859 -2685 36871 -2651
rect 37247 -2685 37259 -2651
rect 36859 -2697 37259 -2685
rect 37477 -2651 37877 -2639
rect 37477 -2685 37489 -2651
rect 37865 -2685 37877 -2651
rect 37477 -2697 37877 -2685
rect 36859 -2909 37259 -2897
rect 36859 -2943 36871 -2909
rect 37247 -2943 37259 -2909
rect 36859 -2955 37259 -2943
rect 37477 -2909 37877 -2897
rect 37477 -2943 37489 -2909
rect 37865 -2943 37877 -2909
rect 37477 -2955 37877 -2943
rect 59 -3305 459 -3293
rect 59 -3339 71 -3305
rect 447 -3339 459 -3305
rect 59 -3351 459 -3339
rect 677 -3305 1077 -3293
rect 677 -3339 689 -3305
rect 1065 -3339 1077 -3305
rect 677 -3351 1077 -3339
rect 59 -4163 459 -4151
rect 59 -4197 71 -4163
rect 447 -4197 459 -4163
rect 59 -4209 459 -4197
rect 677 -4163 1077 -4151
rect 677 -4197 689 -4163
rect 1065 -4197 1077 -4163
rect 677 -4209 1077 -4197
rect 59 -4451 459 -4439
rect 59 -4485 71 -4451
rect 447 -4485 459 -4451
rect 59 -4497 459 -4485
rect 677 -4451 1077 -4439
rect 677 -4485 689 -4451
rect 1065 -4485 1077 -4451
rect 677 -4497 1077 -4485
rect 59 -4709 459 -4697
rect 59 -4743 71 -4709
rect 447 -4743 459 -4709
rect 59 -4755 459 -4743
rect 677 -4709 1077 -4697
rect 677 -4743 689 -4709
rect 1065 -4743 1077 -4709
rect 677 -4755 1077 -4743
rect 1659 -3305 2059 -3293
rect 1659 -3339 1671 -3305
rect 2047 -3339 2059 -3305
rect 1659 -3351 2059 -3339
rect 2277 -3305 2677 -3293
rect 2277 -3339 2289 -3305
rect 2665 -3339 2677 -3305
rect 2277 -3351 2677 -3339
rect 1659 -4163 2059 -4151
rect 1659 -4197 1671 -4163
rect 2047 -4197 2059 -4163
rect 1659 -4209 2059 -4197
rect 2277 -4163 2677 -4151
rect 2277 -4197 2289 -4163
rect 2665 -4197 2677 -4163
rect 2277 -4209 2677 -4197
rect 1659 -4451 2059 -4439
rect 1659 -4485 1671 -4451
rect 2047 -4485 2059 -4451
rect 1659 -4497 2059 -4485
rect 2277 -4451 2677 -4439
rect 2277 -4485 2289 -4451
rect 2665 -4485 2677 -4451
rect 2277 -4497 2677 -4485
rect 1659 -4709 2059 -4697
rect 1659 -4743 1671 -4709
rect 2047 -4743 2059 -4709
rect 1659 -4755 2059 -4743
rect 2277 -4709 2677 -4697
rect 2277 -4743 2289 -4709
rect 2665 -4743 2677 -4709
rect 2277 -4755 2677 -4743
rect 3259 -3305 3659 -3293
rect 3259 -3339 3271 -3305
rect 3647 -3339 3659 -3305
rect 3259 -3351 3659 -3339
rect 3877 -3305 4277 -3293
rect 3877 -3339 3889 -3305
rect 4265 -3339 4277 -3305
rect 3877 -3351 4277 -3339
rect 3259 -4163 3659 -4151
rect 3259 -4197 3271 -4163
rect 3647 -4197 3659 -4163
rect 3259 -4209 3659 -4197
rect 3877 -4163 4277 -4151
rect 3877 -4197 3889 -4163
rect 4265 -4197 4277 -4163
rect 3877 -4209 4277 -4197
rect 3259 -4451 3659 -4439
rect 3259 -4485 3271 -4451
rect 3647 -4485 3659 -4451
rect 3259 -4497 3659 -4485
rect 3877 -4451 4277 -4439
rect 3877 -4485 3889 -4451
rect 4265 -4485 4277 -4451
rect 3877 -4497 4277 -4485
rect 3259 -4709 3659 -4697
rect 3259 -4743 3271 -4709
rect 3647 -4743 3659 -4709
rect 3259 -4755 3659 -4743
rect 3877 -4709 4277 -4697
rect 3877 -4743 3889 -4709
rect 4265 -4743 4277 -4709
rect 3877 -4755 4277 -4743
rect 4859 -3305 5259 -3293
rect 4859 -3339 4871 -3305
rect 5247 -3339 5259 -3305
rect 4859 -3351 5259 -3339
rect 5477 -3305 5877 -3293
rect 5477 -3339 5489 -3305
rect 5865 -3339 5877 -3305
rect 5477 -3351 5877 -3339
rect 4859 -4163 5259 -4151
rect 4859 -4197 4871 -4163
rect 5247 -4197 5259 -4163
rect 4859 -4209 5259 -4197
rect 5477 -4163 5877 -4151
rect 5477 -4197 5489 -4163
rect 5865 -4197 5877 -4163
rect 5477 -4209 5877 -4197
rect 4859 -4451 5259 -4439
rect 4859 -4485 4871 -4451
rect 5247 -4485 5259 -4451
rect 4859 -4497 5259 -4485
rect 5477 -4451 5877 -4439
rect 5477 -4485 5489 -4451
rect 5865 -4485 5877 -4451
rect 5477 -4497 5877 -4485
rect 4859 -4709 5259 -4697
rect 4859 -4743 4871 -4709
rect 5247 -4743 5259 -4709
rect 4859 -4755 5259 -4743
rect 5477 -4709 5877 -4697
rect 5477 -4743 5489 -4709
rect 5865 -4743 5877 -4709
rect 5477 -4755 5877 -4743
rect 6459 -3305 6859 -3293
rect 6459 -3339 6471 -3305
rect 6847 -3339 6859 -3305
rect 6459 -3351 6859 -3339
rect 7077 -3305 7477 -3293
rect 7077 -3339 7089 -3305
rect 7465 -3339 7477 -3305
rect 7077 -3351 7477 -3339
rect 6459 -4163 6859 -4151
rect 6459 -4197 6471 -4163
rect 6847 -4197 6859 -4163
rect 6459 -4209 6859 -4197
rect 7077 -4163 7477 -4151
rect 7077 -4197 7089 -4163
rect 7465 -4197 7477 -4163
rect 7077 -4209 7477 -4197
rect 6459 -4451 6859 -4439
rect 6459 -4485 6471 -4451
rect 6847 -4485 6859 -4451
rect 6459 -4497 6859 -4485
rect 7077 -4451 7477 -4439
rect 7077 -4485 7089 -4451
rect 7465 -4485 7477 -4451
rect 7077 -4497 7477 -4485
rect 6459 -4709 6859 -4697
rect 6459 -4743 6471 -4709
rect 6847 -4743 6859 -4709
rect 6459 -4755 6859 -4743
rect 7077 -4709 7477 -4697
rect 7077 -4743 7089 -4709
rect 7465 -4743 7477 -4709
rect 7077 -4755 7477 -4743
rect 8059 -3305 8459 -3293
rect 8059 -3339 8071 -3305
rect 8447 -3339 8459 -3305
rect 8059 -3351 8459 -3339
rect 8677 -3305 9077 -3293
rect 8677 -3339 8689 -3305
rect 9065 -3339 9077 -3305
rect 8677 -3351 9077 -3339
rect 8059 -4163 8459 -4151
rect 8059 -4197 8071 -4163
rect 8447 -4197 8459 -4163
rect 8059 -4209 8459 -4197
rect 8677 -4163 9077 -4151
rect 8677 -4197 8689 -4163
rect 9065 -4197 9077 -4163
rect 8677 -4209 9077 -4197
rect 8059 -4451 8459 -4439
rect 8059 -4485 8071 -4451
rect 8447 -4485 8459 -4451
rect 8059 -4497 8459 -4485
rect 8677 -4451 9077 -4439
rect 8677 -4485 8689 -4451
rect 9065 -4485 9077 -4451
rect 8677 -4497 9077 -4485
rect 8059 -4709 8459 -4697
rect 8059 -4743 8071 -4709
rect 8447 -4743 8459 -4709
rect 8059 -4755 8459 -4743
rect 8677 -4709 9077 -4697
rect 8677 -4743 8689 -4709
rect 9065 -4743 9077 -4709
rect 8677 -4755 9077 -4743
rect 9659 -3305 10059 -3293
rect 9659 -3339 9671 -3305
rect 10047 -3339 10059 -3305
rect 9659 -3351 10059 -3339
rect 10277 -3305 10677 -3293
rect 10277 -3339 10289 -3305
rect 10665 -3339 10677 -3305
rect 10277 -3351 10677 -3339
rect 9659 -4163 10059 -4151
rect 9659 -4197 9671 -4163
rect 10047 -4197 10059 -4163
rect 9659 -4209 10059 -4197
rect 10277 -4163 10677 -4151
rect 10277 -4197 10289 -4163
rect 10665 -4197 10677 -4163
rect 10277 -4209 10677 -4197
rect 9659 -4451 10059 -4439
rect 9659 -4485 9671 -4451
rect 10047 -4485 10059 -4451
rect 9659 -4497 10059 -4485
rect 10277 -4451 10677 -4439
rect 10277 -4485 10289 -4451
rect 10665 -4485 10677 -4451
rect 10277 -4497 10677 -4485
rect 9659 -4709 10059 -4697
rect 9659 -4743 9671 -4709
rect 10047 -4743 10059 -4709
rect 9659 -4755 10059 -4743
rect 10277 -4709 10677 -4697
rect 10277 -4743 10289 -4709
rect 10665 -4743 10677 -4709
rect 10277 -4755 10677 -4743
rect 11259 -3305 11659 -3293
rect 11259 -3339 11271 -3305
rect 11647 -3339 11659 -3305
rect 11259 -3351 11659 -3339
rect 11877 -3305 12277 -3293
rect 11877 -3339 11889 -3305
rect 12265 -3339 12277 -3305
rect 11877 -3351 12277 -3339
rect 11259 -4163 11659 -4151
rect 11259 -4197 11271 -4163
rect 11647 -4197 11659 -4163
rect 11259 -4209 11659 -4197
rect 11877 -4163 12277 -4151
rect 11877 -4197 11889 -4163
rect 12265 -4197 12277 -4163
rect 11877 -4209 12277 -4197
rect 11259 -4451 11659 -4439
rect 11259 -4485 11271 -4451
rect 11647 -4485 11659 -4451
rect 11259 -4497 11659 -4485
rect 11877 -4451 12277 -4439
rect 11877 -4485 11889 -4451
rect 12265 -4485 12277 -4451
rect 11877 -4497 12277 -4485
rect 11259 -4709 11659 -4697
rect 11259 -4743 11271 -4709
rect 11647 -4743 11659 -4709
rect 11259 -4755 11659 -4743
rect 11877 -4709 12277 -4697
rect 11877 -4743 11889 -4709
rect 12265 -4743 12277 -4709
rect 11877 -4755 12277 -4743
rect 12859 -3305 13259 -3293
rect 12859 -3339 12871 -3305
rect 13247 -3339 13259 -3305
rect 12859 -3351 13259 -3339
rect 13477 -3305 13877 -3293
rect 13477 -3339 13489 -3305
rect 13865 -3339 13877 -3305
rect 13477 -3351 13877 -3339
rect 12859 -4163 13259 -4151
rect 12859 -4197 12871 -4163
rect 13247 -4197 13259 -4163
rect 12859 -4209 13259 -4197
rect 13477 -4163 13877 -4151
rect 13477 -4197 13489 -4163
rect 13865 -4197 13877 -4163
rect 13477 -4209 13877 -4197
rect 12859 -4451 13259 -4439
rect 12859 -4485 12871 -4451
rect 13247 -4485 13259 -4451
rect 12859 -4497 13259 -4485
rect 13477 -4451 13877 -4439
rect 13477 -4485 13489 -4451
rect 13865 -4485 13877 -4451
rect 13477 -4497 13877 -4485
rect 12859 -4709 13259 -4697
rect 12859 -4743 12871 -4709
rect 13247 -4743 13259 -4709
rect 12859 -4755 13259 -4743
rect 13477 -4709 13877 -4697
rect 13477 -4743 13489 -4709
rect 13865 -4743 13877 -4709
rect 13477 -4755 13877 -4743
rect 14459 -3305 14859 -3293
rect 14459 -3339 14471 -3305
rect 14847 -3339 14859 -3305
rect 14459 -3351 14859 -3339
rect 15077 -3305 15477 -3293
rect 15077 -3339 15089 -3305
rect 15465 -3339 15477 -3305
rect 15077 -3351 15477 -3339
rect 14459 -4163 14859 -4151
rect 14459 -4197 14471 -4163
rect 14847 -4197 14859 -4163
rect 14459 -4209 14859 -4197
rect 15077 -4163 15477 -4151
rect 15077 -4197 15089 -4163
rect 15465 -4197 15477 -4163
rect 15077 -4209 15477 -4197
rect 14459 -4451 14859 -4439
rect 14459 -4485 14471 -4451
rect 14847 -4485 14859 -4451
rect 14459 -4497 14859 -4485
rect 15077 -4451 15477 -4439
rect 15077 -4485 15089 -4451
rect 15465 -4485 15477 -4451
rect 15077 -4497 15477 -4485
rect 14459 -4709 14859 -4697
rect 14459 -4743 14471 -4709
rect 14847 -4743 14859 -4709
rect 14459 -4755 14859 -4743
rect 15077 -4709 15477 -4697
rect 15077 -4743 15089 -4709
rect 15465 -4743 15477 -4709
rect 15077 -4755 15477 -4743
rect 16059 -3305 16459 -3293
rect 16059 -3339 16071 -3305
rect 16447 -3339 16459 -3305
rect 16059 -3351 16459 -3339
rect 16677 -3305 17077 -3293
rect 16677 -3339 16689 -3305
rect 17065 -3339 17077 -3305
rect 16677 -3351 17077 -3339
rect 16059 -4163 16459 -4151
rect 16059 -4197 16071 -4163
rect 16447 -4197 16459 -4163
rect 16059 -4209 16459 -4197
rect 16677 -4163 17077 -4151
rect 16677 -4197 16689 -4163
rect 17065 -4197 17077 -4163
rect 16677 -4209 17077 -4197
rect 16059 -4451 16459 -4439
rect 16059 -4485 16071 -4451
rect 16447 -4485 16459 -4451
rect 16059 -4497 16459 -4485
rect 16677 -4451 17077 -4439
rect 16677 -4485 16689 -4451
rect 17065 -4485 17077 -4451
rect 16677 -4497 17077 -4485
rect 16059 -4709 16459 -4697
rect 16059 -4743 16071 -4709
rect 16447 -4743 16459 -4709
rect 16059 -4755 16459 -4743
rect 16677 -4709 17077 -4697
rect 16677 -4743 16689 -4709
rect 17065 -4743 17077 -4709
rect 16677 -4755 17077 -4743
rect 17659 -3305 18059 -3293
rect 17659 -3339 17671 -3305
rect 18047 -3339 18059 -3305
rect 17659 -3351 18059 -3339
rect 18277 -3305 18677 -3293
rect 18277 -3339 18289 -3305
rect 18665 -3339 18677 -3305
rect 18277 -3351 18677 -3339
rect 17659 -4163 18059 -4151
rect 17659 -4197 17671 -4163
rect 18047 -4197 18059 -4163
rect 17659 -4209 18059 -4197
rect 18277 -4163 18677 -4151
rect 18277 -4197 18289 -4163
rect 18665 -4197 18677 -4163
rect 18277 -4209 18677 -4197
rect 17659 -4451 18059 -4439
rect 17659 -4485 17671 -4451
rect 18047 -4485 18059 -4451
rect 17659 -4497 18059 -4485
rect 18277 -4451 18677 -4439
rect 18277 -4485 18289 -4451
rect 18665 -4485 18677 -4451
rect 18277 -4497 18677 -4485
rect 17659 -4709 18059 -4697
rect 17659 -4743 17671 -4709
rect 18047 -4743 18059 -4709
rect 17659 -4755 18059 -4743
rect 18277 -4709 18677 -4697
rect 18277 -4743 18289 -4709
rect 18665 -4743 18677 -4709
rect 18277 -4755 18677 -4743
rect 19259 -3305 19659 -3293
rect 19259 -3339 19271 -3305
rect 19647 -3339 19659 -3305
rect 19259 -3351 19659 -3339
rect 19877 -3305 20277 -3293
rect 19877 -3339 19889 -3305
rect 20265 -3339 20277 -3305
rect 19877 -3351 20277 -3339
rect 19259 -4163 19659 -4151
rect 19259 -4197 19271 -4163
rect 19647 -4197 19659 -4163
rect 19259 -4209 19659 -4197
rect 19877 -4163 20277 -4151
rect 19877 -4197 19889 -4163
rect 20265 -4197 20277 -4163
rect 19877 -4209 20277 -4197
rect 19259 -4451 19659 -4439
rect 19259 -4485 19271 -4451
rect 19647 -4485 19659 -4451
rect 19259 -4497 19659 -4485
rect 19877 -4451 20277 -4439
rect 19877 -4485 19889 -4451
rect 20265 -4485 20277 -4451
rect 19877 -4497 20277 -4485
rect 19259 -4709 19659 -4697
rect 19259 -4743 19271 -4709
rect 19647 -4743 19659 -4709
rect 19259 -4755 19659 -4743
rect 19877 -4709 20277 -4697
rect 19877 -4743 19889 -4709
rect 20265 -4743 20277 -4709
rect 19877 -4755 20277 -4743
rect 20859 -3305 21259 -3293
rect 20859 -3339 20871 -3305
rect 21247 -3339 21259 -3305
rect 20859 -3351 21259 -3339
rect 21477 -3305 21877 -3293
rect 21477 -3339 21489 -3305
rect 21865 -3339 21877 -3305
rect 21477 -3351 21877 -3339
rect 20859 -4163 21259 -4151
rect 20859 -4197 20871 -4163
rect 21247 -4197 21259 -4163
rect 20859 -4209 21259 -4197
rect 21477 -4163 21877 -4151
rect 21477 -4197 21489 -4163
rect 21865 -4197 21877 -4163
rect 21477 -4209 21877 -4197
rect 20859 -4451 21259 -4439
rect 20859 -4485 20871 -4451
rect 21247 -4485 21259 -4451
rect 20859 -4497 21259 -4485
rect 21477 -4451 21877 -4439
rect 21477 -4485 21489 -4451
rect 21865 -4485 21877 -4451
rect 21477 -4497 21877 -4485
rect 20859 -4709 21259 -4697
rect 20859 -4743 20871 -4709
rect 21247 -4743 21259 -4709
rect 20859 -4755 21259 -4743
rect 21477 -4709 21877 -4697
rect 21477 -4743 21489 -4709
rect 21865 -4743 21877 -4709
rect 21477 -4755 21877 -4743
rect 22459 -3305 22859 -3293
rect 22459 -3339 22471 -3305
rect 22847 -3339 22859 -3305
rect 22459 -3351 22859 -3339
rect 23077 -3305 23477 -3293
rect 23077 -3339 23089 -3305
rect 23465 -3339 23477 -3305
rect 23077 -3351 23477 -3339
rect 22459 -4163 22859 -4151
rect 22459 -4197 22471 -4163
rect 22847 -4197 22859 -4163
rect 22459 -4209 22859 -4197
rect 23077 -4163 23477 -4151
rect 23077 -4197 23089 -4163
rect 23465 -4197 23477 -4163
rect 23077 -4209 23477 -4197
rect 22459 -4451 22859 -4439
rect 22459 -4485 22471 -4451
rect 22847 -4485 22859 -4451
rect 22459 -4497 22859 -4485
rect 23077 -4451 23477 -4439
rect 23077 -4485 23089 -4451
rect 23465 -4485 23477 -4451
rect 23077 -4497 23477 -4485
rect 22459 -4709 22859 -4697
rect 22459 -4743 22471 -4709
rect 22847 -4743 22859 -4709
rect 22459 -4755 22859 -4743
rect 23077 -4709 23477 -4697
rect 23077 -4743 23089 -4709
rect 23465 -4743 23477 -4709
rect 23077 -4755 23477 -4743
rect 24059 -3305 24459 -3293
rect 24059 -3339 24071 -3305
rect 24447 -3339 24459 -3305
rect 24059 -3351 24459 -3339
rect 24677 -3305 25077 -3293
rect 24677 -3339 24689 -3305
rect 25065 -3339 25077 -3305
rect 24677 -3351 25077 -3339
rect 24059 -4163 24459 -4151
rect 24059 -4197 24071 -4163
rect 24447 -4197 24459 -4163
rect 24059 -4209 24459 -4197
rect 24677 -4163 25077 -4151
rect 24677 -4197 24689 -4163
rect 25065 -4197 25077 -4163
rect 24677 -4209 25077 -4197
rect 24059 -4451 24459 -4439
rect 24059 -4485 24071 -4451
rect 24447 -4485 24459 -4451
rect 24059 -4497 24459 -4485
rect 24677 -4451 25077 -4439
rect 24677 -4485 24689 -4451
rect 25065 -4485 25077 -4451
rect 24677 -4497 25077 -4485
rect 24059 -4709 24459 -4697
rect 24059 -4743 24071 -4709
rect 24447 -4743 24459 -4709
rect 24059 -4755 24459 -4743
rect 24677 -4709 25077 -4697
rect 24677 -4743 24689 -4709
rect 25065 -4743 25077 -4709
rect 24677 -4755 25077 -4743
rect 25659 -3305 26059 -3293
rect 25659 -3339 25671 -3305
rect 26047 -3339 26059 -3305
rect 25659 -3351 26059 -3339
rect 26277 -3305 26677 -3293
rect 26277 -3339 26289 -3305
rect 26665 -3339 26677 -3305
rect 26277 -3351 26677 -3339
rect 25659 -4163 26059 -4151
rect 25659 -4197 25671 -4163
rect 26047 -4197 26059 -4163
rect 25659 -4209 26059 -4197
rect 26277 -4163 26677 -4151
rect 26277 -4197 26289 -4163
rect 26665 -4197 26677 -4163
rect 26277 -4209 26677 -4197
rect 25659 -4451 26059 -4439
rect 25659 -4485 25671 -4451
rect 26047 -4485 26059 -4451
rect 25659 -4497 26059 -4485
rect 26277 -4451 26677 -4439
rect 26277 -4485 26289 -4451
rect 26665 -4485 26677 -4451
rect 26277 -4497 26677 -4485
rect 25659 -4709 26059 -4697
rect 25659 -4743 25671 -4709
rect 26047 -4743 26059 -4709
rect 25659 -4755 26059 -4743
rect 26277 -4709 26677 -4697
rect 26277 -4743 26289 -4709
rect 26665 -4743 26677 -4709
rect 26277 -4755 26677 -4743
rect 27259 -3305 27659 -3293
rect 27259 -3339 27271 -3305
rect 27647 -3339 27659 -3305
rect 27259 -3351 27659 -3339
rect 27877 -3305 28277 -3293
rect 27877 -3339 27889 -3305
rect 28265 -3339 28277 -3305
rect 27877 -3351 28277 -3339
rect 27259 -4163 27659 -4151
rect 27259 -4197 27271 -4163
rect 27647 -4197 27659 -4163
rect 27259 -4209 27659 -4197
rect 27877 -4163 28277 -4151
rect 27877 -4197 27889 -4163
rect 28265 -4197 28277 -4163
rect 27877 -4209 28277 -4197
rect 27259 -4451 27659 -4439
rect 27259 -4485 27271 -4451
rect 27647 -4485 27659 -4451
rect 27259 -4497 27659 -4485
rect 27877 -4451 28277 -4439
rect 27877 -4485 27889 -4451
rect 28265 -4485 28277 -4451
rect 27877 -4497 28277 -4485
rect 27259 -4709 27659 -4697
rect 27259 -4743 27271 -4709
rect 27647 -4743 27659 -4709
rect 27259 -4755 27659 -4743
rect 27877 -4709 28277 -4697
rect 27877 -4743 27889 -4709
rect 28265 -4743 28277 -4709
rect 27877 -4755 28277 -4743
rect 28859 -3305 29259 -3293
rect 28859 -3339 28871 -3305
rect 29247 -3339 29259 -3305
rect 28859 -3351 29259 -3339
rect 29477 -3305 29877 -3293
rect 29477 -3339 29489 -3305
rect 29865 -3339 29877 -3305
rect 29477 -3351 29877 -3339
rect 28859 -4163 29259 -4151
rect 28859 -4197 28871 -4163
rect 29247 -4197 29259 -4163
rect 28859 -4209 29259 -4197
rect 29477 -4163 29877 -4151
rect 29477 -4197 29489 -4163
rect 29865 -4197 29877 -4163
rect 29477 -4209 29877 -4197
rect 28859 -4451 29259 -4439
rect 28859 -4485 28871 -4451
rect 29247 -4485 29259 -4451
rect 28859 -4497 29259 -4485
rect 29477 -4451 29877 -4439
rect 29477 -4485 29489 -4451
rect 29865 -4485 29877 -4451
rect 29477 -4497 29877 -4485
rect 28859 -4709 29259 -4697
rect 28859 -4743 28871 -4709
rect 29247 -4743 29259 -4709
rect 28859 -4755 29259 -4743
rect 29477 -4709 29877 -4697
rect 29477 -4743 29489 -4709
rect 29865 -4743 29877 -4709
rect 29477 -4755 29877 -4743
rect 30459 -3305 30859 -3293
rect 30459 -3339 30471 -3305
rect 30847 -3339 30859 -3305
rect 30459 -3351 30859 -3339
rect 31077 -3305 31477 -3293
rect 31077 -3339 31089 -3305
rect 31465 -3339 31477 -3305
rect 31077 -3351 31477 -3339
rect 30459 -4163 30859 -4151
rect 30459 -4197 30471 -4163
rect 30847 -4197 30859 -4163
rect 30459 -4209 30859 -4197
rect 31077 -4163 31477 -4151
rect 31077 -4197 31089 -4163
rect 31465 -4197 31477 -4163
rect 31077 -4209 31477 -4197
rect 30459 -4451 30859 -4439
rect 30459 -4485 30471 -4451
rect 30847 -4485 30859 -4451
rect 30459 -4497 30859 -4485
rect 31077 -4451 31477 -4439
rect 31077 -4485 31089 -4451
rect 31465 -4485 31477 -4451
rect 31077 -4497 31477 -4485
rect 30459 -4709 30859 -4697
rect 30459 -4743 30471 -4709
rect 30847 -4743 30859 -4709
rect 30459 -4755 30859 -4743
rect 31077 -4709 31477 -4697
rect 31077 -4743 31089 -4709
rect 31465 -4743 31477 -4709
rect 31077 -4755 31477 -4743
rect 32059 -3305 32459 -3293
rect 32059 -3339 32071 -3305
rect 32447 -3339 32459 -3305
rect 32059 -3351 32459 -3339
rect 32677 -3305 33077 -3293
rect 32677 -3339 32689 -3305
rect 33065 -3339 33077 -3305
rect 32677 -3351 33077 -3339
rect 32059 -4163 32459 -4151
rect 32059 -4197 32071 -4163
rect 32447 -4197 32459 -4163
rect 32059 -4209 32459 -4197
rect 32677 -4163 33077 -4151
rect 32677 -4197 32689 -4163
rect 33065 -4197 33077 -4163
rect 32677 -4209 33077 -4197
rect 32059 -4451 32459 -4439
rect 32059 -4485 32071 -4451
rect 32447 -4485 32459 -4451
rect 32059 -4497 32459 -4485
rect 32677 -4451 33077 -4439
rect 32677 -4485 32689 -4451
rect 33065 -4485 33077 -4451
rect 32677 -4497 33077 -4485
rect 32059 -4709 32459 -4697
rect 32059 -4743 32071 -4709
rect 32447 -4743 32459 -4709
rect 32059 -4755 32459 -4743
rect 32677 -4709 33077 -4697
rect 32677 -4743 32689 -4709
rect 33065 -4743 33077 -4709
rect 32677 -4755 33077 -4743
rect 33659 -3305 34059 -3293
rect 33659 -3339 33671 -3305
rect 34047 -3339 34059 -3305
rect 33659 -3351 34059 -3339
rect 34277 -3305 34677 -3293
rect 34277 -3339 34289 -3305
rect 34665 -3339 34677 -3305
rect 34277 -3351 34677 -3339
rect 33659 -4163 34059 -4151
rect 33659 -4197 33671 -4163
rect 34047 -4197 34059 -4163
rect 33659 -4209 34059 -4197
rect 34277 -4163 34677 -4151
rect 34277 -4197 34289 -4163
rect 34665 -4197 34677 -4163
rect 34277 -4209 34677 -4197
rect 33659 -4451 34059 -4439
rect 33659 -4485 33671 -4451
rect 34047 -4485 34059 -4451
rect 33659 -4497 34059 -4485
rect 34277 -4451 34677 -4439
rect 34277 -4485 34289 -4451
rect 34665 -4485 34677 -4451
rect 34277 -4497 34677 -4485
rect 33659 -4709 34059 -4697
rect 33659 -4743 33671 -4709
rect 34047 -4743 34059 -4709
rect 33659 -4755 34059 -4743
rect 34277 -4709 34677 -4697
rect 34277 -4743 34289 -4709
rect 34665 -4743 34677 -4709
rect 34277 -4755 34677 -4743
rect 35259 -3305 35659 -3293
rect 35259 -3339 35271 -3305
rect 35647 -3339 35659 -3305
rect 35259 -3351 35659 -3339
rect 35877 -3305 36277 -3293
rect 35877 -3339 35889 -3305
rect 36265 -3339 36277 -3305
rect 35877 -3351 36277 -3339
rect 35259 -4163 35659 -4151
rect 35259 -4197 35271 -4163
rect 35647 -4197 35659 -4163
rect 35259 -4209 35659 -4197
rect 35877 -4163 36277 -4151
rect 35877 -4197 35889 -4163
rect 36265 -4197 36277 -4163
rect 35877 -4209 36277 -4197
rect 35259 -4451 35659 -4439
rect 35259 -4485 35271 -4451
rect 35647 -4485 35659 -4451
rect 35259 -4497 35659 -4485
rect 35877 -4451 36277 -4439
rect 35877 -4485 35889 -4451
rect 36265 -4485 36277 -4451
rect 35877 -4497 36277 -4485
rect 35259 -4709 35659 -4697
rect 35259 -4743 35271 -4709
rect 35647 -4743 35659 -4709
rect 35259 -4755 35659 -4743
rect 35877 -4709 36277 -4697
rect 35877 -4743 35889 -4709
rect 36265 -4743 36277 -4709
rect 35877 -4755 36277 -4743
rect 36859 -3305 37259 -3293
rect 36859 -3339 36871 -3305
rect 37247 -3339 37259 -3305
rect 36859 -3351 37259 -3339
rect 37477 -3305 37877 -3293
rect 37477 -3339 37489 -3305
rect 37865 -3339 37877 -3305
rect 37477 -3351 37877 -3339
rect 36859 -4163 37259 -4151
rect 36859 -4197 36871 -4163
rect 37247 -4197 37259 -4163
rect 36859 -4209 37259 -4197
rect 37477 -4163 37877 -4151
rect 37477 -4197 37489 -4163
rect 37865 -4197 37877 -4163
rect 37477 -4209 37877 -4197
rect 36859 -4451 37259 -4439
rect 36859 -4485 36871 -4451
rect 37247 -4485 37259 -4451
rect 36859 -4497 37259 -4485
rect 37477 -4451 37877 -4439
rect 37477 -4485 37489 -4451
rect 37865 -4485 37877 -4451
rect 37477 -4497 37877 -4485
rect 36859 -4709 37259 -4697
rect 36859 -4743 36871 -4709
rect 37247 -4743 37259 -4709
rect 36859 -4755 37259 -4743
rect 37477 -4709 37877 -4697
rect 37477 -4743 37489 -4709
rect 37865 -4743 37877 -4709
rect 37477 -4755 37877 -4743
rect 27910 -24724 27968 -24712
rect 27910 -25100 27922 -24724
rect 27956 -25100 27968 -24724
rect 27910 -25112 27968 -25100
rect 28768 -24724 28826 -24712
rect 28768 -25100 28780 -24724
rect 28814 -25100 28826 -24724
rect 28768 -25112 28826 -25100
rect 27936 -25542 28736 -25530
rect 27936 -25576 27948 -25542
rect 28724 -25576 28736 -25542
rect 27936 -25588 28736 -25576
rect 27936 -25700 28736 -25688
rect 27936 -25734 27948 -25700
rect 28724 -25734 28736 -25700
rect 27936 -25746 28736 -25734
rect 27936 -25858 28736 -25846
rect 27936 -25892 27948 -25858
rect 28724 -25892 28736 -25858
rect 27936 -25904 28736 -25892
rect 27936 -26016 28736 -26004
rect 27936 -26050 27948 -26016
rect 28724 -26050 28736 -26016
rect 27936 -26062 28736 -26050
rect 27936 -26174 28736 -26162
rect 27936 -26208 27948 -26174
rect 28724 -26208 28736 -26174
rect 27936 -26220 28736 -26208
rect 27936 -26582 28736 -26570
rect 27936 -26616 27948 -26582
rect 28724 -26616 28736 -26582
rect 27936 -26628 28736 -26616
rect 27936 -26740 28736 -26728
rect 27936 -26774 27948 -26740
rect 28724 -26774 28736 -26740
rect 27936 -26786 28736 -26774
rect 27936 -26898 28736 -26886
rect 27936 -26932 27948 -26898
rect 28724 -26932 28736 -26898
rect 27936 -26944 28736 -26932
rect 27936 -27056 28736 -27044
rect 27936 -27090 27948 -27056
rect 28724 -27090 28736 -27056
rect 27936 -27102 28736 -27090
rect 27936 -27214 28736 -27202
rect 27936 -27248 27948 -27214
rect 28724 -27248 28736 -27214
rect 27936 -27260 28736 -27248
rect 27936 -27622 28736 -27610
rect 27936 -27656 27948 -27622
rect 28724 -27656 28736 -27622
rect 27936 -27668 28736 -27656
rect 27936 -27780 28736 -27768
rect 27936 -27814 27948 -27780
rect 28724 -27814 28736 -27780
rect 27936 -27826 28736 -27814
rect 27936 -27938 28736 -27926
rect 27936 -27972 27948 -27938
rect 28724 -27972 28736 -27938
rect 27936 -27984 28736 -27972
rect 27936 -28096 28736 -28084
rect 27936 -28130 27948 -28096
rect 28724 -28130 28736 -28096
rect 27936 -28142 28736 -28130
rect 27936 -28254 28736 -28242
rect 27936 -28288 27948 -28254
rect 28724 -28288 28736 -28254
rect 27936 -28300 28736 -28288
rect 27936 -28662 28736 -28650
rect 27936 -28696 27948 -28662
rect 28724 -28696 28736 -28662
rect 27936 -28708 28736 -28696
rect 27936 -28820 28736 -28808
rect 27936 -28854 27948 -28820
rect 28724 -28854 28736 -28820
rect 27936 -28866 28736 -28854
rect 27936 -28978 28736 -28966
rect 27936 -29012 27948 -28978
rect 28724 -29012 28736 -28978
rect 27936 -29024 28736 -29012
rect 27936 -29136 28736 -29124
rect 27936 -29170 27948 -29136
rect 28724 -29170 28736 -29136
rect 27936 -29182 28736 -29170
rect 27936 -29294 28736 -29282
rect 27936 -29328 27948 -29294
rect 28724 -29328 28736 -29294
rect 27936 -29340 28736 -29328
rect 27936 -29702 28736 -29690
rect 27936 -29736 27948 -29702
rect 28724 -29736 28736 -29702
rect 27936 -29748 28736 -29736
rect 27936 -29860 28736 -29848
rect 27936 -29894 27948 -29860
rect 28724 -29894 28736 -29860
rect 27936 -29906 28736 -29894
rect 27936 -30018 28736 -30006
rect 27936 -30052 27948 -30018
rect 28724 -30052 28736 -30018
rect 27936 -30064 28736 -30052
rect 27936 -30176 28736 -30164
rect 27936 -30210 27948 -30176
rect 28724 -30210 28736 -30176
rect 27936 -30222 28736 -30210
rect 27936 -30334 28736 -30322
rect 27936 -30368 27948 -30334
rect 28724 -30368 28736 -30334
rect 27936 -30380 28736 -30368
rect 31801 -29553 31859 -29541
rect 31801 -29729 31813 -29553
rect 31847 -29729 31859 -29553
rect 31801 -29741 31859 -29729
rect 31959 -29553 32017 -29541
rect 31959 -29729 31971 -29553
rect 32005 -29729 32017 -29553
rect 31959 -29741 32017 -29729
rect 32241 -29553 32299 -29541
rect 32241 -29729 32253 -29553
rect 32287 -29729 32299 -29553
rect 32241 -29741 32299 -29729
rect 32399 -29553 32457 -29541
rect 32399 -29729 32411 -29553
rect 32445 -29729 32457 -29553
rect 32399 -29741 32457 -29729
rect 32681 -29553 32739 -29541
rect 32681 -29729 32693 -29553
rect 32727 -29729 32739 -29553
rect 32681 -29741 32739 -29729
rect 32839 -29553 32897 -29541
rect 32839 -29729 32851 -29553
rect 32885 -29729 32897 -29553
rect 32839 -29741 32897 -29729
rect 33120 -29553 33178 -29541
rect 33120 -29729 33132 -29553
rect 33166 -29729 33178 -29553
rect 33120 -29741 33178 -29729
rect 33278 -29553 33336 -29541
rect 33278 -29729 33290 -29553
rect 33324 -29729 33336 -29553
rect 33278 -29741 33336 -29729
rect 33436 -29553 33494 -29541
rect 33436 -29729 33448 -29553
rect 33482 -29729 33494 -29553
rect 33436 -29741 33494 -29729
rect 33594 -29553 33652 -29541
rect 33594 -29729 33606 -29553
rect 33640 -29729 33652 -29553
rect 33594 -29741 33652 -29729
rect 34001 -29553 34059 -29541
rect 34001 -29729 34013 -29553
rect 34047 -29729 34059 -29553
rect 34001 -29741 34059 -29729
rect 34159 -29553 34217 -29541
rect 34159 -29729 34171 -29553
rect 34205 -29729 34217 -29553
rect 34159 -29741 34217 -29729
rect 34441 -29553 34499 -29541
rect 34441 -29729 34453 -29553
rect 34487 -29729 34499 -29553
rect 34441 -29741 34499 -29729
rect 34599 -29553 34657 -29541
rect 34599 -29729 34611 -29553
rect 34645 -29729 34657 -29553
rect 34599 -29741 34657 -29729
rect 34881 -29553 34939 -29541
rect 34881 -29729 34893 -29553
rect 34927 -29729 34939 -29553
rect 34881 -29741 34939 -29729
rect 35039 -29553 35097 -29541
rect 35039 -29729 35051 -29553
rect 35085 -29729 35097 -29553
rect 35039 -29741 35097 -29729
rect 35320 -29553 35378 -29541
rect 35320 -29729 35332 -29553
rect 35366 -29729 35378 -29553
rect 35320 -29741 35378 -29729
rect 35478 -29553 35536 -29541
rect 35478 -29729 35490 -29553
rect 35524 -29729 35536 -29553
rect 35478 -29741 35536 -29729
rect 35636 -29553 35694 -29541
rect 35636 -29729 35648 -29553
rect 35682 -29729 35694 -29553
rect 35636 -29741 35694 -29729
rect 35794 -29553 35852 -29541
rect 35794 -29729 35806 -29553
rect 35840 -29729 35852 -29553
rect 35794 -29741 35852 -29729
rect 36201 -29553 36259 -29541
rect 36201 -29729 36213 -29553
rect 36247 -29729 36259 -29553
rect 36201 -29741 36259 -29729
rect 36359 -29553 36417 -29541
rect 36359 -29729 36371 -29553
rect 36405 -29729 36417 -29553
rect 36359 -29741 36417 -29729
rect 36641 -29553 36699 -29541
rect 36641 -29729 36653 -29553
rect 36687 -29729 36699 -29553
rect 36641 -29741 36699 -29729
rect 36799 -29553 36857 -29541
rect 36799 -29729 36811 -29553
rect 36845 -29729 36857 -29553
rect 36799 -29741 36857 -29729
rect 37081 -29553 37139 -29541
rect 37081 -29729 37093 -29553
rect 37127 -29729 37139 -29553
rect 37081 -29741 37139 -29729
rect 37239 -29553 37297 -29541
rect 37239 -29729 37251 -29553
rect 37285 -29729 37297 -29553
rect 37239 -29741 37297 -29729
rect 37520 -29553 37578 -29541
rect 37520 -29729 37532 -29553
rect 37566 -29729 37578 -29553
rect 37520 -29741 37578 -29729
rect 37678 -29553 37736 -29541
rect 37678 -29729 37690 -29553
rect 37724 -29729 37736 -29553
rect 37678 -29741 37736 -29729
rect 37836 -29553 37894 -29541
rect 37836 -29729 37848 -29553
rect 37882 -29729 37894 -29553
rect 37836 -29741 37894 -29729
rect 37994 -29553 38052 -29541
rect 37994 -29729 38006 -29553
rect 38040 -29729 38052 -29553
rect 37994 -29741 38052 -29729
rect 27936 -30742 28736 -30730
rect 27936 -30776 27948 -30742
rect 28724 -30776 28736 -30742
rect 27936 -30788 28736 -30776
rect 27936 -30900 28736 -30888
rect 27936 -30934 27948 -30900
rect 28724 -30934 28736 -30900
rect 27936 -30946 28736 -30934
rect 27936 -31058 28736 -31046
rect 27936 -31092 27948 -31058
rect 28724 -31092 28736 -31058
rect 27936 -31104 28736 -31092
rect 27936 -31216 28736 -31204
rect 27936 -31250 27948 -31216
rect 28724 -31250 28736 -31216
rect 27936 -31262 28736 -31250
rect 27936 -31374 28736 -31362
rect 27936 -31408 27948 -31374
rect 28724 -31408 28736 -31374
rect 27936 -31420 28736 -31408
rect 31770 -30295 31828 -30283
rect 31770 -30471 31782 -30295
rect 31816 -30471 31828 -30295
rect 31770 -30483 31828 -30471
rect 31928 -30295 31986 -30283
rect 31928 -30471 31940 -30295
rect 31974 -30471 31986 -30295
rect 31928 -30483 31986 -30471
rect 32086 -30295 32144 -30283
rect 32086 -30471 32098 -30295
rect 32132 -30471 32144 -30295
rect 32086 -30483 32144 -30471
rect 32244 -30295 32302 -30283
rect 32244 -30471 32256 -30295
rect 32290 -30471 32302 -30295
rect 32244 -30483 32302 -30471
rect 32525 -30295 32583 -30283
rect 32525 -30471 32537 -30295
rect 32571 -30471 32583 -30295
rect 32525 -30483 32583 -30471
rect 32683 -30295 32741 -30283
rect 32683 -30471 32695 -30295
rect 32729 -30471 32741 -30295
rect 32683 -30483 32741 -30471
rect 32965 -30295 33023 -30283
rect 32965 -30471 32977 -30295
rect 33011 -30471 33023 -30295
rect 32965 -30483 33023 -30471
rect 33123 -30295 33181 -30283
rect 33123 -30471 33135 -30295
rect 33169 -30471 33181 -30295
rect 33123 -30483 33181 -30471
rect 33405 -30295 33463 -30283
rect 33405 -30471 33417 -30295
rect 33451 -30471 33463 -30295
rect 33405 -30483 33463 -30471
rect 33563 -30295 33621 -30283
rect 33563 -30471 33575 -30295
rect 33609 -30471 33621 -30295
rect 33563 -30483 33621 -30471
rect 33970 -30295 34028 -30283
rect 33970 -30471 33982 -30295
rect 34016 -30471 34028 -30295
rect 33970 -30483 34028 -30471
rect 34128 -30295 34186 -30283
rect 34128 -30471 34140 -30295
rect 34174 -30471 34186 -30295
rect 34128 -30483 34186 -30471
rect 34286 -30295 34344 -30283
rect 34286 -30471 34298 -30295
rect 34332 -30471 34344 -30295
rect 34286 -30483 34344 -30471
rect 34444 -30295 34502 -30283
rect 34444 -30471 34456 -30295
rect 34490 -30471 34502 -30295
rect 34444 -30483 34502 -30471
rect 34725 -30295 34783 -30283
rect 34725 -30471 34737 -30295
rect 34771 -30471 34783 -30295
rect 34725 -30483 34783 -30471
rect 34883 -30295 34941 -30283
rect 34883 -30471 34895 -30295
rect 34929 -30471 34941 -30295
rect 34883 -30483 34941 -30471
rect 35165 -30295 35223 -30283
rect 35165 -30471 35177 -30295
rect 35211 -30471 35223 -30295
rect 35165 -30483 35223 -30471
rect 35323 -30295 35381 -30283
rect 35323 -30471 35335 -30295
rect 35369 -30471 35381 -30295
rect 35323 -30483 35381 -30471
rect 35605 -30295 35663 -30283
rect 35605 -30471 35617 -30295
rect 35651 -30471 35663 -30295
rect 35605 -30483 35663 -30471
rect 35763 -30295 35821 -30283
rect 35763 -30471 35775 -30295
rect 35809 -30471 35821 -30295
rect 35763 -30483 35821 -30471
rect 36170 -30295 36228 -30283
rect 36170 -30471 36182 -30295
rect 36216 -30471 36228 -30295
rect 36170 -30483 36228 -30471
rect 36328 -30295 36386 -30283
rect 36328 -30471 36340 -30295
rect 36374 -30471 36386 -30295
rect 36328 -30483 36386 -30471
rect 36486 -30295 36544 -30283
rect 36486 -30471 36498 -30295
rect 36532 -30471 36544 -30295
rect 36486 -30483 36544 -30471
rect 36644 -30295 36702 -30283
rect 36644 -30471 36656 -30295
rect 36690 -30471 36702 -30295
rect 36644 -30483 36702 -30471
rect 36925 -30295 36983 -30283
rect 36925 -30471 36937 -30295
rect 36971 -30471 36983 -30295
rect 36925 -30483 36983 -30471
rect 37083 -30295 37141 -30283
rect 37083 -30471 37095 -30295
rect 37129 -30471 37141 -30295
rect 37083 -30483 37141 -30471
rect 37365 -30295 37423 -30283
rect 37365 -30471 37377 -30295
rect 37411 -30471 37423 -30295
rect 37365 -30483 37423 -30471
rect 37523 -30295 37581 -30283
rect 37523 -30471 37535 -30295
rect 37569 -30471 37581 -30295
rect 37523 -30483 37581 -30471
rect 37805 -30295 37863 -30283
rect 37805 -30471 37817 -30295
rect 37851 -30471 37863 -30295
rect 37805 -30483 37863 -30471
rect 37963 -30295 38021 -30283
rect 37963 -30471 37975 -30295
rect 38009 -30471 38021 -30295
rect 37963 -30483 38021 -30471
<< mvpdiff >>
rect 27926 11458 28726 11470
rect 27926 11424 27938 11458
rect 28714 11424 28726 11458
rect 27926 11412 28726 11424
rect 27926 11300 28726 11312
rect 27926 11266 27938 11300
rect 28714 11266 28726 11300
rect 27926 11254 28726 11266
rect 27926 11142 28726 11154
rect 27926 11108 27938 11142
rect 28714 11108 28726 11142
rect 27926 11096 28726 11108
rect 27926 10984 28726 10996
rect 27926 10950 27938 10984
rect 28714 10950 28726 10984
rect 27926 10938 28726 10950
rect 27926 10826 28726 10838
rect 27926 10792 27938 10826
rect 28714 10792 28726 10826
rect 27926 10780 28726 10792
rect 30132 10895 30190 10907
rect 30132 10819 30144 10895
rect 30178 10819 30190 10895
rect 30132 10807 30190 10819
rect 30590 10895 30648 10907
rect 30590 10819 30602 10895
rect 30636 10819 30648 10895
rect 30590 10807 30648 10819
rect 30846 10895 30904 10907
rect 27926 10418 28726 10430
rect 27926 10384 27938 10418
rect 28714 10384 28726 10418
rect 27926 10372 28726 10384
rect 27926 10260 28726 10272
rect 27926 10226 27938 10260
rect 28714 10226 28726 10260
rect 27926 10214 28726 10226
rect 27926 10102 28726 10114
rect 27926 10068 27938 10102
rect 28714 10068 28726 10102
rect 27926 10056 28726 10068
rect 27926 9944 28726 9956
rect 27926 9910 27938 9944
rect 28714 9910 28726 9944
rect 27926 9898 28726 9910
rect 27926 9786 28726 9798
rect 27926 9752 27938 9786
rect 28714 9752 28726 9786
rect 27926 9740 28726 9752
rect 30846 10519 30858 10895
rect 30892 10519 30904 10895
rect 30846 10507 30904 10519
rect 31004 10895 31062 10907
rect 31004 10519 31016 10895
rect 31050 10519 31062 10895
rect 31004 10507 31062 10519
rect 31286 10895 31344 10907
rect 31286 10519 31298 10895
rect 31332 10519 31344 10895
rect 31286 10507 31344 10519
rect 31444 10895 31502 10907
rect 31444 10519 31456 10895
rect 31490 10519 31502 10895
rect 31444 10507 31502 10519
rect 31726 10895 31784 10907
rect 31726 10519 31738 10895
rect 31772 10519 31784 10895
rect 31726 10507 31784 10519
rect 31884 10895 31942 10907
rect 31884 10519 31896 10895
rect 31930 10519 31942 10895
rect 31884 10507 31942 10519
rect 32332 10895 32390 10907
rect 32332 10819 32344 10895
rect 32378 10819 32390 10895
rect 32332 10807 32390 10819
rect 32790 10895 32848 10907
rect 32790 10819 32802 10895
rect 32836 10819 32848 10895
rect 32790 10807 32848 10819
rect 33046 10895 33104 10907
rect 33046 10519 33058 10895
rect 33092 10519 33104 10895
rect 33046 10507 33104 10519
rect 33204 10895 33262 10907
rect 33204 10519 33216 10895
rect 33250 10519 33262 10895
rect 33204 10507 33262 10519
rect 33486 10895 33544 10907
rect 33486 10519 33498 10895
rect 33532 10519 33544 10895
rect 33486 10507 33544 10519
rect 33644 10895 33702 10907
rect 33644 10519 33656 10895
rect 33690 10519 33702 10895
rect 33644 10507 33702 10519
rect 33926 10895 33984 10907
rect 33926 10519 33938 10895
rect 33972 10519 33984 10895
rect 33926 10507 33984 10519
rect 34084 10895 34142 10907
rect 34084 10519 34096 10895
rect 34130 10519 34142 10895
rect 34084 10507 34142 10519
rect 34532 10895 34590 10907
rect 34532 10819 34544 10895
rect 34578 10819 34590 10895
rect 34532 10807 34590 10819
rect 34990 10895 35048 10907
rect 34990 10819 35002 10895
rect 35036 10819 35048 10895
rect 34990 10807 35048 10819
rect 35246 10895 35304 10907
rect 35246 10519 35258 10895
rect 35292 10519 35304 10895
rect 35246 10507 35304 10519
rect 35404 10895 35462 10907
rect 35404 10519 35416 10895
rect 35450 10519 35462 10895
rect 35404 10507 35462 10519
rect 35686 10895 35744 10907
rect 35686 10519 35698 10895
rect 35732 10519 35744 10895
rect 35686 10507 35744 10519
rect 35844 10895 35902 10907
rect 35844 10519 35856 10895
rect 35890 10519 35902 10895
rect 35844 10507 35902 10519
rect 36126 10895 36184 10907
rect 36126 10519 36138 10895
rect 36172 10519 36184 10895
rect 36126 10507 36184 10519
rect 36284 10895 36342 10907
rect 36284 10519 36296 10895
rect 36330 10519 36342 10895
rect 36284 10507 36342 10519
rect 27926 9378 28726 9390
rect 27926 9344 27938 9378
rect 28714 9344 28726 9378
rect 27926 9332 28726 9344
rect 27926 9220 28726 9232
rect 27926 9186 27938 9220
rect 28714 9186 28726 9220
rect 27926 9174 28726 9186
rect 27926 9062 28726 9074
rect 27926 9028 27938 9062
rect 28714 9028 28726 9062
rect 27926 9016 28726 9028
rect 27926 8904 28726 8916
rect 27926 8870 27938 8904
rect 28714 8870 28726 8904
rect 27926 8858 28726 8870
rect 27926 8746 28726 8758
rect 27926 8712 27938 8746
rect 28714 8712 28726 8746
rect 27926 8700 28726 8712
rect 29720 9585 29778 9597
rect 29720 9209 29732 9585
rect 29766 9209 29778 9585
rect 29720 9197 29778 9209
rect 30578 9585 30636 9597
rect 30578 9209 30590 9585
rect 30624 9209 30636 9585
rect 30578 9197 30636 9209
rect 31436 9585 31494 9597
rect 31436 9209 31448 9585
rect 31482 9209 31494 9585
rect 31436 9197 31494 9209
rect 27926 8338 28726 8350
rect 27926 8304 27938 8338
rect 28714 8304 28726 8338
rect 27926 8292 28726 8304
rect 27926 8180 28726 8192
rect 27926 8146 27938 8180
rect 28714 8146 28726 8180
rect 27926 8134 28726 8146
rect 27926 8022 28726 8034
rect 27926 7988 27938 8022
rect 28714 7988 28726 8022
rect 27926 7976 28726 7988
rect 27926 7864 28726 7876
rect 27926 7830 27938 7864
rect 28714 7830 28726 7864
rect 27926 7818 28726 7830
rect 27926 7706 28726 7718
rect 27926 7672 27938 7706
rect 28714 7672 28726 7706
rect 27926 7660 28726 7672
rect 27926 7298 28726 7310
rect 27926 7264 27938 7298
rect 28714 7264 28726 7298
rect 27926 7252 28726 7264
rect 27926 7140 28726 7152
rect 27926 7106 27938 7140
rect 28714 7106 28726 7140
rect 27926 7094 28726 7106
rect 27926 6982 28726 6994
rect 27926 6948 27938 6982
rect 28714 6948 28726 6982
rect 27926 6936 28726 6948
rect 27926 6824 28726 6836
rect 27926 6790 27938 6824
rect 28714 6790 28726 6824
rect 27926 6778 28726 6790
rect 27926 6666 28726 6678
rect 27926 6632 27938 6666
rect 28714 6632 28726 6666
rect 27926 6620 28726 6632
rect 29720 8581 29778 8593
rect 29720 8205 29732 8581
rect 29766 8205 29778 8581
rect 29720 8193 29778 8205
rect 30578 8581 30636 8593
rect 30578 8205 30590 8581
rect 30624 8205 30636 8581
rect 30578 8193 30636 8205
rect 31436 8581 31494 8593
rect 31436 8205 31448 8581
rect 31482 8205 31494 8581
rect 31436 8193 31494 8205
rect 29720 7945 29778 7957
rect 29720 7569 29732 7945
rect 29766 7569 29778 7945
rect 29720 7557 29778 7569
rect 30578 7945 30636 7957
rect 30578 7569 30590 7945
rect 30624 7569 30636 7945
rect 30578 7557 30636 7569
rect 31436 7945 31494 7957
rect 31436 7569 31448 7945
rect 31482 7569 31494 7945
rect 31436 7557 31494 7569
rect 29757 7064 30557 7076
rect 29757 7030 29769 7064
rect 30545 7030 30557 7064
rect 29757 7018 30557 7030
rect 29757 6806 30557 6818
rect 29757 6772 29769 6806
rect 30545 6772 30557 6806
rect 29757 6760 30557 6772
rect 31097 7064 31897 7076
rect 31097 7030 31109 7064
rect 31885 7030 31897 7064
rect 31097 7018 31897 7030
rect 31097 6806 31897 6818
rect 31097 6772 31109 6806
rect 31885 6772 31897 6806
rect 31097 6760 31897 6772
rect 27926 6258 28726 6270
rect 27926 6224 27938 6258
rect 28714 6224 28726 6258
rect 27926 6212 28726 6224
rect 27926 6100 28726 6112
rect 27926 6066 27938 6100
rect 28714 6066 28726 6100
rect 27926 6054 28726 6066
rect 27926 5942 28726 5954
rect 27926 5908 27938 5942
rect 28714 5908 28726 5942
rect 27926 5896 28726 5908
rect 27926 5784 28726 5796
rect 27926 5750 27938 5784
rect 28714 5750 28726 5784
rect 27926 5738 28726 5750
rect 27926 5626 28726 5638
rect 27926 5592 27938 5626
rect 28714 5592 28726 5626
rect 27926 5580 28726 5592
rect 27900 5145 27958 5157
rect 27900 4369 27912 5145
rect 27946 4369 27958 5145
rect 27900 4357 27958 4369
rect 28758 5145 28816 5157
rect 28758 4369 28770 5145
rect 28804 4369 28816 5145
rect 28758 4357 28816 4369
rect 57 -8170 457 -8158
rect 57 -8204 69 -8170
rect 445 -8204 457 -8170
rect 57 -8216 457 -8204
rect 693 -8170 1093 -8158
rect 693 -8204 705 -8170
rect 1081 -8204 1093 -8170
rect 693 -8216 1093 -8204
rect 57 -8428 457 -8416
rect 57 -8462 69 -8428
rect 445 -8462 457 -8428
rect 57 -8474 457 -8462
rect 693 -8428 1093 -8416
rect 693 -8462 705 -8428
rect 1081 -8462 1093 -8428
rect 693 -8474 1093 -8462
rect 57 -8696 457 -8684
rect 57 -8730 69 -8696
rect 445 -8730 457 -8696
rect 57 -8742 457 -8730
rect 693 -8696 1093 -8684
rect 693 -8730 705 -8696
rect 1081 -8730 1093 -8696
rect 693 -8742 1093 -8730
rect 57 -9554 457 -9542
rect 57 -9588 69 -9554
rect 445 -9588 457 -9554
rect 57 -9600 457 -9588
rect 693 -9554 1093 -9542
rect 693 -9588 705 -9554
rect 1081 -9588 1093 -9554
rect 693 -9600 1093 -9588
rect 1657 -8170 2057 -8158
rect 1657 -8204 1669 -8170
rect 2045 -8204 2057 -8170
rect 1657 -8216 2057 -8204
rect 2293 -8170 2693 -8158
rect 2293 -8204 2305 -8170
rect 2681 -8204 2693 -8170
rect 2293 -8216 2693 -8204
rect 1657 -8428 2057 -8416
rect 1657 -8462 1669 -8428
rect 2045 -8462 2057 -8428
rect 1657 -8474 2057 -8462
rect 2293 -8428 2693 -8416
rect 2293 -8462 2305 -8428
rect 2681 -8462 2693 -8428
rect 2293 -8474 2693 -8462
rect 1657 -8696 2057 -8684
rect 1657 -8730 1669 -8696
rect 2045 -8730 2057 -8696
rect 1657 -8742 2057 -8730
rect 2293 -8696 2693 -8684
rect 2293 -8730 2305 -8696
rect 2681 -8730 2693 -8696
rect 2293 -8742 2693 -8730
rect 1657 -9554 2057 -9542
rect 1657 -9588 1669 -9554
rect 2045 -9588 2057 -9554
rect 1657 -9600 2057 -9588
rect 2293 -9554 2693 -9542
rect 2293 -9588 2305 -9554
rect 2681 -9588 2693 -9554
rect 2293 -9600 2693 -9588
rect 3257 -8170 3657 -8158
rect 3257 -8204 3269 -8170
rect 3645 -8204 3657 -8170
rect 3257 -8216 3657 -8204
rect 3893 -8170 4293 -8158
rect 3893 -8204 3905 -8170
rect 4281 -8204 4293 -8170
rect 3893 -8216 4293 -8204
rect 3257 -8428 3657 -8416
rect 3257 -8462 3269 -8428
rect 3645 -8462 3657 -8428
rect 3257 -8474 3657 -8462
rect 3893 -8428 4293 -8416
rect 3893 -8462 3905 -8428
rect 4281 -8462 4293 -8428
rect 3893 -8474 4293 -8462
rect 3257 -8696 3657 -8684
rect 3257 -8730 3269 -8696
rect 3645 -8730 3657 -8696
rect 3257 -8742 3657 -8730
rect 3893 -8696 4293 -8684
rect 3893 -8730 3905 -8696
rect 4281 -8730 4293 -8696
rect 3893 -8742 4293 -8730
rect 3257 -9554 3657 -9542
rect 3257 -9588 3269 -9554
rect 3645 -9588 3657 -9554
rect 3257 -9600 3657 -9588
rect 3893 -9554 4293 -9542
rect 3893 -9588 3905 -9554
rect 4281 -9588 4293 -9554
rect 3893 -9600 4293 -9588
rect 4857 -8170 5257 -8158
rect 4857 -8204 4869 -8170
rect 5245 -8204 5257 -8170
rect 4857 -8216 5257 -8204
rect 5493 -8170 5893 -8158
rect 5493 -8204 5505 -8170
rect 5881 -8204 5893 -8170
rect 5493 -8216 5893 -8204
rect 4857 -8428 5257 -8416
rect 4857 -8462 4869 -8428
rect 5245 -8462 5257 -8428
rect 4857 -8474 5257 -8462
rect 5493 -8428 5893 -8416
rect 5493 -8462 5505 -8428
rect 5881 -8462 5893 -8428
rect 5493 -8474 5893 -8462
rect 4857 -8696 5257 -8684
rect 4857 -8730 4869 -8696
rect 5245 -8730 5257 -8696
rect 4857 -8742 5257 -8730
rect 5493 -8696 5893 -8684
rect 5493 -8730 5505 -8696
rect 5881 -8730 5893 -8696
rect 5493 -8742 5893 -8730
rect 4857 -9554 5257 -9542
rect 4857 -9588 4869 -9554
rect 5245 -9588 5257 -9554
rect 4857 -9600 5257 -9588
rect 5493 -9554 5893 -9542
rect 5493 -9588 5505 -9554
rect 5881 -9588 5893 -9554
rect 5493 -9600 5893 -9588
rect 6457 -8170 6857 -8158
rect 6457 -8204 6469 -8170
rect 6845 -8204 6857 -8170
rect 6457 -8216 6857 -8204
rect 7093 -8170 7493 -8158
rect 7093 -8204 7105 -8170
rect 7481 -8204 7493 -8170
rect 7093 -8216 7493 -8204
rect 6457 -8428 6857 -8416
rect 6457 -8462 6469 -8428
rect 6845 -8462 6857 -8428
rect 6457 -8474 6857 -8462
rect 7093 -8428 7493 -8416
rect 7093 -8462 7105 -8428
rect 7481 -8462 7493 -8428
rect 7093 -8474 7493 -8462
rect 6457 -8696 6857 -8684
rect 6457 -8730 6469 -8696
rect 6845 -8730 6857 -8696
rect 6457 -8742 6857 -8730
rect 7093 -8696 7493 -8684
rect 7093 -8730 7105 -8696
rect 7481 -8730 7493 -8696
rect 7093 -8742 7493 -8730
rect 6457 -9554 6857 -9542
rect 6457 -9588 6469 -9554
rect 6845 -9588 6857 -9554
rect 6457 -9600 6857 -9588
rect 7093 -9554 7493 -9542
rect 7093 -9588 7105 -9554
rect 7481 -9588 7493 -9554
rect 7093 -9600 7493 -9588
rect 8057 -8170 8457 -8158
rect 8057 -8204 8069 -8170
rect 8445 -8204 8457 -8170
rect 8057 -8216 8457 -8204
rect 8693 -8170 9093 -8158
rect 8693 -8204 8705 -8170
rect 9081 -8204 9093 -8170
rect 8693 -8216 9093 -8204
rect 8057 -8428 8457 -8416
rect 8057 -8462 8069 -8428
rect 8445 -8462 8457 -8428
rect 8057 -8474 8457 -8462
rect 8693 -8428 9093 -8416
rect 8693 -8462 8705 -8428
rect 9081 -8462 9093 -8428
rect 8693 -8474 9093 -8462
rect 8057 -8696 8457 -8684
rect 8057 -8730 8069 -8696
rect 8445 -8730 8457 -8696
rect 8057 -8742 8457 -8730
rect 8693 -8696 9093 -8684
rect 8693 -8730 8705 -8696
rect 9081 -8730 9093 -8696
rect 8693 -8742 9093 -8730
rect 8057 -9554 8457 -9542
rect 8057 -9588 8069 -9554
rect 8445 -9588 8457 -9554
rect 8057 -9600 8457 -9588
rect 8693 -9554 9093 -9542
rect 8693 -9588 8705 -9554
rect 9081 -9588 9093 -9554
rect 8693 -9600 9093 -9588
rect 9657 -8170 10057 -8158
rect 9657 -8204 9669 -8170
rect 10045 -8204 10057 -8170
rect 9657 -8216 10057 -8204
rect 10293 -8170 10693 -8158
rect 10293 -8204 10305 -8170
rect 10681 -8204 10693 -8170
rect 10293 -8216 10693 -8204
rect 9657 -8428 10057 -8416
rect 9657 -8462 9669 -8428
rect 10045 -8462 10057 -8428
rect 9657 -8474 10057 -8462
rect 10293 -8428 10693 -8416
rect 10293 -8462 10305 -8428
rect 10681 -8462 10693 -8428
rect 10293 -8474 10693 -8462
rect 9657 -8696 10057 -8684
rect 9657 -8730 9669 -8696
rect 10045 -8730 10057 -8696
rect 9657 -8742 10057 -8730
rect 10293 -8696 10693 -8684
rect 10293 -8730 10305 -8696
rect 10681 -8730 10693 -8696
rect 10293 -8742 10693 -8730
rect 9657 -9554 10057 -9542
rect 9657 -9588 9669 -9554
rect 10045 -9588 10057 -9554
rect 9657 -9600 10057 -9588
rect 10293 -9554 10693 -9542
rect 10293 -9588 10305 -9554
rect 10681 -9588 10693 -9554
rect 10293 -9600 10693 -9588
rect 11257 -8170 11657 -8158
rect 11257 -8204 11269 -8170
rect 11645 -8204 11657 -8170
rect 11257 -8216 11657 -8204
rect 11893 -8170 12293 -8158
rect 11893 -8204 11905 -8170
rect 12281 -8204 12293 -8170
rect 11893 -8216 12293 -8204
rect 11257 -8428 11657 -8416
rect 11257 -8462 11269 -8428
rect 11645 -8462 11657 -8428
rect 11257 -8474 11657 -8462
rect 11893 -8428 12293 -8416
rect 11893 -8462 11905 -8428
rect 12281 -8462 12293 -8428
rect 11893 -8474 12293 -8462
rect 11257 -8696 11657 -8684
rect 11257 -8730 11269 -8696
rect 11645 -8730 11657 -8696
rect 11257 -8742 11657 -8730
rect 11893 -8696 12293 -8684
rect 11893 -8730 11905 -8696
rect 12281 -8730 12293 -8696
rect 11893 -8742 12293 -8730
rect 11257 -9554 11657 -9542
rect 11257 -9588 11269 -9554
rect 11645 -9588 11657 -9554
rect 11257 -9600 11657 -9588
rect 11893 -9554 12293 -9542
rect 11893 -9588 11905 -9554
rect 12281 -9588 12293 -9554
rect 11893 -9600 12293 -9588
rect 12857 -8170 13257 -8158
rect 12857 -8204 12869 -8170
rect 13245 -8204 13257 -8170
rect 12857 -8216 13257 -8204
rect 13493 -8170 13893 -8158
rect 13493 -8204 13505 -8170
rect 13881 -8204 13893 -8170
rect 13493 -8216 13893 -8204
rect 12857 -8428 13257 -8416
rect 12857 -8462 12869 -8428
rect 13245 -8462 13257 -8428
rect 12857 -8474 13257 -8462
rect 13493 -8428 13893 -8416
rect 13493 -8462 13505 -8428
rect 13881 -8462 13893 -8428
rect 13493 -8474 13893 -8462
rect 12857 -8696 13257 -8684
rect 12857 -8730 12869 -8696
rect 13245 -8730 13257 -8696
rect 12857 -8742 13257 -8730
rect 13493 -8696 13893 -8684
rect 13493 -8730 13505 -8696
rect 13881 -8730 13893 -8696
rect 13493 -8742 13893 -8730
rect 12857 -9554 13257 -9542
rect 12857 -9588 12869 -9554
rect 13245 -9588 13257 -9554
rect 12857 -9600 13257 -9588
rect 13493 -9554 13893 -9542
rect 13493 -9588 13505 -9554
rect 13881 -9588 13893 -9554
rect 13493 -9600 13893 -9588
rect 14457 -8170 14857 -8158
rect 14457 -8204 14469 -8170
rect 14845 -8204 14857 -8170
rect 14457 -8216 14857 -8204
rect 15093 -8170 15493 -8158
rect 15093 -8204 15105 -8170
rect 15481 -8204 15493 -8170
rect 15093 -8216 15493 -8204
rect 14457 -8428 14857 -8416
rect 14457 -8462 14469 -8428
rect 14845 -8462 14857 -8428
rect 14457 -8474 14857 -8462
rect 15093 -8428 15493 -8416
rect 15093 -8462 15105 -8428
rect 15481 -8462 15493 -8428
rect 15093 -8474 15493 -8462
rect 14457 -8696 14857 -8684
rect 14457 -8730 14469 -8696
rect 14845 -8730 14857 -8696
rect 14457 -8742 14857 -8730
rect 15093 -8696 15493 -8684
rect 15093 -8730 15105 -8696
rect 15481 -8730 15493 -8696
rect 15093 -8742 15493 -8730
rect 14457 -9554 14857 -9542
rect 14457 -9588 14469 -9554
rect 14845 -9588 14857 -9554
rect 14457 -9600 14857 -9588
rect 15093 -9554 15493 -9542
rect 15093 -9588 15105 -9554
rect 15481 -9588 15493 -9554
rect 15093 -9600 15493 -9588
rect 16057 -8170 16457 -8158
rect 16057 -8204 16069 -8170
rect 16445 -8204 16457 -8170
rect 16057 -8216 16457 -8204
rect 16693 -8170 17093 -8158
rect 16693 -8204 16705 -8170
rect 17081 -8204 17093 -8170
rect 16693 -8216 17093 -8204
rect 16057 -8428 16457 -8416
rect 16057 -8462 16069 -8428
rect 16445 -8462 16457 -8428
rect 16057 -8474 16457 -8462
rect 16693 -8428 17093 -8416
rect 16693 -8462 16705 -8428
rect 17081 -8462 17093 -8428
rect 16693 -8474 17093 -8462
rect 16057 -8696 16457 -8684
rect 16057 -8730 16069 -8696
rect 16445 -8730 16457 -8696
rect 16057 -8742 16457 -8730
rect 16693 -8696 17093 -8684
rect 16693 -8730 16705 -8696
rect 17081 -8730 17093 -8696
rect 16693 -8742 17093 -8730
rect 16057 -9554 16457 -9542
rect 16057 -9588 16069 -9554
rect 16445 -9588 16457 -9554
rect 16057 -9600 16457 -9588
rect 16693 -9554 17093 -9542
rect 16693 -9588 16705 -9554
rect 17081 -9588 17093 -9554
rect 16693 -9600 17093 -9588
rect 17657 -8170 18057 -8158
rect 17657 -8204 17669 -8170
rect 18045 -8204 18057 -8170
rect 17657 -8216 18057 -8204
rect 18293 -8170 18693 -8158
rect 18293 -8204 18305 -8170
rect 18681 -8204 18693 -8170
rect 18293 -8216 18693 -8204
rect 17657 -8428 18057 -8416
rect 17657 -8462 17669 -8428
rect 18045 -8462 18057 -8428
rect 17657 -8474 18057 -8462
rect 18293 -8428 18693 -8416
rect 18293 -8462 18305 -8428
rect 18681 -8462 18693 -8428
rect 18293 -8474 18693 -8462
rect 17657 -8696 18057 -8684
rect 17657 -8730 17669 -8696
rect 18045 -8730 18057 -8696
rect 17657 -8742 18057 -8730
rect 18293 -8696 18693 -8684
rect 18293 -8730 18305 -8696
rect 18681 -8730 18693 -8696
rect 18293 -8742 18693 -8730
rect 17657 -9554 18057 -9542
rect 17657 -9588 17669 -9554
rect 18045 -9588 18057 -9554
rect 17657 -9600 18057 -9588
rect 18293 -9554 18693 -9542
rect 18293 -9588 18305 -9554
rect 18681 -9588 18693 -9554
rect 18293 -9600 18693 -9588
rect 19257 -8170 19657 -8158
rect 19257 -8204 19269 -8170
rect 19645 -8204 19657 -8170
rect 19257 -8216 19657 -8204
rect 19893 -8170 20293 -8158
rect 19893 -8204 19905 -8170
rect 20281 -8204 20293 -8170
rect 19893 -8216 20293 -8204
rect 19257 -8428 19657 -8416
rect 19257 -8462 19269 -8428
rect 19645 -8462 19657 -8428
rect 19257 -8474 19657 -8462
rect 19893 -8428 20293 -8416
rect 19893 -8462 19905 -8428
rect 20281 -8462 20293 -8428
rect 19893 -8474 20293 -8462
rect 19257 -8696 19657 -8684
rect 19257 -8730 19269 -8696
rect 19645 -8730 19657 -8696
rect 19257 -8742 19657 -8730
rect 19893 -8696 20293 -8684
rect 19893 -8730 19905 -8696
rect 20281 -8730 20293 -8696
rect 19893 -8742 20293 -8730
rect 19257 -9554 19657 -9542
rect 19257 -9588 19269 -9554
rect 19645 -9588 19657 -9554
rect 19257 -9600 19657 -9588
rect 19893 -9554 20293 -9542
rect 19893 -9588 19905 -9554
rect 20281 -9588 20293 -9554
rect 19893 -9600 20293 -9588
rect 20857 -8170 21257 -8158
rect 20857 -8204 20869 -8170
rect 21245 -8204 21257 -8170
rect 20857 -8216 21257 -8204
rect 21493 -8170 21893 -8158
rect 21493 -8204 21505 -8170
rect 21881 -8204 21893 -8170
rect 21493 -8216 21893 -8204
rect 20857 -8428 21257 -8416
rect 20857 -8462 20869 -8428
rect 21245 -8462 21257 -8428
rect 20857 -8474 21257 -8462
rect 21493 -8428 21893 -8416
rect 21493 -8462 21505 -8428
rect 21881 -8462 21893 -8428
rect 21493 -8474 21893 -8462
rect 20857 -8696 21257 -8684
rect 20857 -8730 20869 -8696
rect 21245 -8730 21257 -8696
rect 20857 -8742 21257 -8730
rect 21493 -8696 21893 -8684
rect 21493 -8730 21505 -8696
rect 21881 -8730 21893 -8696
rect 21493 -8742 21893 -8730
rect 20857 -9554 21257 -9542
rect 20857 -9588 20869 -9554
rect 21245 -9588 21257 -9554
rect 20857 -9600 21257 -9588
rect 21493 -9554 21893 -9542
rect 21493 -9588 21505 -9554
rect 21881 -9588 21893 -9554
rect 21493 -9600 21893 -9588
rect 22457 -8170 22857 -8158
rect 22457 -8204 22469 -8170
rect 22845 -8204 22857 -8170
rect 22457 -8216 22857 -8204
rect 23093 -8170 23493 -8158
rect 23093 -8204 23105 -8170
rect 23481 -8204 23493 -8170
rect 23093 -8216 23493 -8204
rect 22457 -8428 22857 -8416
rect 22457 -8462 22469 -8428
rect 22845 -8462 22857 -8428
rect 22457 -8474 22857 -8462
rect 23093 -8428 23493 -8416
rect 23093 -8462 23105 -8428
rect 23481 -8462 23493 -8428
rect 23093 -8474 23493 -8462
rect 22457 -8696 22857 -8684
rect 22457 -8730 22469 -8696
rect 22845 -8730 22857 -8696
rect 22457 -8742 22857 -8730
rect 23093 -8696 23493 -8684
rect 23093 -8730 23105 -8696
rect 23481 -8730 23493 -8696
rect 23093 -8742 23493 -8730
rect 22457 -9554 22857 -9542
rect 22457 -9588 22469 -9554
rect 22845 -9588 22857 -9554
rect 22457 -9600 22857 -9588
rect 23093 -9554 23493 -9542
rect 23093 -9588 23105 -9554
rect 23481 -9588 23493 -9554
rect 23093 -9600 23493 -9588
rect 24057 -8170 24457 -8158
rect 24057 -8204 24069 -8170
rect 24445 -8204 24457 -8170
rect 24057 -8216 24457 -8204
rect 24693 -8170 25093 -8158
rect 24693 -8204 24705 -8170
rect 25081 -8204 25093 -8170
rect 24693 -8216 25093 -8204
rect 24057 -8428 24457 -8416
rect 24057 -8462 24069 -8428
rect 24445 -8462 24457 -8428
rect 24057 -8474 24457 -8462
rect 24693 -8428 25093 -8416
rect 24693 -8462 24705 -8428
rect 25081 -8462 25093 -8428
rect 24693 -8474 25093 -8462
rect 24057 -8696 24457 -8684
rect 24057 -8730 24069 -8696
rect 24445 -8730 24457 -8696
rect 24057 -8742 24457 -8730
rect 24693 -8696 25093 -8684
rect 24693 -8730 24705 -8696
rect 25081 -8730 25093 -8696
rect 24693 -8742 25093 -8730
rect 24057 -9554 24457 -9542
rect 24057 -9588 24069 -9554
rect 24445 -9588 24457 -9554
rect 24057 -9600 24457 -9588
rect 24693 -9554 25093 -9542
rect 24693 -9588 24705 -9554
rect 25081 -9588 25093 -9554
rect 24693 -9600 25093 -9588
rect 25657 -8170 26057 -8158
rect 25657 -8204 25669 -8170
rect 26045 -8204 26057 -8170
rect 25657 -8216 26057 -8204
rect 26293 -8170 26693 -8158
rect 26293 -8204 26305 -8170
rect 26681 -8204 26693 -8170
rect 26293 -8216 26693 -8204
rect 25657 -8428 26057 -8416
rect 25657 -8462 25669 -8428
rect 26045 -8462 26057 -8428
rect 25657 -8474 26057 -8462
rect 26293 -8428 26693 -8416
rect 26293 -8462 26305 -8428
rect 26681 -8462 26693 -8428
rect 26293 -8474 26693 -8462
rect 25657 -8696 26057 -8684
rect 25657 -8730 25669 -8696
rect 26045 -8730 26057 -8696
rect 25657 -8742 26057 -8730
rect 26293 -8696 26693 -8684
rect 26293 -8730 26305 -8696
rect 26681 -8730 26693 -8696
rect 26293 -8742 26693 -8730
rect 25657 -9554 26057 -9542
rect 25657 -9588 25669 -9554
rect 26045 -9588 26057 -9554
rect 25657 -9600 26057 -9588
rect 26293 -9554 26693 -9542
rect 26293 -9588 26305 -9554
rect 26681 -9588 26693 -9554
rect 26293 -9600 26693 -9588
rect 27257 -8170 27657 -8158
rect 27257 -8204 27269 -8170
rect 27645 -8204 27657 -8170
rect 27257 -8216 27657 -8204
rect 27893 -8170 28293 -8158
rect 27893 -8204 27905 -8170
rect 28281 -8204 28293 -8170
rect 27893 -8216 28293 -8204
rect 27257 -8428 27657 -8416
rect 27257 -8462 27269 -8428
rect 27645 -8462 27657 -8428
rect 27257 -8474 27657 -8462
rect 27893 -8428 28293 -8416
rect 27893 -8462 27905 -8428
rect 28281 -8462 28293 -8428
rect 27893 -8474 28293 -8462
rect 27257 -8696 27657 -8684
rect 27257 -8730 27269 -8696
rect 27645 -8730 27657 -8696
rect 27257 -8742 27657 -8730
rect 27893 -8696 28293 -8684
rect 27893 -8730 27905 -8696
rect 28281 -8730 28293 -8696
rect 27893 -8742 28293 -8730
rect 27257 -9554 27657 -9542
rect 27257 -9588 27269 -9554
rect 27645 -9588 27657 -9554
rect 27257 -9600 27657 -9588
rect 27893 -9554 28293 -9542
rect 27893 -9588 27905 -9554
rect 28281 -9588 28293 -9554
rect 27893 -9600 28293 -9588
rect 28857 -8170 29257 -8158
rect 28857 -8204 28869 -8170
rect 29245 -8204 29257 -8170
rect 28857 -8216 29257 -8204
rect 29493 -8170 29893 -8158
rect 29493 -8204 29505 -8170
rect 29881 -8204 29893 -8170
rect 29493 -8216 29893 -8204
rect 28857 -8428 29257 -8416
rect 28857 -8462 28869 -8428
rect 29245 -8462 29257 -8428
rect 28857 -8474 29257 -8462
rect 29493 -8428 29893 -8416
rect 29493 -8462 29505 -8428
rect 29881 -8462 29893 -8428
rect 29493 -8474 29893 -8462
rect 28857 -8696 29257 -8684
rect 28857 -8730 28869 -8696
rect 29245 -8730 29257 -8696
rect 28857 -8742 29257 -8730
rect 29493 -8696 29893 -8684
rect 29493 -8730 29505 -8696
rect 29881 -8730 29893 -8696
rect 29493 -8742 29893 -8730
rect 28857 -9554 29257 -9542
rect 28857 -9588 28869 -9554
rect 29245 -9588 29257 -9554
rect 28857 -9600 29257 -9588
rect 29493 -9554 29893 -9542
rect 29493 -9588 29505 -9554
rect 29881 -9588 29893 -9554
rect 29493 -9600 29893 -9588
rect 30457 -8170 30857 -8158
rect 30457 -8204 30469 -8170
rect 30845 -8204 30857 -8170
rect 30457 -8216 30857 -8204
rect 31093 -8170 31493 -8158
rect 31093 -8204 31105 -8170
rect 31481 -8204 31493 -8170
rect 31093 -8216 31493 -8204
rect 30457 -8428 30857 -8416
rect 30457 -8462 30469 -8428
rect 30845 -8462 30857 -8428
rect 30457 -8474 30857 -8462
rect 31093 -8428 31493 -8416
rect 31093 -8462 31105 -8428
rect 31481 -8462 31493 -8428
rect 31093 -8474 31493 -8462
rect 30457 -8696 30857 -8684
rect 30457 -8730 30469 -8696
rect 30845 -8730 30857 -8696
rect 30457 -8742 30857 -8730
rect 31093 -8696 31493 -8684
rect 31093 -8730 31105 -8696
rect 31481 -8730 31493 -8696
rect 31093 -8742 31493 -8730
rect 30457 -9554 30857 -9542
rect 30457 -9588 30469 -9554
rect 30845 -9588 30857 -9554
rect 30457 -9600 30857 -9588
rect 31093 -9554 31493 -9542
rect 31093 -9588 31105 -9554
rect 31481 -9588 31493 -9554
rect 31093 -9600 31493 -9588
rect 32057 -8170 32457 -8158
rect 32057 -8204 32069 -8170
rect 32445 -8204 32457 -8170
rect 32057 -8216 32457 -8204
rect 32693 -8170 33093 -8158
rect 32693 -8204 32705 -8170
rect 33081 -8204 33093 -8170
rect 32693 -8216 33093 -8204
rect 32057 -8428 32457 -8416
rect 32057 -8462 32069 -8428
rect 32445 -8462 32457 -8428
rect 32057 -8474 32457 -8462
rect 32693 -8428 33093 -8416
rect 32693 -8462 32705 -8428
rect 33081 -8462 33093 -8428
rect 32693 -8474 33093 -8462
rect 32057 -8696 32457 -8684
rect 32057 -8730 32069 -8696
rect 32445 -8730 32457 -8696
rect 32057 -8742 32457 -8730
rect 32693 -8696 33093 -8684
rect 32693 -8730 32705 -8696
rect 33081 -8730 33093 -8696
rect 32693 -8742 33093 -8730
rect 32057 -9554 32457 -9542
rect 32057 -9588 32069 -9554
rect 32445 -9588 32457 -9554
rect 32057 -9600 32457 -9588
rect 32693 -9554 33093 -9542
rect 32693 -9588 32705 -9554
rect 33081 -9588 33093 -9554
rect 32693 -9600 33093 -9588
rect 33657 -8170 34057 -8158
rect 33657 -8204 33669 -8170
rect 34045 -8204 34057 -8170
rect 33657 -8216 34057 -8204
rect 34293 -8170 34693 -8158
rect 34293 -8204 34305 -8170
rect 34681 -8204 34693 -8170
rect 34293 -8216 34693 -8204
rect 33657 -8428 34057 -8416
rect 33657 -8462 33669 -8428
rect 34045 -8462 34057 -8428
rect 33657 -8474 34057 -8462
rect 34293 -8428 34693 -8416
rect 34293 -8462 34305 -8428
rect 34681 -8462 34693 -8428
rect 34293 -8474 34693 -8462
rect 33657 -8696 34057 -8684
rect 33657 -8730 33669 -8696
rect 34045 -8730 34057 -8696
rect 33657 -8742 34057 -8730
rect 34293 -8696 34693 -8684
rect 34293 -8730 34305 -8696
rect 34681 -8730 34693 -8696
rect 34293 -8742 34693 -8730
rect 33657 -9554 34057 -9542
rect 33657 -9588 33669 -9554
rect 34045 -9588 34057 -9554
rect 33657 -9600 34057 -9588
rect 34293 -9554 34693 -9542
rect 34293 -9588 34305 -9554
rect 34681 -9588 34693 -9554
rect 34293 -9600 34693 -9588
rect 35257 -8170 35657 -8158
rect 35257 -8204 35269 -8170
rect 35645 -8204 35657 -8170
rect 35257 -8216 35657 -8204
rect 35893 -8170 36293 -8158
rect 35893 -8204 35905 -8170
rect 36281 -8204 36293 -8170
rect 35893 -8216 36293 -8204
rect 35257 -8428 35657 -8416
rect 35257 -8462 35269 -8428
rect 35645 -8462 35657 -8428
rect 35257 -8474 35657 -8462
rect 35893 -8428 36293 -8416
rect 35893 -8462 35905 -8428
rect 36281 -8462 36293 -8428
rect 35893 -8474 36293 -8462
rect 35257 -8696 35657 -8684
rect 35257 -8730 35269 -8696
rect 35645 -8730 35657 -8696
rect 35257 -8742 35657 -8730
rect 35893 -8696 36293 -8684
rect 35893 -8730 35905 -8696
rect 36281 -8730 36293 -8696
rect 35893 -8742 36293 -8730
rect 35257 -9554 35657 -9542
rect 35257 -9588 35269 -9554
rect 35645 -9588 35657 -9554
rect 35257 -9600 35657 -9588
rect 35893 -9554 36293 -9542
rect 35893 -9588 35905 -9554
rect 36281 -9588 36293 -9554
rect 35893 -9600 36293 -9588
rect 36857 -8170 37257 -8158
rect 36857 -8204 36869 -8170
rect 37245 -8204 37257 -8170
rect 36857 -8216 37257 -8204
rect 37493 -8170 37893 -8158
rect 37493 -8204 37505 -8170
rect 37881 -8204 37893 -8170
rect 37493 -8216 37893 -8204
rect 36857 -8428 37257 -8416
rect 36857 -8462 36869 -8428
rect 37245 -8462 37257 -8428
rect 36857 -8474 37257 -8462
rect 37493 -8428 37893 -8416
rect 37493 -8462 37505 -8428
rect 37881 -8462 37893 -8428
rect 37493 -8474 37893 -8462
rect 36857 -8696 37257 -8684
rect 36857 -8730 36869 -8696
rect 37245 -8730 37257 -8696
rect 36857 -8742 37257 -8730
rect 37493 -8696 37893 -8684
rect 37493 -8730 37505 -8696
rect 37881 -8730 37893 -8696
rect 37493 -8742 37893 -8730
rect 36857 -9554 37257 -9542
rect 36857 -9588 36869 -9554
rect 37245 -9588 37257 -9554
rect 36857 -9600 37257 -9588
rect 37493 -9554 37893 -9542
rect 37493 -9588 37505 -9554
rect 37881 -9588 37893 -9554
rect 37493 -9600 37893 -9588
rect 57 -9970 457 -9958
rect 57 -10004 69 -9970
rect 445 -10004 457 -9970
rect 57 -10016 457 -10004
rect 693 -9970 1093 -9958
rect 693 -10004 705 -9970
rect 1081 -10004 1093 -9970
rect 693 -10016 1093 -10004
rect 57 -10228 457 -10216
rect 57 -10262 69 -10228
rect 445 -10262 457 -10228
rect 57 -10274 457 -10262
rect 693 -10228 1093 -10216
rect 693 -10262 705 -10228
rect 1081 -10262 1093 -10228
rect 693 -10274 1093 -10262
rect 57 -10496 457 -10484
rect 57 -10530 69 -10496
rect 445 -10530 457 -10496
rect 57 -10542 457 -10530
rect 693 -10496 1093 -10484
rect 693 -10530 705 -10496
rect 1081 -10530 1093 -10496
rect 693 -10542 1093 -10530
rect 57 -11354 457 -11342
rect 57 -11388 69 -11354
rect 445 -11388 457 -11354
rect 57 -11400 457 -11388
rect 693 -11354 1093 -11342
rect 693 -11388 705 -11354
rect 1081 -11388 1093 -11354
rect 693 -11400 1093 -11388
rect 1657 -9970 2057 -9958
rect 1657 -10004 1669 -9970
rect 2045 -10004 2057 -9970
rect 1657 -10016 2057 -10004
rect 2293 -9970 2693 -9958
rect 2293 -10004 2305 -9970
rect 2681 -10004 2693 -9970
rect 2293 -10016 2693 -10004
rect 1657 -10228 2057 -10216
rect 1657 -10262 1669 -10228
rect 2045 -10262 2057 -10228
rect 1657 -10274 2057 -10262
rect 2293 -10228 2693 -10216
rect 2293 -10262 2305 -10228
rect 2681 -10262 2693 -10228
rect 2293 -10274 2693 -10262
rect 1657 -10496 2057 -10484
rect 1657 -10530 1669 -10496
rect 2045 -10530 2057 -10496
rect 1657 -10542 2057 -10530
rect 2293 -10496 2693 -10484
rect 2293 -10530 2305 -10496
rect 2681 -10530 2693 -10496
rect 2293 -10542 2693 -10530
rect 1657 -11354 2057 -11342
rect 1657 -11388 1669 -11354
rect 2045 -11388 2057 -11354
rect 1657 -11400 2057 -11388
rect 2293 -11354 2693 -11342
rect 2293 -11388 2305 -11354
rect 2681 -11388 2693 -11354
rect 2293 -11400 2693 -11388
rect 3257 -9970 3657 -9958
rect 3257 -10004 3269 -9970
rect 3645 -10004 3657 -9970
rect 3257 -10016 3657 -10004
rect 3893 -9970 4293 -9958
rect 3893 -10004 3905 -9970
rect 4281 -10004 4293 -9970
rect 3893 -10016 4293 -10004
rect 3257 -10228 3657 -10216
rect 3257 -10262 3269 -10228
rect 3645 -10262 3657 -10228
rect 3257 -10274 3657 -10262
rect 3893 -10228 4293 -10216
rect 3893 -10262 3905 -10228
rect 4281 -10262 4293 -10228
rect 3893 -10274 4293 -10262
rect 3257 -10496 3657 -10484
rect 3257 -10530 3269 -10496
rect 3645 -10530 3657 -10496
rect 3257 -10542 3657 -10530
rect 3893 -10496 4293 -10484
rect 3893 -10530 3905 -10496
rect 4281 -10530 4293 -10496
rect 3893 -10542 4293 -10530
rect 3257 -11354 3657 -11342
rect 3257 -11388 3269 -11354
rect 3645 -11388 3657 -11354
rect 3257 -11400 3657 -11388
rect 3893 -11354 4293 -11342
rect 3893 -11388 3905 -11354
rect 4281 -11388 4293 -11354
rect 3893 -11400 4293 -11388
rect 4857 -9970 5257 -9958
rect 4857 -10004 4869 -9970
rect 5245 -10004 5257 -9970
rect 4857 -10016 5257 -10004
rect 5493 -9970 5893 -9958
rect 5493 -10004 5505 -9970
rect 5881 -10004 5893 -9970
rect 5493 -10016 5893 -10004
rect 4857 -10228 5257 -10216
rect 4857 -10262 4869 -10228
rect 5245 -10262 5257 -10228
rect 4857 -10274 5257 -10262
rect 5493 -10228 5893 -10216
rect 5493 -10262 5505 -10228
rect 5881 -10262 5893 -10228
rect 5493 -10274 5893 -10262
rect 4857 -10496 5257 -10484
rect 4857 -10530 4869 -10496
rect 5245 -10530 5257 -10496
rect 4857 -10542 5257 -10530
rect 5493 -10496 5893 -10484
rect 5493 -10530 5505 -10496
rect 5881 -10530 5893 -10496
rect 5493 -10542 5893 -10530
rect 4857 -11354 5257 -11342
rect 4857 -11388 4869 -11354
rect 5245 -11388 5257 -11354
rect 4857 -11400 5257 -11388
rect 5493 -11354 5893 -11342
rect 5493 -11388 5505 -11354
rect 5881 -11388 5893 -11354
rect 5493 -11400 5893 -11388
rect 6457 -9970 6857 -9958
rect 6457 -10004 6469 -9970
rect 6845 -10004 6857 -9970
rect 6457 -10016 6857 -10004
rect 7093 -9970 7493 -9958
rect 7093 -10004 7105 -9970
rect 7481 -10004 7493 -9970
rect 7093 -10016 7493 -10004
rect 6457 -10228 6857 -10216
rect 6457 -10262 6469 -10228
rect 6845 -10262 6857 -10228
rect 6457 -10274 6857 -10262
rect 7093 -10228 7493 -10216
rect 7093 -10262 7105 -10228
rect 7481 -10262 7493 -10228
rect 7093 -10274 7493 -10262
rect 6457 -10496 6857 -10484
rect 6457 -10530 6469 -10496
rect 6845 -10530 6857 -10496
rect 6457 -10542 6857 -10530
rect 7093 -10496 7493 -10484
rect 7093 -10530 7105 -10496
rect 7481 -10530 7493 -10496
rect 7093 -10542 7493 -10530
rect 6457 -11354 6857 -11342
rect 6457 -11388 6469 -11354
rect 6845 -11388 6857 -11354
rect 6457 -11400 6857 -11388
rect 7093 -11354 7493 -11342
rect 7093 -11388 7105 -11354
rect 7481 -11388 7493 -11354
rect 7093 -11400 7493 -11388
rect 8057 -9970 8457 -9958
rect 8057 -10004 8069 -9970
rect 8445 -10004 8457 -9970
rect 8057 -10016 8457 -10004
rect 8693 -9970 9093 -9958
rect 8693 -10004 8705 -9970
rect 9081 -10004 9093 -9970
rect 8693 -10016 9093 -10004
rect 8057 -10228 8457 -10216
rect 8057 -10262 8069 -10228
rect 8445 -10262 8457 -10228
rect 8057 -10274 8457 -10262
rect 8693 -10228 9093 -10216
rect 8693 -10262 8705 -10228
rect 9081 -10262 9093 -10228
rect 8693 -10274 9093 -10262
rect 8057 -10496 8457 -10484
rect 8057 -10530 8069 -10496
rect 8445 -10530 8457 -10496
rect 8057 -10542 8457 -10530
rect 8693 -10496 9093 -10484
rect 8693 -10530 8705 -10496
rect 9081 -10530 9093 -10496
rect 8693 -10542 9093 -10530
rect 8057 -11354 8457 -11342
rect 8057 -11388 8069 -11354
rect 8445 -11388 8457 -11354
rect 8057 -11400 8457 -11388
rect 8693 -11354 9093 -11342
rect 8693 -11388 8705 -11354
rect 9081 -11388 9093 -11354
rect 8693 -11400 9093 -11388
rect 9657 -9970 10057 -9958
rect 9657 -10004 9669 -9970
rect 10045 -10004 10057 -9970
rect 9657 -10016 10057 -10004
rect 10293 -9970 10693 -9958
rect 10293 -10004 10305 -9970
rect 10681 -10004 10693 -9970
rect 10293 -10016 10693 -10004
rect 9657 -10228 10057 -10216
rect 9657 -10262 9669 -10228
rect 10045 -10262 10057 -10228
rect 9657 -10274 10057 -10262
rect 10293 -10228 10693 -10216
rect 10293 -10262 10305 -10228
rect 10681 -10262 10693 -10228
rect 10293 -10274 10693 -10262
rect 9657 -10496 10057 -10484
rect 9657 -10530 9669 -10496
rect 10045 -10530 10057 -10496
rect 9657 -10542 10057 -10530
rect 10293 -10496 10693 -10484
rect 10293 -10530 10305 -10496
rect 10681 -10530 10693 -10496
rect 10293 -10542 10693 -10530
rect 9657 -11354 10057 -11342
rect 9657 -11388 9669 -11354
rect 10045 -11388 10057 -11354
rect 9657 -11400 10057 -11388
rect 10293 -11354 10693 -11342
rect 10293 -11388 10305 -11354
rect 10681 -11388 10693 -11354
rect 10293 -11400 10693 -11388
rect 11257 -9970 11657 -9958
rect 11257 -10004 11269 -9970
rect 11645 -10004 11657 -9970
rect 11257 -10016 11657 -10004
rect 11893 -9970 12293 -9958
rect 11893 -10004 11905 -9970
rect 12281 -10004 12293 -9970
rect 11893 -10016 12293 -10004
rect 11257 -10228 11657 -10216
rect 11257 -10262 11269 -10228
rect 11645 -10262 11657 -10228
rect 11257 -10274 11657 -10262
rect 11893 -10228 12293 -10216
rect 11893 -10262 11905 -10228
rect 12281 -10262 12293 -10228
rect 11893 -10274 12293 -10262
rect 11257 -10496 11657 -10484
rect 11257 -10530 11269 -10496
rect 11645 -10530 11657 -10496
rect 11257 -10542 11657 -10530
rect 11893 -10496 12293 -10484
rect 11893 -10530 11905 -10496
rect 12281 -10530 12293 -10496
rect 11893 -10542 12293 -10530
rect 11257 -11354 11657 -11342
rect 11257 -11388 11269 -11354
rect 11645 -11388 11657 -11354
rect 11257 -11400 11657 -11388
rect 11893 -11354 12293 -11342
rect 11893 -11388 11905 -11354
rect 12281 -11388 12293 -11354
rect 11893 -11400 12293 -11388
rect 12857 -9970 13257 -9958
rect 12857 -10004 12869 -9970
rect 13245 -10004 13257 -9970
rect 12857 -10016 13257 -10004
rect 13493 -9970 13893 -9958
rect 13493 -10004 13505 -9970
rect 13881 -10004 13893 -9970
rect 13493 -10016 13893 -10004
rect 12857 -10228 13257 -10216
rect 12857 -10262 12869 -10228
rect 13245 -10262 13257 -10228
rect 12857 -10274 13257 -10262
rect 13493 -10228 13893 -10216
rect 13493 -10262 13505 -10228
rect 13881 -10262 13893 -10228
rect 13493 -10274 13893 -10262
rect 12857 -10496 13257 -10484
rect 12857 -10530 12869 -10496
rect 13245 -10530 13257 -10496
rect 12857 -10542 13257 -10530
rect 13493 -10496 13893 -10484
rect 13493 -10530 13505 -10496
rect 13881 -10530 13893 -10496
rect 13493 -10542 13893 -10530
rect 12857 -11354 13257 -11342
rect 12857 -11388 12869 -11354
rect 13245 -11388 13257 -11354
rect 12857 -11400 13257 -11388
rect 13493 -11354 13893 -11342
rect 13493 -11388 13505 -11354
rect 13881 -11388 13893 -11354
rect 13493 -11400 13893 -11388
rect 14457 -9970 14857 -9958
rect 14457 -10004 14469 -9970
rect 14845 -10004 14857 -9970
rect 14457 -10016 14857 -10004
rect 15093 -9970 15493 -9958
rect 15093 -10004 15105 -9970
rect 15481 -10004 15493 -9970
rect 15093 -10016 15493 -10004
rect 14457 -10228 14857 -10216
rect 14457 -10262 14469 -10228
rect 14845 -10262 14857 -10228
rect 14457 -10274 14857 -10262
rect 15093 -10228 15493 -10216
rect 15093 -10262 15105 -10228
rect 15481 -10262 15493 -10228
rect 15093 -10274 15493 -10262
rect 14457 -10496 14857 -10484
rect 14457 -10530 14469 -10496
rect 14845 -10530 14857 -10496
rect 14457 -10542 14857 -10530
rect 15093 -10496 15493 -10484
rect 15093 -10530 15105 -10496
rect 15481 -10530 15493 -10496
rect 15093 -10542 15493 -10530
rect 14457 -11354 14857 -11342
rect 14457 -11388 14469 -11354
rect 14845 -11388 14857 -11354
rect 14457 -11400 14857 -11388
rect 15093 -11354 15493 -11342
rect 15093 -11388 15105 -11354
rect 15481 -11388 15493 -11354
rect 15093 -11400 15493 -11388
rect 16057 -9970 16457 -9958
rect 16057 -10004 16069 -9970
rect 16445 -10004 16457 -9970
rect 16057 -10016 16457 -10004
rect 16693 -9970 17093 -9958
rect 16693 -10004 16705 -9970
rect 17081 -10004 17093 -9970
rect 16693 -10016 17093 -10004
rect 16057 -10228 16457 -10216
rect 16057 -10262 16069 -10228
rect 16445 -10262 16457 -10228
rect 16057 -10274 16457 -10262
rect 16693 -10228 17093 -10216
rect 16693 -10262 16705 -10228
rect 17081 -10262 17093 -10228
rect 16693 -10274 17093 -10262
rect 16057 -10496 16457 -10484
rect 16057 -10530 16069 -10496
rect 16445 -10530 16457 -10496
rect 16057 -10542 16457 -10530
rect 16693 -10496 17093 -10484
rect 16693 -10530 16705 -10496
rect 17081 -10530 17093 -10496
rect 16693 -10542 17093 -10530
rect 16057 -11354 16457 -11342
rect 16057 -11388 16069 -11354
rect 16445 -11388 16457 -11354
rect 16057 -11400 16457 -11388
rect 16693 -11354 17093 -11342
rect 16693 -11388 16705 -11354
rect 17081 -11388 17093 -11354
rect 16693 -11400 17093 -11388
rect 17657 -9970 18057 -9958
rect 17657 -10004 17669 -9970
rect 18045 -10004 18057 -9970
rect 17657 -10016 18057 -10004
rect 18293 -9970 18693 -9958
rect 18293 -10004 18305 -9970
rect 18681 -10004 18693 -9970
rect 18293 -10016 18693 -10004
rect 17657 -10228 18057 -10216
rect 17657 -10262 17669 -10228
rect 18045 -10262 18057 -10228
rect 17657 -10274 18057 -10262
rect 18293 -10228 18693 -10216
rect 18293 -10262 18305 -10228
rect 18681 -10262 18693 -10228
rect 18293 -10274 18693 -10262
rect 17657 -10496 18057 -10484
rect 17657 -10530 17669 -10496
rect 18045 -10530 18057 -10496
rect 17657 -10542 18057 -10530
rect 18293 -10496 18693 -10484
rect 18293 -10530 18305 -10496
rect 18681 -10530 18693 -10496
rect 18293 -10542 18693 -10530
rect 17657 -11354 18057 -11342
rect 17657 -11388 17669 -11354
rect 18045 -11388 18057 -11354
rect 17657 -11400 18057 -11388
rect 18293 -11354 18693 -11342
rect 18293 -11388 18305 -11354
rect 18681 -11388 18693 -11354
rect 18293 -11400 18693 -11388
rect 19257 -9970 19657 -9958
rect 19257 -10004 19269 -9970
rect 19645 -10004 19657 -9970
rect 19257 -10016 19657 -10004
rect 19893 -9970 20293 -9958
rect 19893 -10004 19905 -9970
rect 20281 -10004 20293 -9970
rect 19893 -10016 20293 -10004
rect 19257 -10228 19657 -10216
rect 19257 -10262 19269 -10228
rect 19645 -10262 19657 -10228
rect 19257 -10274 19657 -10262
rect 19893 -10228 20293 -10216
rect 19893 -10262 19905 -10228
rect 20281 -10262 20293 -10228
rect 19893 -10274 20293 -10262
rect 19257 -10496 19657 -10484
rect 19257 -10530 19269 -10496
rect 19645 -10530 19657 -10496
rect 19257 -10542 19657 -10530
rect 19893 -10496 20293 -10484
rect 19893 -10530 19905 -10496
rect 20281 -10530 20293 -10496
rect 19893 -10542 20293 -10530
rect 19257 -11354 19657 -11342
rect 19257 -11388 19269 -11354
rect 19645 -11388 19657 -11354
rect 19257 -11400 19657 -11388
rect 19893 -11354 20293 -11342
rect 19893 -11388 19905 -11354
rect 20281 -11388 20293 -11354
rect 19893 -11400 20293 -11388
rect 20857 -9970 21257 -9958
rect 20857 -10004 20869 -9970
rect 21245 -10004 21257 -9970
rect 20857 -10016 21257 -10004
rect 21493 -9970 21893 -9958
rect 21493 -10004 21505 -9970
rect 21881 -10004 21893 -9970
rect 21493 -10016 21893 -10004
rect 20857 -10228 21257 -10216
rect 20857 -10262 20869 -10228
rect 21245 -10262 21257 -10228
rect 20857 -10274 21257 -10262
rect 21493 -10228 21893 -10216
rect 21493 -10262 21505 -10228
rect 21881 -10262 21893 -10228
rect 21493 -10274 21893 -10262
rect 20857 -10496 21257 -10484
rect 20857 -10530 20869 -10496
rect 21245 -10530 21257 -10496
rect 20857 -10542 21257 -10530
rect 21493 -10496 21893 -10484
rect 21493 -10530 21505 -10496
rect 21881 -10530 21893 -10496
rect 21493 -10542 21893 -10530
rect 20857 -11354 21257 -11342
rect 20857 -11388 20869 -11354
rect 21245 -11388 21257 -11354
rect 20857 -11400 21257 -11388
rect 21493 -11354 21893 -11342
rect 21493 -11388 21505 -11354
rect 21881 -11388 21893 -11354
rect 21493 -11400 21893 -11388
rect 22457 -9970 22857 -9958
rect 22457 -10004 22469 -9970
rect 22845 -10004 22857 -9970
rect 22457 -10016 22857 -10004
rect 23093 -9970 23493 -9958
rect 23093 -10004 23105 -9970
rect 23481 -10004 23493 -9970
rect 23093 -10016 23493 -10004
rect 22457 -10228 22857 -10216
rect 22457 -10262 22469 -10228
rect 22845 -10262 22857 -10228
rect 22457 -10274 22857 -10262
rect 23093 -10228 23493 -10216
rect 23093 -10262 23105 -10228
rect 23481 -10262 23493 -10228
rect 23093 -10274 23493 -10262
rect 22457 -10496 22857 -10484
rect 22457 -10530 22469 -10496
rect 22845 -10530 22857 -10496
rect 22457 -10542 22857 -10530
rect 23093 -10496 23493 -10484
rect 23093 -10530 23105 -10496
rect 23481 -10530 23493 -10496
rect 23093 -10542 23493 -10530
rect 22457 -11354 22857 -11342
rect 22457 -11388 22469 -11354
rect 22845 -11388 22857 -11354
rect 22457 -11400 22857 -11388
rect 23093 -11354 23493 -11342
rect 23093 -11388 23105 -11354
rect 23481 -11388 23493 -11354
rect 23093 -11400 23493 -11388
rect 24057 -9970 24457 -9958
rect 24057 -10004 24069 -9970
rect 24445 -10004 24457 -9970
rect 24057 -10016 24457 -10004
rect 24693 -9970 25093 -9958
rect 24693 -10004 24705 -9970
rect 25081 -10004 25093 -9970
rect 24693 -10016 25093 -10004
rect 24057 -10228 24457 -10216
rect 24057 -10262 24069 -10228
rect 24445 -10262 24457 -10228
rect 24057 -10274 24457 -10262
rect 24693 -10228 25093 -10216
rect 24693 -10262 24705 -10228
rect 25081 -10262 25093 -10228
rect 24693 -10274 25093 -10262
rect 24057 -10496 24457 -10484
rect 24057 -10530 24069 -10496
rect 24445 -10530 24457 -10496
rect 24057 -10542 24457 -10530
rect 24693 -10496 25093 -10484
rect 24693 -10530 24705 -10496
rect 25081 -10530 25093 -10496
rect 24693 -10542 25093 -10530
rect 24057 -11354 24457 -11342
rect 24057 -11388 24069 -11354
rect 24445 -11388 24457 -11354
rect 24057 -11400 24457 -11388
rect 24693 -11354 25093 -11342
rect 24693 -11388 24705 -11354
rect 25081 -11388 25093 -11354
rect 24693 -11400 25093 -11388
rect 25657 -9970 26057 -9958
rect 25657 -10004 25669 -9970
rect 26045 -10004 26057 -9970
rect 25657 -10016 26057 -10004
rect 26293 -9970 26693 -9958
rect 26293 -10004 26305 -9970
rect 26681 -10004 26693 -9970
rect 26293 -10016 26693 -10004
rect 25657 -10228 26057 -10216
rect 25657 -10262 25669 -10228
rect 26045 -10262 26057 -10228
rect 25657 -10274 26057 -10262
rect 26293 -10228 26693 -10216
rect 26293 -10262 26305 -10228
rect 26681 -10262 26693 -10228
rect 26293 -10274 26693 -10262
rect 25657 -10496 26057 -10484
rect 25657 -10530 25669 -10496
rect 26045 -10530 26057 -10496
rect 25657 -10542 26057 -10530
rect 26293 -10496 26693 -10484
rect 26293 -10530 26305 -10496
rect 26681 -10530 26693 -10496
rect 26293 -10542 26693 -10530
rect 25657 -11354 26057 -11342
rect 25657 -11388 25669 -11354
rect 26045 -11388 26057 -11354
rect 25657 -11400 26057 -11388
rect 26293 -11354 26693 -11342
rect 26293 -11388 26305 -11354
rect 26681 -11388 26693 -11354
rect 26293 -11400 26693 -11388
rect 27257 -9970 27657 -9958
rect 27257 -10004 27269 -9970
rect 27645 -10004 27657 -9970
rect 27257 -10016 27657 -10004
rect 27893 -9970 28293 -9958
rect 27893 -10004 27905 -9970
rect 28281 -10004 28293 -9970
rect 27893 -10016 28293 -10004
rect 27257 -10228 27657 -10216
rect 27257 -10262 27269 -10228
rect 27645 -10262 27657 -10228
rect 27257 -10274 27657 -10262
rect 27893 -10228 28293 -10216
rect 27893 -10262 27905 -10228
rect 28281 -10262 28293 -10228
rect 27893 -10274 28293 -10262
rect 27257 -10496 27657 -10484
rect 27257 -10530 27269 -10496
rect 27645 -10530 27657 -10496
rect 27257 -10542 27657 -10530
rect 27893 -10496 28293 -10484
rect 27893 -10530 27905 -10496
rect 28281 -10530 28293 -10496
rect 27893 -10542 28293 -10530
rect 27257 -11354 27657 -11342
rect 27257 -11388 27269 -11354
rect 27645 -11388 27657 -11354
rect 27257 -11400 27657 -11388
rect 27893 -11354 28293 -11342
rect 27893 -11388 27905 -11354
rect 28281 -11388 28293 -11354
rect 27893 -11400 28293 -11388
rect 28857 -9970 29257 -9958
rect 28857 -10004 28869 -9970
rect 29245 -10004 29257 -9970
rect 28857 -10016 29257 -10004
rect 29493 -9970 29893 -9958
rect 29493 -10004 29505 -9970
rect 29881 -10004 29893 -9970
rect 29493 -10016 29893 -10004
rect 28857 -10228 29257 -10216
rect 28857 -10262 28869 -10228
rect 29245 -10262 29257 -10228
rect 28857 -10274 29257 -10262
rect 29493 -10228 29893 -10216
rect 29493 -10262 29505 -10228
rect 29881 -10262 29893 -10228
rect 29493 -10274 29893 -10262
rect 28857 -10496 29257 -10484
rect 28857 -10530 28869 -10496
rect 29245 -10530 29257 -10496
rect 28857 -10542 29257 -10530
rect 29493 -10496 29893 -10484
rect 29493 -10530 29505 -10496
rect 29881 -10530 29893 -10496
rect 29493 -10542 29893 -10530
rect 28857 -11354 29257 -11342
rect 28857 -11388 28869 -11354
rect 29245 -11388 29257 -11354
rect 28857 -11400 29257 -11388
rect 29493 -11354 29893 -11342
rect 29493 -11388 29505 -11354
rect 29881 -11388 29893 -11354
rect 29493 -11400 29893 -11388
rect 30457 -9970 30857 -9958
rect 30457 -10004 30469 -9970
rect 30845 -10004 30857 -9970
rect 30457 -10016 30857 -10004
rect 31093 -9970 31493 -9958
rect 31093 -10004 31105 -9970
rect 31481 -10004 31493 -9970
rect 31093 -10016 31493 -10004
rect 30457 -10228 30857 -10216
rect 30457 -10262 30469 -10228
rect 30845 -10262 30857 -10228
rect 30457 -10274 30857 -10262
rect 31093 -10228 31493 -10216
rect 31093 -10262 31105 -10228
rect 31481 -10262 31493 -10228
rect 31093 -10274 31493 -10262
rect 30457 -10496 30857 -10484
rect 30457 -10530 30469 -10496
rect 30845 -10530 30857 -10496
rect 30457 -10542 30857 -10530
rect 31093 -10496 31493 -10484
rect 31093 -10530 31105 -10496
rect 31481 -10530 31493 -10496
rect 31093 -10542 31493 -10530
rect 30457 -11354 30857 -11342
rect 30457 -11388 30469 -11354
rect 30845 -11388 30857 -11354
rect 30457 -11400 30857 -11388
rect 31093 -11354 31493 -11342
rect 31093 -11388 31105 -11354
rect 31481 -11388 31493 -11354
rect 31093 -11400 31493 -11388
rect 32057 -9970 32457 -9958
rect 32057 -10004 32069 -9970
rect 32445 -10004 32457 -9970
rect 32057 -10016 32457 -10004
rect 32693 -9970 33093 -9958
rect 32693 -10004 32705 -9970
rect 33081 -10004 33093 -9970
rect 32693 -10016 33093 -10004
rect 32057 -10228 32457 -10216
rect 32057 -10262 32069 -10228
rect 32445 -10262 32457 -10228
rect 32057 -10274 32457 -10262
rect 32693 -10228 33093 -10216
rect 32693 -10262 32705 -10228
rect 33081 -10262 33093 -10228
rect 32693 -10274 33093 -10262
rect 32057 -10496 32457 -10484
rect 32057 -10530 32069 -10496
rect 32445 -10530 32457 -10496
rect 32057 -10542 32457 -10530
rect 32693 -10496 33093 -10484
rect 32693 -10530 32705 -10496
rect 33081 -10530 33093 -10496
rect 32693 -10542 33093 -10530
rect 32057 -11354 32457 -11342
rect 32057 -11388 32069 -11354
rect 32445 -11388 32457 -11354
rect 32057 -11400 32457 -11388
rect 32693 -11354 33093 -11342
rect 32693 -11388 32705 -11354
rect 33081 -11388 33093 -11354
rect 32693 -11400 33093 -11388
rect 33657 -9970 34057 -9958
rect 33657 -10004 33669 -9970
rect 34045 -10004 34057 -9970
rect 33657 -10016 34057 -10004
rect 34293 -9970 34693 -9958
rect 34293 -10004 34305 -9970
rect 34681 -10004 34693 -9970
rect 34293 -10016 34693 -10004
rect 33657 -10228 34057 -10216
rect 33657 -10262 33669 -10228
rect 34045 -10262 34057 -10228
rect 33657 -10274 34057 -10262
rect 34293 -10228 34693 -10216
rect 34293 -10262 34305 -10228
rect 34681 -10262 34693 -10228
rect 34293 -10274 34693 -10262
rect 33657 -10496 34057 -10484
rect 33657 -10530 33669 -10496
rect 34045 -10530 34057 -10496
rect 33657 -10542 34057 -10530
rect 34293 -10496 34693 -10484
rect 34293 -10530 34305 -10496
rect 34681 -10530 34693 -10496
rect 34293 -10542 34693 -10530
rect 33657 -11354 34057 -11342
rect 33657 -11388 33669 -11354
rect 34045 -11388 34057 -11354
rect 33657 -11400 34057 -11388
rect 34293 -11354 34693 -11342
rect 34293 -11388 34305 -11354
rect 34681 -11388 34693 -11354
rect 34293 -11400 34693 -11388
rect 35257 -9970 35657 -9958
rect 35257 -10004 35269 -9970
rect 35645 -10004 35657 -9970
rect 35257 -10016 35657 -10004
rect 35893 -9970 36293 -9958
rect 35893 -10004 35905 -9970
rect 36281 -10004 36293 -9970
rect 35893 -10016 36293 -10004
rect 35257 -10228 35657 -10216
rect 35257 -10262 35269 -10228
rect 35645 -10262 35657 -10228
rect 35257 -10274 35657 -10262
rect 35893 -10228 36293 -10216
rect 35893 -10262 35905 -10228
rect 36281 -10262 36293 -10228
rect 35893 -10274 36293 -10262
rect 35257 -10496 35657 -10484
rect 35257 -10530 35269 -10496
rect 35645 -10530 35657 -10496
rect 35257 -10542 35657 -10530
rect 35893 -10496 36293 -10484
rect 35893 -10530 35905 -10496
rect 36281 -10530 36293 -10496
rect 35893 -10542 36293 -10530
rect 35257 -11354 35657 -11342
rect 35257 -11388 35269 -11354
rect 35645 -11388 35657 -11354
rect 35257 -11400 35657 -11388
rect 35893 -11354 36293 -11342
rect 35893 -11388 35905 -11354
rect 36281 -11388 36293 -11354
rect 35893 -11400 36293 -11388
rect 36857 -9970 37257 -9958
rect 36857 -10004 36869 -9970
rect 37245 -10004 37257 -9970
rect 36857 -10016 37257 -10004
rect 37493 -9970 37893 -9958
rect 37493 -10004 37505 -9970
rect 37881 -10004 37893 -9970
rect 37493 -10016 37893 -10004
rect 36857 -10228 37257 -10216
rect 36857 -10262 36869 -10228
rect 37245 -10262 37257 -10228
rect 36857 -10274 37257 -10262
rect 37493 -10228 37893 -10216
rect 37493 -10262 37505 -10228
rect 37881 -10262 37893 -10228
rect 37493 -10274 37893 -10262
rect 36857 -10496 37257 -10484
rect 36857 -10530 36869 -10496
rect 37245 -10530 37257 -10496
rect 36857 -10542 37257 -10530
rect 37493 -10496 37893 -10484
rect 37493 -10530 37505 -10496
rect 37881 -10530 37893 -10496
rect 37493 -10542 37893 -10530
rect 36857 -11354 37257 -11342
rect 36857 -11388 36869 -11354
rect 37245 -11388 37257 -11354
rect 36857 -11400 37257 -11388
rect 37493 -11354 37893 -11342
rect 37493 -11388 37505 -11354
rect 37881 -11388 37893 -11354
rect 37493 -11400 37893 -11388
rect 57 -11770 457 -11758
rect 57 -11804 69 -11770
rect 445 -11804 457 -11770
rect 57 -11816 457 -11804
rect 693 -11770 1093 -11758
rect 693 -11804 705 -11770
rect 1081 -11804 1093 -11770
rect 693 -11816 1093 -11804
rect 57 -12028 457 -12016
rect 57 -12062 69 -12028
rect 445 -12062 457 -12028
rect 57 -12074 457 -12062
rect 693 -12028 1093 -12016
rect 693 -12062 705 -12028
rect 1081 -12062 1093 -12028
rect 693 -12074 1093 -12062
rect 57 -12296 457 -12284
rect 57 -12330 69 -12296
rect 445 -12330 457 -12296
rect 57 -12342 457 -12330
rect 693 -12296 1093 -12284
rect 693 -12330 705 -12296
rect 1081 -12330 1093 -12296
rect 693 -12342 1093 -12330
rect 57 -13154 457 -13142
rect 57 -13188 69 -13154
rect 445 -13188 457 -13154
rect 57 -13200 457 -13188
rect 693 -13154 1093 -13142
rect 693 -13188 705 -13154
rect 1081 -13188 1093 -13154
rect 693 -13200 1093 -13188
rect 1657 -11770 2057 -11758
rect 1657 -11804 1669 -11770
rect 2045 -11804 2057 -11770
rect 1657 -11816 2057 -11804
rect 2293 -11770 2693 -11758
rect 2293 -11804 2305 -11770
rect 2681 -11804 2693 -11770
rect 2293 -11816 2693 -11804
rect 1657 -12028 2057 -12016
rect 1657 -12062 1669 -12028
rect 2045 -12062 2057 -12028
rect 1657 -12074 2057 -12062
rect 2293 -12028 2693 -12016
rect 2293 -12062 2305 -12028
rect 2681 -12062 2693 -12028
rect 2293 -12074 2693 -12062
rect 1657 -12296 2057 -12284
rect 1657 -12330 1669 -12296
rect 2045 -12330 2057 -12296
rect 1657 -12342 2057 -12330
rect 2293 -12296 2693 -12284
rect 2293 -12330 2305 -12296
rect 2681 -12330 2693 -12296
rect 2293 -12342 2693 -12330
rect 1657 -13154 2057 -13142
rect 1657 -13188 1669 -13154
rect 2045 -13188 2057 -13154
rect 1657 -13200 2057 -13188
rect 2293 -13154 2693 -13142
rect 2293 -13188 2305 -13154
rect 2681 -13188 2693 -13154
rect 2293 -13200 2693 -13188
rect 3257 -11770 3657 -11758
rect 3257 -11804 3269 -11770
rect 3645 -11804 3657 -11770
rect 3257 -11816 3657 -11804
rect 3893 -11770 4293 -11758
rect 3893 -11804 3905 -11770
rect 4281 -11804 4293 -11770
rect 3893 -11816 4293 -11804
rect 3257 -12028 3657 -12016
rect 3257 -12062 3269 -12028
rect 3645 -12062 3657 -12028
rect 3257 -12074 3657 -12062
rect 3893 -12028 4293 -12016
rect 3893 -12062 3905 -12028
rect 4281 -12062 4293 -12028
rect 3893 -12074 4293 -12062
rect 3257 -12296 3657 -12284
rect 3257 -12330 3269 -12296
rect 3645 -12330 3657 -12296
rect 3257 -12342 3657 -12330
rect 3893 -12296 4293 -12284
rect 3893 -12330 3905 -12296
rect 4281 -12330 4293 -12296
rect 3893 -12342 4293 -12330
rect 3257 -13154 3657 -13142
rect 3257 -13188 3269 -13154
rect 3645 -13188 3657 -13154
rect 3257 -13200 3657 -13188
rect 3893 -13154 4293 -13142
rect 3893 -13188 3905 -13154
rect 4281 -13188 4293 -13154
rect 3893 -13200 4293 -13188
rect 4857 -11770 5257 -11758
rect 4857 -11804 4869 -11770
rect 5245 -11804 5257 -11770
rect 4857 -11816 5257 -11804
rect 5493 -11770 5893 -11758
rect 5493 -11804 5505 -11770
rect 5881 -11804 5893 -11770
rect 5493 -11816 5893 -11804
rect 4857 -12028 5257 -12016
rect 4857 -12062 4869 -12028
rect 5245 -12062 5257 -12028
rect 4857 -12074 5257 -12062
rect 5493 -12028 5893 -12016
rect 5493 -12062 5505 -12028
rect 5881 -12062 5893 -12028
rect 5493 -12074 5893 -12062
rect 4857 -12296 5257 -12284
rect 4857 -12330 4869 -12296
rect 5245 -12330 5257 -12296
rect 4857 -12342 5257 -12330
rect 5493 -12296 5893 -12284
rect 5493 -12330 5505 -12296
rect 5881 -12330 5893 -12296
rect 5493 -12342 5893 -12330
rect 4857 -13154 5257 -13142
rect 4857 -13188 4869 -13154
rect 5245 -13188 5257 -13154
rect 4857 -13200 5257 -13188
rect 5493 -13154 5893 -13142
rect 5493 -13188 5505 -13154
rect 5881 -13188 5893 -13154
rect 5493 -13200 5893 -13188
rect 6457 -11770 6857 -11758
rect 6457 -11804 6469 -11770
rect 6845 -11804 6857 -11770
rect 6457 -11816 6857 -11804
rect 7093 -11770 7493 -11758
rect 7093 -11804 7105 -11770
rect 7481 -11804 7493 -11770
rect 7093 -11816 7493 -11804
rect 6457 -12028 6857 -12016
rect 6457 -12062 6469 -12028
rect 6845 -12062 6857 -12028
rect 6457 -12074 6857 -12062
rect 7093 -12028 7493 -12016
rect 7093 -12062 7105 -12028
rect 7481 -12062 7493 -12028
rect 7093 -12074 7493 -12062
rect 6457 -12296 6857 -12284
rect 6457 -12330 6469 -12296
rect 6845 -12330 6857 -12296
rect 6457 -12342 6857 -12330
rect 7093 -12296 7493 -12284
rect 7093 -12330 7105 -12296
rect 7481 -12330 7493 -12296
rect 7093 -12342 7493 -12330
rect 6457 -13154 6857 -13142
rect 6457 -13188 6469 -13154
rect 6845 -13188 6857 -13154
rect 6457 -13200 6857 -13188
rect 7093 -13154 7493 -13142
rect 7093 -13188 7105 -13154
rect 7481 -13188 7493 -13154
rect 7093 -13200 7493 -13188
rect 8057 -11770 8457 -11758
rect 8057 -11804 8069 -11770
rect 8445 -11804 8457 -11770
rect 8057 -11816 8457 -11804
rect 8693 -11770 9093 -11758
rect 8693 -11804 8705 -11770
rect 9081 -11804 9093 -11770
rect 8693 -11816 9093 -11804
rect 8057 -12028 8457 -12016
rect 8057 -12062 8069 -12028
rect 8445 -12062 8457 -12028
rect 8057 -12074 8457 -12062
rect 8693 -12028 9093 -12016
rect 8693 -12062 8705 -12028
rect 9081 -12062 9093 -12028
rect 8693 -12074 9093 -12062
rect 8057 -12296 8457 -12284
rect 8057 -12330 8069 -12296
rect 8445 -12330 8457 -12296
rect 8057 -12342 8457 -12330
rect 8693 -12296 9093 -12284
rect 8693 -12330 8705 -12296
rect 9081 -12330 9093 -12296
rect 8693 -12342 9093 -12330
rect 8057 -13154 8457 -13142
rect 8057 -13188 8069 -13154
rect 8445 -13188 8457 -13154
rect 8057 -13200 8457 -13188
rect 8693 -13154 9093 -13142
rect 8693 -13188 8705 -13154
rect 9081 -13188 9093 -13154
rect 8693 -13200 9093 -13188
rect 9657 -11770 10057 -11758
rect 9657 -11804 9669 -11770
rect 10045 -11804 10057 -11770
rect 9657 -11816 10057 -11804
rect 10293 -11770 10693 -11758
rect 10293 -11804 10305 -11770
rect 10681 -11804 10693 -11770
rect 10293 -11816 10693 -11804
rect 9657 -12028 10057 -12016
rect 9657 -12062 9669 -12028
rect 10045 -12062 10057 -12028
rect 9657 -12074 10057 -12062
rect 10293 -12028 10693 -12016
rect 10293 -12062 10305 -12028
rect 10681 -12062 10693 -12028
rect 10293 -12074 10693 -12062
rect 9657 -12296 10057 -12284
rect 9657 -12330 9669 -12296
rect 10045 -12330 10057 -12296
rect 9657 -12342 10057 -12330
rect 10293 -12296 10693 -12284
rect 10293 -12330 10305 -12296
rect 10681 -12330 10693 -12296
rect 10293 -12342 10693 -12330
rect 9657 -13154 10057 -13142
rect 9657 -13188 9669 -13154
rect 10045 -13188 10057 -13154
rect 9657 -13200 10057 -13188
rect 10293 -13154 10693 -13142
rect 10293 -13188 10305 -13154
rect 10681 -13188 10693 -13154
rect 10293 -13200 10693 -13188
rect 11257 -11770 11657 -11758
rect 11257 -11804 11269 -11770
rect 11645 -11804 11657 -11770
rect 11257 -11816 11657 -11804
rect 11893 -11770 12293 -11758
rect 11893 -11804 11905 -11770
rect 12281 -11804 12293 -11770
rect 11893 -11816 12293 -11804
rect 11257 -12028 11657 -12016
rect 11257 -12062 11269 -12028
rect 11645 -12062 11657 -12028
rect 11257 -12074 11657 -12062
rect 11893 -12028 12293 -12016
rect 11893 -12062 11905 -12028
rect 12281 -12062 12293 -12028
rect 11893 -12074 12293 -12062
rect 11257 -12296 11657 -12284
rect 11257 -12330 11269 -12296
rect 11645 -12330 11657 -12296
rect 11257 -12342 11657 -12330
rect 11893 -12296 12293 -12284
rect 11893 -12330 11905 -12296
rect 12281 -12330 12293 -12296
rect 11893 -12342 12293 -12330
rect 11257 -13154 11657 -13142
rect 11257 -13188 11269 -13154
rect 11645 -13188 11657 -13154
rect 11257 -13200 11657 -13188
rect 11893 -13154 12293 -13142
rect 11893 -13188 11905 -13154
rect 12281 -13188 12293 -13154
rect 11893 -13200 12293 -13188
rect 12857 -11770 13257 -11758
rect 12857 -11804 12869 -11770
rect 13245 -11804 13257 -11770
rect 12857 -11816 13257 -11804
rect 13493 -11770 13893 -11758
rect 13493 -11804 13505 -11770
rect 13881 -11804 13893 -11770
rect 13493 -11816 13893 -11804
rect 12857 -12028 13257 -12016
rect 12857 -12062 12869 -12028
rect 13245 -12062 13257 -12028
rect 12857 -12074 13257 -12062
rect 13493 -12028 13893 -12016
rect 13493 -12062 13505 -12028
rect 13881 -12062 13893 -12028
rect 13493 -12074 13893 -12062
rect 12857 -12296 13257 -12284
rect 12857 -12330 12869 -12296
rect 13245 -12330 13257 -12296
rect 12857 -12342 13257 -12330
rect 13493 -12296 13893 -12284
rect 13493 -12330 13505 -12296
rect 13881 -12330 13893 -12296
rect 13493 -12342 13893 -12330
rect 12857 -13154 13257 -13142
rect 12857 -13188 12869 -13154
rect 13245 -13188 13257 -13154
rect 12857 -13200 13257 -13188
rect 13493 -13154 13893 -13142
rect 13493 -13188 13505 -13154
rect 13881 -13188 13893 -13154
rect 13493 -13200 13893 -13188
rect 14457 -11770 14857 -11758
rect 14457 -11804 14469 -11770
rect 14845 -11804 14857 -11770
rect 14457 -11816 14857 -11804
rect 15093 -11770 15493 -11758
rect 15093 -11804 15105 -11770
rect 15481 -11804 15493 -11770
rect 15093 -11816 15493 -11804
rect 14457 -12028 14857 -12016
rect 14457 -12062 14469 -12028
rect 14845 -12062 14857 -12028
rect 14457 -12074 14857 -12062
rect 15093 -12028 15493 -12016
rect 15093 -12062 15105 -12028
rect 15481 -12062 15493 -12028
rect 15093 -12074 15493 -12062
rect 14457 -12296 14857 -12284
rect 14457 -12330 14469 -12296
rect 14845 -12330 14857 -12296
rect 14457 -12342 14857 -12330
rect 15093 -12296 15493 -12284
rect 15093 -12330 15105 -12296
rect 15481 -12330 15493 -12296
rect 15093 -12342 15493 -12330
rect 14457 -13154 14857 -13142
rect 14457 -13188 14469 -13154
rect 14845 -13188 14857 -13154
rect 14457 -13200 14857 -13188
rect 15093 -13154 15493 -13142
rect 15093 -13188 15105 -13154
rect 15481 -13188 15493 -13154
rect 15093 -13200 15493 -13188
rect 16057 -11770 16457 -11758
rect 16057 -11804 16069 -11770
rect 16445 -11804 16457 -11770
rect 16057 -11816 16457 -11804
rect 16693 -11770 17093 -11758
rect 16693 -11804 16705 -11770
rect 17081 -11804 17093 -11770
rect 16693 -11816 17093 -11804
rect 16057 -12028 16457 -12016
rect 16057 -12062 16069 -12028
rect 16445 -12062 16457 -12028
rect 16057 -12074 16457 -12062
rect 16693 -12028 17093 -12016
rect 16693 -12062 16705 -12028
rect 17081 -12062 17093 -12028
rect 16693 -12074 17093 -12062
rect 16057 -12296 16457 -12284
rect 16057 -12330 16069 -12296
rect 16445 -12330 16457 -12296
rect 16057 -12342 16457 -12330
rect 16693 -12296 17093 -12284
rect 16693 -12330 16705 -12296
rect 17081 -12330 17093 -12296
rect 16693 -12342 17093 -12330
rect 16057 -13154 16457 -13142
rect 16057 -13188 16069 -13154
rect 16445 -13188 16457 -13154
rect 16057 -13200 16457 -13188
rect 16693 -13154 17093 -13142
rect 16693 -13188 16705 -13154
rect 17081 -13188 17093 -13154
rect 16693 -13200 17093 -13188
rect 17657 -11770 18057 -11758
rect 17657 -11804 17669 -11770
rect 18045 -11804 18057 -11770
rect 17657 -11816 18057 -11804
rect 18293 -11770 18693 -11758
rect 18293 -11804 18305 -11770
rect 18681 -11804 18693 -11770
rect 18293 -11816 18693 -11804
rect 17657 -12028 18057 -12016
rect 17657 -12062 17669 -12028
rect 18045 -12062 18057 -12028
rect 17657 -12074 18057 -12062
rect 18293 -12028 18693 -12016
rect 18293 -12062 18305 -12028
rect 18681 -12062 18693 -12028
rect 18293 -12074 18693 -12062
rect 17657 -12296 18057 -12284
rect 17657 -12330 17669 -12296
rect 18045 -12330 18057 -12296
rect 17657 -12342 18057 -12330
rect 18293 -12296 18693 -12284
rect 18293 -12330 18305 -12296
rect 18681 -12330 18693 -12296
rect 18293 -12342 18693 -12330
rect 17657 -13154 18057 -13142
rect 17657 -13188 17669 -13154
rect 18045 -13188 18057 -13154
rect 17657 -13200 18057 -13188
rect 18293 -13154 18693 -13142
rect 18293 -13188 18305 -13154
rect 18681 -13188 18693 -13154
rect 18293 -13200 18693 -13188
rect 19257 -11770 19657 -11758
rect 19257 -11804 19269 -11770
rect 19645 -11804 19657 -11770
rect 19257 -11816 19657 -11804
rect 19893 -11770 20293 -11758
rect 19893 -11804 19905 -11770
rect 20281 -11804 20293 -11770
rect 19893 -11816 20293 -11804
rect 19257 -12028 19657 -12016
rect 19257 -12062 19269 -12028
rect 19645 -12062 19657 -12028
rect 19257 -12074 19657 -12062
rect 19893 -12028 20293 -12016
rect 19893 -12062 19905 -12028
rect 20281 -12062 20293 -12028
rect 19893 -12074 20293 -12062
rect 19257 -12296 19657 -12284
rect 19257 -12330 19269 -12296
rect 19645 -12330 19657 -12296
rect 19257 -12342 19657 -12330
rect 19893 -12296 20293 -12284
rect 19893 -12330 19905 -12296
rect 20281 -12330 20293 -12296
rect 19893 -12342 20293 -12330
rect 19257 -13154 19657 -13142
rect 19257 -13188 19269 -13154
rect 19645 -13188 19657 -13154
rect 19257 -13200 19657 -13188
rect 19893 -13154 20293 -13142
rect 19893 -13188 19905 -13154
rect 20281 -13188 20293 -13154
rect 19893 -13200 20293 -13188
rect 20857 -11770 21257 -11758
rect 20857 -11804 20869 -11770
rect 21245 -11804 21257 -11770
rect 20857 -11816 21257 -11804
rect 21493 -11770 21893 -11758
rect 21493 -11804 21505 -11770
rect 21881 -11804 21893 -11770
rect 21493 -11816 21893 -11804
rect 20857 -12028 21257 -12016
rect 20857 -12062 20869 -12028
rect 21245 -12062 21257 -12028
rect 20857 -12074 21257 -12062
rect 21493 -12028 21893 -12016
rect 21493 -12062 21505 -12028
rect 21881 -12062 21893 -12028
rect 21493 -12074 21893 -12062
rect 20857 -12296 21257 -12284
rect 20857 -12330 20869 -12296
rect 21245 -12330 21257 -12296
rect 20857 -12342 21257 -12330
rect 21493 -12296 21893 -12284
rect 21493 -12330 21505 -12296
rect 21881 -12330 21893 -12296
rect 21493 -12342 21893 -12330
rect 20857 -13154 21257 -13142
rect 20857 -13188 20869 -13154
rect 21245 -13188 21257 -13154
rect 20857 -13200 21257 -13188
rect 21493 -13154 21893 -13142
rect 21493 -13188 21505 -13154
rect 21881 -13188 21893 -13154
rect 21493 -13200 21893 -13188
rect 22457 -11770 22857 -11758
rect 22457 -11804 22469 -11770
rect 22845 -11804 22857 -11770
rect 22457 -11816 22857 -11804
rect 23093 -11770 23493 -11758
rect 23093 -11804 23105 -11770
rect 23481 -11804 23493 -11770
rect 23093 -11816 23493 -11804
rect 22457 -12028 22857 -12016
rect 22457 -12062 22469 -12028
rect 22845 -12062 22857 -12028
rect 22457 -12074 22857 -12062
rect 23093 -12028 23493 -12016
rect 23093 -12062 23105 -12028
rect 23481 -12062 23493 -12028
rect 23093 -12074 23493 -12062
rect 22457 -12296 22857 -12284
rect 22457 -12330 22469 -12296
rect 22845 -12330 22857 -12296
rect 22457 -12342 22857 -12330
rect 23093 -12296 23493 -12284
rect 23093 -12330 23105 -12296
rect 23481 -12330 23493 -12296
rect 23093 -12342 23493 -12330
rect 22457 -13154 22857 -13142
rect 22457 -13188 22469 -13154
rect 22845 -13188 22857 -13154
rect 22457 -13200 22857 -13188
rect 23093 -13154 23493 -13142
rect 23093 -13188 23105 -13154
rect 23481 -13188 23493 -13154
rect 23093 -13200 23493 -13188
rect 24057 -11770 24457 -11758
rect 24057 -11804 24069 -11770
rect 24445 -11804 24457 -11770
rect 24057 -11816 24457 -11804
rect 24693 -11770 25093 -11758
rect 24693 -11804 24705 -11770
rect 25081 -11804 25093 -11770
rect 24693 -11816 25093 -11804
rect 24057 -12028 24457 -12016
rect 24057 -12062 24069 -12028
rect 24445 -12062 24457 -12028
rect 24057 -12074 24457 -12062
rect 24693 -12028 25093 -12016
rect 24693 -12062 24705 -12028
rect 25081 -12062 25093 -12028
rect 24693 -12074 25093 -12062
rect 24057 -12296 24457 -12284
rect 24057 -12330 24069 -12296
rect 24445 -12330 24457 -12296
rect 24057 -12342 24457 -12330
rect 24693 -12296 25093 -12284
rect 24693 -12330 24705 -12296
rect 25081 -12330 25093 -12296
rect 24693 -12342 25093 -12330
rect 24057 -13154 24457 -13142
rect 24057 -13188 24069 -13154
rect 24445 -13188 24457 -13154
rect 24057 -13200 24457 -13188
rect 24693 -13154 25093 -13142
rect 24693 -13188 24705 -13154
rect 25081 -13188 25093 -13154
rect 24693 -13200 25093 -13188
rect 25657 -11770 26057 -11758
rect 25657 -11804 25669 -11770
rect 26045 -11804 26057 -11770
rect 25657 -11816 26057 -11804
rect 26293 -11770 26693 -11758
rect 26293 -11804 26305 -11770
rect 26681 -11804 26693 -11770
rect 26293 -11816 26693 -11804
rect 25657 -12028 26057 -12016
rect 25657 -12062 25669 -12028
rect 26045 -12062 26057 -12028
rect 25657 -12074 26057 -12062
rect 26293 -12028 26693 -12016
rect 26293 -12062 26305 -12028
rect 26681 -12062 26693 -12028
rect 26293 -12074 26693 -12062
rect 25657 -12296 26057 -12284
rect 25657 -12330 25669 -12296
rect 26045 -12330 26057 -12296
rect 25657 -12342 26057 -12330
rect 26293 -12296 26693 -12284
rect 26293 -12330 26305 -12296
rect 26681 -12330 26693 -12296
rect 26293 -12342 26693 -12330
rect 25657 -13154 26057 -13142
rect 25657 -13188 25669 -13154
rect 26045 -13188 26057 -13154
rect 25657 -13200 26057 -13188
rect 26293 -13154 26693 -13142
rect 26293 -13188 26305 -13154
rect 26681 -13188 26693 -13154
rect 26293 -13200 26693 -13188
rect 27257 -11770 27657 -11758
rect 27257 -11804 27269 -11770
rect 27645 -11804 27657 -11770
rect 27257 -11816 27657 -11804
rect 27893 -11770 28293 -11758
rect 27893 -11804 27905 -11770
rect 28281 -11804 28293 -11770
rect 27893 -11816 28293 -11804
rect 27257 -12028 27657 -12016
rect 27257 -12062 27269 -12028
rect 27645 -12062 27657 -12028
rect 27257 -12074 27657 -12062
rect 27893 -12028 28293 -12016
rect 27893 -12062 27905 -12028
rect 28281 -12062 28293 -12028
rect 27893 -12074 28293 -12062
rect 27257 -12296 27657 -12284
rect 27257 -12330 27269 -12296
rect 27645 -12330 27657 -12296
rect 27257 -12342 27657 -12330
rect 27893 -12296 28293 -12284
rect 27893 -12330 27905 -12296
rect 28281 -12330 28293 -12296
rect 27893 -12342 28293 -12330
rect 27257 -13154 27657 -13142
rect 27257 -13188 27269 -13154
rect 27645 -13188 27657 -13154
rect 27257 -13200 27657 -13188
rect 27893 -13154 28293 -13142
rect 27893 -13188 27905 -13154
rect 28281 -13188 28293 -13154
rect 27893 -13200 28293 -13188
rect 28857 -11770 29257 -11758
rect 28857 -11804 28869 -11770
rect 29245 -11804 29257 -11770
rect 28857 -11816 29257 -11804
rect 29493 -11770 29893 -11758
rect 29493 -11804 29505 -11770
rect 29881 -11804 29893 -11770
rect 29493 -11816 29893 -11804
rect 28857 -12028 29257 -12016
rect 28857 -12062 28869 -12028
rect 29245 -12062 29257 -12028
rect 28857 -12074 29257 -12062
rect 29493 -12028 29893 -12016
rect 29493 -12062 29505 -12028
rect 29881 -12062 29893 -12028
rect 29493 -12074 29893 -12062
rect 28857 -12296 29257 -12284
rect 28857 -12330 28869 -12296
rect 29245 -12330 29257 -12296
rect 28857 -12342 29257 -12330
rect 29493 -12296 29893 -12284
rect 29493 -12330 29505 -12296
rect 29881 -12330 29893 -12296
rect 29493 -12342 29893 -12330
rect 28857 -13154 29257 -13142
rect 28857 -13188 28869 -13154
rect 29245 -13188 29257 -13154
rect 28857 -13200 29257 -13188
rect 29493 -13154 29893 -13142
rect 29493 -13188 29505 -13154
rect 29881 -13188 29893 -13154
rect 29493 -13200 29893 -13188
rect 30457 -11770 30857 -11758
rect 30457 -11804 30469 -11770
rect 30845 -11804 30857 -11770
rect 30457 -11816 30857 -11804
rect 31093 -11770 31493 -11758
rect 31093 -11804 31105 -11770
rect 31481 -11804 31493 -11770
rect 31093 -11816 31493 -11804
rect 30457 -12028 30857 -12016
rect 30457 -12062 30469 -12028
rect 30845 -12062 30857 -12028
rect 30457 -12074 30857 -12062
rect 31093 -12028 31493 -12016
rect 31093 -12062 31105 -12028
rect 31481 -12062 31493 -12028
rect 31093 -12074 31493 -12062
rect 30457 -12296 30857 -12284
rect 30457 -12330 30469 -12296
rect 30845 -12330 30857 -12296
rect 30457 -12342 30857 -12330
rect 31093 -12296 31493 -12284
rect 31093 -12330 31105 -12296
rect 31481 -12330 31493 -12296
rect 31093 -12342 31493 -12330
rect 30457 -13154 30857 -13142
rect 30457 -13188 30469 -13154
rect 30845 -13188 30857 -13154
rect 30457 -13200 30857 -13188
rect 31093 -13154 31493 -13142
rect 31093 -13188 31105 -13154
rect 31481 -13188 31493 -13154
rect 31093 -13200 31493 -13188
rect 32057 -11770 32457 -11758
rect 32057 -11804 32069 -11770
rect 32445 -11804 32457 -11770
rect 32057 -11816 32457 -11804
rect 32693 -11770 33093 -11758
rect 32693 -11804 32705 -11770
rect 33081 -11804 33093 -11770
rect 32693 -11816 33093 -11804
rect 32057 -12028 32457 -12016
rect 32057 -12062 32069 -12028
rect 32445 -12062 32457 -12028
rect 32057 -12074 32457 -12062
rect 32693 -12028 33093 -12016
rect 32693 -12062 32705 -12028
rect 33081 -12062 33093 -12028
rect 32693 -12074 33093 -12062
rect 32057 -12296 32457 -12284
rect 32057 -12330 32069 -12296
rect 32445 -12330 32457 -12296
rect 32057 -12342 32457 -12330
rect 32693 -12296 33093 -12284
rect 32693 -12330 32705 -12296
rect 33081 -12330 33093 -12296
rect 32693 -12342 33093 -12330
rect 32057 -13154 32457 -13142
rect 32057 -13188 32069 -13154
rect 32445 -13188 32457 -13154
rect 32057 -13200 32457 -13188
rect 32693 -13154 33093 -13142
rect 32693 -13188 32705 -13154
rect 33081 -13188 33093 -13154
rect 32693 -13200 33093 -13188
rect 33657 -11770 34057 -11758
rect 33657 -11804 33669 -11770
rect 34045 -11804 34057 -11770
rect 33657 -11816 34057 -11804
rect 34293 -11770 34693 -11758
rect 34293 -11804 34305 -11770
rect 34681 -11804 34693 -11770
rect 34293 -11816 34693 -11804
rect 33657 -12028 34057 -12016
rect 33657 -12062 33669 -12028
rect 34045 -12062 34057 -12028
rect 33657 -12074 34057 -12062
rect 34293 -12028 34693 -12016
rect 34293 -12062 34305 -12028
rect 34681 -12062 34693 -12028
rect 34293 -12074 34693 -12062
rect 33657 -12296 34057 -12284
rect 33657 -12330 33669 -12296
rect 34045 -12330 34057 -12296
rect 33657 -12342 34057 -12330
rect 34293 -12296 34693 -12284
rect 34293 -12330 34305 -12296
rect 34681 -12330 34693 -12296
rect 34293 -12342 34693 -12330
rect 33657 -13154 34057 -13142
rect 33657 -13188 33669 -13154
rect 34045 -13188 34057 -13154
rect 33657 -13200 34057 -13188
rect 34293 -13154 34693 -13142
rect 34293 -13188 34305 -13154
rect 34681 -13188 34693 -13154
rect 34293 -13200 34693 -13188
rect 35257 -11770 35657 -11758
rect 35257 -11804 35269 -11770
rect 35645 -11804 35657 -11770
rect 35257 -11816 35657 -11804
rect 35893 -11770 36293 -11758
rect 35893 -11804 35905 -11770
rect 36281 -11804 36293 -11770
rect 35893 -11816 36293 -11804
rect 35257 -12028 35657 -12016
rect 35257 -12062 35269 -12028
rect 35645 -12062 35657 -12028
rect 35257 -12074 35657 -12062
rect 35893 -12028 36293 -12016
rect 35893 -12062 35905 -12028
rect 36281 -12062 36293 -12028
rect 35893 -12074 36293 -12062
rect 35257 -12296 35657 -12284
rect 35257 -12330 35269 -12296
rect 35645 -12330 35657 -12296
rect 35257 -12342 35657 -12330
rect 35893 -12296 36293 -12284
rect 35893 -12330 35905 -12296
rect 36281 -12330 36293 -12296
rect 35893 -12342 36293 -12330
rect 35257 -13154 35657 -13142
rect 35257 -13188 35269 -13154
rect 35645 -13188 35657 -13154
rect 35257 -13200 35657 -13188
rect 35893 -13154 36293 -13142
rect 35893 -13188 35905 -13154
rect 36281 -13188 36293 -13154
rect 35893 -13200 36293 -13188
rect 36857 -11770 37257 -11758
rect 36857 -11804 36869 -11770
rect 37245 -11804 37257 -11770
rect 36857 -11816 37257 -11804
rect 37493 -11770 37893 -11758
rect 37493 -11804 37505 -11770
rect 37881 -11804 37893 -11770
rect 37493 -11816 37893 -11804
rect 36857 -12028 37257 -12016
rect 36857 -12062 36869 -12028
rect 37245 -12062 37257 -12028
rect 36857 -12074 37257 -12062
rect 37493 -12028 37893 -12016
rect 37493 -12062 37505 -12028
rect 37881 -12062 37893 -12028
rect 37493 -12074 37893 -12062
rect 36857 -12296 37257 -12284
rect 36857 -12330 36869 -12296
rect 37245 -12330 37257 -12296
rect 36857 -12342 37257 -12330
rect 37493 -12296 37893 -12284
rect 37493 -12330 37505 -12296
rect 37881 -12330 37893 -12296
rect 37493 -12342 37893 -12330
rect 36857 -13154 37257 -13142
rect 36857 -13188 36869 -13154
rect 37245 -13188 37257 -13154
rect 36857 -13200 37257 -13188
rect 37493 -13154 37893 -13142
rect 37493 -13188 37505 -13154
rect 37881 -13188 37893 -13154
rect 37493 -13200 37893 -13188
rect 57 -13570 457 -13558
rect 57 -13604 69 -13570
rect 445 -13604 457 -13570
rect 57 -13616 457 -13604
rect 693 -13570 1093 -13558
rect 693 -13604 705 -13570
rect 1081 -13604 1093 -13570
rect 693 -13616 1093 -13604
rect 57 -13828 457 -13816
rect 57 -13862 69 -13828
rect 445 -13862 457 -13828
rect 57 -13874 457 -13862
rect 693 -13828 1093 -13816
rect 693 -13862 705 -13828
rect 1081 -13862 1093 -13828
rect 693 -13874 1093 -13862
rect 57 -14096 457 -14084
rect 57 -14130 69 -14096
rect 445 -14130 457 -14096
rect 57 -14142 457 -14130
rect 693 -14096 1093 -14084
rect 693 -14130 705 -14096
rect 1081 -14130 1093 -14096
rect 693 -14142 1093 -14130
rect 57 -14954 457 -14942
rect 57 -14988 69 -14954
rect 445 -14988 457 -14954
rect 57 -15000 457 -14988
rect 693 -14954 1093 -14942
rect 693 -14988 705 -14954
rect 1081 -14988 1093 -14954
rect 693 -15000 1093 -14988
rect 1657 -13570 2057 -13558
rect 1657 -13604 1669 -13570
rect 2045 -13604 2057 -13570
rect 1657 -13616 2057 -13604
rect 2293 -13570 2693 -13558
rect 2293 -13604 2305 -13570
rect 2681 -13604 2693 -13570
rect 2293 -13616 2693 -13604
rect 1657 -13828 2057 -13816
rect 1657 -13862 1669 -13828
rect 2045 -13862 2057 -13828
rect 1657 -13874 2057 -13862
rect 2293 -13828 2693 -13816
rect 2293 -13862 2305 -13828
rect 2681 -13862 2693 -13828
rect 2293 -13874 2693 -13862
rect 1657 -14096 2057 -14084
rect 1657 -14130 1669 -14096
rect 2045 -14130 2057 -14096
rect 1657 -14142 2057 -14130
rect 2293 -14096 2693 -14084
rect 2293 -14130 2305 -14096
rect 2681 -14130 2693 -14096
rect 2293 -14142 2693 -14130
rect 1657 -14954 2057 -14942
rect 1657 -14988 1669 -14954
rect 2045 -14988 2057 -14954
rect 1657 -15000 2057 -14988
rect 2293 -14954 2693 -14942
rect 2293 -14988 2305 -14954
rect 2681 -14988 2693 -14954
rect 2293 -15000 2693 -14988
rect 3257 -13570 3657 -13558
rect 3257 -13604 3269 -13570
rect 3645 -13604 3657 -13570
rect 3257 -13616 3657 -13604
rect 3893 -13570 4293 -13558
rect 3893 -13604 3905 -13570
rect 4281 -13604 4293 -13570
rect 3893 -13616 4293 -13604
rect 3257 -13828 3657 -13816
rect 3257 -13862 3269 -13828
rect 3645 -13862 3657 -13828
rect 3257 -13874 3657 -13862
rect 3893 -13828 4293 -13816
rect 3893 -13862 3905 -13828
rect 4281 -13862 4293 -13828
rect 3893 -13874 4293 -13862
rect 3257 -14096 3657 -14084
rect 3257 -14130 3269 -14096
rect 3645 -14130 3657 -14096
rect 3257 -14142 3657 -14130
rect 3893 -14096 4293 -14084
rect 3893 -14130 3905 -14096
rect 4281 -14130 4293 -14096
rect 3893 -14142 4293 -14130
rect 3257 -14954 3657 -14942
rect 3257 -14988 3269 -14954
rect 3645 -14988 3657 -14954
rect 3257 -15000 3657 -14988
rect 3893 -14954 4293 -14942
rect 3893 -14988 3905 -14954
rect 4281 -14988 4293 -14954
rect 3893 -15000 4293 -14988
rect 4857 -13570 5257 -13558
rect 4857 -13604 4869 -13570
rect 5245 -13604 5257 -13570
rect 4857 -13616 5257 -13604
rect 5493 -13570 5893 -13558
rect 5493 -13604 5505 -13570
rect 5881 -13604 5893 -13570
rect 5493 -13616 5893 -13604
rect 4857 -13828 5257 -13816
rect 4857 -13862 4869 -13828
rect 5245 -13862 5257 -13828
rect 4857 -13874 5257 -13862
rect 5493 -13828 5893 -13816
rect 5493 -13862 5505 -13828
rect 5881 -13862 5893 -13828
rect 5493 -13874 5893 -13862
rect 4857 -14096 5257 -14084
rect 4857 -14130 4869 -14096
rect 5245 -14130 5257 -14096
rect 4857 -14142 5257 -14130
rect 5493 -14096 5893 -14084
rect 5493 -14130 5505 -14096
rect 5881 -14130 5893 -14096
rect 5493 -14142 5893 -14130
rect 4857 -14954 5257 -14942
rect 4857 -14988 4869 -14954
rect 5245 -14988 5257 -14954
rect 4857 -15000 5257 -14988
rect 5493 -14954 5893 -14942
rect 5493 -14988 5505 -14954
rect 5881 -14988 5893 -14954
rect 5493 -15000 5893 -14988
rect 6457 -13570 6857 -13558
rect 6457 -13604 6469 -13570
rect 6845 -13604 6857 -13570
rect 6457 -13616 6857 -13604
rect 7093 -13570 7493 -13558
rect 7093 -13604 7105 -13570
rect 7481 -13604 7493 -13570
rect 7093 -13616 7493 -13604
rect 6457 -13828 6857 -13816
rect 6457 -13862 6469 -13828
rect 6845 -13862 6857 -13828
rect 6457 -13874 6857 -13862
rect 7093 -13828 7493 -13816
rect 7093 -13862 7105 -13828
rect 7481 -13862 7493 -13828
rect 7093 -13874 7493 -13862
rect 6457 -14096 6857 -14084
rect 6457 -14130 6469 -14096
rect 6845 -14130 6857 -14096
rect 6457 -14142 6857 -14130
rect 7093 -14096 7493 -14084
rect 7093 -14130 7105 -14096
rect 7481 -14130 7493 -14096
rect 7093 -14142 7493 -14130
rect 6457 -14954 6857 -14942
rect 6457 -14988 6469 -14954
rect 6845 -14988 6857 -14954
rect 6457 -15000 6857 -14988
rect 7093 -14954 7493 -14942
rect 7093 -14988 7105 -14954
rect 7481 -14988 7493 -14954
rect 7093 -15000 7493 -14988
rect 8057 -13570 8457 -13558
rect 8057 -13604 8069 -13570
rect 8445 -13604 8457 -13570
rect 8057 -13616 8457 -13604
rect 8693 -13570 9093 -13558
rect 8693 -13604 8705 -13570
rect 9081 -13604 9093 -13570
rect 8693 -13616 9093 -13604
rect 8057 -13828 8457 -13816
rect 8057 -13862 8069 -13828
rect 8445 -13862 8457 -13828
rect 8057 -13874 8457 -13862
rect 8693 -13828 9093 -13816
rect 8693 -13862 8705 -13828
rect 9081 -13862 9093 -13828
rect 8693 -13874 9093 -13862
rect 8057 -14096 8457 -14084
rect 8057 -14130 8069 -14096
rect 8445 -14130 8457 -14096
rect 8057 -14142 8457 -14130
rect 8693 -14096 9093 -14084
rect 8693 -14130 8705 -14096
rect 9081 -14130 9093 -14096
rect 8693 -14142 9093 -14130
rect 8057 -14954 8457 -14942
rect 8057 -14988 8069 -14954
rect 8445 -14988 8457 -14954
rect 8057 -15000 8457 -14988
rect 8693 -14954 9093 -14942
rect 8693 -14988 8705 -14954
rect 9081 -14988 9093 -14954
rect 8693 -15000 9093 -14988
rect 9657 -13570 10057 -13558
rect 9657 -13604 9669 -13570
rect 10045 -13604 10057 -13570
rect 9657 -13616 10057 -13604
rect 10293 -13570 10693 -13558
rect 10293 -13604 10305 -13570
rect 10681 -13604 10693 -13570
rect 10293 -13616 10693 -13604
rect 9657 -13828 10057 -13816
rect 9657 -13862 9669 -13828
rect 10045 -13862 10057 -13828
rect 9657 -13874 10057 -13862
rect 10293 -13828 10693 -13816
rect 10293 -13862 10305 -13828
rect 10681 -13862 10693 -13828
rect 10293 -13874 10693 -13862
rect 9657 -14096 10057 -14084
rect 9657 -14130 9669 -14096
rect 10045 -14130 10057 -14096
rect 9657 -14142 10057 -14130
rect 10293 -14096 10693 -14084
rect 10293 -14130 10305 -14096
rect 10681 -14130 10693 -14096
rect 10293 -14142 10693 -14130
rect 9657 -14954 10057 -14942
rect 9657 -14988 9669 -14954
rect 10045 -14988 10057 -14954
rect 9657 -15000 10057 -14988
rect 10293 -14954 10693 -14942
rect 10293 -14988 10305 -14954
rect 10681 -14988 10693 -14954
rect 10293 -15000 10693 -14988
rect 11257 -13570 11657 -13558
rect 11257 -13604 11269 -13570
rect 11645 -13604 11657 -13570
rect 11257 -13616 11657 -13604
rect 11893 -13570 12293 -13558
rect 11893 -13604 11905 -13570
rect 12281 -13604 12293 -13570
rect 11893 -13616 12293 -13604
rect 11257 -13828 11657 -13816
rect 11257 -13862 11269 -13828
rect 11645 -13862 11657 -13828
rect 11257 -13874 11657 -13862
rect 11893 -13828 12293 -13816
rect 11893 -13862 11905 -13828
rect 12281 -13862 12293 -13828
rect 11893 -13874 12293 -13862
rect 11257 -14096 11657 -14084
rect 11257 -14130 11269 -14096
rect 11645 -14130 11657 -14096
rect 11257 -14142 11657 -14130
rect 11893 -14096 12293 -14084
rect 11893 -14130 11905 -14096
rect 12281 -14130 12293 -14096
rect 11893 -14142 12293 -14130
rect 11257 -14954 11657 -14942
rect 11257 -14988 11269 -14954
rect 11645 -14988 11657 -14954
rect 11257 -15000 11657 -14988
rect 11893 -14954 12293 -14942
rect 11893 -14988 11905 -14954
rect 12281 -14988 12293 -14954
rect 11893 -15000 12293 -14988
rect 12857 -13570 13257 -13558
rect 12857 -13604 12869 -13570
rect 13245 -13604 13257 -13570
rect 12857 -13616 13257 -13604
rect 13493 -13570 13893 -13558
rect 13493 -13604 13505 -13570
rect 13881 -13604 13893 -13570
rect 13493 -13616 13893 -13604
rect 12857 -13828 13257 -13816
rect 12857 -13862 12869 -13828
rect 13245 -13862 13257 -13828
rect 12857 -13874 13257 -13862
rect 13493 -13828 13893 -13816
rect 13493 -13862 13505 -13828
rect 13881 -13862 13893 -13828
rect 13493 -13874 13893 -13862
rect 12857 -14096 13257 -14084
rect 12857 -14130 12869 -14096
rect 13245 -14130 13257 -14096
rect 12857 -14142 13257 -14130
rect 13493 -14096 13893 -14084
rect 13493 -14130 13505 -14096
rect 13881 -14130 13893 -14096
rect 13493 -14142 13893 -14130
rect 12857 -14954 13257 -14942
rect 12857 -14988 12869 -14954
rect 13245 -14988 13257 -14954
rect 12857 -15000 13257 -14988
rect 13493 -14954 13893 -14942
rect 13493 -14988 13505 -14954
rect 13881 -14988 13893 -14954
rect 13493 -15000 13893 -14988
rect 14457 -13570 14857 -13558
rect 14457 -13604 14469 -13570
rect 14845 -13604 14857 -13570
rect 14457 -13616 14857 -13604
rect 15093 -13570 15493 -13558
rect 15093 -13604 15105 -13570
rect 15481 -13604 15493 -13570
rect 15093 -13616 15493 -13604
rect 14457 -13828 14857 -13816
rect 14457 -13862 14469 -13828
rect 14845 -13862 14857 -13828
rect 14457 -13874 14857 -13862
rect 15093 -13828 15493 -13816
rect 15093 -13862 15105 -13828
rect 15481 -13862 15493 -13828
rect 15093 -13874 15493 -13862
rect 14457 -14096 14857 -14084
rect 14457 -14130 14469 -14096
rect 14845 -14130 14857 -14096
rect 14457 -14142 14857 -14130
rect 15093 -14096 15493 -14084
rect 15093 -14130 15105 -14096
rect 15481 -14130 15493 -14096
rect 15093 -14142 15493 -14130
rect 14457 -14954 14857 -14942
rect 14457 -14988 14469 -14954
rect 14845 -14988 14857 -14954
rect 14457 -15000 14857 -14988
rect 15093 -14954 15493 -14942
rect 15093 -14988 15105 -14954
rect 15481 -14988 15493 -14954
rect 15093 -15000 15493 -14988
rect 16057 -13570 16457 -13558
rect 16057 -13604 16069 -13570
rect 16445 -13604 16457 -13570
rect 16057 -13616 16457 -13604
rect 16693 -13570 17093 -13558
rect 16693 -13604 16705 -13570
rect 17081 -13604 17093 -13570
rect 16693 -13616 17093 -13604
rect 16057 -13828 16457 -13816
rect 16057 -13862 16069 -13828
rect 16445 -13862 16457 -13828
rect 16057 -13874 16457 -13862
rect 16693 -13828 17093 -13816
rect 16693 -13862 16705 -13828
rect 17081 -13862 17093 -13828
rect 16693 -13874 17093 -13862
rect 16057 -14096 16457 -14084
rect 16057 -14130 16069 -14096
rect 16445 -14130 16457 -14096
rect 16057 -14142 16457 -14130
rect 16693 -14096 17093 -14084
rect 16693 -14130 16705 -14096
rect 17081 -14130 17093 -14096
rect 16693 -14142 17093 -14130
rect 16057 -14954 16457 -14942
rect 16057 -14988 16069 -14954
rect 16445 -14988 16457 -14954
rect 16057 -15000 16457 -14988
rect 16693 -14954 17093 -14942
rect 16693 -14988 16705 -14954
rect 17081 -14988 17093 -14954
rect 16693 -15000 17093 -14988
rect 17657 -13570 18057 -13558
rect 17657 -13604 17669 -13570
rect 18045 -13604 18057 -13570
rect 17657 -13616 18057 -13604
rect 18293 -13570 18693 -13558
rect 18293 -13604 18305 -13570
rect 18681 -13604 18693 -13570
rect 18293 -13616 18693 -13604
rect 17657 -13828 18057 -13816
rect 17657 -13862 17669 -13828
rect 18045 -13862 18057 -13828
rect 17657 -13874 18057 -13862
rect 18293 -13828 18693 -13816
rect 18293 -13862 18305 -13828
rect 18681 -13862 18693 -13828
rect 18293 -13874 18693 -13862
rect 17657 -14096 18057 -14084
rect 17657 -14130 17669 -14096
rect 18045 -14130 18057 -14096
rect 17657 -14142 18057 -14130
rect 18293 -14096 18693 -14084
rect 18293 -14130 18305 -14096
rect 18681 -14130 18693 -14096
rect 18293 -14142 18693 -14130
rect 17657 -14954 18057 -14942
rect 17657 -14988 17669 -14954
rect 18045 -14988 18057 -14954
rect 17657 -15000 18057 -14988
rect 18293 -14954 18693 -14942
rect 18293 -14988 18305 -14954
rect 18681 -14988 18693 -14954
rect 18293 -15000 18693 -14988
rect 19257 -13570 19657 -13558
rect 19257 -13604 19269 -13570
rect 19645 -13604 19657 -13570
rect 19257 -13616 19657 -13604
rect 19893 -13570 20293 -13558
rect 19893 -13604 19905 -13570
rect 20281 -13604 20293 -13570
rect 19893 -13616 20293 -13604
rect 19257 -13828 19657 -13816
rect 19257 -13862 19269 -13828
rect 19645 -13862 19657 -13828
rect 19257 -13874 19657 -13862
rect 19893 -13828 20293 -13816
rect 19893 -13862 19905 -13828
rect 20281 -13862 20293 -13828
rect 19893 -13874 20293 -13862
rect 19257 -14096 19657 -14084
rect 19257 -14130 19269 -14096
rect 19645 -14130 19657 -14096
rect 19257 -14142 19657 -14130
rect 19893 -14096 20293 -14084
rect 19893 -14130 19905 -14096
rect 20281 -14130 20293 -14096
rect 19893 -14142 20293 -14130
rect 19257 -14954 19657 -14942
rect 19257 -14988 19269 -14954
rect 19645 -14988 19657 -14954
rect 19257 -15000 19657 -14988
rect 19893 -14954 20293 -14942
rect 19893 -14988 19905 -14954
rect 20281 -14988 20293 -14954
rect 19893 -15000 20293 -14988
rect 20857 -13570 21257 -13558
rect 20857 -13604 20869 -13570
rect 21245 -13604 21257 -13570
rect 20857 -13616 21257 -13604
rect 21493 -13570 21893 -13558
rect 21493 -13604 21505 -13570
rect 21881 -13604 21893 -13570
rect 21493 -13616 21893 -13604
rect 20857 -13828 21257 -13816
rect 20857 -13862 20869 -13828
rect 21245 -13862 21257 -13828
rect 20857 -13874 21257 -13862
rect 21493 -13828 21893 -13816
rect 21493 -13862 21505 -13828
rect 21881 -13862 21893 -13828
rect 21493 -13874 21893 -13862
rect 20857 -14096 21257 -14084
rect 20857 -14130 20869 -14096
rect 21245 -14130 21257 -14096
rect 20857 -14142 21257 -14130
rect 21493 -14096 21893 -14084
rect 21493 -14130 21505 -14096
rect 21881 -14130 21893 -14096
rect 21493 -14142 21893 -14130
rect 20857 -14954 21257 -14942
rect 20857 -14988 20869 -14954
rect 21245 -14988 21257 -14954
rect 20857 -15000 21257 -14988
rect 21493 -14954 21893 -14942
rect 21493 -14988 21505 -14954
rect 21881 -14988 21893 -14954
rect 21493 -15000 21893 -14988
rect 22457 -13570 22857 -13558
rect 22457 -13604 22469 -13570
rect 22845 -13604 22857 -13570
rect 22457 -13616 22857 -13604
rect 23093 -13570 23493 -13558
rect 23093 -13604 23105 -13570
rect 23481 -13604 23493 -13570
rect 23093 -13616 23493 -13604
rect 22457 -13828 22857 -13816
rect 22457 -13862 22469 -13828
rect 22845 -13862 22857 -13828
rect 22457 -13874 22857 -13862
rect 23093 -13828 23493 -13816
rect 23093 -13862 23105 -13828
rect 23481 -13862 23493 -13828
rect 23093 -13874 23493 -13862
rect 22457 -14096 22857 -14084
rect 22457 -14130 22469 -14096
rect 22845 -14130 22857 -14096
rect 22457 -14142 22857 -14130
rect 23093 -14096 23493 -14084
rect 23093 -14130 23105 -14096
rect 23481 -14130 23493 -14096
rect 23093 -14142 23493 -14130
rect 22457 -14954 22857 -14942
rect 22457 -14988 22469 -14954
rect 22845 -14988 22857 -14954
rect 22457 -15000 22857 -14988
rect 23093 -14954 23493 -14942
rect 23093 -14988 23105 -14954
rect 23481 -14988 23493 -14954
rect 23093 -15000 23493 -14988
rect 24057 -13570 24457 -13558
rect 24057 -13604 24069 -13570
rect 24445 -13604 24457 -13570
rect 24057 -13616 24457 -13604
rect 24693 -13570 25093 -13558
rect 24693 -13604 24705 -13570
rect 25081 -13604 25093 -13570
rect 24693 -13616 25093 -13604
rect 24057 -13828 24457 -13816
rect 24057 -13862 24069 -13828
rect 24445 -13862 24457 -13828
rect 24057 -13874 24457 -13862
rect 24693 -13828 25093 -13816
rect 24693 -13862 24705 -13828
rect 25081 -13862 25093 -13828
rect 24693 -13874 25093 -13862
rect 24057 -14096 24457 -14084
rect 24057 -14130 24069 -14096
rect 24445 -14130 24457 -14096
rect 24057 -14142 24457 -14130
rect 24693 -14096 25093 -14084
rect 24693 -14130 24705 -14096
rect 25081 -14130 25093 -14096
rect 24693 -14142 25093 -14130
rect 24057 -14954 24457 -14942
rect 24057 -14988 24069 -14954
rect 24445 -14988 24457 -14954
rect 24057 -15000 24457 -14988
rect 24693 -14954 25093 -14942
rect 24693 -14988 24705 -14954
rect 25081 -14988 25093 -14954
rect 24693 -15000 25093 -14988
rect 25657 -13570 26057 -13558
rect 25657 -13604 25669 -13570
rect 26045 -13604 26057 -13570
rect 25657 -13616 26057 -13604
rect 26293 -13570 26693 -13558
rect 26293 -13604 26305 -13570
rect 26681 -13604 26693 -13570
rect 26293 -13616 26693 -13604
rect 25657 -13828 26057 -13816
rect 25657 -13862 25669 -13828
rect 26045 -13862 26057 -13828
rect 25657 -13874 26057 -13862
rect 26293 -13828 26693 -13816
rect 26293 -13862 26305 -13828
rect 26681 -13862 26693 -13828
rect 26293 -13874 26693 -13862
rect 25657 -14096 26057 -14084
rect 25657 -14130 25669 -14096
rect 26045 -14130 26057 -14096
rect 25657 -14142 26057 -14130
rect 26293 -14096 26693 -14084
rect 26293 -14130 26305 -14096
rect 26681 -14130 26693 -14096
rect 26293 -14142 26693 -14130
rect 25657 -14954 26057 -14942
rect 25657 -14988 25669 -14954
rect 26045 -14988 26057 -14954
rect 25657 -15000 26057 -14988
rect 26293 -14954 26693 -14942
rect 26293 -14988 26305 -14954
rect 26681 -14988 26693 -14954
rect 26293 -15000 26693 -14988
rect 27257 -13570 27657 -13558
rect 27257 -13604 27269 -13570
rect 27645 -13604 27657 -13570
rect 27257 -13616 27657 -13604
rect 27893 -13570 28293 -13558
rect 27893 -13604 27905 -13570
rect 28281 -13604 28293 -13570
rect 27893 -13616 28293 -13604
rect 27257 -13828 27657 -13816
rect 27257 -13862 27269 -13828
rect 27645 -13862 27657 -13828
rect 27257 -13874 27657 -13862
rect 27893 -13828 28293 -13816
rect 27893 -13862 27905 -13828
rect 28281 -13862 28293 -13828
rect 27893 -13874 28293 -13862
rect 27257 -14096 27657 -14084
rect 27257 -14130 27269 -14096
rect 27645 -14130 27657 -14096
rect 27257 -14142 27657 -14130
rect 27893 -14096 28293 -14084
rect 27893 -14130 27905 -14096
rect 28281 -14130 28293 -14096
rect 27893 -14142 28293 -14130
rect 27257 -14954 27657 -14942
rect 27257 -14988 27269 -14954
rect 27645 -14988 27657 -14954
rect 27257 -15000 27657 -14988
rect 27893 -14954 28293 -14942
rect 27893 -14988 27905 -14954
rect 28281 -14988 28293 -14954
rect 27893 -15000 28293 -14988
rect 28857 -13570 29257 -13558
rect 28857 -13604 28869 -13570
rect 29245 -13604 29257 -13570
rect 28857 -13616 29257 -13604
rect 29493 -13570 29893 -13558
rect 29493 -13604 29505 -13570
rect 29881 -13604 29893 -13570
rect 29493 -13616 29893 -13604
rect 28857 -13828 29257 -13816
rect 28857 -13862 28869 -13828
rect 29245 -13862 29257 -13828
rect 28857 -13874 29257 -13862
rect 29493 -13828 29893 -13816
rect 29493 -13862 29505 -13828
rect 29881 -13862 29893 -13828
rect 29493 -13874 29893 -13862
rect 28857 -14096 29257 -14084
rect 28857 -14130 28869 -14096
rect 29245 -14130 29257 -14096
rect 28857 -14142 29257 -14130
rect 29493 -14096 29893 -14084
rect 29493 -14130 29505 -14096
rect 29881 -14130 29893 -14096
rect 29493 -14142 29893 -14130
rect 28857 -14954 29257 -14942
rect 28857 -14988 28869 -14954
rect 29245 -14988 29257 -14954
rect 28857 -15000 29257 -14988
rect 29493 -14954 29893 -14942
rect 29493 -14988 29505 -14954
rect 29881 -14988 29893 -14954
rect 29493 -15000 29893 -14988
rect 30457 -13570 30857 -13558
rect 30457 -13604 30469 -13570
rect 30845 -13604 30857 -13570
rect 30457 -13616 30857 -13604
rect 31093 -13570 31493 -13558
rect 31093 -13604 31105 -13570
rect 31481 -13604 31493 -13570
rect 31093 -13616 31493 -13604
rect 30457 -13828 30857 -13816
rect 30457 -13862 30469 -13828
rect 30845 -13862 30857 -13828
rect 30457 -13874 30857 -13862
rect 31093 -13828 31493 -13816
rect 31093 -13862 31105 -13828
rect 31481 -13862 31493 -13828
rect 31093 -13874 31493 -13862
rect 30457 -14096 30857 -14084
rect 30457 -14130 30469 -14096
rect 30845 -14130 30857 -14096
rect 30457 -14142 30857 -14130
rect 31093 -14096 31493 -14084
rect 31093 -14130 31105 -14096
rect 31481 -14130 31493 -14096
rect 31093 -14142 31493 -14130
rect 30457 -14954 30857 -14942
rect 30457 -14988 30469 -14954
rect 30845 -14988 30857 -14954
rect 30457 -15000 30857 -14988
rect 31093 -14954 31493 -14942
rect 31093 -14988 31105 -14954
rect 31481 -14988 31493 -14954
rect 31093 -15000 31493 -14988
rect 32057 -13570 32457 -13558
rect 32057 -13604 32069 -13570
rect 32445 -13604 32457 -13570
rect 32057 -13616 32457 -13604
rect 32693 -13570 33093 -13558
rect 32693 -13604 32705 -13570
rect 33081 -13604 33093 -13570
rect 32693 -13616 33093 -13604
rect 32057 -13828 32457 -13816
rect 32057 -13862 32069 -13828
rect 32445 -13862 32457 -13828
rect 32057 -13874 32457 -13862
rect 32693 -13828 33093 -13816
rect 32693 -13862 32705 -13828
rect 33081 -13862 33093 -13828
rect 32693 -13874 33093 -13862
rect 32057 -14096 32457 -14084
rect 32057 -14130 32069 -14096
rect 32445 -14130 32457 -14096
rect 32057 -14142 32457 -14130
rect 32693 -14096 33093 -14084
rect 32693 -14130 32705 -14096
rect 33081 -14130 33093 -14096
rect 32693 -14142 33093 -14130
rect 32057 -14954 32457 -14942
rect 32057 -14988 32069 -14954
rect 32445 -14988 32457 -14954
rect 32057 -15000 32457 -14988
rect 32693 -14954 33093 -14942
rect 32693 -14988 32705 -14954
rect 33081 -14988 33093 -14954
rect 32693 -15000 33093 -14988
rect 33657 -13570 34057 -13558
rect 33657 -13604 33669 -13570
rect 34045 -13604 34057 -13570
rect 33657 -13616 34057 -13604
rect 34293 -13570 34693 -13558
rect 34293 -13604 34305 -13570
rect 34681 -13604 34693 -13570
rect 34293 -13616 34693 -13604
rect 33657 -13828 34057 -13816
rect 33657 -13862 33669 -13828
rect 34045 -13862 34057 -13828
rect 33657 -13874 34057 -13862
rect 34293 -13828 34693 -13816
rect 34293 -13862 34305 -13828
rect 34681 -13862 34693 -13828
rect 34293 -13874 34693 -13862
rect 33657 -14096 34057 -14084
rect 33657 -14130 33669 -14096
rect 34045 -14130 34057 -14096
rect 33657 -14142 34057 -14130
rect 34293 -14096 34693 -14084
rect 34293 -14130 34305 -14096
rect 34681 -14130 34693 -14096
rect 34293 -14142 34693 -14130
rect 33657 -14954 34057 -14942
rect 33657 -14988 33669 -14954
rect 34045 -14988 34057 -14954
rect 33657 -15000 34057 -14988
rect 34293 -14954 34693 -14942
rect 34293 -14988 34305 -14954
rect 34681 -14988 34693 -14954
rect 34293 -15000 34693 -14988
rect 35257 -13570 35657 -13558
rect 35257 -13604 35269 -13570
rect 35645 -13604 35657 -13570
rect 35257 -13616 35657 -13604
rect 35893 -13570 36293 -13558
rect 35893 -13604 35905 -13570
rect 36281 -13604 36293 -13570
rect 35893 -13616 36293 -13604
rect 35257 -13828 35657 -13816
rect 35257 -13862 35269 -13828
rect 35645 -13862 35657 -13828
rect 35257 -13874 35657 -13862
rect 35893 -13828 36293 -13816
rect 35893 -13862 35905 -13828
rect 36281 -13862 36293 -13828
rect 35893 -13874 36293 -13862
rect 35257 -14096 35657 -14084
rect 35257 -14130 35269 -14096
rect 35645 -14130 35657 -14096
rect 35257 -14142 35657 -14130
rect 35893 -14096 36293 -14084
rect 35893 -14130 35905 -14096
rect 36281 -14130 36293 -14096
rect 35893 -14142 36293 -14130
rect 35257 -14954 35657 -14942
rect 35257 -14988 35269 -14954
rect 35645 -14988 35657 -14954
rect 35257 -15000 35657 -14988
rect 35893 -14954 36293 -14942
rect 35893 -14988 35905 -14954
rect 36281 -14988 36293 -14954
rect 35893 -15000 36293 -14988
rect 36857 -13570 37257 -13558
rect 36857 -13604 36869 -13570
rect 37245 -13604 37257 -13570
rect 36857 -13616 37257 -13604
rect 37493 -13570 37893 -13558
rect 37493 -13604 37505 -13570
rect 37881 -13604 37893 -13570
rect 37493 -13616 37893 -13604
rect 36857 -13828 37257 -13816
rect 36857 -13862 36869 -13828
rect 37245 -13862 37257 -13828
rect 36857 -13874 37257 -13862
rect 37493 -13828 37893 -13816
rect 37493 -13862 37505 -13828
rect 37881 -13862 37893 -13828
rect 37493 -13874 37893 -13862
rect 36857 -14096 37257 -14084
rect 36857 -14130 36869 -14096
rect 37245 -14130 37257 -14096
rect 36857 -14142 37257 -14130
rect 37493 -14096 37893 -14084
rect 37493 -14130 37505 -14096
rect 37881 -14130 37893 -14096
rect 37493 -14142 37893 -14130
rect 36857 -14954 37257 -14942
rect 36857 -14988 36869 -14954
rect 37245 -14988 37257 -14954
rect 36857 -15000 37257 -14988
rect 37493 -14954 37893 -14942
rect 37493 -14988 37505 -14954
rect 37881 -14988 37893 -14954
rect 37493 -15000 37893 -14988
rect 57 -15370 457 -15358
rect 57 -15404 69 -15370
rect 445 -15404 457 -15370
rect 57 -15416 457 -15404
rect 693 -15370 1093 -15358
rect 693 -15404 705 -15370
rect 1081 -15404 1093 -15370
rect 693 -15416 1093 -15404
rect 57 -15628 457 -15616
rect 57 -15662 69 -15628
rect 445 -15662 457 -15628
rect 57 -15674 457 -15662
rect 693 -15628 1093 -15616
rect 693 -15662 705 -15628
rect 1081 -15662 1093 -15628
rect 693 -15674 1093 -15662
rect 57 -15896 457 -15884
rect 57 -15930 69 -15896
rect 445 -15930 457 -15896
rect 57 -15942 457 -15930
rect 693 -15896 1093 -15884
rect 693 -15930 705 -15896
rect 1081 -15930 1093 -15896
rect 693 -15942 1093 -15930
rect 57 -16754 457 -16742
rect 57 -16788 69 -16754
rect 445 -16788 457 -16754
rect 57 -16800 457 -16788
rect 693 -16754 1093 -16742
rect 693 -16788 705 -16754
rect 1081 -16788 1093 -16754
rect 693 -16800 1093 -16788
rect 1657 -15370 2057 -15358
rect 1657 -15404 1669 -15370
rect 2045 -15404 2057 -15370
rect 1657 -15416 2057 -15404
rect 2293 -15370 2693 -15358
rect 2293 -15404 2305 -15370
rect 2681 -15404 2693 -15370
rect 2293 -15416 2693 -15404
rect 1657 -15628 2057 -15616
rect 1657 -15662 1669 -15628
rect 2045 -15662 2057 -15628
rect 1657 -15674 2057 -15662
rect 2293 -15628 2693 -15616
rect 2293 -15662 2305 -15628
rect 2681 -15662 2693 -15628
rect 2293 -15674 2693 -15662
rect 1657 -15896 2057 -15884
rect 1657 -15930 1669 -15896
rect 2045 -15930 2057 -15896
rect 1657 -15942 2057 -15930
rect 2293 -15896 2693 -15884
rect 2293 -15930 2305 -15896
rect 2681 -15930 2693 -15896
rect 2293 -15942 2693 -15930
rect 1657 -16754 2057 -16742
rect 1657 -16788 1669 -16754
rect 2045 -16788 2057 -16754
rect 1657 -16800 2057 -16788
rect 2293 -16754 2693 -16742
rect 2293 -16788 2305 -16754
rect 2681 -16788 2693 -16754
rect 2293 -16800 2693 -16788
rect 3257 -15370 3657 -15358
rect 3257 -15404 3269 -15370
rect 3645 -15404 3657 -15370
rect 3257 -15416 3657 -15404
rect 3893 -15370 4293 -15358
rect 3893 -15404 3905 -15370
rect 4281 -15404 4293 -15370
rect 3893 -15416 4293 -15404
rect 3257 -15628 3657 -15616
rect 3257 -15662 3269 -15628
rect 3645 -15662 3657 -15628
rect 3257 -15674 3657 -15662
rect 3893 -15628 4293 -15616
rect 3893 -15662 3905 -15628
rect 4281 -15662 4293 -15628
rect 3893 -15674 4293 -15662
rect 3257 -15896 3657 -15884
rect 3257 -15930 3269 -15896
rect 3645 -15930 3657 -15896
rect 3257 -15942 3657 -15930
rect 3893 -15896 4293 -15884
rect 3893 -15930 3905 -15896
rect 4281 -15930 4293 -15896
rect 3893 -15942 4293 -15930
rect 3257 -16754 3657 -16742
rect 3257 -16788 3269 -16754
rect 3645 -16788 3657 -16754
rect 3257 -16800 3657 -16788
rect 3893 -16754 4293 -16742
rect 3893 -16788 3905 -16754
rect 4281 -16788 4293 -16754
rect 3893 -16800 4293 -16788
rect 4857 -15370 5257 -15358
rect 4857 -15404 4869 -15370
rect 5245 -15404 5257 -15370
rect 4857 -15416 5257 -15404
rect 5493 -15370 5893 -15358
rect 5493 -15404 5505 -15370
rect 5881 -15404 5893 -15370
rect 5493 -15416 5893 -15404
rect 4857 -15628 5257 -15616
rect 4857 -15662 4869 -15628
rect 5245 -15662 5257 -15628
rect 4857 -15674 5257 -15662
rect 5493 -15628 5893 -15616
rect 5493 -15662 5505 -15628
rect 5881 -15662 5893 -15628
rect 5493 -15674 5893 -15662
rect 4857 -15896 5257 -15884
rect 4857 -15930 4869 -15896
rect 5245 -15930 5257 -15896
rect 4857 -15942 5257 -15930
rect 5493 -15896 5893 -15884
rect 5493 -15930 5505 -15896
rect 5881 -15930 5893 -15896
rect 5493 -15942 5893 -15930
rect 4857 -16754 5257 -16742
rect 4857 -16788 4869 -16754
rect 5245 -16788 5257 -16754
rect 4857 -16800 5257 -16788
rect 5493 -16754 5893 -16742
rect 5493 -16788 5505 -16754
rect 5881 -16788 5893 -16754
rect 5493 -16800 5893 -16788
rect 6457 -15370 6857 -15358
rect 6457 -15404 6469 -15370
rect 6845 -15404 6857 -15370
rect 6457 -15416 6857 -15404
rect 7093 -15370 7493 -15358
rect 7093 -15404 7105 -15370
rect 7481 -15404 7493 -15370
rect 7093 -15416 7493 -15404
rect 6457 -15628 6857 -15616
rect 6457 -15662 6469 -15628
rect 6845 -15662 6857 -15628
rect 6457 -15674 6857 -15662
rect 7093 -15628 7493 -15616
rect 7093 -15662 7105 -15628
rect 7481 -15662 7493 -15628
rect 7093 -15674 7493 -15662
rect 6457 -15896 6857 -15884
rect 6457 -15930 6469 -15896
rect 6845 -15930 6857 -15896
rect 6457 -15942 6857 -15930
rect 7093 -15896 7493 -15884
rect 7093 -15930 7105 -15896
rect 7481 -15930 7493 -15896
rect 7093 -15942 7493 -15930
rect 6457 -16754 6857 -16742
rect 6457 -16788 6469 -16754
rect 6845 -16788 6857 -16754
rect 6457 -16800 6857 -16788
rect 7093 -16754 7493 -16742
rect 7093 -16788 7105 -16754
rect 7481 -16788 7493 -16754
rect 7093 -16800 7493 -16788
rect 8057 -15370 8457 -15358
rect 8057 -15404 8069 -15370
rect 8445 -15404 8457 -15370
rect 8057 -15416 8457 -15404
rect 8693 -15370 9093 -15358
rect 8693 -15404 8705 -15370
rect 9081 -15404 9093 -15370
rect 8693 -15416 9093 -15404
rect 8057 -15628 8457 -15616
rect 8057 -15662 8069 -15628
rect 8445 -15662 8457 -15628
rect 8057 -15674 8457 -15662
rect 8693 -15628 9093 -15616
rect 8693 -15662 8705 -15628
rect 9081 -15662 9093 -15628
rect 8693 -15674 9093 -15662
rect 8057 -15896 8457 -15884
rect 8057 -15930 8069 -15896
rect 8445 -15930 8457 -15896
rect 8057 -15942 8457 -15930
rect 8693 -15896 9093 -15884
rect 8693 -15930 8705 -15896
rect 9081 -15930 9093 -15896
rect 8693 -15942 9093 -15930
rect 8057 -16754 8457 -16742
rect 8057 -16788 8069 -16754
rect 8445 -16788 8457 -16754
rect 8057 -16800 8457 -16788
rect 8693 -16754 9093 -16742
rect 8693 -16788 8705 -16754
rect 9081 -16788 9093 -16754
rect 8693 -16800 9093 -16788
rect 9657 -15370 10057 -15358
rect 9657 -15404 9669 -15370
rect 10045 -15404 10057 -15370
rect 9657 -15416 10057 -15404
rect 10293 -15370 10693 -15358
rect 10293 -15404 10305 -15370
rect 10681 -15404 10693 -15370
rect 10293 -15416 10693 -15404
rect 9657 -15628 10057 -15616
rect 9657 -15662 9669 -15628
rect 10045 -15662 10057 -15628
rect 9657 -15674 10057 -15662
rect 10293 -15628 10693 -15616
rect 10293 -15662 10305 -15628
rect 10681 -15662 10693 -15628
rect 10293 -15674 10693 -15662
rect 9657 -15896 10057 -15884
rect 9657 -15930 9669 -15896
rect 10045 -15930 10057 -15896
rect 9657 -15942 10057 -15930
rect 10293 -15896 10693 -15884
rect 10293 -15930 10305 -15896
rect 10681 -15930 10693 -15896
rect 10293 -15942 10693 -15930
rect 9657 -16754 10057 -16742
rect 9657 -16788 9669 -16754
rect 10045 -16788 10057 -16754
rect 9657 -16800 10057 -16788
rect 10293 -16754 10693 -16742
rect 10293 -16788 10305 -16754
rect 10681 -16788 10693 -16754
rect 10293 -16800 10693 -16788
rect 11257 -15370 11657 -15358
rect 11257 -15404 11269 -15370
rect 11645 -15404 11657 -15370
rect 11257 -15416 11657 -15404
rect 11893 -15370 12293 -15358
rect 11893 -15404 11905 -15370
rect 12281 -15404 12293 -15370
rect 11893 -15416 12293 -15404
rect 11257 -15628 11657 -15616
rect 11257 -15662 11269 -15628
rect 11645 -15662 11657 -15628
rect 11257 -15674 11657 -15662
rect 11893 -15628 12293 -15616
rect 11893 -15662 11905 -15628
rect 12281 -15662 12293 -15628
rect 11893 -15674 12293 -15662
rect 11257 -15896 11657 -15884
rect 11257 -15930 11269 -15896
rect 11645 -15930 11657 -15896
rect 11257 -15942 11657 -15930
rect 11893 -15896 12293 -15884
rect 11893 -15930 11905 -15896
rect 12281 -15930 12293 -15896
rect 11893 -15942 12293 -15930
rect 11257 -16754 11657 -16742
rect 11257 -16788 11269 -16754
rect 11645 -16788 11657 -16754
rect 11257 -16800 11657 -16788
rect 11893 -16754 12293 -16742
rect 11893 -16788 11905 -16754
rect 12281 -16788 12293 -16754
rect 11893 -16800 12293 -16788
rect 12857 -15370 13257 -15358
rect 12857 -15404 12869 -15370
rect 13245 -15404 13257 -15370
rect 12857 -15416 13257 -15404
rect 13493 -15370 13893 -15358
rect 13493 -15404 13505 -15370
rect 13881 -15404 13893 -15370
rect 13493 -15416 13893 -15404
rect 12857 -15628 13257 -15616
rect 12857 -15662 12869 -15628
rect 13245 -15662 13257 -15628
rect 12857 -15674 13257 -15662
rect 13493 -15628 13893 -15616
rect 13493 -15662 13505 -15628
rect 13881 -15662 13893 -15628
rect 13493 -15674 13893 -15662
rect 12857 -15896 13257 -15884
rect 12857 -15930 12869 -15896
rect 13245 -15930 13257 -15896
rect 12857 -15942 13257 -15930
rect 13493 -15896 13893 -15884
rect 13493 -15930 13505 -15896
rect 13881 -15930 13893 -15896
rect 13493 -15942 13893 -15930
rect 12857 -16754 13257 -16742
rect 12857 -16788 12869 -16754
rect 13245 -16788 13257 -16754
rect 12857 -16800 13257 -16788
rect 13493 -16754 13893 -16742
rect 13493 -16788 13505 -16754
rect 13881 -16788 13893 -16754
rect 13493 -16800 13893 -16788
rect 14457 -15370 14857 -15358
rect 14457 -15404 14469 -15370
rect 14845 -15404 14857 -15370
rect 14457 -15416 14857 -15404
rect 15093 -15370 15493 -15358
rect 15093 -15404 15105 -15370
rect 15481 -15404 15493 -15370
rect 15093 -15416 15493 -15404
rect 14457 -15628 14857 -15616
rect 14457 -15662 14469 -15628
rect 14845 -15662 14857 -15628
rect 14457 -15674 14857 -15662
rect 15093 -15628 15493 -15616
rect 15093 -15662 15105 -15628
rect 15481 -15662 15493 -15628
rect 15093 -15674 15493 -15662
rect 14457 -15896 14857 -15884
rect 14457 -15930 14469 -15896
rect 14845 -15930 14857 -15896
rect 14457 -15942 14857 -15930
rect 15093 -15896 15493 -15884
rect 15093 -15930 15105 -15896
rect 15481 -15930 15493 -15896
rect 15093 -15942 15493 -15930
rect 14457 -16754 14857 -16742
rect 14457 -16788 14469 -16754
rect 14845 -16788 14857 -16754
rect 14457 -16800 14857 -16788
rect 15093 -16754 15493 -16742
rect 15093 -16788 15105 -16754
rect 15481 -16788 15493 -16754
rect 15093 -16800 15493 -16788
rect 16057 -15370 16457 -15358
rect 16057 -15404 16069 -15370
rect 16445 -15404 16457 -15370
rect 16057 -15416 16457 -15404
rect 16693 -15370 17093 -15358
rect 16693 -15404 16705 -15370
rect 17081 -15404 17093 -15370
rect 16693 -15416 17093 -15404
rect 16057 -15628 16457 -15616
rect 16057 -15662 16069 -15628
rect 16445 -15662 16457 -15628
rect 16057 -15674 16457 -15662
rect 16693 -15628 17093 -15616
rect 16693 -15662 16705 -15628
rect 17081 -15662 17093 -15628
rect 16693 -15674 17093 -15662
rect 16057 -15896 16457 -15884
rect 16057 -15930 16069 -15896
rect 16445 -15930 16457 -15896
rect 16057 -15942 16457 -15930
rect 16693 -15896 17093 -15884
rect 16693 -15930 16705 -15896
rect 17081 -15930 17093 -15896
rect 16693 -15942 17093 -15930
rect 16057 -16754 16457 -16742
rect 16057 -16788 16069 -16754
rect 16445 -16788 16457 -16754
rect 16057 -16800 16457 -16788
rect 16693 -16754 17093 -16742
rect 16693 -16788 16705 -16754
rect 17081 -16788 17093 -16754
rect 16693 -16800 17093 -16788
rect 17657 -15370 18057 -15358
rect 17657 -15404 17669 -15370
rect 18045 -15404 18057 -15370
rect 17657 -15416 18057 -15404
rect 18293 -15370 18693 -15358
rect 18293 -15404 18305 -15370
rect 18681 -15404 18693 -15370
rect 18293 -15416 18693 -15404
rect 17657 -15628 18057 -15616
rect 17657 -15662 17669 -15628
rect 18045 -15662 18057 -15628
rect 17657 -15674 18057 -15662
rect 18293 -15628 18693 -15616
rect 18293 -15662 18305 -15628
rect 18681 -15662 18693 -15628
rect 18293 -15674 18693 -15662
rect 17657 -15896 18057 -15884
rect 17657 -15930 17669 -15896
rect 18045 -15930 18057 -15896
rect 17657 -15942 18057 -15930
rect 18293 -15896 18693 -15884
rect 18293 -15930 18305 -15896
rect 18681 -15930 18693 -15896
rect 18293 -15942 18693 -15930
rect 17657 -16754 18057 -16742
rect 17657 -16788 17669 -16754
rect 18045 -16788 18057 -16754
rect 17657 -16800 18057 -16788
rect 18293 -16754 18693 -16742
rect 18293 -16788 18305 -16754
rect 18681 -16788 18693 -16754
rect 18293 -16800 18693 -16788
rect 19257 -15370 19657 -15358
rect 19257 -15404 19269 -15370
rect 19645 -15404 19657 -15370
rect 19257 -15416 19657 -15404
rect 19893 -15370 20293 -15358
rect 19893 -15404 19905 -15370
rect 20281 -15404 20293 -15370
rect 19893 -15416 20293 -15404
rect 19257 -15628 19657 -15616
rect 19257 -15662 19269 -15628
rect 19645 -15662 19657 -15628
rect 19257 -15674 19657 -15662
rect 19893 -15628 20293 -15616
rect 19893 -15662 19905 -15628
rect 20281 -15662 20293 -15628
rect 19893 -15674 20293 -15662
rect 19257 -15896 19657 -15884
rect 19257 -15930 19269 -15896
rect 19645 -15930 19657 -15896
rect 19257 -15942 19657 -15930
rect 19893 -15896 20293 -15884
rect 19893 -15930 19905 -15896
rect 20281 -15930 20293 -15896
rect 19893 -15942 20293 -15930
rect 19257 -16754 19657 -16742
rect 19257 -16788 19269 -16754
rect 19645 -16788 19657 -16754
rect 19257 -16800 19657 -16788
rect 19893 -16754 20293 -16742
rect 19893 -16788 19905 -16754
rect 20281 -16788 20293 -16754
rect 19893 -16800 20293 -16788
rect 20857 -15370 21257 -15358
rect 20857 -15404 20869 -15370
rect 21245 -15404 21257 -15370
rect 20857 -15416 21257 -15404
rect 21493 -15370 21893 -15358
rect 21493 -15404 21505 -15370
rect 21881 -15404 21893 -15370
rect 21493 -15416 21893 -15404
rect 20857 -15628 21257 -15616
rect 20857 -15662 20869 -15628
rect 21245 -15662 21257 -15628
rect 20857 -15674 21257 -15662
rect 21493 -15628 21893 -15616
rect 21493 -15662 21505 -15628
rect 21881 -15662 21893 -15628
rect 21493 -15674 21893 -15662
rect 20857 -15896 21257 -15884
rect 20857 -15930 20869 -15896
rect 21245 -15930 21257 -15896
rect 20857 -15942 21257 -15930
rect 21493 -15896 21893 -15884
rect 21493 -15930 21505 -15896
rect 21881 -15930 21893 -15896
rect 21493 -15942 21893 -15930
rect 20857 -16754 21257 -16742
rect 20857 -16788 20869 -16754
rect 21245 -16788 21257 -16754
rect 20857 -16800 21257 -16788
rect 21493 -16754 21893 -16742
rect 21493 -16788 21505 -16754
rect 21881 -16788 21893 -16754
rect 21493 -16800 21893 -16788
rect 22457 -15370 22857 -15358
rect 22457 -15404 22469 -15370
rect 22845 -15404 22857 -15370
rect 22457 -15416 22857 -15404
rect 23093 -15370 23493 -15358
rect 23093 -15404 23105 -15370
rect 23481 -15404 23493 -15370
rect 23093 -15416 23493 -15404
rect 22457 -15628 22857 -15616
rect 22457 -15662 22469 -15628
rect 22845 -15662 22857 -15628
rect 22457 -15674 22857 -15662
rect 23093 -15628 23493 -15616
rect 23093 -15662 23105 -15628
rect 23481 -15662 23493 -15628
rect 23093 -15674 23493 -15662
rect 22457 -15896 22857 -15884
rect 22457 -15930 22469 -15896
rect 22845 -15930 22857 -15896
rect 22457 -15942 22857 -15930
rect 23093 -15896 23493 -15884
rect 23093 -15930 23105 -15896
rect 23481 -15930 23493 -15896
rect 23093 -15942 23493 -15930
rect 22457 -16754 22857 -16742
rect 22457 -16788 22469 -16754
rect 22845 -16788 22857 -16754
rect 22457 -16800 22857 -16788
rect 23093 -16754 23493 -16742
rect 23093 -16788 23105 -16754
rect 23481 -16788 23493 -16754
rect 23093 -16800 23493 -16788
rect 24057 -15370 24457 -15358
rect 24057 -15404 24069 -15370
rect 24445 -15404 24457 -15370
rect 24057 -15416 24457 -15404
rect 24693 -15370 25093 -15358
rect 24693 -15404 24705 -15370
rect 25081 -15404 25093 -15370
rect 24693 -15416 25093 -15404
rect 24057 -15628 24457 -15616
rect 24057 -15662 24069 -15628
rect 24445 -15662 24457 -15628
rect 24057 -15674 24457 -15662
rect 24693 -15628 25093 -15616
rect 24693 -15662 24705 -15628
rect 25081 -15662 25093 -15628
rect 24693 -15674 25093 -15662
rect 24057 -15896 24457 -15884
rect 24057 -15930 24069 -15896
rect 24445 -15930 24457 -15896
rect 24057 -15942 24457 -15930
rect 24693 -15896 25093 -15884
rect 24693 -15930 24705 -15896
rect 25081 -15930 25093 -15896
rect 24693 -15942 25093 -15930
rect 24057 -16754 24457 -16742
rect 24057 -16788 24069 -16754
rect 24445 -16788 24457 -16754
rect 24057 -16800 24457 -16788
rect 24693 -16754 25093 -16742
rect 24693 -16788 24705 -16754
rect 25081 -16788 25093 -16754
rect 24693 -16800 25093 -16788
rect 25657 -15370 26057 -15358
rect 25657 -15404 25669 -15370
rect 26045 -15404 26057 -15370
rect 25657 -15416 26057 -15404
rect 26293 -15370 26693 -15358
rect 26293 -15404 26305 -15370
rect 26681 -15404 26693 -15370
rect 26293 -15416 26693 -15404
rect 25657 -15628 26057 -15616
rect 25657 -15662 25669 -15628
rect 26045 -15662 26057 -15628
rect 25657 -15674 26057 -15662
rect 26293 -15628 26693 -15616
rect 26293 -15662 26305 -15628
rect 26681 -15662 26693 -15628
rect 26293 -15674 26693 -15662
rect 25657 -15896 26057 -15884
rect 25657 -15930 25669 -15896
rect 26045 -15930 26057 -15896
rect 25657 -15942 26057 -15930
rect 26293 -15896 26693 -15884
rect 26293 -15930 26305 -15896
rect 26681 -15930 26693 -15896
rect 26293 -15942 26693 -15930
rect 25657 -16754 26057 -16742
rect 25657 -16788 25669 -16754
rect 26045 -16788 26057 -16754
rect 25657 -16800 26057 -16788
rect 26293 -16754 26693 -16742
rect 26293 -16788 26305 -16754
rect 26681 -16788 26693 -16754
rect 26293 -16800 26693 -16788
rect 27257 -15370 27657 -15358
rect 27257 -15404 27269 -15370
rect 27645 -15404 27657 -15370
rect 27257 -15416 27657 -15404
rect 27893 -15370 28293 -15358
rect 27893 -15404 27905 -15370
rect 28281 -15404 28293 -15370
rect 27893 -15416 28293 -15404
rect 27257 -15628 27657 -15616
rect 27257 -15662 27269 -15628
rect 27645 -15662 27657 -15628
rect 27257 -15674 27657 -15662
rect 27893 -15628 28293 -15616
rect 27893 -15662 27905 -15628
rect 28281 -15662 28293 -15628
rect 27893 -15674 28293 -15662
rect 27257 -15896 27657 -15884
rect 27257 -15930 27269 -15896
rect 27645 -15930 27657 -15896
rect 27257 -15942 27657 -15930
rect 27893 -15896 28293 -15884
rect 27893 -15930 27905 -15896
rect 28281 -15930 28293 -15896
rect 27893 -15942 28293 -15930
rect 27257 -16754 27657 -16742
rect 27257 -16788 27269 -16754
rect 27645 -16788 27657 -16754
rect 27257 -16800 27657 -16788
rect 27893 -16754 28293 -16742
rect 27893 -16788 27905 -16754
rect 28281 -16788 28293 -16754
rect 27893 -16800 28293 -16788
rect 28857 -15370 29257 -15358
rect 28857 -15404 28869 -15370
rect 29245 -15404 29257 -15370
rect 28857 -15416 29257 -15404
rect 29493 -15370 29893 -15358
rect 29493 -15404 29505 -15370
rect 29881 -15404 29893 -15370
rect 29493 -15416 29893 -15404
rect 28857 -15628 29257 -15616
rect 28857 -15662 28869 -15628
rect 29245 -15662 29257 -15628
rect 28857 -15674 29257 -15662
rect 29493 -15628 29893 -15616
rect 29493 -15662 29505 -15628
rect 29881 -15662 29893 -15628
rect 29493 -15674 29893 -15662
rect 28857 -15896 29257 -15884
rect 28857 -15930 28869 -15896
rect 29245 -15930 29257 -15896
rect 28857 -15942 29257 -15930
rect 29493 -15896 29893 -15884
rect 29493 -15930 29505 -15896
rect 29881 -15930 29893 -15896
rect 29493 -15942 29893 -15930
rect 28857 -16754 29257 -16742
rect 28857 -16788 28869 -16754
rect 29245 -16788 29257 -16754
rect 28857 -16800 29257 -16788
rect 29493 -16754 29893 -16742
rect 29493 -16788 29505 -16754
rect 29881 -16788 29893 -16754
rect 29493 -16800 29893 -16788
rect 30457 -15370 30857 -15358
rect 30457 -15404 30469 -15370
rect 30845 -15404 30857 -15370
rect 30457 -15416 30857 -15404
rect 31093 -15370 31493 -15358
rect 31093 -15404 31105 -15370
rect 31481 -15404 31493 -15370
rect 31093 -15416 31493 -15404
rect 30457 -15628 30857 -15616
rect 30457 -15662 30469 -15628
rect 30845 -15662 30857 -15628
rect 30457 -15674 30857 -15662
rect 31093 -15628 31493 -15616
rect 31093 -15662 31105 -15628
rect 31481 -15662 31493 -15628
rect 31093 -15674 31493 -15662
rect 30457 -15896 30857 -15884
rect 30457 -15930 30469 -15896
rect 30845 -15930 30857 -15896
rect 30457 -15942 30857 -15930
rect 31093 -15896 31493 -15884
rect 31093 -15930 31105 -15896
rect 31481 -15930 31493 -15896
rect 31093 -15942 31493 -15930
rect 30457 -16754 30857 -16742
rect 30457 -16788 30469 -16754
rect 30845 -16788 30857 -16754
rect 30457 -16800 30857 -16788
rect 31093 -16754 31493 -16742
rect 31093 -16788 31105 -16754
rect 31481 -16788 31493 -16754
rect 31093 -16800 31493 -16788
rect 32057 -15370 32457 -15358
rect 32057 -15404 32069 -15370
rect 32445 -15404 32457 -15370
rect 32057 -15416 32457 -15404
rect 32693 -15370 33093 -15358
rect 32693 -15404 32705 -15370
rect 33081 -15404 33093 -15370
rect 32693 -15416 33093 -15404
rect 32057 -15628 32457 -15616
rect 32057 -15662 32069 -15628
rect 32445 -15662 32457 -15628
rect 32057 -15674 32457 -15662
rect 32693 -15628 33093 -15616
rect 32693 -15662 32705 -15628
rect 33081 -15662 33093 -15628
rect 32693 -15674 33093 -15662
rect 32057 -15896 32457 -15884
rect 32057 -15930 32069 -15896
rect 32445 -15930 32457 -15896
rect 32057 -15942 32457 -15930
rect 32693 -15896 33093 -15884
rect 32693 -15930 32705 -15896
rect 33081 -15930 33093 -15896
rect 32693 -15942 33093 -15930
rect 32057 -16754 32457 -16742
rect 32057 -16788 32069 -16754
rect 32445 -16788 32457 -16754
rect 32057 -16800 32457 -16788
rect 32693 -16754 33093 -16742
rect 32693 -16788 32705 -16754
rect 33081 -16788 33093 -16754
rect 32693 -16800 33093 -16788
rect 33657 -15370 34057 -15358
rect 33657 -15404 33669 -15370
rect 34045 -15404 34057 -15370
rect 33657 -15416 34057 -15404
rect 34293 -15370 34693 -15358
rect 34293 -15404 34305 -15370
rect 34681 -15404 34693 -15370
rect 34293 -15416 34693 -15404
rect 33657 -15628 34057 -15616
rect 33657 -15662 33669 -15628
rect 34045 -15662 34057 -15628
rect 33657 -15674 34057 -15662
rect 34293 -15628 34693 -15616
rect 34293 -15662 34305 -15628
rect 34681 -15662 34693 -15628
rect 34293 -15674 34693 -15662
rect 33657 -15896 34057 -15884
rect 33657 -15930 33669 -15896
rect 34045 -15930 34057 -15896
rect 33657 -15942 34057 -15930
rect 34293 -15896 34693 -15884
rect 34293 -15930 34305 -15896
rect 34681 -15930 34693 -15896
rect 34293 -15942 34693 -15930
rect 33657 -16754 34057 -16742
rect 33657 -16788 33669 -16754
rect 34045 -16788 34057 -16754
rect 33657 -16800 34057 -16788
rect 34293 -16754 34693 -16742
rect 34293 -16788 34305 -16754
rect 34681 -16788 34693 -16754
rect 34293 -16800 34693 -16788
rect 35257 -15370 35657 -15358
rect 35257 -15404 35269 -15370
rect 35645 -15404 35657 -15370
rect 35257 -15416 35657 -15404
rect 35893 -15370 36293 -15358
rect 35893 -15404 35905 -15370
rect 36281 -15404 36293 -15370
rect 35893 -15416 36293 -15404
rect 35257 -15628 35657 -15616
rect 35257 -15662 35269 -15628
rect 35645 -15662 35657 -15628
rect 35257 -15674 35657 -15662
rect 35893 -15628 36293 -15616
rect 35893 -15662 35905 -15628
rect 36281 -15662 36293 -15628
rect 35893 -15674 36293 -15662
rect 35257 -15896 35657 -15884
rect 35257 -15930 35269 -15896
rect 35645 -15930 35657 -15896
rect 35257 -15942 35657 -15930
rect 35893 -15896 36293 -15884
rect 35893 -15930 35905 -15896
rect 36281 -15930 36293 -15896
rect 35893 -15942 36293 -15930
rect 35257 -16754 35657 -16742
rect 35257 -16788 35269 -16754
rect 35645 -16788 35657 -16754
rect 35257 -16800 35657 -16788
rect 35893 -16754 36293 -16742
rect 35893 -16788 35905 -16754
rect 36281 -16788 36293 -16754
rect 35893 -16800 36293 -16788
rect 36857 -15370 37257 -15358
rect 36857 -15404 36869 -15370
rect 37245 -15404 37257 -15370
rect 36857 -15416 37257 -15404
rect 37493 -15370 37893 -15358
rect 37493 -15404 37505 -15370
rect 37881 -15404 37893 -15370
rect 37493 -15416 37893 -15404
rect 36857 -15628 37257 -15616
rect 36857 -15662 36869 -15628
rect 37245 -15662 37257 -15628
rect 36857 -15674 37257 -15662
rect 37493 -15628 37893 -15616
rect 37493 -15662 37505 -15628
rect 37881 -15662 37893 -15628
rect 37493 -15674 37893 -15662
rect 36857 -15896 37257 -15884
rect 36857 -15930 36869 -15896
rect 37245 -15930 37257 -15896
rect 36857 -15942 37257 -15930
rect 37493 -15896 37893 -15884
rect 37493 -15930 37505 -15896
rect 37881 -15930 37893 -15896
rect 37493 -15942 37893 -15930
rect 36857 -16754 37257 -16742
rect 36857 -16788 36869 -16754
rect 37245 -16788 37257 -16754
rect 36857 -16800 37257 -16788
rect 37493 -16754 37893 -16742
rect 37493 -16788 37505 -16754
rect 37881 -16788 37893 -16754
rect 37493 -16800 37893 -16788
rect 57 -17170 457 -17158
rect 57 -17204 69 -17170
rect 445 -17204 457 -17170
rect 57 -17216 457 -17204
rect 693 -17170 1093 -17158
rect 693 -17204 705 -17170
rect 1081 -17204 1093 -17170
rect 693 -17216 1093 -17204
rect 57 -17428 457 -17416
rect 57 -17462 69 -17428
rect 445 -17462 457 -17428
rect 57 -17474 457 -17462
rect 693 -17428 1093 -17416
rect 693 -17462 705 -17428
rect 1081 -17462 1093 -17428
rect 693 -17474 1093 -17462
rect 57 -17696 457 -17684
rect 57 -17730 69 -17696
rect 445 -17730 457 -17696
rect 57 -17742 457 -17730
rect 693 -17696 1093 -17684
rect 693 -17730 705 -17696
rect 1081 -17730 1093 -17696
rect 693 -17742 1093 -17730
rect 57 -18554 457 -18542
rect 57 -18588 69 -18554
rect 445 -18588 457 -18554
rect 57 -18600 457 -18588
rect 693 -18554 1093 -18542
rect 693 -18588 705 -18554
rect 1081 -18588 1093 -18554
rect 693 -18600 1093 -18588
rect 1657 -17170 2057 -17158
rect 1657 -17204 1669 -17170
rect 2045 -17204 2057 -17170
rect 1657 -17216 2057 -17204
rect 2293 -17170 2693 -17158
rect 2293 -17204 2305 -17170
rect 2681 -17204 2693 -17170
rect 2293 -17216 2693 -17204
rect 1657 -17428 2057 -17416
rect 1657 -17462 1669 -17428
rect 2045 -17462 2057 -17428
rect 1657 -17474 2057 -17462
rect 2293 -17428 2693 -17416
rect 2293 -17462 2305 -17428
rect 2681 -17462 2693 -17428
rect 2293 -17474 2693 -17462
rect 1657 -17696 2057 -17684
rect 1657 -17730 1669 -17696
rect 2045 -17730 2057 -17696
rect 1657 -17742 2057 -17730
rect 2293 -17696 2693 -17684
rect 2293 -17730 2305 -17696
rect 2681 -17730 2693 -17696
rect 2293 -17742 2693 -17730
rect 1657 -18554 2057 -18542
rect 1657 -18588 1669 -18554
rect 2045 -18588 2057 -18554
rect 1657 -18600 2057 -18588
rect 2293 -18554 2693 -18542
rect 2293 -18588 2305 -18554
rect 2681 -18588 2693 -18554
rect 2293 -18600 2693 -18588
rect 3257 -17170 3657 -17158
rect 3257 -17204 3269 -17170
rect 3645 -17204 3657 -17170
rect 3257 -17216 3657 -17204
rect 3893 -17170 4293 -17158
rect 3893 -17204 3905 -17170
rect 4281 -17204 4293 -17170
rect 3893 -17216 4293 -17204
rect 3257 -17428 3657 -17416
rect 3257 -17462 3269 -17428
rect 3645 -17462 3657 -17428
rect 3257 -17474 3657 -17462
rect 3893 -17428 4293 -17416
rect 3893 -17462 3905 -17428
rect 4281 -17462 4293 -17428
rect 3893 -17474 4293 -17462
rect 3257 -17696 3657 -17684
rect 3257 -17730 3269 -17696
rect 3645 -17730 3657 -17696
rect 3257 -17742 3657 -17730
rect 3893 -17696 4293 -17684
rect 3893 -17730 3905 -17696
rect 4281 -17730 4293 -17696
rect 3893 -17742 4293 -17730
rect 3257 -18554 3657 -18542
rect 3257 -18588 3269 -18554
rect 3645 -18588 3657 -18554
rect 3257 -18600 3657 -18588
rect 3893 -18554 4293 -18542
rect 3893 -18588 3905 -18554
rect 4281 -18588 4293 -18554
rect 3893 -18600 4293 -18588
rect 4857 -17170 5257 -17158
rect 4857 -17204 4869 -17170
rect 5245 -17204 5257 -17170
rect 4857 -17216 5257 -17204
rect 5493 -17170 5893 -17158
rect 5493 -17204 5505 -17170
rect 5881 -17204 5893 -17170
rect 5493 -17216 5893 -17204
rect 4857 -17428 5257 -17416
rect 4857 -17462 4869 -17428
rect 5245 -17462 5257 -17428
rect 4857 -17474 5257 -17462
rect 5493 -17428 5893 -17416
rect 5493 -17462 5505 -17428
rect 5881 -17462 5893 -17428
rect 5493 -17474 5893 -17462
rect 4857 -17696 5257 -17684
rect 4857 -17730 4869 -17696
rect 5245 -17730 5257 -17696
rect 4857 -17742 5257 -17730
rect 5493 -17696 5893 -17684
rect 5493 -17730 5505 -17696
rect 5881 -17730 5893 -17696
rect 5493 -17742 5893 -17730
rect 4857 -18554 5257 -18542
rect 4857 -18588 4869 -18554
rect 5245 -18588 5257 -18554
rect 4857 -18600 5257 -18588
rect 5493 -18554 5893 -18542
rect 5493 -18588 5505 -18554
rect 5881 -18588 5893 -18554
rect 5493 -18600 5893 -18588
rect 6457 -17170 6857 -17158
rect 6457 -17204 6469 -17170
rect 6845 -17204 6857 -17170
rect 6457 -17216 6857 -17204
rect 7093 -17170 7493 -17158
rect 7093 -17204 7105 -17170
rect 7481 -17204 7493 -17170
rect 7093 -17216 7493 -17204
rect 6457 -17428 6857 -17416
rect 6457 -17462 6469 -17428
rect 6845 -17462 6857 -17428
rect 6457 -17474 6857 -17462
rect 7093 -17428 7493 -17416
rect 7093 -17462 7105 -17428
rect 7481 -17462 7493 -17428
rect 7093 -17474 7493 -17462
rect 6457 -17696 6857 -17684
rect 6457 -17730 6469 -17696
rect 6845 -17730 6857 -17696
rect 6457 -17742 6857 -17730
rect 7093 -17696 7493 -17684
rect 7093 -17730 7105 -17696
rect 7481 -17730 7493 -17696
rect 7093 -17742 7493 -17730
rect 6457 -18554 6857 -18542
rect 6457 -18588 6469 -18554
rect 6845 -18588 6857 -18554
rect 6457 -18600 6857 -18588
rect 7093 -18554 7493 -18542
rect 7093 -18588 7105 -18554
rect 7481 -18588 7493 -18554
rect 7093 -18600 7493 -18588
rect 8057 -17170 8457 -17158
rect 8057 -17204 8069 -17170
rect 8445 -17204 8457 -17170
rect 8057 -17216 8457 -17204
rect 8693 -17170 9093 -17158
rect 8693 -17204 8705 -17170
rect 9081 -17204 9093 -17170
rect 8693 -17216 9093 -17204
rect 8057 -17428 8457 -17416
rect 8057 -17462 8069 -17428
rect 8445 -17462 8457 -17428
rect 8057 -17474 8457 -17462
rect 8693 -17428 9093 -17416
rect 8693 -17462 8705 -17428
rect 9081 -17462 9093 -17428
rect 8693 -17474 9093 -17462
rect 8057 -17696 8457 -17684
rect 8057 -17730 8069 -17696
rect 8445 -17730 8457 -17696
rect 8057 -17742 8457 -17730
rect 8693 -17696 9093 -17684
rect 8693 -17730 8705 -17696
rect 9081 -17730 9093 -17696
rect 8693 -17742 9093 -17730
rect 8057 -18554 8457 -18542
rect 8057 -18588 8069 -18554
rect 8445 -18588 8457 -18554
rect 8057 -18600 8457 -18588
rect 8693 -18554 9093 -18542
rect 8693 -18588 8705 -18554
rect 9081 -18588 9093 -18554
rect 8693 -18600 9093 -18588
rect 9657 -17170 10057 -17158
rect 9657 -17204 9669 -17170
rect 10045 -17204 10057 -17170
rect 9657 -17216 10057 -17204
rect 10293 -17170 10693 -17158
rect 10293 -17204 10305 -17170
rect 10681 -17204 10693 -17170
rect 10293 -17216 10693 -17204
rect 9657 -17428 10057 -17416
rect 9657 -17462 9669 -17428
rect 10045 -17462 10057 -17428
rect 9657 -17474 10057 -17462
rect 10293 -17428 10693 -17416
rect 10293 -17462 10305 -17428
rect 10681 -17462 10693 -17428
rect 10293 -17474 10693 -17462
rect 9657 -17696 10057 -17684
rect 9657 -17730 9669 -17696
rect 10045 -17730 10057 -17696
rect 9657 -17742 10057 -17730
rect 10293 -17696 10693 -17684
rect 10293 -17730 10305 -17696
rect 10681 -17730 10693 -17696
rect 10293 -17742 10693 -17730
rect 9657 -18554 10057 -18542
rect 9657 -18588 9669 -18554
rect 10045 -18588 10057 -18554
rect 9657 -18600 10057 -18588
rect 10293 -18554 10693 -18542
rect 10293 -18588 10305 -18554
rect 10681 -18588 10693 -18554
rect 10293 -18600 10693 -18588
rect 11257 -17170 11657 -17158
rect 11257 -17204 11269 -17170
rect 11645 -17204 11657 -17170
rect 11257 -17216 11657 -17204
rect 11893 -17170 12293 -17158
rect 11893 -17204 11905 -17170
rect 12281 -17204 12293 -17170
rect 11893 -17216 12293 -17204
rect 11257 -17428 11657 -17416
rect 11257 -17462 11269 -17428
rect 11645 -17462 11657 -17428
rect 11257 -17474 11657 -17462
rect 11893 -17428 12293 -17416
rect 11893 -17462 11905 -17428
rect 12281 -17462 12293 -17428
rect 11893 -17474 12293 -17462
rect 11257 -17696 11657 -17684
rect 11257 -17730 11269 -17696
rect 11645 -17730 11657 -17696
rect 11257 -17742 11657 -17730
rect 11893 -17696 12293 -17684
rect 11893 -17730 11905 -17696
rect 12281 -17730 12293 -17696
rect 11893 -17742 12293 -17730
rect 11257 -18554 11657 -18542
rect 11257 -18588 11269 -18554
rect 11645 -18588 11657 -18554
rect 11257 -18600 11657 -18588
rect 11893 -18554 12293 -18542
rect 11893 -18588 11905 -18554
rect 12281 -18588 12293 -18554
rect 11893 -18600 12293 -18588
rect 12857 -17170 13257 -17158
rect 12857 -17204 12869 -17170
rect 13245 -17204 13257 -17170
rect 12857 -17216 13257 -17204
rect 13493 -17170 13893 -17158
rect 13493 -17204 13505 -17170
rect 13881 -17204 13893 -17170
rect 13493 -17216 13893 -17204
rect 12857 -17428 13257 -17416
rect 12857 -17462 12869 -17428
rect 13245 -17462 13257 -17428
rect 12857 -17474 13257 -17462
rect 13493 -17428 13893 -17416
rect 13493 -17462 13505 -17428
rect 13881 -17462 13893 -17428
rect 13493 -17474 13893 -17462
rect 12857 -17696 13257 -17684
rect 12857 -17730 12869 -17696
rect 13245 -17730 13257 -17696
rect 12857 -17742 13257 -17730
rect 13493 -17696 13893 -17684
rect 13493 -17730 13505 -17696
rect 13881 -17730 13893 -17696
rect 13493 -17742 13893 -17730
rect 12857 -18554 13257 -18542
rect 12857 -18588 12869 -18554
rect 13245 -18588 13257 -18554
rect 12857 -18600 13257 -18588
rect 13493 -18554 13893 -18542
rect 13493 -18588 13505 -18554
rect 13881 -18588 13893 -18554
rect 13493 -18600 13893 -18588
rect 14457 -17170 14857 -17158
rect 14457 -17204 14469 -17170
rect 14845 -17204 14857 -17170
rect 14457 -17216 14857 -17204
rect 15093 -17170 15493 -17158
rect 15093 -17204 15105 -17170
rect 15481 -17204 15493 -17170
rect 15093 -17216 15493 -17204
rect 14457 -17428 14857 -17416
rect 14457 -17462 14469 -17428
rect 14845 -17462 14857 -17428
rect 14457 -17474 14857 -17462
rect 15093 -17428 15493 -17416
rect 15093 -17462 15105 -17428
rect 15481 -17462 15493 -17428
rect 15093 -17474 15493 -17462
rect 14457 -17696 14857 -17684
rect 14457 -17730 14469 -17696
rect 14845 -17730 14857 -17696
rect 14457 -17742 14857 -17730
rect 15093 -17696 15493 -17684
rect 15093 -17730 15105 -17696
rect 15481 -17730 15493 -17696
rect 15093 -17742 15493 -17730
rect 14457 -18554 14857 -18542
rect 14457 -18588 14469 -18554
rect 14845 -18588 14857 -18554
rect 14457 -18600 14857 -18588
rect 15093 -18554 15493 -18542
rect 15093 -18588 15105 -18554
rect 15481 -18588 15493 -18554
rect 15093 -18600 15493 -18588
rect 16057 -17170 16457 -17158
rect 16057 -17204 16069 -17170
rect 16445 -17204 16457 -17170
rect 16057 -17216 16457 -17204
rect 16693 -17170 17093 -17158
rect 16693 -17204 16705 -17170
rect 17081 -17204 17093 -17170
rect 16693 -17216 17093 -17204
rect 16057 -17428 16457 -17416
rect 16057 -17462 16069 -17428
rect 16445 -17462 16457 -17428
rect 16057 -17474 16457 -17462
rect 16693 -17428 17093 -17416
rect 16693 -17462 16705 -17428
rect 17081 -17462 17093 -17428
rect 16693 -17474 17093 -17462
rect 16057 -17696 16457 -17684
rect 16057 -17730 16069 -17696
rect 16445 -17730 16457 -17696
rect 16057 -17742 16457 -17730
rect 16693 -17696 17093 -17684
rect 16693 -17730 16705 -17696
rect 17081 -17730 17093 -17696
rect 16693 -17742 17093 -17730
rect 16057 -18554 16457 -18542
rect 16057 -18588 16069 -18554
rect 16445 -18588 16457 -18554
rect 16057 -18600 16457 -18588
rect 16693 -18554 17093 -18542
rect 16693 -18588 16705 -18554
rect 17081 -18588 17093 -18554
rect 16693 -18600 17093 -18588
rect 17657 -17170 18057 -17158
rect 17657 -17204 17669 -17170
rect 18045 -17204 18057 -17170
rect 17657 -17216 18057 -17204
rect 18293 -17170 18693 -17158
rect 18293 -17204 18305 -17170
rect 18681 -17204 18693 -17170
rect 18293 -17216 18693 -17204
rect 17657 -17428 18057 -17416
rect 17657 -17462 17669 -17428
rect 18045 -17462 18057 -17428
rect 17657 -17474 18057 -17462
rect 18293 -17428 18693 -17416
rect 18293 -17462 18305 -17428
rect 18681 -17462 18693 -17428
rect 18293 -17474 18693 -17462
rect 17657 -17696 18057 -17684
rect 17657 -17730 17669 -17696
rect 18045 -17730 18057 -17696
rect 17657 -17742 18057 -17730
rect 18293 -17696 18693 -17684
rect 18293 -17730 18305 -17696
rect 18681 -17730 18693 -17696
rect 18293 -17742 18693 -17730
rect 17657 -18554 18057 -18542
rect 17657 -18588 17669 -18554
rect 18045 -18588 18057 -18554
rect 17657 -18600 18057 -18588
rect 18293 -18554 18693 -18542
rect 18293 -18588 18305 -18554
rect 18681 -18588 18693 -18554
rect 18293 -18600 18693 -18588
rect 19257 -17170 19657 -17158
rect 19257 -17204 19269 -17170
rect 19645 -17204 19657 -17170
rect 19257 -17216 19657 -17204
rect 19893 -17170 20293 -17158
rect 19893 -17204 19905 -17170
rect 20281 -17204 20293 -17170
rect 19893 -17216 20293 -17204
rect 19257 -17428 19657 -17416
rect 19257 -17462 19269 -17428
rect 19645 -17462 19657 -17428
rect 19257 -17474 19657 -17462
rect 19893 -17428 20293 -17416
rect 19893 -17462 19905 -17428
rect 20281 -17462 20293 -17428
rect 19893 -17474 20293 -17462
rect 19257 -17696 19657 -17684
rect 19257 -17730 19269 -17696
rect 19645 -17730 19657 -17696
rect 19257 -17742 19657 -17730
rect 19893 -17696 20293 -17684
rect 19893 -17730 19905 -17696
rect 20281 -17730 20293 -17696
rect 19893 -17742 20293 -17730
rect 19257 -18554 19657 -18542
rect 19257 -18588 19269 -18554
rect 19645 -18588 19657 -18554
rect 19257 -18600 19657 -18588
rect 19893 -18554 20293 -18542
rect 19893 -18588 19905 -18554
rect 20281 -18588 20293 -18554
rect 19893 -18600 20293 -18588
rect 20857 -17170 21257 -17158
rect 20857 -17204 20869 -17170
rect 21245 -17204 21257 -17170
rect 20857 -17216 21257 -17204
rect 21493 -17170 21893 -17158
rect 21493 -17204 21505 -17170
rect 21881 -17204 21893 -17170
rect 21493 -17216 21893 -17204
rect 20857 -17428 21257 -17416
rect 20857 -17462 20869 -17428
rect 21245 -17462 21257 -17428
rect 20857 -17474 21257 -17462
rect 21493 -17428 21893 -17416
rect 21493 -17462 21505 -17428
rect 21881 -17462 21893 -17428
rect 21493 -17474 21893 -17462
rect 20857 -17696 21257 -17684
rect 20857 -17730 20869 -17696
rect 21245 -17730 21257 -17696
rect 20857 -17742 21257 -17730
rect 21493 -17696 21893 -17684
rect 21493 -17730 21505 -17696
rect 21881 -17730 21893 -17696
rect 21493 -17742 21893 -17730
rect 20857 -18554 21257 -18542
rect 20857 -18588 20869 -18554
rect 21245 -18588 21257 -18554
rect 20857 -18600 21257 -18588
rect 21493 -18554 21893 -18542
rect 21493 -18588 21505 -18554
rect 21881 -18588 21893 -18554
rect 21493 -18600 21893 -18588
rect 22457 -17170 22857 -17158
rect 22457 -17204 22469 -17170
rect 22845 -17204 22857 -17170
rect 22457 -17216 22857 -17204
rect 23093 -17170 23493 -17158
rect 23093 -17204 23105 -17170
rect 23481 -17204 23493 -17170
rect 23093 -17216 23493 -17204
rect 22457 -17428 22857 -17416
rect 22457 -17462 22469 -17428
rect 22845 -17462 22857 -17428
rect 22457 -17474 22857 -17462
rect 23093 -17428 23493 -17416
rect 23093 -17462 23105 -17428
rect 23481 -17462 23493 -17428
rect 23093 -17474 23493 -17462
rect 22457 -17696 22857 -17684
rect 22457 -17730 22469 -17696
rect 22845 -17730 22857 -17696
rect 22457 -17742 22857 -17730
rect 23093 -17696 23493 -17684
rect 23093 -17730 23105 -17696
rect 23481 -17730 23493 -17696
rect 23093 -17742 23493 -17730
rect 22457 -18554 22857 -18542
rect 22457 -18588 22469 -18554
rect 22845 -18588 22857 -18554
rect 22457 -18600 22857 -18588
rect 23093 -18554 23493 -18542
rect 23093 -18588 23105 -18554
rect 23481 -18588 23493 -18554
rect 23093 -18600 23493 -18588
rect 24057 -17170 24457 -17158
rect 24057 -17204 24069 -17170
rect 24445 -17204 24457 -17170
rect 24057 -17216 24457 -17204
rect 24693 -17170 25093 -17158
rect 24693 -17204 24705 -17170
rect 25081 -17204 25093 -17170
rect 24693 -17216 25093 -17204
rect 24057 -17428 24457 -17416
rect 24057 -17462 24069 -17428
rect 24445 -17462 24457 -17428
rect 24057 -17474 24457 -17462
rect 24693 -17428 25093 -17416
rect 24693 -17462 24705 -17428
rect 25081 -17462 25093 -17428
rect 24693 -17474 25093 -17462
rect 24057 -17696 24457 -17684
rect 24057 -17730 24069 -17696
rect 24445 -17730 24457 -17696
rect 24057 -17742 24457 -17730
rect 24693 -17696 25093 -17684
rect 24693 -17730 24705 -17696
rect 25081 -17730 25093 -17696
rect 24693 -17742 25093 -17730
rect 24057 -18554 24457 -18542
rect 24057 -18588 24069 -18554
rect 24445 -18588 24457 -18554
rect 24057 -18600 24457 -18588
rect 24693 -18554 25093 -18542
rect 24693 -18588 24705 -18554
rect 25081 -18588 25093 -18554
rect 24693 -18600 25093 -18588
rect 25657 -17170 26057 -17158
rect 25657 -17204 25669 -17170
rect 26045 -17204 26057 -17170
rect 25657 -17216 26057 -17204
rect 26293 -17170 26693 -17158
rect 26293 -17204 26305 -17170
rect 26681 -17204 26693 -17170
rect 26293 -17216 26693 -17204
rect 25657 -17428 26057 -17416
rect 25657 -17462 25669 -17428
rect 26045 -17462 26057 -17428
rect 25657 -17474 26057 -17462
rect 26293 -17428 26693 -17416
rect 26293 -17462 26305 -17428
rect 26681 -17462 26693 -17428
rect 26293 -17474 26693 -17462
rect 25657 -17696 26057 -17684
rect 25657 -17730 25669 -17696
rect 26045 -17730 26057 -17696
rect 25657 -17742 26057 -17730
rect 26293 -17696 26693 -17684
rect 26293 -17730 26305 -17696
rect 26681 -17730 26693 -17696
rect 26293 -17742 26693 -17730
rect 25657 -18554 26057 -18542
rect 25657 -18588 25669 -18554
rect 26045 -18588 26057 -18554
rect 25657 -18600 26057 -18588
rect 26293 -18554 26693 -18542
rect 26293 -18588 26305 -18554
rect 26681 -18588 26693 -18554
rect 26293 -18600 26693 -18588
rect 27257 -17170 27657 -17158
rect 27257 -17204 27269 -17170
rect 27645 -17204 27657 -17170
rect 27257 -17216 27657 -17204
rect 27893 -17170 28293 -17158
rect 27893 -17204 27905 -17170
rect 28281 -17204 28293 -17170
rect 27893 -17216 28293 -17204
rect 27257 -17428 27657 -17416
rect 27257 -17462 27269 -17428
rect 27645 -17462 27657 -17428
rect 27257 -17474 27657 -17462
rect 27893 -17428 28293 -17416
rect 27893 -17462 27905 -17428
rect 28281 -17462 28293 -17428
rect 27893 -17474 28293 -17462
rect 27257 -17696 27657 -17684
rect 27257 -17730 27269 -17696
rect 27645 -17730 27657 -17696
rect 27257 -17742 27657 -17730
rect 27893 -17696 28293 -17684
rect 27893 -17730 27905 -17696
rect 28281 -17730 28293 -17696
rect 27893 -17742 28293 -17730
rect 27257 -18554 27657 -18542
rect 27257 -18588 27269 -18554
rect 27645 -18588 27657 -18554
rect 27257 -18600 27657 -18588
rect 27893 -18554 28293 -18542
rect 27893 -18588 27905 -18554
rect 28281 -18588 28293 -18554
rect 27893 -18600 28293 -18588
rect 28857 -17170 29257 -17158
rect 28857 -17204 28869 -17170
rect 29245 -17204 29257 -17170
rect 28857 -17216 29257 -17204
rect 29493 -17170 29893 -17158
rect 29493 -17204 29505 -17170
rect 29881 -17204 29893 -17170
rect 29493 -17216 29893 -17204
rect 28857 -17428 29257 -17416
rect 28857 -17462 28869 -17428
rect 29245 -17462 29257 -17428
rect 28857 -17474 29257 -17462
rect 29493 -17428 29893 -17416
rect 29493 -17462 29505 -17428
rect 29881 -17462 29893 -17428
rect 29493 -17474 29893 -17462
rect 28857 -17696 29257 -17684
rect 28857 -17730 28869 -17696
rect 29245 -17730 29257 -17696
rect 28857 -17742 29257 -17730
rect 29493 -17696 29893 -17684
rect 29493 -17730 29505 -17696
rect 29881 -17730 29893 -17696
rect 29493 -17742 29893 -17730
rect 28857 -18554 29257 -18542
rect 28857 -18588 28869 -18554
rect 29245 -18588 29257 -18554
rect 28857 -18600 29257 -18588
rect 29493 -18554 29893 -18542
rect 29493 -18588 29505 -18554
rect 29881 -18588 29893 -18554
rect 29493 -18600 29893 -18588
rect 30457 -17170 30857 -17158
rect 30457 -17204 30469 -17170
rect 30845 -17204 30857 -17170
rect 30457 -17216 30857 -17204
rect 31093 -17170 31493 -17158
rect 31093 -17204 31105 -17170
rect 31481 -17204 31493 -17170
rect 31093 -17216 31493 -17204
rect 30457 -17428 30857 -17416
rect 30457 -17462 30469 -17428
rect 30845 -17462 30857 -17428
rect 30457 -17474 30857 -17462
rect 31093 -17428 31493 -17416
rect 31093 -17462 31105 -17428
rect 31481 -17462 31493 -17428
rect 31093 -17474 31493 -17462
rect 30457 -17696 30857 -17684
rect 30457 -17730 30469 -17696
rect 30845 -17730 30857 -17696
rect 30457 -17742 30857 -17730
rect 31093 -17696 31493 -17684
rect 31093 -17730 31105 -17696
rect 31481 -17730 31493 -17696
rect 31093 -17742 31493 -17730
rect 30457 -18554 30857 -18542
rect 30457 -18588 30469 -18554
rect 30845 -18588 30857 -18554
rect 30457 -18600 30857 -18588
rect 31093 -18554 31493 -18542
rect 31093 -18588 31105 -18554
rect 31481 -18588 31493 -18554
rect 31093 -18600 31493 -18588
rect 32057 -17170 32457 -17158
rect 32057 -17204 32069 -17170
rect 32445 -17204 32457 -17170
rect 32057 -17216 32457 -17204
rect 32693 -17170 33093 -17158
rect 32693 -17204 32705 -17170
rect 33081 -17204 33093 -17170
rect 32693 -17216 33093 -17204
rect 32057 -17428 32457 -17416
rect 32057 -17462 32069 -17428
rect 32445 -17462 32457 -17428
rect 32057 -17474 32457 -17462
rect 32693 -17428 33093 -17416
rect 32693 -17462 32705 -17428
rect 33081 -17462 33093 -17428
rect 32693 -17474 33093 -17462
rect 32057 -17696 32457 -17684
rect 32057 -17730 32069 -17696
rect 32445 -17730 32457 -17696
rect 32057 -17742 32457 -17730
rect 32693 -17696 33093 -17684
rect 32693 -17730 32705 -17696
rect 33081 -17730 33093 -17696
rect 32693 -17742 33093 -17730
rect 32057 -18554 32457 -18542
rect 32057 -18588 32069 -18554
rect 32445 -18588 32457 -18554
rect 32057 -18600 32457 -18588
rect 32693 -18554 33093 -18542
rect 32693 -18588 32705 -18554
rect 33081 -18588 33093 -18554
rect 32693 -18600 33093 -18588
rect 33657 -17170 34057 -17158
rect 33657 -17204 33669 -17170
rect 34045 -17204 34057 -17170
rect 33657 -17216 34057 -17204
rect 34293 -17170 34693 -17158
rect 34293 -17204 34305 -17170
rect 34681 -17204 34693 -17170
rect 34293 -17216 34693 -17204
rect 33657 -17428 34057 -17416
rect 33657 -17462 33669 -17428
rect 34045 -17462 34057 -17428
rect 33657 -17474 34057 -17462
rect 34293 -17428 34693 -17416
rect 34293 -17462 34305 -17428
rect 34681 -17462 34693 -17428
rect 34293 -17474 34693 -17462
rect 33657 -17696 34057 -17684
rect 33657 -17730 33669 -17696
rect 34045 -17730 34057 -17696
rect 33657 -17742 34057 -17730
rect 34293 -17696 34693 -17684
rect 34293 -17730 34305 -17696
rect 34681 -17730 34693 -17696
rect 34293 -17742 34693 -17730
rect 33657 -18554 34057 -18542
rect 33657 -18588 33669 -18554
rect 34045 -18588 34057 -18554
rect 33657 -18600 34057 -18588
rect 34293 -18554 34693 -18542
rect 34293 -18588 34305 -18554
rect 34681 -18588 34693 -18554
rect 34293 -18600 34693 -18588
rect 35257 -17170 35657 -17158
rect 35257 -17204 35269 -17170
rect 35645 -17204 35657 -17170
rect 35257 -17216 35657 -17204
rect 35893 -17170 36293 -17158
rect 35893 -17204 35905 -17170
rect 36281 -17204 36293 -17170
rect 35893 -17216 36293 -17204
rect 35257 -17428 35657 -17416
rect 35257 -17462 35269 -17428
rect 35645 -17462 35657 -17428
rect 35257 -17474 35657 -17462
rect 35893 -17428 36293 -17416
rect 35893 -17462 35905 -17428
rect 36281 -17462 36293 -17428
rect 35893 -17474 36293 -17462
rect 35257 -17696 35657 -17684
rect 35257 -17730 35269 -17696
rect 35645 -17730 35657 -17696
rect 35257 -17742 35657 -17730
rect 35893 -17696 36293 -17684
rect 35893 -17730 35905 -17696
rect 36281 -17730 36293 -17696
rect 35893 -17742 36293 -17730
rect 35257 -18554 35657 -18542
rect 35257 -18588 35269 -18554
rect 35645 -18588 35657 -18554
rect 35257 -18600 35657 -18588
rect 35893 -18554 36293 -18542
rect 35893 -18588 35905 -18554
rect 36281 -18588 36293 -18554
rect 35893 -18600 36293 -18588
rect 36857 -17170 37257 -17158
rect 36857 -17204 36869 -17170
rect 37245 -17204 37257 -17170
rect 36857 -17216 37257 -17204
rect 37493 -17170 37893 -17158
rect 37493 -17204 37505 -17170
rect 37881 -17204 37893 -17170
rect 37493 -17216 37893 -17204
rect 36857 -17428 37257 -17416
rect 36857 -17462 36869 -17428
rect 37245 -17462 37257 -17428
rect 36857 -17474 37257 -17462
rect 37493 -17428 37893 -17416
rect 37493 -17462 37505 -17428
rect 37881 -17462 37893 -17428
rect 37493 -17474 37893 -17462
rect 36857 -17696 37257 -17684
rect 36857 -17730 36869 -17696
rect 37245 -17730 37257 -17696
rect 36857 -17742 37257 -17730
rect 37493 -17696 37893 -17684
rect 37493 -17730 37505 -17696
rect 37881 -17730 37893 -17696
rect 37493 -17742 37893 -17730
rect 36857 -18554 37257 -18542
rect 36857 -18588 36869 -18554
rect 37245 -18588 37257 -18554
rect 36857 -18600 37257 -18588
rect 37493 -18554 37893 -18542
rect 37493 -18588 37505 -18554
rect 37881 -18588 37893 -18554
rect 37493 -18600 37893 -18588
rect 57 -18970 457 -18958
rect 57 -19004 69 -18970
rect 445 -19004 457 -18970
rect 57 -19016 457 -19004
rect 693 -18970 1093 -18958
rect 693 -19004 705 -18970
rect 1081 -19004 1093 -18970
rect 693 -19016 1093 -19004
rect 57 -19228 457 -19216
rect 57 -19262 69 -19228
rect 445 -19262 457 -19228
rect 57 -19274 457 -19262
rect 693 -19228 1093 -19216
rect 693 -19262 705 -19228
rect 1081 -19262 1093 -19228
rect 693 -19274 1093 -19262
rect 57 -19496 457 -19484
rect 57 -19530 69 -19496
rect 445 -19530 457 -19496
rect 57 -19542 457 -19530
rect 693 -19496 1093 -19484
rect 693 -19530 705 -19496
rect 1081 -19530 1093 -19496
rect 693 -19542 1093 -19530
rect 57 -20354 457 -20342
rect 57 -20388 69 -20354
rect 445 -20388 457 -20354
rect 57 -20400 457 -20388
rect 693 -20354 1093 -20342
rect 693 -20388 705 -20354
rect 1081 -20388 1093 -20354
rect 693 -20400 1093 -20388
rect 1657 -18970 2057 -18958
rect 1657 -19004 1669 -18970
rect 2045 -19004 2057 -18970
rect 1657 -19016 2057 -19004
rect 2293 -18970 2693 -18958
rect 2293 -19004 2305 -18970
rect 2681 -19004 2693 -18970
rect 2293 -19016 2693 -19004
rect 1657 -19228 2057 -19216
rect 1657 -19262 1669 -19228
rect 2045 -19262 2057 -19228
rect 1657 -19274 2057 -19262
rect 2293 -19228 2693 -19216
rect 2293 -19262 2305 -19228
rect 2681 -19262 2693 -19228
rect 2293 -19274 2693 -19262
rect 1657 -19496 2057 -19484
rect 1657 -19530 1669 -19496
rect 2045 -19530 2057 -19496
rect 1657 -19542 2057 -19530
rect 2293 -19496 2693 -19484
rect 2293 -19530 2305 -19496
rect 2681 -19530 2693 -19496
rect 2293 -19542 2693 -19530
rect 1657 -20354 2057 -20342
rect 1657 -20388 1669 -20354
rect 2045 -20388 2057 -20354
rect 1657 -20400 2057 -20388
rect 2293 -20354 2693 -20342
rect 2293 -20388 2305 -20354
rect 2681 -20388 2693 -20354
rect 2293 -20400 2693 -20388
rect 3257 -18970 3657 -18958
rect 3257 -19004 3269 -18970
rect 3645 -19004 3657 -18970
rect 3257 -19016 3657 -19004
rect 3893 -18970 4293 -18958
rect 3893 -19004 3905 -18970
rect 4281 -19004 4293 -18970
rect 3893 -19016 4293 -19004
rect 3257 -19228 3657 -19216
rect 3257 -19262 3269 -19228
rect 3645 -19262 3657 -19228
rect 3257 -19274 3657 -19262
rect 3893 -19228 4293 -19216
rect 3893 -19262 3905 -19228
rect 4281 -19262 4293 -19228
rect 3893 -19274 4293 -19262
rect 3257 -19496 3657 -19484
rect 3257 -19530 3269 -19496
rect 3645 -19530 3657 -19496
rect 3257 -19542 3657 -19530
rect 3893 -19496 4293 -19484
rect 3893 -19530 3905 -19496
rect 4281 -19530 4293 -19496
rect 3893 -19542 4293 -19530
rect 3257 -20354 3657 -20342
rect 3257 -20388 3269 -20354
rect 3645 -20388 3657 -20354
rect 3257 -20400 3657 -20388
rect 3893 -20354 4293 -20342
rect 3893 -20388 3905 -20354
rect 4281 -20388 4293 -20354
rect 3893 -20400 4293 -20388
rect 4857 -18970 5257 -18958
rect 4857 -19004 4869 -18970
rect 5245 -19004 5257 -18970
rect 4857 -19016 5257 -19004
rect 5493 -18970 5893 -18958
rect 5493 -19004 5505 -18970
rect 5881 -19004 5893 -18970
rect 5493 -19016 5893 -19004
rect 4857 -19228 5257 -19216
rect 4857 -19262 4869 -19228
rect 5245 -19262 5257 -19228
rect 4857 -19274 5257 -19262
rect 5493 -19228 5893 -19216
rect 5493 -19262 5505 -19228
rect 5881 -19262 5893 -19228
rect 5493 -19274 5893 -19262
rect 4857 -19496 5257 -19484
rect 4857 -19530 4869 -19496
rect 5245 -19530 5257 -19496
rect 4857 -19542 5257 -19530
rect 5493 -19496 5893 -19484
rect 5493 -19530 5505 -19496
rect 5881 -19530 5893 -19496
rect 5493 -19542 5893 -19530
rect 4857 -20354 5257 -20342
rect 4857 -20388 4869 -20354
rect 5245 -20388 5257 -20354
rect 4857 -20400 5257 -20388
rect 5493 -20354 5893 -20342
rect 5493 -20388 5505 -20354
rect 5881 -20388 5893 -20354
rect 5493 -20400 5893 -20388
rect 6457 -18970 6857 -18958
rect 6457 -19004 6469 -18970
rect 6845 -19004 6857 -18970
rect 6457 -19016 6857 -19004
rect 7093 -18970 7493 -18958
rect 7093 -19004 7105 -18970
rect 7481 -19004 7493 -18970
rect 7093 -19016 7493 -19004
rect 6457 -19228 6857 -19216
rect 6457 -19262 6469 -19228
rect 6845 -19262 6857 -19228
rect 6457 -19274 6857 -19262
rect 7093 -19228 7493 -19216
rect 7093 -19262 7105 -19228
rect 7481 -19262 7493 -19228
rect 7093 -19274 7493 -19262
rect 6457 -19496 6857 -19484
rect 6457 -19530 6469 -19496
rect 6845 -19530 6857 -19496
rect 6457 -19542 6857 -19530
rect 7093 -19496 7493 -19484
rect 7093 -19530 7105 -19496
rect 7481 -19530 7493 -19496
rect 7093 -19542 7493 -19530
rect 6457 -20354 6857 -20342
rect 6457 -20388 6469 -20354
rect 6845 -20388 6857 -20354
rect 6457 -20400 6857 -20388
rect 7093 -20354 7493 -20342
rect 7093 -20388 7105 -20354
rect 7481 -20388 7493 -20354
rect 7093 -20400 7493 -20388
rect 8057 -18970 8457 -18958
rect 8057 -19004 8069 -18970
rect 8445 -19004 8457 -18970
rect 8057 -19016 8457 -19004
rect 8693 -18970 9093 -18958
rect 8693 -19004 8705 -18970
rect 9081 -19004 9093 -18970
rect 8693 -19016 9093 -19004
rect 8057 -19228 8457 -19216
rect 8057 -19262 8069 -19228
rect 8445 -19262 8457 -19228
rect 8057 -19274 8457 -19262
rect 8693 -19228 9093 -19216
rect 8693 -19262 8705 -19228
rect 9081 -19262 9093 -19228
rect 8693 -19274 9093 -19262
rect 8057 -19496 8457 -19484
rect 8057 -19530 8069 -19496
rect 8445 -19530 8457 -19496
rect 8057 -19542 8457 -19530
rect 8693 -19496 9093 -19484
rect 8693 -19530 8705 -19496
rect 9081 -19530 9093 -19496
rect 8693 -19542 9093 -19530
rect 8057 -20354 8457 -20342
rect 8057 -20388 8069 -20354
rect 8445 -20388 8457 -20354
rect 8057 -20400 8457 -20388
rect 8693 -20354 9093 -20342
rect 8693 -20388 8705 -20354
rect 9081 -20388 9093 -20354
rect 8693 -20400 9093 -20388
rect 9657 -18970 10057 -18958
rect 9657 -19004 9669 -18970
rect 10045 -19004 10057 -18970
rect 9657 -19016 10057 -19004
rect 10293 -18970 10693 -18958
rect 10293 -19004 10305 -18970
rect 10681 -19004 10693 -18970
rect 10293 -19016 10693 -19004
rect 9657 -19228 10057 -19216
rect 9657 -19262 9669 -19228
rect 10045 -19262 10057 -19228
rect 9657 -19274 10057 -19262
rect 10293 -19228 10693 -19216
rect 10293 -19262 10305 -19228
rect 10681 -19262 10693 -19228
rect 10293 -19274 10693 -19262
rect 9657 -19496 10057 -19484
rect 9657 -19530 9669 -19496
rect 10045 -19530 10057 -19496
rect 9657 -19542 10057 -19530
rect 10293 -19496 10693 -19484
rect 10293 -19530 10305 -19496
rect 10681 -19530 10693 -19496
rect 10293 -19542 10693 -19530
rect 9657 -20354 10057 -20342
rect 9657 -20388 9669 -20354
rect 10045 -20388 10057 -20354
rect 9657 -20400 10057 -20388
rect 10293 -20354 10693 -20342
rect 10293 -20388 10305 -20354
rect 10681 -20388 10693 -20354
rect 10293 -20400 10693 -20388
rect 11257 -18970 11657 -18958
rect 11257 -19004 11269 -18970
rect 11645 -19004 11657 -18970
rect 11257 -19016 11657 -19004
rect 11893 -18970 12293 -18958
rect 11893 -19004 11905 -18970
rect 12281 -19004 12293 -18970
rect 11893 -19016 12293 -19004
rect 11257 -19228 11657 -19216
rect 11257 -19262 11269 -19228
rect 11645 -19262 11657 -19228
rect 11257 -19274 11657 -19262
rect 11893 -19228 12293 -19216
rect 11893 -19262 11905 -19228
rect 12281 -19262 12293 -19228
rect 11893 -19274 12293 -19262
rect 11257 -19496 11657 -19484
rect 11257 -19530 11269 -19496
rect 11645 -19530 11657 -19496
rect 11257 -19542 11657 -19530
rect 11893 -19496 12293 -19484
rect 11893 -19530 11905 -19496
rect 12281 -19530 12293 -19496
rect 11893 -19542 12293 -19530
rect 11257 -20354 11657 -20342
rect 11257 -20388 11269 -20354
rect 11645 -20388 11657 -20354
rect 11257 -20400 11657 -20388
rect 11893 -20354 12293 -20342
rect 11893 -20388 11905 -20354
rect 12281 -20388 12293 -20354
rect 11893 -20400 12293 -20388
rect 12857 -18970 13257 -18958
rect 12857 -19004 12869 -18970
rect 13245 -19004 13257 -18970
rect 12857 -19016 13257 -19004
rect 13493 -18970 13893 -18958
rect 13493 -19004 13505 -18970
rect 13881 -19004 13893 -18970
rect 13493 -19016 13893 -19004
rect 12857 -19228 13257 -19216
rect 12857 -19262 12869 -19228
rect 13245 -19262 13257 -19228
rect 12857 -19274 13257 -19262
rect 13493 -19228 13893 -19216
rect 13493 -19262 13505 -19228
rect 13881 -19262 13893 -19228
rect 13493 -19274 13893 -19262
rect 12857 -19496 13257 -19484
rect 12857 -19530 12869 -19496
rect 13245 -19530 13257 -19496
rect 12857 -19542 13257 -19530
rect 13493 -19496 13893 -19484
rect 13493 -19530 13505 -19496
rect 13881 -19530 13893 -19496
rect 13493 -19542 13893 -19530
rect 12857 -20354 13257 -20342
rect 12857 -20388 12869 -20354
rect 13245 -20388 13257 -20354
rect 12857 -20400 13257 -20388
rect 13493 -20354 13893 -20342
rect 13493 -20388 13505 -20354
rect 13881 -20388 13893 -20354
rect 13493 -20400 13893 -20388
rect 14457 -18970 14857 -18958
rect 14457 -19004 14469 -18970
rect 14845 -19004 14857 -18970
rect 14457 -19016 14857 -19004
rect 15093 -18970 15493 -18958
rect 15093 -19004 15105 -18970
rect 15481 -19004 15493 -18970
rect 15093 -19016 15493 -19004
rect 14457 -19228 14857 -19216
rect 14457 -19262 14469 -19228
rect 14845 -19262 14857 -19228
rect 14457 -19274 14857 -19262
rect 15093 -19228 15493 -19216
rect 15093 -19262 15105 -19228
rect 15481 -19262 15493 -19228
rect 15093 -19274 15493 -19262
rect 14457 -19496 14857 -19484
rect 14457 -19530 14469 -19496
rect 14845 -19530 14857 -19496
rect 14457 -19542 14857 -19530
rect 15093 -19496 15493 -19484
rect 15093 -19530 15105 -19496
rect 15481 -19530 15493 -19496
rect 15093 -19542 15493 -19530
rect 14457 -20354 14857 -20342
rect 14457 -20388 14469 -20354
rect 14845 -20388 14857 -20354
rect 14457 -20400 14857 -20388
rect 15093 -20354 15493 -20342
rect 15093 -20388 15105 -20354
rect 15481 -20388 15493 -20354
rect 15093 -20400 15493 -20388
rect 16057 -18970 16457 -18958
rect 16057 -19004 16069 -18970
rect 16445 -19004 16457 -18970
rect 16057 -19016 16457 -19004
rect 16693 -18970 17093 -18958
rect 16693 -19004 16705 -18970
rect 17081 -19004 17093 -18970
rect 16693 -19016 17093 -19004
rect 16057 -19228 16457 -19216
rect 16057 -19262 16069 -19228
rect 16445 -19262 16457 -19228
rect 16057 -19274 16457 -19262
rect 16693 -19228 17093 -19216
rect 16693 -19262 16705 -19228
rect 17081 -19262 17093 -19228
rect 16693 -19274 17093 -19262
rect 16057 -19496 16457 -19484
rect 16057 -19530 16069 -19496
rect 16445 -19530 16457 -19496
rect 16057 -19542 16457 -19530
rect 16693 -19496 17093 -19484
rect 16693 -19530 16705 -19496
rect 17081 -19530 17093 -19496
rect 16693 -19542 17093 -19530
rect 16057 -20354 16457 -20342
rect 16057 -20388 16069 -20354
rect 16445 -20388 16457 -20354
rect 16057 -20400 16457 -20388
rect 16693 -20354 17093 -20342
rect 16693 -20388 16705 -20354
rect 17081 -20388 17093 -20354
rect 16693 -20400 17093 -20388
rect 17657 -18970 18057 -18958
rect 17657 -19004 17669 -18970
rect 18045 -19004 18057 -18970
rect 17657 -19016 18057 -19004
rect 18293 -18970 18693 -18958
rect 18293 -19004 18305 -18970
rect 18681 -19004 18693 -18970
rect 18293 -19016 18693 -19004
rect 17657 -19228 18057 -19216
rect 17657 -19262 17669 -19228
rect 18045 -19262 18057 -19228
rect 17657 -19274 18057 -19262
rect 18293 -19228 18693 -19216
rect 18293 -19262 18305 -19228
rect 18681 -19262 18693 -19228
rect 18293 -19274 18693 -19262
rect 17657 -19496 18057 -19484
rect 17657 -19530 17669 -19496
rect 18045 -19530 18057 -19496
rect 17657 -19542 18057 -19530
rect 18293 -19496 18693 -19484
rect 18293 -19530 18305 -19496
rect 18681 -19530 18693 -19496
rect 18293 -19542 18693 -19530
rect 17657 -20354 18057 -20342
rect 17657 -20388 17669 -20354
rect 18045 -20388 18057 -20354
rect 17657 -20400 18057 -20388
rect 18293 -20354 18693 -20342
rect 18293 -20388 18305 -20354
rect 18681 -20388 18693 -20354
rect 18293 -20400 18693 -20388
rect 19257 -18970 19657 -18958
rect 19257 -19004 19269 -18970
rect 19645 -19004 19657 -18970
rect 19257 -19016 19657 -19004
rect 19893 -18970 20293 -18958
rect 19893 -19004 19905 -18970
rect 20281 -19004 20293 -18970
rect 19893 -19016 20293 -19004
rect 19257 -19228 19657 -19216
rect 19257 -19262 19269 -19228
rect 19645 -19262 19657 -19228
rect 19257 -19274 19657 -19262
rect 19893 -19228 20293 -19216
rect 19893 -19262 19905 -19228
rect 20281 -19262 20293 -19228
rect 19893 -19274 20293 -19262
rect 19257 -19496 19657 -19484
rect 19257 -19530 19269 -19496
rect 19645 -19530 19657 -19496
rect 19257 -19542 19657 -19530
rect 19893 -19496 20293 -19484
rect 19893 -19530 19905 -19496
rect 20281 -19530 20293 -19496
rect 19893 -19542 20293 -19530
rect 19257 -20354 19657 -20342
rect 19257 -20388 19269 -20354
rect 19645 -20388 19657 -20354
rect 19257 -20400 19657 -20388
rect 19893 -20354 20293 -20342
rect 19893 -20388 19905 -20354
rect 20281 -20388 20293 -20354
rect 19893 -20400 20293 -20388
rect 20857 -18970 21257 -18958
rect 20857 -19004 20869 -18970
rect 21245 -19004 21257 -18970
rect 20857 -19016 21257 -19004
rect 21493 -18970 21893 -18958
rect 21493 -19004 21505 -18970
rect 21881 -19004 21893 -18970
rect 21493 -19016 21893 -19004
rect 20857 -19228 21257 -19216
rect 20857 -19262 20869 -19228
rect 21245 -19262 21257 -19228
rect 20857 -19274 21257 -19262
rect 21493 -19228 21893 -19216
rect 21493 -19262 21505 -19228
rect 21881 -19262 21893 -19228
rect 21493 -19274 21893 -19262
rect 20857 -19496 21257 -19484
rect 20857 -19530 20869 -19496
rect 21245 -19530 21257 -19496
rect 20857 -19542 21257 -19530
rect 21493 -19496 21893 -19484
rect 21493 -19530 21505 -19496
rect 21881 -19530 21893 -19496
rect 21493 -19542 21893 -19530
rect 20857 -20354 21257 -20342
rect 20857 -20388 20869 -20354
rect 21245 -20388 21257 -20354
rect 20857 -20400 21257 -20388
rect 21493 -20354 21893 -20342
rect 21493 -20388 21505 -20354
rect 21881 -20388 21893 -20354
rect 21493 -20400 21893 -20388
rect 22457 -18970 22857 -18958
rect 22457 -19004 22469 -18970
rect 22845 -19004 22857 -18970
rect 22457 -19016 22857 -19004
rect 23093 -18970 23493 -18958
rect 23093 -19004 23105 -18970
rect 23481 -19004 23493 -18970
rect 23093 -19016 23493 -19004
rect 22457 -19228 22857 -19216
rect 22457 -19262 22469 -19228
rect 22845 -19262 22857 -19228
rect 22457 -19274 22857 -19262
rect 23093 -19228 23493 -19216
rect 23093 -19262 23105 -19228
rect 23481 -19262 23493 -19228
rect 23093 -19274 23493 -19262
rect 22457 -19496 22857 -19484
rect 22457 -19530 22469 -19496
rect 22845 -19530 22857 -19496
rect 22457 -19542 22857 -19530
rect 23093 -19496 23493 -19484
rect 23093 -19530 23105 -19496
rect 23481 -19530 23493 -19496
rect 23093 -19542 23493 -19530
rect 22457 -20354 22857 -20342
rect 22457 -20388 22469 -20354
rect 22845 -20388 22857 -20354
rect 22457 -20400 22857 -20388
rect 23093 -20354 23493 -20342
rect 23093 -20388 23105 -20354
rect 23481 -20388 23493 -20354
rect 23093 -20400 23493 -20388
rect 24057 -18970 24457 -18958
rect 24057 -19004 24069 -18970
rect 24445 -19004 24457 -18970
rect 24057 -19016 24457 -19004
rect 24693 -18970 25093 -18958
rect 24693 -19004 24705 -18970
rect 25081 -19004 25093 -18970
rect 24693 -19016 25093 -19004
rect 24057 -19228 24457 -19216
rect 24057 -19262 24069 -19228
rect 24445 -19262 24457 -19228
rect 24057 -19274 24457 -19262
rect 24693 -19228 25093 -19216
rect 24693 -19262 24705 -19228
rect 25081 -19262 25093 -19228
rect 24693 -19274 25093 -19262
rect 24057 -19496 24457 -19484
rect 24057 -19530 24069 -19496
rect 24445 -19530 24457 -19496
rect 24057 -19542 24457 -19530
rect 24693 -19496 25093 -19484
rect 24693 -19530 24705 -19496
rect 25081 -19530 25093 -19496
rect 24693 -19542 25093 -19530
rect 24057 -20354 24457 -20342
rect 24057 -20388 24069 -20354
rect 24445 -20388 24457 -20354
rect 24057 -20400 24457 -20388
rect 24693 -20354 25093 -20342
rect 24693 -20388 24705 -20354
rect 25081 -20388 25093 -20354
rect 24693 -20400 25093 -20388
rect 25657 -18970 26057 -18958
rect 25657 -19004 25669 -18970
rect 26045 -19004 26057 -18970
rect 25657 -19016 26057 -19004
rect 26293 -18970 26693 -18958
rect 26293 -19004 26305 -18970
rect 26681 -19004 26693 -18970
rect 26293 -19016 26693 -19004
rect 25657 -19228 26057 -19216
rect 25657 -19262 25669 -19228
rect 26045 -19262 26057 -19228
rect 25657 -19274 26057 -19262
rect 26293 -19228 26693 -19216
rect 26293 -19262 26305 -19228
rect 26681 -19262 26693 -19228
rect 26293 -19274 26693 -19262
rect 25657 -19496 26057 -19484
rect 25657 -19530 25669 -19496
rect 26045 -19530 26057 -19496
rect 25657 -19542 26057 -19530
rect 26293 -19496 26693 -19484
rect 26293 -19530 26305 -19496
rect 26681 -19530 26693 -19496
rect 26293 -19542 26693 -19530
rect 25657 -20354 26057 -20342
rect 25657 -20388 25669 -20354
rect 26045 -20388 26057 -20354
rect 25657 -20400 26057 -20388
rect 26293 -20354 26693 -20342
rect 26293 -20388 26305 -20354
rect 26681 -20388 26693 -20354
rect 26293 -20400 26693 -20388
rect 27257 -18970 27657 -18958
rect 27257 -19004 27269 -18970
rect 27645 -19004 27657 -18970
rect 27257 -19016 27657 -19004
rect 27893 -18970 28293 -18958
rect 27893 -19004 27905 -18970
rect 28281 -19004 28293 -18970
rect 27893 -19016 28293 -19004
rect 27257 -19228 27657 -19216
rect 27257 -19262 27269 -19228
rect 27645 -19262 27657 -19228
rect 27257 -19274 27657 -19262
rect 27893 -19228 28293 -19216
rect 27893 -19262 27905 -19228
rect 28281 -19262 28293 -19228
rect 27893 -19274 28293 -19262
rect 27257 -19496 27657 -19484
rect 27257 -19530 27269 -19496
rect 27645 -19530 27657 -19496
rect 27257 -19542 27657 -19530
rect 27893 -19496 28293 -19484
rect 27893 -19530 27905 -19496
rect 28281 -19530 28293 -19496
rect 27893 -19542 28293 -19530
rect 27257 -20354 27657 -20342
rect 27257 -20388 27269 -20354
rect 27645 -20388 27657 -20354
rect 27257 -20400 27657 -20388
rect 27893 -20354 28293 -20342
rect 27893 -20388 27905 -20354
rect 28281 -20388 28293 -20354
rect 27893 -20400 28293 -20388
rect 28857 -18970 29257 -18958
rect 28857 -19004 28869 -18970
rect 29245 -19004 29257 -18970
rect 28857 -19016 29257 -19004
rect 29493 -18970 29893 -18958
rect 29493 -19004 29505 -18970
rect 29881 -19004 29893 -18970
rect 29493 -19016 29893 -19004
rect 28857 -19228 29257 -19216
rect 28857 -19262 28869 -19228
rect 29245 -19262 29257 -19228
rect 28857 -19274 29257 -19262
rect 29493 -19228 29893 -19216
rect 29493 -19262 29505 -19228
rect 29881 -19262 29893 -19228
rect 29493 -19274 29893 -19262
rect 28857 -19496 29257 -19484
rect 28857 -19530 28869 -19496
rect 29245 -19530 29257 -19496
rect 28857 -19542 29257 -19530
rect 29493 -19496 29893 -19484
rect 29493 -19530 29505 -19496
rect 29881 -19530 29893 -19496
rect 29493 -19542 29893 -19530
rect 28857 -20354 29257 -20342
rect 28857 -20388 28869 -20354
rect 29245 -20388 29257 -20354
rect 28857 -20400 29257 -20388
rect 29493 -20354 29893 -20342
rect 29493 -20388 29505 -20354
rect 29881 -20388 29893 -20354
rect 29493 -20400 29893 -20388
rect 30457 -18970 30857 -18958
rect 30457 -19004 30469 -18970
rect 30845 -19004 30857 -18970
rect 30457 -19016 30857 -19004
rect 31093 -18970 31493 -18958
rect 31093 -19004 31105 -18970
rect 31481 -19004 31493 -18970
rect 31093 -19016 31493 -19004
rect 30457 -19228 30857 -19216
rect 30457 -19262 30469 -19228
rect 30845 -19262 30857 -19228
rect 30457 -19274 30857 -19262
rect 31093 -19228 31493 -19216
rect 31093 -19262 31105 -19228
rect 31481 -19262 31493 -19228
rect 31093 -19274 31493 -19262
rect 30457 -19496 30857 -19484
rect 30457 -19530 30469 -19496
rect 30845 -19530 30857 -19496
rect 30457 -19542 30857 -19530
rect 31093 -19496 31493 -19484
rect 31093 -19530 31105 -19496
rect 31481 -19530 31493 -19496
rect 31093 -19542 31493 -19530
rect 30457 -20354 30857 -20342
rect 30457 -20388 30469 -20354
rect 30845 -20388 30857 -20354
rect 30457 -20400 30857 -20388
rect 31093 -20354 31493 -20342
rect 31093 -20388 31105 -20354
rect 31481 -20388 31493 -20354
rect 31093 -20400 31493 -20388
rect 32057 -18970 32457 -18958
rect 32057 -19004 32069 -18970
rect 32445 -19004 32457 -18970
rect 32057 -19016 32457 -19004
rect 32693 -18970 33093 -18958
rect 32693 -19004 32705 -18970
rect 33081 -19004 33093 -18970
rect 32693 -19016 33093 -19004
rect 32057 -19228 32457 -19216
rect 32057 -19262 32069 -19228
rect 32445 -19262 32457 -19228
rect 32057 -19274 32457 -19262
rect 32693 -19228 33093 -19216
rect 32693 -19262 32705 -19228
rect 33081 -19262 33093 -19228
rect 32693 -19274 33093 -19262
rect 32057 -19496 32457 -19484
rect 32057 -19530 32069 -19496
rect 32445 -19530 32457 -19496
rect 32057 -19542 32457 -19530
rect 32693 -19496 33093 -19484
rect 32693 -19530 32705 -19496
rect 33081 -19530 33093 -19496
rect 32693 -19542 33093 -19530
rect 32057 -20354 32457 -20342
rect 32057 -20388 32069 -20354
rect 32445 -20388 32457 -20354
rect 32057 -20400 32457 -20388
rect 32693 -20354 33093 -20342
rect 32693 -20388 32705 -20354
rect 33081 -20388 33093 -20354
rect 32693 -20400 33093 -20388
rect 33657 -18970 34057 -18958
rect 33657 -19004 33669 -18970
rect 34045 -19004 34057 -18970
rect 33657 -19016 34057 -19004
rect 34293 -18970 34693 -18958
rect 34293 -19004 34305 -18970
rect 34681 -19004 34693 -18970
rect 34293 -19016 34693 -19004
rect 33657 -19228 34057 -19216
rect 33657 -19262 33669 -19228
rect 34045 -19262 34057 -19228
rect 33657 -19274 34057 -19262
rect 34293 -19228 34693 -19216
rect 34293 -19262 34305 -19228
rect 34681 -19262 34693 -19228
rect 34293 -19274 34693 -19262
rect 33657 -19496 34057 -19484
rect 33657 -19530 33669 -19496
rect 34045 -19530 34057 -19496
rect 33657 -19542 34057 -19530
rect 34293 -19496 34693 -19484
rect 34293 -19530 34305 -19496
rect 34681 -19530 34693 -19496
rect 34293 -19542 34693 -19530
rect 33657 -20354 34057 -20342
rect 33657 -20388 33669 -20354
rect 34045 -20388 34057 -20354
rect 33657 -20400 34057 -20388
rect 34293 -20354 34693 -20342
rect 34293 -20388 34305 -20354
rect 34681 -20388 34693 -20354
rect 34293 -20400 34693 -20388
rect 35257 -18970 35657 -18958
rect 35257 -19004 35269 -18970
rect 35645 -19004 35657 -18970
rect 35257 -19016 35657 -19004
rect 35893 -18970 36293 -18958
rect 35893 -19004 35905 -18970
rect 36281 -19004 36293 -18970
rect 35893 -19016 36293 -19004
rect 35257 -19228 35657 -19216
rect 35257 -19262 35269 -19228
rect 35645 -19262 35657 -19228
rect 35257 -19274 35657 -19262
rect 35893 -19228 36293 -19216
rect 35893 -19262 35905 -19228
rect 36281 -19262 36293 -19228
rect 35893 -19274 36293 -19262
rect 35257 -19496 35657 -19484
rect 35257 -19530 35269 -19496
rect 35645 -19530 35657 -19496
rect 35257 -19542 35657 -19530
rect 35893 -19496 36293 -19484
rect 35893 -19530 35905 -19496
rect 36281 -19530 36293 -19496
rect 35893 -19542 36293 -19530
rect 35257 -20354 35657 -20342
rect 35257 -20388 35269 -20354
rect 35645 -20388 35657 -20354
rect 35257 -20400 35657 -20388
rect 35893 -20354 36293 -20342
rect 35893 -20388 35905 -20354
rect 36281 -20388 36293 -20354
rect 35893 -20400 36293 -20388
rect 36857 -18970 37257 -18958
rect 36857 -19004 36869 -18970
rect 37245 -19004 37257 -18970
rect 36857 -19016 37257 -19004
rect 37493 -18970 37893 -18958
rect 37493 -19004 37505 -18970
rect 37881 -19004 37893 -18970
rect 37493 -19016 37893 -19004
rect 36857 -19228 37257 -19216
rect 36857 -19262 36869 -19228
rect 37245 -19262 37257 -19228
rect 36857 -19274 37257 -19262
rect 37493 -19228 37893 -19216
rect 37493 -19262 37505 -19228
rect 37881 -19262 37893 -19228
rect 37493 -19274 37893 -19262
rect 36857 -19496 37257 -19484
rect 36857 -19530 36869 -19496
rect 37245 -19530 37257 -19496
rect 36857 -19542 37257 -19530
rect 37493 -19496 37893 -19484
rect 37493 -19530 37505 -19496
rect 37881 -19530 37893 -19496
rect 37493 -19542 37893 -19530
rect 36857 -20354 37257 -20342
rect 36857 -20388 36869 -20354
rect 37245 -20388 37257 -20354
rect 36857 -20400 37257 -20388
rect 37493 -20354 37893 -20342
rect 37493 -20388 37505 -20354
rect 37881 -20388 37893 -20354
rect 37493 -20400 37893 -20388
rect 57 -20770 457 -20758
rect 57 -20804 69 -20770
rect 445 -20804 457 -20770
rect 57 -20816 457 -20804
rect 693 -20770 1093 -20758
rect 693 -20804 705 -20770
rect 1081 -20804 1093 -20770
rect 693 -20816 1093 -20804
rect 57 -21028 457 -21016
rect 57 -21062 69 -21028
rect 445 -21062 457 -21028
rect 57 -21074 457 -21062
rect 693 -21028 1093 -21016
rect 693 -21062 705 -21028
rect 1081 -21062 1093 -21028
rect 693 -21074 1093 -21062
rect 57 -21296 457 -21284
rect 57 -21330 69 -21296
rect 445 -21330 457 -21296
rect 57 -21342 457 -21330
rect 693 -21296 1093 -21284
rect 693 -21330 705 -21296
rect 1081 -21330 1093 -21296
rect 693 -21342 1093 -21330
rect 57 -22154 457 -22142
rect 57 -22188 69 -22154
rect 445 -22188 457 -22154
rect 57 -22200 457 -22188
rect 693 -22154 1093 -22142
rect 693 -22188 705 -22154
rect 1081 -22188 1093 -22154
rect 693 -22200 1093 -22188
rect 1657 -20770 2057 -20758
rect 1657 -20804 1669 -20770
rect 2045 -20804 2057 -20770
rect 1657 -20816 2057 -20804
rect 2293 -20770 2693 -20758
rect 2293 -20804 2305 -20770
rect 2681 -20804 2693 -20770
rect 2293 -20816 2693 -20804
rect 1657 -21028 2057 -21016
rect 1657 -21062 1669 -21028
rect 2045 -21062 2057 -21028
rect 1657 -21074 2057 -21062
rect 2293 -21028 2693 -21016
rect 2293 -21062 2305 -21028
rect 2681 -21062 2693 -21028
rect 2293 -21074 2693 -21062
rect 1657 -21296 2057 -21284
rect 1657 -21330 1669 -21296
rect 2045 -21330 2057 -21296
rect 1657 -21342 2057 -21330
rect 2293 -21296 2693 -21284
rect 2293 -21330 2305 -21296
rect 2681 -21330 2693 -21296
rect 2293 -21342 2693 -21330
rect 1657 -22154 2057 -22142
rect 1657 -22188 1669 -22154
rect 2045 -22188 2057 -22154
rect 1657 -22200 2057 -22188
rect 2293 -22154 2693 -22142
rect 2293 -22188 2305 -22154
rect 2681 -22188 2693 -22154
rect 2293 -22200 2693 -22188
rect 3257 -20770 3657 -20758
rect 3257 -20804 3269 -20770
rect 3645 -20804 3657 -20770
rect 3257 -20816 3657 -20804
rect 3893 -20770 4293 -20758
rect 3893 -20804 3905 -20770
rect 4281 -20804 4293 -20770
rect 3893 -20816 4293 -20804
rect 3257 -21028 3657 -21016
rect 3257 -21062 3269 -21028
rect 3645 -21062 3657 -21028
rect 3257 -21074 3657 -21062
rect 3893 -21028 4293 -21016
rect 3893 -21062 3905 -21028
rect 4281 -21062 4293 -21028
rect 3893 -21074 4293 -21062
rect 3257 -21296 3657 -21284
rect 3257 -21330 3269 -21296
rect 3645 -21330 3657 -21296
rect 3257 -21342 3657 -21330
rect 3893 -21296 4293 -21284
rect 3893 -21330 3905 -21296
rect 4281 -21330 4293 -21296
rect 3893 -21342 4293 -21330
rect 3257 -22154 3657 -22142
rect 3257 -22188 3269 -22154
rect 3645 -22188 3657 -22154
rect 3257 -22200 3657 -22188
rect 3893 -22154 4293 -22142
rect 3893 -22188 3905 -22154
rect 4281 -22188 4293 -22154
rect 3893 -22200 4293 -22188
rect 4857 -20770 5257 -20758
rect 4857 -20804 4869 -20770
rect 5245 -20804 5257 -20770
rect 4857 -20816 5257 -20804
rect 5493 -20770 5893 -20758
rect 5493 -20804 5505 -20770
rect 5881 -20804 5893 -20770
rect 5493 -20816 5893 -20804
rect 4857 -21028 5257 -21016
rect 4857 -21062 4869 -21028
rect 5245 -21062 5257 -21028
rect 4857 -21074 5257 -21062
rect 5493 -21028 5893 -21016
rect 5493 -21062 5505 -21028
rect 5881 -21062 5893 -21028
rect 5493 -21074 5893 -21062
rect 4857 -21296 5257 -21284
rect 4857 -21330 4869 -21296
rect 5245 -21330 5257 -21296
rect 4857 -21342 5257 -21330
rect 5493 -21296 5893 -21284
rect 5493 -21330 5505 -21296
rect 5881 -21330 5893 -21296
rect 5493 -21342 5893 -21330
rect 4857 -22154 5257 -22142
rect 4857 -22188 4869 -22154
rect 5245 -22188 5257 -22154
rect 4857 -22200 5257 -22188
rect 5493 -22154 5893 -22142
rect 5493 -22188 5505 -22154
rect 5881 -22188 5893 -22154
rect 5493 -22200 5893 -22188
rect 6457 -20770 6857 -20758
rect 6457 -20804 6469 -20770
rect 6845 -20804 6857 -20770
rect 6457 -20816 6857 -20804
rect 7093 -20770 7493 -20758
rect 7093 -20804 7105 -20770
rect 7481 -20804 7493 -20770
rect 7093 -20816 7493 -20804
rect 6457 -21028 6857 -21016
rect 6457 -21062 6469 -21028
rect 6845 -21062 6857 -21028
rect 6457 -21074 6857 -21062
rect 7093 -21028 7493 -21016
rect 7093 -21062 7105 -21028
rect 7481 -21062 7493 -21028
rect 7093 -21074 7493 -21062
rect 6457 -21296 6857 -21284
rect 6457 -21330 6469 -21296
rect 6845 -21330 6857 -21296
rect 6457 -21342 6857 -21330
rect 7093 -21296 7493 -21284
rect 7093 -21330 7105 -21296
rect 7481 -21330 7493 -21296
rect 7093 -21342 7493 -21330
rect 6457 -22154 6857 -22142
rect 6457 -22188 6469 -22154
rect 6845 -22188 6857 -22154
rect 6457 -22200 6857 -22188
rect 7093 -22154 7493 -22142
rect 7093 -22188 7105 -22154
rect 7481 -22188 7493 -22154
rect 7093 -22200 7493 -22188
rect 8057 -20770 8457 -20758
rect 8057 -20804 8069 -20770
rect 8445 -20804 8457 -20770
rect 8057 -20816 8457 -20804
rect 8693 -20770 9093 -20758
rect 8693 -20804 8705 -20770
rect 9081 -20804 9093 -20770
rect 8693 -20816 9093 -20804
rect 8057 -21028 8457 -21016
rect 8057 -21062 8069 -21028
rect 8445 -21062 8457 -21028
rect 8057 -21074 8457 -21062
rect 8693 -21028 9093 -21016
rect 8693 -21062 8705 -21028
rect 9081 -21062 9093 -21028
rect 8693 -21074 9093 -21062
rect 8057 -21296 8457 -21284
rect 8057 -21330 8069 -21296
rect 8445 -21330 8457 -21296
rect 8057 -21342 8457 -21330
rect 8693 -21296 9093 -21284
rect 8693 -21330 8705 -21296
rect 9081 -21330 9093 -21296
rect 8693 -21342 9093 -21330
rect 8057 -22154 8457 -22142
rect 8057 -22188 8069 -22154
rect 8445 -22188 8457 -22154
rect 8057 -22200 8457 -22188
rect 8693 -22154 9093 -22142
rect 8693 -22188 8705 -22154
rect 9081 -22188 9093 -22154
rect 8693 -22200 9093 -22188
rect 9657 -20770 10057 -20758
rect 9657 -20804 9669 -20770
rect 10045 -20804 10057 -20770
rect 9657 -20816 10057 -20804
rect 10293 -20770 10693 -20758
rect 10293 -20804 10305 -20770
rect 10681 -20804 10693 -20770
rect 10293 -20816 10693 -20804
rect 9657 -21028 10057 -21016
rect 9657 -21062 9669 -21028
rect 10045 -21062 10057 -21028
rect 9657 -21074 10057 -21062
rect 10293 -21028 10693 -21016
rect 10293 -21062 10305 -21028
rect 10681 -21062 10693 -21028
rect 10293 -21074 10693 -21062
rect 9657 -21296 10057 -21284
rect 9657 -21330 9669 -21296
rect 10045 -21330 10057 -21296
rect 9657 -21342 10057 -21330
rect 10293 -21296 10693 -21284
rect 10293 -21330 10305 -21296
rect 10681 -21330 10693 -21296
rect 10293 -21342 10693 -21330
rect 9657 -22154 10057 -22142
rect 9657 -22188 9669 -22154
rect 10045 -22188 10057 -22154
rect 9657 -22200 10057 -22188
rect 10293 -22154 10693 -22142
rect 10293 -22188 10305 -22154
rect 10681 -22188 10693 -22154
rect 10293 -22200 10693 -22188
rect 11257 -20770 11657 -20758
rect 11257 -20804 11269 -20770
rect 11645 -20804 11657 -20770
rect 11257 -20816 11657 -20804
rect 11893 -20770 12293 -20758
rect 11893 -20804 11905 -20770
rect 12281 -20804 12293 -20770
rect 11893 -20816 12293 -20804
rect 11257 -21028 11657 -21016
rect 11257 -21062 11269 -21028
rect 11645 -21062 11657 -21028
rect 11257 -21074 11657 -21062
rect 11893 -21028 12293 -21016
rect 11893 -21062 11905 -21028
rect 12281 -21062 12293 -21028
rect 11893 -21074 12293 -21062
rect 11257 -21296 11657 -21284
rect 11257 -21330 11269 -21296
rect 11645 -21330 11657 -21296
rect 11257 -21342 11657 -21330
rect 11893 -21296 12293 -21284
rect 11893 -21330 11905 -21296
rect 12281 -21330 12293 -21296
rect 11893 -21342 12293 -21330
rect 11257 -22154 11657 -22142
rect 11257 -22188 11269 -22154
rect 11645 -22188 11657 -22154
rect 11257 -22200 11657 -22188
rect 11893 -22154 12293 -22142
rect 11893 -22188 11905 -22154
rect 12281 -22188 12293 -22154
rect 11893 -22200 12293 -22188
rect 12857 -20770 13257 -20758
rect 12857 -20804 12869 -20770
rect 13245 -20804 13257 -20770
rect 12857 -20816 13257 -20804
rect 13493 -20770 13893 -20758
rect 13493 -20804 13505 -20770
rect 13881 -20804 13893 -20770
rect 13493 -20816 13893 -20804
rect 12857 -21028 13257 -21016
rect 12857 -21062 12869 -21028
rect 13245 -21062 13257 -21028
rect 12857 -21074 13257 -21062
rect 13493 -21028 13893 -21016
rect 13493 -21062 13505 -21028
rect 13881 -21062 13893 -21028
rect 13493 -21074 13893 -21062
rect 12857 -21296 13257 -21284
rect 12857 -21330 12869 -21296
rect 13245 -21330 13257 -21296
rect 12857 -21342 13257 -21330
rect 13493 -21296 13893 -21284
rect 13493 -21330 13505 -21296
rect 13881 -21330 13893 -21296
rect 13493 -21342 13893 -21330
rect 12857 -22154 13257 -22142
rect 12857 -22188 12869 -22154
rect 13245 -22188 13257 -22154
rect 12857 -22200 13257 -22188
rect 13493 -22154 13893 -22142
rect 13493 -22188 13505 -22154
rect 13881 -22188 13893 -22154
rect 13493 -22200 13893 -22188
rect 14457 -20770 14857 -20758
rect 14457 -20804 14469 -20770
rect 14845 -20804 14857 -20770
rect 14457 -20816 14857 -20804
rect 15093 -20770 15493 -20758
rect 15093 -20804 15105 -20770
rect 15481 -20804 15493 -20770
rect 15093 -20816 15493 -20804
rect 14457 -21028 14857 -21016
rect 14457 -21062 14469 -21028
rect 14845 -21062 14857 -21028
rect 14457 -21074 14857 -21062
rect 15093 -21028 15493 -21016
rect 15093 -21062 15105 -21028
rect 15481 -21062 15493 -21028
rect 15093 -21074 15493 -21062
rect 14457 -21296 14857 -21284
rect 14457 -21330 14469 -21296
rect 14845 -21330 14857 -21296
rect 14457 -21342 14857 -21330
rect 15093 -21296 15493 -21284
rect 15093 -21330 15105 -21296
rect 15481 -21330 15493 -21296
rect 15093 -21342 15493 -21330
rect 14457 -22154 14857 -22142
rect 14457 -22188 14469 -22154
rect 14845 -22188 14857 -22154
rect 14457 -22200 14857 -22188
rect 15093 -22154 15493 -22142
rect 15093 -22188 15105 -22154
rect 15481 -22188 15493 -22154
rect 15093 -22200 15493 -22188
rect 16057 -20770 16457 -20758
rect 16057 -20804 16069 -20770
rect 16445 -20804 16457 -20770
rect 16057 -20816 16457 -20804
rect 16693 -20770 17093 -20758
rect 16693 -20804 16705 -20770
rect 17081 -20804 17093 -20770
rect 16693 -20816 17093 -20804
rect 16057 -21028 16457 -21016
rect 16057 -21062 16069 -21028
rect 16445 -21062 16457 -21028
rect 16057 -21074 16457 -21062
rect 16693 -21028 17093 -21016
rect 16693 -21062 16705 -21028
rect 17081 -21062 17093 -21028
rect 16693 -21074 17093 -21062
rect 16057 -21296 16457 -21284
rect 16057 -21330 16069 -21296
rect 16445 -21330 16457 -21296
rect 16057 -21342 16457 -21330
rect 16693 -21296 17093 -21284
rect 16693 -21330 16705 -21296
rect 17081 -21330 17093 -21296
rect 16693 -21342 17093 -21330
rect 16057 -22154 16457 -22142
rect 16057 -22188 16069 -22154
rect 16445 -22188 16457 -22154
rect 16057 -22200 16457 -22188
rect 16693 -22154 17093 -22142
rect 16693 -22188 16705 -22154
rect 17081 -22188 17093 -22154
rect 16693 -22200 17093 -22188
rect 17657 -20770 18057 -20758
rect 17657 -20804 17669 -20770
rect 18045 -20804 18057 -20770
rect 17657 -20816 18057 -20804
rect 18293 -20770 18693 -20758
rect 18293 -20804 18305 -20770
rect 18681 -20804 18693 -20770
rect 18293 -20816 18693 -20804
rect 17657 -21028 18057 -21016
rect 17657 -21062 17669 -21028
rect 18045 -21062 18057 -21028
rect 17657 -21074 18057 -21062
rect 18293 -21028 18693 -21016
rect 18293 -21062 18305 -21028
rect 18681 -21062 18693 -21028
rect 18293 -21074 18693 -21062
rect 17657 -21296 18057 -21284
rect 17657 -21330 17669 -21296
rect 18045 -21330 18057 -21296
rect 17657 -21342 18057 -21330
rect 18293 -21296 18693 -21284
rect 18293 -21330 18305 -21296
rect 18681 -21330 18693 -21296
rect 18293 -21342 18693 -21330
rect 17657 -22154 18057 -22142
rect 17657 -22188 17669 -22154
rect 18045 -22188 18057 -22154
rect 17657 -22200 18057 -22188
rect 18293 -22154 18693 -22142
rect 18293 -22188 18305 -22154
rect 18681 -22188 18693 -22154
rect 18293 -22200 18693 -22188
rect 19257 -20770 19657 -20758
rect 19257 -20804 19269 -20770
rect 19645 -20804 19657 -20770
rect 19257 -20816 19657 -20804
rect 19893 -20770 20293 -20758
rect 19893 -20804 19905 -20770
rect 20281 -20804 20293 -20770
rect 19893 -20816 20293 -20804
rect 19257 -21028 19657 -21016
rect 19257 -21062 19269 -21028
rect 19645 -21062 19657 -21028
rect 19257 -21074 19657 -21062
rect 19893 -21028 20293 -21016
rect 19893 -21062 19905 -21028
rect 20281 -21062 20293 -21028
rect 19893 -21074 20293 -21062
rect 19257 -21296 19657 -21284
rect 19257 -21330 19269 -21296
rect 19645 -21330 19657 -21296
rect 19257 -21342 19657 -21330
rect 19893 -21296 20293 -21284
rect 19893 -21330 19905 -21296
rect 20281 -21330 20293 -21296
rect 19893 -21342 20293 -21330
rect 19257 -22154 19657 -22142
rect 19257 -22188 19269 -22154
rect 19645 -22188 19657 -22154
rect 19257 -22200 19657 -22188
rect 19893 -22154 20293 -22142
rect 19893 -22188 19905 -22154
rect 20281 -22188 20293 -22154
rect 19893 -22200 20293 -22188
rect 20857 -20770 21257 -20758
rect 20857 -20804 20869 -20770
rect 21245 -20804 21257 -20770
rect 20857 -20816 21257 -20804
rect 21493 -20770 21893 -20758
rect 21493 -20804 21505 -20770
rect 21881 -20804 21893 -20770
rect 21493 -20816 21893 -20804
rect 20857 -21028 21257 -21016
rect 20857 -21062 20869 -21028
rect 21245 -21062 21257 -21028
rect 20857 -21074 21257 -21062
rect 21493 -21028 21893 -21016
rect 21493 -21062 21505 -21028
rect 21881 -21062 21893 -21028
rect 21493 -21074 21893 -21062
rect 20857 -21296 21257 -21284
rect 20857 -21330 20869 -21296
rect 21245 -21330 21257 -21296
rect 20857 -21342 21257 -21330
rect 21493 -21296 21893 -21284
rect 21493 -21330 21505 -21296
rect 21881 -21330 21893 -21296
rect 21493 -21342 21893 -21330
rect 20857 -22154 21257 -22142
rect 20857 -22188 20869 -22154
rect 21245 -22188 21257 -22154
rect 20857 -22200 21257 -22188
rect 21493 -22154 21893 -22142
rect 21493 -22188 21505 -22154
rect 21881 -22188 21893 -22154
rect 21493 -22200 21893 -22188
rect 22457 -20770 22857 -20758
rect 22457 -20804 22469 -20770
rect 22845 -20804 22857 -20770
rect 22457 -20816 22857 -20804
rect 23093 -20770 23493 -20758
rect 23093 -20804 23105 -20770
rect 23481 -20804 23493 -20770
rect 23093 -20816 23493 -20804
rect 22457 -21028 22857 -21016
rect 22457 -21062 22469 -21028
rect 22845 -21062 22857 -21028
rect 22457 -21074 22857 -21062
rect 23093 -21028 23493 -21016
rect 23093 -21062 23105 -21028
rect 23481 -21062 23493 -21028
rect 23093 -21074 23493 -21062
rect 22457 -21296 22857 -21284
rect 22457 -21330 22469 -21296
rect 22845 -21330 22857 -21296
rect 22457 -21342 22857 -21330
rect 23093 -21296 23493 -21284
rect 23093 -21330 23105 -21296
rect 23481 -21330 23493 -21296
rect 23093 -21342 23493 -21330
rect 22457 -22154 22857 -22142
rect 22457 -22188 22469 -22154
rect 22845 -22188 22857 -22154
rect 22457 -22200 22857 -22188
rect 23093 -22154 23493 -22142
rect 23093 -22188 23105 -22154
rect 23481 -22188 23493 -22154
rect 23093 -22200 23493 -22188
rect 24057 -20770 24457 -20758
rect 24057 -20804 24069 -20770
rect 24445 -20804 24457 -20770
rect 24057 -20816 24457 -20804
rect 24693 -20770 25093 -20758
rect 24693 -20804 24705 -20770
rect 25081 -20804 25093 -20770
rect 24693 -20816 25093 -20804
rect 24057 -21028 24457 -21016
rect 24057 -21062 24069 -21028
rect 24445 -21062 24457 -21028
rect 24057 -21074 24457 -21062
rect 24693 -21028 25093 -21016
rect 24693 -21062 24705 -21028
rect 25081 -21062 25093 -21028
rect 24693 -21074 25093 -21062
rect 24057 -21296 24457 -21284
rect 24057 -21330 24069 -21296
rect 24445 -21330 24457 -21296
rect 24057 -21342 24457 -21330
rect 24693 -21296 25093 -21284
rect 24693 -21330 24705 -21296
rect 25081 -21330 25093 -21296
rect 24693 -21342 25093 -21330
rect 24057 -22154 24457 -22142
rect 24057 -22188 24069 -22154
rect 24445 -22188 24457 -22154
rect 24057 -22200 24457 -22188
rect 24693 -22154 25093 -22142
rect 24693 -22188 24705 -22154
rect 25081 -22188 25093 -22154
rect 24693 -22200 25093 -22188
rect 25657 -20770 26057 -20758
rect 25657 -20804 25669 -20770
rect 26045 -20804 26057 -20770
rect 25657 -20816 26057 -20804
rect 26293 -20770 26693 -20758
rect 26293 -20804 26305 -20770
rect 26681 -20804 26693 -20770
rect 26293 -20816 26693 -20804
rect 25657 -21028 26057 -21016
rect 25657 -21062 25669 -21028
rect 26045 -21062 26057 -21028
rect 25657 -21074 26057 -21062
rect 26293 -21028 26693 -21016
rect 26293 -21062 26305 -21028
rect 26681 -21062 26693 -21028
rect 26293 -21074 26693 -21062
rect 25657 -21296 26057 -21284
rect 25657 -21330 25669 -21296
rect 26045 -21330 26057 -21296
rect 25657 -21342 26057 -21330
rect 26293 -21296 26693 -21284
rect 26293 -21330 26305 -21296
rect 26681 -21330 26693 -21296
rect 26293 -21342 26693 -21330
rect 25657 -22154 26057 -22142
rect 25657 -22188 25669 -22154
rect 26045 -22188 26057 -22154
rect 25657 -22200 26057 -22188
rect 26293 -22154 26693 -22142
rect 26293 -22188 26305 -22154
rect 26681 -22188 26693 -22154
rect 26293 -22200 26693 -22188
rect 27257 -20770 27657 -20758
rect 27257 -20804 27269 -20770
rect 27645 -20804 27657 -20770
rect 27257 -20816 27657 -20804
rect 27893 -20770 28293 -20758
rect 27893 -20804 27905 -20770
rect 28281 -20804 28293 -20770
rect 27893 -20816 28293 -20804
rect 27257 -21028 27657 -21016
rect 27257 -21062 27269 -21028
rect 27645 -21062 27657 -21028
rect 27257 -21074 27657 -21062
rect 27893 -21028 28293 -21016
rect 27893 -21062 27905 -21028
rect 28281 -21062 28293 -21028
rect 27893 -21074 28293 -21062
rect 27257 -21296 27657 -21284
rect 27257 -21330 27269 -21296
rect 27645 -21330 27657 -21296
rect 27257 -21342 27657 -21330
rect 27893 -21296 28293 -21284
rect 27893 -21330 27905 -21296
rect 28281 -21330 28293 -21296
rect 27893 -21342 28293 -21330
rect 27257 -22154 27657 -22142
rect 27257 -22188 27269 -22154
rect 27645 -22188 27657 -22154
rect 27257 -22200 27657 -22188
rect 27893 -22154 28293 -22142
rect 27893 -22188 27905 -22154
rect 28281 -22188 28293 -22154
rect 27893 -22200 28293 -22188
rect 28857 -20770 29257 -20758
rect 28857 -20804 28869 -20770
rect 29245 -20804 29257 -20770
rect 28857 -20816 29257 -20804
rect 29493 -20770 29893 -20758
rect 29493 -20804 29505 -20770
rect 29881 -20804 29893 -20770
rect 29493 -20816 29893 -20804
rect 28857 -21028 29257 -21016
rect 28857 -21062 28869 -21028
rect 29245 -21062 29257 -21028
rect 28857 -21074 29257 -21062
rect 29493 -21028 29893 -21016
rect 29493 -21062 29505 -21028
rect 29881 -21062 29893 -21028
rect 29493 -21074 29893 -21062
rect 28857 -21296 29257 -21284
rect 28857 -21330 28869 -21296
rect 29245 -21330 29257 -21296
rect 28857 -21342 29257 -21330
rect 29493 -21296 29893 -21284
rect 29493 -21330 29505 -21296
rect 29881 -21330 29893 -21296
rect 29493 -21342 29893 -21330
rect 28857 -22154 29257 -22142
rect 28857 -22188 28869 -22154
rect 29245 -22188 29257 -22154
rect 28857 -22200 29257 -22188
rect 29493 -22154 29893 -22142
rect 29493 -22188 29505 -22154
rect 29881 -22188 29893 -22154
rect 29493 -22200 29893 -22188
rect 30457 -20770 30857 -20758
rect 30457 -20804 30469 -20770
rect 30845 -20804 30857 -20770
rect 30457 -20816 30857 -20804
rect 31093 -20770 31493 -20758
rect 31093 -20804 31105 -20770
rect 31481 -20804 31493 -20770
rect 31093 -20816 31493 -20804
rect 30457 -21028 30857 -21016
rect 30457 -21062 30469 -21028
rect 30845 -21062 30857 -21028
rect 30457 -21074 30857 -21062
rect 31093 -21028 31493 -21016
rect 31093 -21062 31105 -21028
rect 31481 -21062 31493 -21028
rect 31093 -21074 31493 -21062
rect 30457 -21296 30857 -21284
rect 30457 -21330 30469 -21296
rect 30845 -21330 30857 -21296
rect 30457 -21342 30857 -21330
rect 31093 -21296 31493 -21284
rect 31093 -21330 31105 -21296
rect 31481 -21330 31493 -21296
rect 31093 -21342 31493 -21330
rect 30457 -22154 30857 -22142
rect 30457 -22188 30469 -22154
rect 30845 -22188 30857 -22154
rect 30457 -22200 30857 -22188
rect 31093 -22154 31493 -22142
rect 31093 -22188 31105 -22154
rect 31481 -22188 31493 -22154
rect 31093 -22200 31493 -22188
rect 32057 -20770 32457 -20758
rect 32057 -20804 32069 -20770
rect 32445 -20804 32457 -20770
rect 32057 -20816 32457 -20804
rect 32693 -20770 33093 -20758
rect 32693 -20804 32705 -20770
rect 33081 -20804 33093 -20770
rect 32693 -20816 33093 -20804
rect 32057 -21028 32457 -21016
rect 32057 -21062 32069 -21028
rect 32445 -21062 32457 -21028
rect 32057 -21074 32457 -21062
rect 32693 -21028 33093 -21016
rect 32693 -21062 32705 -21028
rect 33081 -21062 33093 -21028
rect 32693 -21074 33093 -21062
rect 32057 -21296 32457 -21284
rect 32057 -21330 32069 -21296
rect 32445 -21330 32457 -21296
rect 32057 -21342 32457 -21330
rect 32693 -21296 33093 -21284
rect 32693 -21330 32705 -21296
rect 33081 -21330 33093 -21296
rect 32693 -21342 33093 -21330
rect 32057 -22154 32457 -22142
rect 32057 -22188 32069 -22154
rect 32445 -22188 32457 -22154
rect 32057 -22200 32457 -22188
rect 32693 -22154 33093 -22142
rect 32693 -22188 32705 -22154
rect 33081 -22188 33093 -22154
rect 32693 -22200 33093 -22188
rect 33657 -20770 34057 -20758
rect 33657 -20804 33669 -20770
rect 34045 -20804 34057 -20770
rect 33657 -20816 34057 -20804
rect 34293 -20770 34693 -20758
rect 34293 -20804 34305 -20770
rect 34681 -20804 34693 -20770
rect 34293 -20816 34693 -20804
rect 33657 -21028 34057 -21016
rect 33657 -21062 33669 -21028
rect 34045 -21062 34057 -21028
rect 33657 -21074 34057 -21062
rect 34293 -21028 34693 -21016
rect 34293 -21062 34305 -21028
rect 34681 -21062 34693 -21028
rect 34293 -21074 34693 -21062
rect 33657 -21296 34057 -21284
rect 33657 -21330 33669 -21296
rect 34045 -21330 34057 -21296
rect 33657 -21342 34057 -21330
rect 34293 -21296 34693 -21284
rect 34293 -21330 34305 -21296
rect 34681 -21330 34693 -21296
rect 34293 -21342 34693 -21330
rect 33657 -22154 34057 -22142
rect 33657 -22188 33669 -22154
rect 34045 -22188 34057 -22154
rect 33657 -22200 34057 -22188
rect 34293 -22154 34693 -22142
rect 34293 -22188 34305 -22154
rect 34681 -22188 34693 -22154
rect 34293 -22200 34693 -22188
rect 35257 -20770 35657 -20758
rect 35257 -20804 35269 -20770
rect 35645 -20804 35657 -20770
rect 35257 -20816 35657 -20804
rect 35893 -20770 36293 -20758
rect 35893 -20804 35905 -20770
rect 36281 -20804 36293 -20770
rect 35893 -20816 36293 -20804
rect 35257 -21028 35657 -21016
rect 35257 -21062 35269 -21028
rect 35645 -21062 35657 -21028
rect 35257 -21074 35657 -21062
rect 35893 -21028 36293 -21016
rect 35893 -21062 35905 -21028
rect 36281 -21062 36293 -21028
rect 35893 -21074 36293 -21062
rect 35257 -21296 35657 -21284
rect 35257 -21330 35269 -21296
rect 35645 -21330 35657 -21296
rect 35257 -21342 35657 -21330
rect 35893 -21296 36293 -21284
rect 35893 -21330 35905 -21296
rect 36281 -21330 36293 -21296
rect 35893 -21342 36293 -21330
rect 35257 -22154 35657 -22142
rect 35257 -22188 35269 -22154
rect 35645 -22188 35657 -22154
rect 35257 -22200 35657 -22188
rect 35893 -22154 36293 -22142
rect 35893 -22188 35905 -22154
rect 36281 -22188 36293 -22154
rect 35893 -22200 36293 -22188
rect 36857 -20770 37257 -20758
rect 36857 -20804 36869 -20770
rect 37245 -20804 37257 -20770
rect 36857 -20816 37257 -20804
rect 37493 -20770 37893 -20758
rect 37493 -20804 37505 -20770
rect 37881 -20804 37893 -20770
rect 37493 -20816 37893 -20804
rect 36857 -21028 37257 -21016
rect 36857 -21062 36869 -21028
rect 37245 -21062 37257 -21028
rect 36857 -21074 37257 -21062
rect 37493 -21028 37893 -21016
rect 37493 -21062 37505 -21028
rect 37881 -21062 37893 -21028
rect 37493 -21074 37893 -21062
rect 36857 -21296 37257 -21284
rect 36857 -21330 36869 -21296
rect 37245 -21330 37257 -21296
rect 36857 -21342 37257 -21330
rect 37493 -21296 37893 -21284
rect 37493 -21330 37505 -21296
rect 37881 -21330 37893 -21296
rect 37493 -21342 37893 -21330
rect 36857 -22154 37257 -22142
rect 36857 -22188 36869 -22154
rect 37245 -22188 37257 -22154
rect 36857 -22200 37257 -22188
rect 37493 -22154 37893 -22142
rect 37493 -22188 37505 -22154
rect 37881 -22188 37893 -22154
rect 37493 -22200 37893 -22188
rect 28340 -22684 28398 -22672
rect 28340 -23460 28352 -22684
rect 28386 -23460 28398 -22684
rect 28340 -23472 28398 -23460
rect 28498 -22684 28556 -22672
rect 28498 -23460 28510 -22684
rect 28544 -23460 28556 -22684
rect 28498 -23472 28556 -23460
rect 28656 -22684 28714 -22672
rect 28656 -23460 28668 -22684
rect 28702 -23460 28714 -22684
rect 28656 -23472 28714 -23460
rect 28814 -22684 28872 -22672
rect 28814 -23460 28826 -22684
rect 28860 -23460 28872 -22684
rect 28814 -23472 28872 -23460
rect 28972 -22684 29030 -22672
rect 28972 -23460 28984 -22684
rect 29018 -23460 29030 -22684
rect 28972 -23472 29030 -23460
rect 32620 -22635 32678 -22623
rect 32620 -23011 32632 -22635
rect 32666 -23011 32678 -22635
rect 32620 -23023 32678 -23011
rect 32778 -22635 32836 -22623
rect 32778 -23011 32790 -22635
rect 32824 -23011 32836 -22635
rect 32778 -23023 32836 -23011
rect 32936 -22635 32994 -22623
rect 32936 -23011 32948 -22635
rect 32982 -23011 32994 -22635
rect 32936 -23023 32994 -23011
rect 33094 -22635 33152 -22623
rect 33094 -23011 33106 -22635
rect 33140 -23011 33152 -22635
rect 33094 -23023 33152 -23011
rect 33252 -22635 33310 -22623
rect 33252 -23011 33264 -22635
rect 33298 -23011 33310 -22635
rect 33252 -23023 33310 -23011
rect 33990 -22655 34048 -22643
rect 33990 -23031 34002 -22655
rect 34036 -23031 34048 -22655
rect 33990 -23043 34048 -23031
rect 34148 -22655 34206 -22643
rect 34148 -23031 34160 -22655
rect 34194 -23031 34206 -22655
rect 34148 -23043 34206 -23031
rect 34306 -22655 34364 -22643
rect 34306 -23031 34318 -22655
rect 34352 -23031 34364 -22655
rect 34306 -23043 34364 -23031
rect 267 -24306 1867 -24294
rect 267 -24340 279 -24306
rect 1855 -24340 1867 -24306
rect 267 -24352 1867 -24340
rect 267 -24664 1867 -24652
rect 267 -24698 279 -24664
rect 1855 -24698 1867 -24664
rect 267 -24710 1867 -24698
rect 2467 -24306 4067 -24294
rect 2467 -24340 2479 -24306
rect 4055 -24340 4067 -24306
rect 2467 -24352 4067 -24340
rect 2467 -24664 4067 -24652
rect 2467 -24698 2479 -24664
rect 4055 -24698 4067 -24664
rect 2467 -24710 4067 -24698
rect 4667 -24306 6267 -24294
rect 4667 -24340 4679 -24306
rect 6255 -24340 6267 -24306
rect 4667 -24352 6267 -24340
rect 4667 -24664 6267 -24652
rect 4667 -24698 4679 -24664
rect 6255 -24698 6267 -24664
rect 4667 -24710 6267 -24698
rect 6867 -24306 8467 -24294
rect 6867 -24340 6879 -24306
rect 8455 -24340 8467 -24306
rect 6867 -24352 8467 -24340
rect 6867 -24664 8467 -24652
rect 6867 -24698 6879 -24664
rect 8455 -24698 8467 -24664
rect 6867 -24710 8467 -24698
rect 9067 -24306 10667 -24294
rect 9067 -24340 9079 -24306
rect 10655 -24340 10667 -24306
rect 9067 -24352 10667 -24340
rect 9067 -24664 10667 -24652
rect 9067 -24698 9079 -24664
rect 10655 -24698 10667 -24664
rect 9067 -24710 10667 -24698
rect 11267 -24306 12867 -24294
rect 11267 -24340 11279 -24306
rect 12855 -24340 12867 -24306
rect 11267 -24352 12867 -24340
rect 11267 -24664 12867 -24652
rect 11267 -24698 11279 -24664
rect 12855 -24698 12867 -24664
rect 11267 -24710 12867 -24698
rect 13467 -24306 15067 -24294
rect 13467 -24340 13479 -24306
rect 15055 -24340 15067 -24306
rect 13467 -24352 15067 -24340
rect 13467 -24664 15067 -24652
rect 13467 -24698 13479 -24664
rect 15055 -24698 15067 -24664
rect 13467 -24710 15067 -24698
rect 15667 -24306 17267 -24294
rect 15667 -24340 15679 -24306
rect 17255 -24340 17267 -24306
rect 15667 -24352 17267 -24340
rect 15667 -24664 17267 -24652
rect 15667 -24698 15679 -24664
rect 17255 -24698 17267 -24664
rect 15667 -24710 17267 -24698
rect 17867 -24306 19467 -24294
rect 17867 -24340 17879 -24306
rect 19455 -24340 19467 -24306
rect 17867 -24352 19467 -24340
rect 17867 -24664 19467 -24652
rect 17867 -24698 17879 -24664
rect 19455 -24698 19467 -24664
rect 17867 -24710 19467 -24698
rect 20067 -24306 21667 -24294
rect 20067 -24340 20079 -24306
rect 21655 -24340 21667 -24306
rect 20067 -24352 21667 -24340
rect 20067 -24664 21667 -24652
rect 20067 -24698 20079 -24664
rect 21655 -24698 21667 -24664
rect 20067 -24710 21667 -24698
rect 33158 -23777 33216 -23765
rect 33158 -24153 33170 -23777
rect 33204 -24153 33216 -23777
rect 33158 -24165 33216 -24153
rect 33316 -23777 33374 -23765
rect 33316 -24153 33328 -23777
rect 33362 -24153 33374 -23777
rect 33316 -24165 33374 -24153
rect 33474 -23777 33532 -23765
rect 33474 -24153 33486 -23777
rect 33520 -24153 33532 -23777
rect 33474 -24165 33532 -24153
rect 33632 -23777 33690 -23765
rect 33632 -24153 33644 -23777
rect 33678 -24153 33690 -23777
rect 33632 -24165 33690 -24153
rect 33790 -23777 33848 -23765
rect 33790 -24153 33802 -23777
rect 33836 -24153 33848 -23777
rect 33790 -24165 33848 -24153
rect 33948 -23777 34006 -23765
rect 33948 -24153 33960 -23777
rect 33994 -24153 34006 -23777
rect 33948 -24165 34006 -24153
rect 34106 -23777 34164 -23765
rect 34106 -24153 34118 -23777
rect 34152 -24153 34164 -23777
rect 34106 -24165 34164 -24153
rect 34530 -23775 34588 -23763
rect 34530 -24151 34542 -23775
rect 34576 -24151 34588 -23775
rect 34530 -24163 34588 -24151
rect 34688 -23775 34746 -23763
rect 34688 -24151 34700 -23775
rect 34734 -24151 34746 -23775
rect 34688 -24163 34746 -24151
rect 34846 -23775 34904 -23763
rect 34846 -24151 34858 -23775
rect 34892 -24151 34904 -23775
rect 34846 -24163 34904 -24151
rect 35004 -23775 35062 -23763
rect 35004 -24151 35016 -23775
rect 35050 -24151 35062 -23775
rect 35004 -24163 35062 -24151
rect 35162 -23775 35220 -23763
rect 35162 -24151 35174 -23775
rect 35208 -24151 35220 -23775
rect 35162 -24163 35220 -24151
rect 35320 -23775 35378 -23763
rect 35320 -24151 35332 -23775
rect 35366 -24151 35378 -23775
rect 35320 -24163 35378 -24151
rect 35478 -23775 35536 -23763
rect 35478 -24151 35490 -23775
rect 35524 -24151 35536 -23775
rect 35478 -24163 35536 -24151
rect 35636 -23775 35694 -23763
rect 35636 -24151 35648 -23775
rect 35682 -24151 35694 -23775
rect 35636 -24163 35694 -24151
rect 35794 -23775 35852 -23763
rect 35794 -24151 35806 -23775
rect 35840 -24151 35852 -23775
rect 35794 -24163 35852 -24151
rect 35952 -23775 36010 -23763
rect 35952 -24151 35964 -23775
rect 35998 -24151 36010 -23775
rect 35952 -24163 36010 -24151
rect 36110 -23775 36168 -23763
rect 36110 -24151 36122 -23775
rect 36156 -24151 36168 -23775
rect 36110 -24163 36168 -24151
rect 36268 -23775 36326 -23763
rect 36268 -24151 36280 -23775
rect 36314 -24151 36326 -23775
rect 36268 -24163 36326 -24151
rect 36426 -23775 36484 -23763
rect 36426 -24151 36438 -23775
rect 36472 -24151 36484 -23775
rect 36426 -24163 36484 -24151
rect 36584 -23775 36642 -23763
rect 36584 -24151 36596 -23775
rect 36630 -24151 36642 -23775
rect 36584 -24163 36642 -24151
rect 36742 -23775 36800 -23763
rect 36742 -24151 36754 -23775
rect 36788 -24151 36800 -23775
rect 36742 -24163 36800 -24151
rect 36900 -23775 36958 -23763
rect 36900 -24151 36912 -23775
rect 36946 -24151 36958 -23775
rect 36900 -24163 36958 -24151
rect 37058 -23775 37116 -23763
rect 37058 -24151 37070 -23775
rect 37104 -24151 37116 -23775
rect 37058 -24163 37116 -24151
rect 267 -25106 1867 -25094
rect 267 -25140 279 -25106
rect 1855 -25140 1867 -25106
rect 267 -25152 1867 -25140
rect 267 -25464 1867 -25452
rect 267 -25498 279 -25464
rect 1855 -25498 1867 -25464
rect 267 -25510 1867 -25498
rect 2467 -25106 4067 -25094
rect 2467 -25140 2479 -25106
rect 4055 -25140 4067 -25106
rect 2467 -25152 4067 -25140
rect 2467 -25464 4067 -25452
rect 2467 -25498 2479 -25464
rect 4055 -25498 4067 -25464
rect 2467 -25510 4067 -25498
rect 4667 -25106 6267 -25094
rect 4667 -25140 4679 -25106
rect 6255 -25140 6267 -25106
rect 4667 -25152 6267 -25140
rect 4667 -25464 6267 -25452
rect 4667 -25498 4679 -25464
rect 6255 -25498 6267 -25464
rect 4667 -25510 6267 -25498
rect 6867 -25106 8467 -25094
rect 6867 -25140 6879 -25106
rect 8455 -25140 8467 -25106
rect 6867 -25152 8467 -25140
rect 6867 -25464 8467 -25452
rect 6867 -25498 6879 -25464
rect 8455 -25498 8467 -25464
rect 6867 -25510 8467 -25498
rect 9067 -25106 10667 -25094
rect 9067 -25140 9079 -25106
rect 10655 -25140 10667 -25106
rect 9067 -25152 10667 -25140
rect 9067 -25464 10667 -25452
rect 9067 -25498 9079 -25464
rect 10655 -25498 10667 -25464
rect 9067 -25510 10667 -25498
rect 11267 -25106 12867 -25094
rect 11267 -25140 11279 -25106
rect 12855 -25140 12867 -25106
rect 11267 -25152 12867 -25140
rect 11267 -25464 12867 -25452
rect 11267 -25498 11279 -25464
rect 12855 -25498 12867 -25464
rect 11267 -25510 12867 -25498
rect 13467 -25106 15067 -25094
rect 13467 -25140 13479 -25106
rect 15055 -25140 15067 -25106
rect 13467 -25152 15067 -25140
rect 13467 -25464 15067 -25452
rect 13467 -25498 13479 -25464
rect 15055 -25498 15067 -25464
rect 13467 -25510 15067 -25498
rect 15667 -25106 17267 -25094
rect 15667 -25140 15679 -25106
rect 17255 -25140 17267 -25106
rect 15667 -25152 17267 -25140
rect 15667 -25464 17267 -25452
rect 15667 -25498 15679 -25464
rect 17255 -25498 17267 -25464
rect 15667 -25510 17267 -25498
rect 17867 -25106 19467 -25094
rect 17867 -25140 17879 -25106
rect 19455 -25140 19467 -25106
rect 17867 -25152 19467 -25140
rect 17867 -25464 19467 -25452
rect 17867 -25498 17879 -25464
rect 19455 -25498 19467 -25464
rect 17867 -25510 19467 -25498
rect 20067 -25106 21667 -25094
rect 20067 -25140 20079 -25106
rect 21655 -25140 21667 -25106
rect 20067 -25152 21667 -25140
rect 20067 -25464 21667 -25452
rect 20067 -25498 20079 -25464
rect 21655 -25498 21667 -25464
rect 20067 -25510 21667 -25498
rect 267 -25906 1867 -25894
rect 267 -25940 279 -25906
rect 1855 -25940 1867 -25906
rect 267 -25952 1867 -25940
rect 267 -26264 1867 -26252
rect 267 -26298 279 -26264
rect 1855 -26298 1867 -26264
rect 267 -26310 1867 -26298
rect 2467 -25906 4067 -25894
rect 2467 -25940 2479 -25906
rect 4055 -25940 4067 -25906
rect 2467 -25952 4067 -25940
rect 2467 -26264 4067 -26252
rect 2467 -26298 2479 -26264
rect 4055 -26298 4067 -26264
rect 2467 -26310 4067 -26298
rect 4667 -25906 6267 -25894
rect 4667 -25940 4679 -25906
rect 6255 -25940 6267 -25906
rect 4667 -25952 6267 -25940
rect 4667 -26264 6267 -26252
rect 4667 -26298 4679 -26264
rect 6255 -26298 6267 -26264
rect 4667 -26310 6267 -26298
rect 6867 -25906 8467 -25894
rect 6867 -25940 6879 -25906
rect 8455 -25940 8467 -25906
rect 6867 -25952 8467 -25940
rect 6867 -26264 8467 -26252
rect 6867 -26298 6879 -26264
rect 8455 -26298 8467 -26264
rect 6867 -26310 8467 -26298
rect 9067 -25906 10667 -25894
rect 9067 -25940 9079 -25906
rect 10655 -25940 10667 -25906
rect 9067 -25952 10667 -25940
rect 9067 -26264 10667 -26252
rect 9067 -26298 9079 -26264
rect 10655 -26298 10667 -26264
rect 9067 -26310 10667 -26298
rect 11267 -25906 12867 -25894
rect 11267 -25940 11279 -25906
rect 12855 -25940 12867 -25906
rect 11267 -25952 12867 -25940
rect 11267 -26264 12867 -26252
rect 11267 -26298 11279 -26264
rect 12855 -26298 12867 -26264
rect 11267 -26310 12867 -26298
rect 13467 -25906 15067 -25894
rect 13467 -25940 13479 -25906
rect 15055 -25940 15067 -25906
rect 13467 -25952 15067 -25940
rect 13467 -26264 15067 -26252
rect 13467 -26298 13479 -26264
rect 15055 -26298 15067 -26264
rect 13467 -26310 15067 -26298
rect 15667 -25906 17267 -25894
rect 15667 -25940 15679 -25906
rect 17255 -25940 17267 -25906
rect 15667 -25952 17267 -25940
rect 15667 -26264 17267 -26252
rect 15667 -26298 15679 -26264
rect 17255 -26298 17267 -26264
rect 15667 -26310 17267 -26298
rect 17867 -25906 19467 -25894
rect 17867 -25940 17879 -25906
rect 19455 -25940 19467 -25906
rect 17867 -25952 19467 -25940
rect 17867 -26264 19467 -26252
rect 17867 -26298 17879 -26264
rect 19455 -26298 19467 -26264
rect 17867 -26310 19467 -26298
rect 20067 -25906 21667 -25894
rect 20067 -25940 20079 -25906
rect 21655 -25940 21667 -25906
rect 20067 -25952 21667 -25940
rect 20067 -26264 21667 -26252
rect 20067 -26298 20079 -26264
rect 21655 -26298 21667 -26264
rect 20067 -26310 21667 -26298
rect 267 -26706 1867 -26694
rect 267 -26740 279 -26706
rect 1855 -26740 1867 -26706
rect 267 -26752 1867 -26740
rect 267 -27064 1867 -27052
rect 267 -27098 279 -27064
rect 1855 -27098 1867 -27064
rect 267 -27110 1867 -27098
rect 2467 -26706 4067 -26694
rect 2467 -26740 2479 -26706
rect 4055 -26740 4067 -26706
rect 2467 -26752 4067 -26740
rect 2467 -27064 4067 -27052
rect 2467 -27098 2479 -27064
rect 4055 -27098 4067 -27064
rect 2467 -27110 4067 -27098
rect 4667 -26706 6267 -26694
rect 4667 -26740 4679 -26706
rect 6255 -26740 6267 -26706
rect 4667 -26752 6267 -26740
rect 4667 -27064 6267 -27052
rect 4667 -27098 4679 -27064
rect 6255 -27098 6267 -27064
rect 4667 -27110 6267 -27098
rect 6867 -26706 8467 -26694
rect 6867 -26740 6879 -26706
rect 8455 -26740 8467 -26706
rect 6867 -26752 8467 -26740
rect 6867 -27064 8467 -27052
rect 6867 -27098 6879 -27064
rect 8455 -27098 8467 -27064
rect 6867 -27110 8467 -27098
rect 9067 -26706 10667 -26694
rect 9067 -26740 9079 -26706
rect 10655 -26740 10667 -26706
rect 9067 -26752 10667 -26740
rect 9067 -27064 10667 -27052
rect 9067 -27098 9079 -27064
rect 10655 -27098 10667 -27064
rect 9067 -27110 10667 -27098
rect 11267 -26706 12867 -26694
rect 11267 -26740 11279 -26706
rect 12855 -26740 12867 -26706
rect 11267 -26752 12867 -26740
rect 11267 -27064 12867 -27052
rect 11267 -27098 11279 -27064
rect 12855 -27098 12867 -27064
rect 11267 -27110 12867 -27098
rect 13467 -26706 15067 -26694
rect 13467 -26740 13479 -26706
rect 15055 -26740 15067 -26706
rect 13467 -26752 15067 -26740
rect 13467 -27064 15067 -27052
rect 13467 -27098 13479 -27064
rect 15055 -27098 15067 -27064
rect 13467 -27110 15067 -27098
rect 15667 -26706 17267 -26694
rect 15667 -26740 15679 -26706
rect 17255 -26740 17267 -26706
rect 15667 -26752 17267 -26740
rect 15667 -27064 17267 -27052
rect 15667 -27098 15679 -27064
rect 17255 -27098 17267 -27064
rect 15667 -27110 17267 -27098
rect 17867 -26706 19467 -26694
rect 17867 -26740 17879 -26706
rect 19455 -26740 19467 -26706
rect 17867 -26752 19467 -26740
rect 17867 -27064 19467 -27052
rect 17867 -27098 17879 -27064
rect 19455 -27098 19467 -27064
rect 17867 -27110 19467 -27098
rect 20067 -26706 21667 -26694
rect 20067 -26740 20079 -26706
rect 21655 -26740 21667 -26706
rect 20067 -26752 21667 -26740
rect 20067 -27064 21667 -27052
rect 20067 -27098 20079 -27064
rect 21655 -27098 21667 -27064
rect 20067 -27110 21667 -27098
rect 267 -27506 1867 -27494
rect 267 -27540 279 -27506
rect 1855 -27540 1867 -27506
rect 267 -27552 1867 -27540
rect 267 -27864 1867 -27852
rect 267 -27898 279 -27864
rect 1855 -27898 1867 -27864
rect 267 -27910 1867 -27898
rect 2467 -27506 4067 -27494
rect 2467 -27540 2479 -27506
rect 4055 -27540 4067 -27506
rect 2467 -27552 4067 -27540
rect 2467 -27864 4067 -27852
rect 2467 -27898 2479 -27864
rect 4055 -27898 4067 -27864
rect 2467 -27910 4067 -27898
rect 4667 -27506 6267 -27494
rect 4667 -27540 4679 -27506
rect 6255 -27540 6267 -27506
rect 4667 -27552 6267 -27540
rect 4667 -27864 6267 -27852
rect 4667 -27898 4679 -27864
rect 6255 -27898 6267 -27864
rect 4667 -27910 6267 -27898
rect 6867 -27506 8467 -27494
rect 6867 -27540 6879 -27506
rect 8455 -27540 8467 -27506
rect 6867 -27552 8467 -27540
rect 6867 -27864 8467 -27852
rect 6867 -27898 6879 -27864
rect 8455 -27898 8467 -27864
rect 6867 -27910 8467 -27898
rect 9067 -27506 10667 -27494
rect 9067 -27540 9079 -27506
rect 10655 -27540 10667 -27506
rect 9067 -27552 10667 -27540
rect 9067 -27864 10667 -27852
rect 9067 -27898 9079 -27864
rect 10655 -27898 10667 -27864
rect 9067 -27910 10667 -27898
rect 11267 -27506 12867 -27494
rect 11267 -27540 11279 -27506
rect 12855 -27540 12867 -27506
rect 11267 -27552 12867 -27540
rect 11267 -27864 12867 -27852
rect 11267 -27898 11279 -27864
rect 12855 -27898 12867 -27864
rect 11267 -27910 12867 -27898
rect 13467 -27506 15067 -27494
rect 13467 -27540 13479 -27506
rect 15055 -27540 15067 -27506
rect 13467 -27552 15067 -27540
rect 13467 -27864 15067 -27852
rect 13467 -27898 13479 -27864
rect 15055 -27898 15067 -27864
rect 13467 -27910 15067 -27898
rect 15667 -27506 17267 -27494
rect 15667 -27540 15679 -27506
rect 17255 -27540 17267 -27506
rect 15667 -27552 17267 -27540
rect 15667 -27864 17267 -27852
rect 15667 -27898 15679 -27864
rect 17255 -27898 17267 -27864
rect 15667 -27910 17267 -27898
rect 17867 -27506 19467 -27494
rect 17867 -27540 17879 -27506
rect 19455 -27540 19467 -27506
rect 17867 -27552 19467 -27540
rect 17867 -27864 19467 -27852
rect 17867 -27898 17879 -27864
rect 19455 -27898 19467 -27864
rect 17867 -27910 19467 -27898
rect 20067 -27506 21667 -27494
rect 20067 -27540 20079 -27506
rect 21655 -27540 21667 -27506
rect 20067 -27552 21667 -27540
rect 20067 -27864 21667 -27852
rect 20067 -27898 20079 -27864
rect 21655 -27898 21667 -27864
rect 20067 -27910 21667 -27898
rect 267 -28306 1867 -28294
rect 267 -28340 279 -28306
rect 1855 -28340 1867 -28306
rect 267 -28352 1867 -28340
rect 267 -28664 1867 -28652
rect 267 -28698 279 -28664
rect 1855 -28698 1867 -28664
rect 267 -28710 1867 -28698
rect 2467 -28306 4067 -28294
rect 2467 -28340 2479 -28306
rect 4055 -28340 4067 -28306
rect 2467 -28352 4067 -28340
rect 2467 -28664 4067 -28652
rect 2467 -28698 2479 -28664
rect 4055 -28698 4067 -28664
rect 2467 -28710 4067 -28698
rect 4667 -28306 6267 -28294
rect 4667 -28340 4679 -28306
rect 6255 -28340 6267 -28306
rect 4667 -28352 6267 -28340
rect 4667 -28664 6267 -28652
rect 4667 -28698 4679 -28664
rect 6255 -28698 6267 -28664
rect 4667 -28710 6267 -28698
rect 6867 -28306 8467 -28294
rect 6867 -28340 6879 -28306
rect 8455 -28340 8467 -28306
rect 6867 -28352 8467 -28340
rect 6867 -28664 8467 -28652
rect 6867 -28698 6879 -28664
rect 8455 -28698 8467 -28664
rect 6867 -28710 8467 -28698
rect 9067 -28306 10667 -28294
rect 9067 -28340 9079 -28306
rect 10655 -28340 10667 -28306
rect 9067 -28352 10667 -28340
rect 9067 -28664 10667 -28652
rect 9067 -28698 9079 -28664
rect 10655 -28698 10667 -28664
rect 9067 -28710 10667 -28698
rect 11267 -28306 12867 -28294
rect 11267 -28340 11279 -28306
rect 12855 -28340 12867 -28306
rect 11267 -28352 12867 -28340
rect 11267 -28664 12867 -28652
rect 11267 -28698 11279 -28664
rect 12855 -28698 12867 -28664
rect 11267 -28710 12867 -28698
rect 13467 -28306 15067 -28294
rect 13467 -28340 13479 -28306
rect 15055 -28340 15067 -28306
rect 13467 -28352 15067 -28340
rect 13467 -28664 15067 -28652
rect 13467 -28698 13479 -28664
rect 15055 -28698 15067 -28664
rect 13467 -28710 15067 -28698
rect 15667 -28306 17267 -28294
rect 15667 -28340 15679 -28306
rect 17255 -28340 17267 -28306
rect 15667 -28352 17267 -28340
rect 15667 -28664 17267 -28652
rect 15667 -28698 15679 -28664
rect 17255 -28698 17267 -28664
rect 15667 -28710 17267 -28698
rect 17867 -28306 19467 -28294
rect 17867 -28340 17879 -28306
rect 19455 -28340 19467 -28306
rect 17867 -28352 19467 -28340
rect 17867 -28664 19467 -28652
rect 17867 -28698 17879 -28664
rect 19455 -28698 19467 -28664
rect 17867 -28710 19467 -28698
rect 20067 -28306 21667 -28294
rect 20067 -28340 20079 -28306
rect 21655 -28340 21667 -28306
rect 20067 -28352 21667 -28340
rect 20067 -28664 21667 -28652
rect 20067 -28698 20079 -28664
rect 21655 -28698 21667 -28664
rect 20067 -28710 21667 -28698
rect 267 -29106 1867 -29094
rect 267 -29140 279 -29106
rect 1855 -29140 1867 -29106
rect 267 -29152 1867 -29140
rect 267 -29464 1867 -29452
rect 267 -29498 279 -29464
rect 1855 -29498 1867 -29464
rect 267 -29510 1867 -29498
rect 2467 -29106 4067 -29094
rect 2467 -29140 2479 -29106
rect 4055 -29140 4067 -29106
rect 2467 -29152 4067 -29140
rect 2467 -29464 4067 -29452
rect 2467 -29498 2479 -29464
rect 4055 -29498 4067 -29464
rect 2467 -29510 4067 -29498
rect 4667 -29106 6267 -29094
rect 4667 -29140 4679 -29106
rect 6255 -29140 6267 -29106
rect 4667 -29152 6267 -29140
rect 4667 -29464 6267 -29452
rect 4667 -29498 4679 -29464
rect 6255 -29498 6267 -29464
rect 4667 -29510 6267 -29498
rect 6867 -29106 8467 -29094
rect 6867 -29140 6879 -29106
rect 8455 -29140 8467 -29106
rect 6867 -29152 8467 -29140
rect 6867 -29464 8467 -29452
rect 6867 -29498 6879 -29464
rect 8455 -29498 8467 -29464
rect 6867 -29510 8467 -29498
rect 9067 -29106 10667 -29094
rect 9067 -29140 9079 -29106
rect 10655 -29140 10667 -29106
rect 9067 -29152 10667 -29140
rect 9067 -29464 10667 -29452
rect 9067 -29498 9079 -29464
rect 10655 -29498 10667 -29464
rect 9067 -29510 10667 -29498
rect 11267 -29106 12867 -29094
rect 11267 -29140 11279 -29106
rect 12855 -29140 12867 -29106
rect 11267 -29152 12867 -29140
rect 11267 -29464 12867 -29452
rect 11267 -29498 11279 -29464
rect 12855 -29498 12867 -29464
rect 11267 -29510 12867 -29498
rect 13467 -29106 15067 -29094
rect 13467 -29140 13479 -29106
rect 15055 -29140 15067 -29106
rect 13467 -29152 15067 -29140
rect 13467 -29464 15067 -29452
rect 13467 -29498 13479 -29464
rect 15055 -29498 15067 -29464
rect 13467 -29510 15067 -29498
rect 15667 -29106 17267 -29094
rect 15667 -29140 15679 -29106
rect 17255 -29140 17267 -29106
rect 15667 -29152 17267 -29140
rect 15667 -29464 17267 -29452
rect 15667 -29498 15679 -29464
rect 17255 -29498 17267 -29464
rect 15667 -29510 17267 -29498
rect 17867 -29106 19467 -29094
rect 17867 -29140 17879 -29106
rect 19455 -29140 19467 -29106
rect 17867 -29152 19467 -29140
rect 17867 -29464 19467 -29452
rect 17867 -29498 17879 -29464
rect 19455 -29498 19467 -29464
rect 17867 -29510 19467 -29498
rect 20067 -29106 21667 -29094
rect 20067 -29140 20079 -29106
rect 21655 -29140 21667 -29106
rect 20067 -29152 21667 -29140
rect 20067 -29464 21667 -29452
rect 20067 -29498 20079 -29464
rect 21655 -29498 21667 -29464
rect 20067 -29510 21667 -29498
rect 267 -29906 1867 -29894
rect 267 -29940 279 -29906
rect 1855 -29940 1867 -29906
rect 267 -29952 1867 -29940
rect 267 -30264 1867 -30252
rect 267 -30298 279 -30264
rect 1855 -30298 1867 -30264
rect 267 -30310 1867 -30298
rect 2467 -29906 4067 -29894
rect 2467 -29940 2479 -29906
rect 4055 -29940 4067 -29906
rect 2467 -29952 4067 -29940
rect 2467 -30264 4067 -30252
rect 2467 -30298 2479 -30264
rect 4055 -30298 4067 -30264
rect 2467 -30310 4067 -30298
rect 4667 -29906 6267 -29894
rect 4667 -29940 4679 -29906
rect 6255 -29940 6267 -29906
rect 4667 -29952 6267 -29940
rect 4667 -30264 6267 -30252
rect 4667 -30298 4679 -30264
rect 6255 -30298 6267 -30264
rect 4667 -30310 6267 -30298
rect 6867 -29906 8467 -29894
rect 6867 -29940 6879 -29906
rect 8455 -29940 8467 -29906
rect 6867 -29952 8467 -29940
rect 6867 -30264 8467 -30252
rect 6867 -30298 6879 -30264
rect 8455 -30298 8467 -30264
rect 6867 -30310 8467 -30298
rect 9067 -29906 10667 -29894
rect 9067 -29940 9079 -29906
rect 10655 -29940 10667 -29906
rect 9067 -29952 10667 -29940
rect 9067 -30264 10667 -30252
rect 9067 -30298 9079 -30264
rect 10655 -30298 10667 -30264
rect 9067 -30310 10667 -30298
rect 11267 -29906 12867 -29894
rect 11267 -29940 11279 -29906
rect 12855 -29940 12867 -29906
rect 11267 -29952 12867 -29940
rect 11267 -30264 12867 -30252
rect 11267 -30298 11279 -30264
rect 12855 -30298 12867 -30264
rect 11267 -30310 12867 -30298
rect 13467 -29906 15067 -29894
rect 13467 -29940 13479 -29906
rect 15055 -29940 15067 -29906
rect 13467 -29952 15067 -29940
rect 13467 -30264 15067 -30252
rect 13467 -30298 13479 -30264
rect 15055 -30298 15067 -30264
rect 13467 -30310 15067 -30298
rect 15667 -29906 17267 -29894
rect 15667 -29940 15679 -29906
rect 17255 -29940 17267 -29906
rect 15667 -29952 17267 -29940
rect 15667 -30264 17267 -30252
rect 15667 -30298 15679 -30264
rect 17255 -30298 17267 -30264
rect 15667 -30310 17267 -30298
rect 17867 -29906 19467 -29894
rect 17867 -29940 17879 -29906
rect 19455 -29940 19467 -29906
rect 17867 -29952 19467 -29940
rect 17867 -30264 19467 -30252
rect 17867 -30298 17879 -30264
rect 19455 -30298 19467 -30264
rect 17867 -30310 19467 -30298
rect 20067 -29906 21667 -29894
rect 20067 -29940 20079 -29906
rect 21655 -29940 21667 -29906
rect 20067 -29952 21667 -29940
rect 20067 -30264 21667 -30252
rect 20067 -30298 20079 -30264
rect 21655 -30298 21667 -30264
rect 20067 -30310 21667 -30298
rect 267 -30706 1867 -30694
rect 267 -30740 279 -30706
rect 1855 -30740 1867 -30706
rect 267 -30752 1867 -30740
rect 267 -31064 1867 -31052
rect 267 -31098 279 -31064
rect 1855 -31098 1867 -31064
rect 267 -31110 1867 -31098
rect 2467 -30706 4067 -30694
rect 2467 -30740 2479 -30706
rect 4055 -30740 4067 -30706
rect 2467 -30752 4067 -30740
rect 2467 -31064 4067 -31052
rect 2467 -31098 2479 -31064
rect 4055 -31098 4067 -31064
rect 2467 -31110 4067 -31098
rect 4667 -30706 6267 -30694
rect 4667 -30740 4679 -30706
rect 6255 -30740 6267 -30706
rect 4667 -30752 6267 -30740
rect 4667 -31064 6267 -31052
rect 4667 -31098 4679 -31064
rect 6255 -31098 6267 -31064
rect 4667 -31110 6267 -31098
rect 6867 -30706 8467 -30694
rect 6867 -30740 6879 -30706
rect 8455 -30740 8467 -30706
rect 6867 -30752 8467 -30740
rect 6867 -31064 8467 -31052
rect 6867 -31098 6879 -31064
rect 8455 -31098 8467 -31064
rect 6867 -31110 8467 -31098
rect 9067 -30706 10667 -30694
rect 9067 -30740 9079 -30706
rect 10655 -30740 10667 -30706
rect 9067 -30752 10667 -30740
rect 9067 -31064 10667 -31052
rect 9067 -31098 9079 -31064
rect 10655 -31098 10667 -31064
rect 9067 -31110 10667 -31098
rect 11267 -30706 12867 -30694
rect 11267 -30740 11279 -30706
rect 12855 -30740 12867 -30706
rect 11267 -30752 12867 -30740
rect 11267 -31064 12867 -31052
rect 11267 -31098 11279 -31064
rect 12855 -31098 12867 -31064
rect 11267 -31110 12867 -31098
rect 13467 -30706 15067 -30694
rect 13467 -30740 13479 -30706
rect 15055 -30740 15067 -30706
rect 13467 -30752 15067 -30740
rect 13467 -31064 15067 -31052
rect 13467 -31098 13479 -31064
rect 15055 -31098 15067 -31064
rect 13467 -31110 15067 -31098
rect 15667 -30706 17267 -30694
rect 15667 -30740 15679 -30706
rect 17255 -30740 17267 -30706
rect 15667 -30752 17267 -30740
rect 15667 -31064 17267 -31052
rect 15667 -31098 15679 -31064
rect 17255 -31098 17267 -31064
rect 15667 -31110 17267 -31098
rect 17867 -30706 19467 -30694
rect 17867 -30740 17879 -30706
rect 19455 -30740 19467 -30706
rect 17867 -30752 19467 -30740
rect 17867 -31064 19467 -31052
rect 17867 -31098 17879 -31064
rect 19455 -31098 19467 -31064
rect 17867 -31110 19467 -31098
rect 20067 -30706 21667 -30694
rect 20067 -30740 20079 -30706
rect 21655 -30740 21667 -30706
rect 20067 -30752 21667 -30740
rect 20067 -31064 21667 -31052
rect 20067 -31098 20079 -31064
rect 21655 -31098 21667 -31064
rect 20067 -31110 21667 -31098
rect 267 -31506 1867 -31494
rect 267 -31540 279 -31506
rect 1855 -31540 1867 -31506
rect 267 -31552 1867 -31540
rect 267 -31864 1867 -31852
rect 267 -31898 279 -31864
rect 1855 -31898 1867 -31864
rect 267 -31910 1867 -31898
rect 2467 -31506 4067 -31494
rect 2467 -31540 2479 -31506
rect 4055 -31540 4067 -31506
rect 2467 -31552 4067 -31540
rect 2467 -31864 4067 -31852
rect 2467 -31898 2479 -31864
rect 4055 -31898 4067 -31864
rect 2467 -31910 4067 -31898
rect 4667 -31506 6267 -31494
rect 4667 -31540 4679 -31506
rect 6255 -31540 6267 -31506
rect 4667 -31552 6267 -31540
rect 4667 -31864 6267 -31852
rect 4667 -31898 4679 -31864
rect 6255 -31898 6267 -31864
rect 4667 -31910 6267 -31898
rect 6867 -31506 8467 -31494
rect 6867 -31540 6879 -31506
rect 8455 -31540 8467 -31506
rect 6867 -31552 8467 -31540
rect 6867 -31864 8467 -31852
rect 6867 -31898 6879 -31864
rect 8455 -31898 8467 -31864
rect 6867 -31910 8467 -31898
rect 9067 -31506 10667 -31494
rect 9067 -31540 9079 -31506
rect 10655 -31540 10667 -31506
rect 9067 -31552 10667 -31540
rect 9067 -31864 10667 -31852
rect 9067 -31898 9079 -31864
rect 10655 -31898 10667 -31864
rect 9067 -31910 10667 -31898
rect 11267 -31506 12867 -31494
rect 11267 -31540 11279 -31506
rect 12855 -31540 12867 -31506
rect 11267 -31552 12867 -31540
rect 11267 -31864 12867 -31852
rect 11267 -31898 11279 -31864
rect 12855 -31898 12867 -31864
rect 11267 -31910 12867 -31898
rect 13467 -31506 15067 -31494
rect 13467 -31540 13479 -31506
rect 15055 -31540 15067 -31506
rect 13467 -31552 15067 -31540
rect 13467 -31864 15067 -31852
rect 13467 -31898 13479 -31864
rect 15055 -31898 15067 -31864
rect 13467 -31910 15067 -31898
rect 15667 -31506 17267 -31494
rect 15667 -31540 15679 -31506
rect 17255 -31540 17267 -31506
rect 15667 -31552 17267 -31540
rect 15667 -31864 17267 -31852
rect 15667 -31898 15679 -31864
rect 17255 -31898 17267 -31864
rect 15667 -31910 17267 -31898
rect 17867 -31506 19467 -31494
rect 17867 -31540 17879 -31506
rect 19455 -31540 19467 -31506
rect 17867 -31552 19467 -31540
rect 17867 -31864 19467 -31852
rect 17867 -31898 17879 -31864
rect 19455 -31898 19467 -31864
rect 17867 -31910 19467 -31898
rect 20067 -31506 21667 -31494
rect 20067 -31540 20079 -31506
rect 21655 -31540 21667 -31506
rect 20067 -31552 21667 -31540
rect 20067 -31864 21667 -31852
rect 20067 -31898 20079 -31864
rect 21655 -31898 21667 -31864
rect 20067 -31910 21667 -31898
rect 34977 -24830 35777 -24818
rect 34977 -24864 34989 -24830
rect 35765 -24864 35777 -24830
rect 34977 -24876 35777 -24864
rect 34977 -25088 35777 -25076
rect 34977 -25122 34989 -25088
rect 35765 -25122 35777 -25088
rect 34977 -25134 35777 -25122
rect 34977 -25346 35777 -25334
rect 34977 -25380 34989 -25346
rect 35765 -25380 35777 -25346
rect 34977 -25392 35777 -25380
rect 34977 -25604 35777 -25592
rect 34977 -25638 34989 -25604
rect 35765 -25638 35777 -25604
rect 34977 -25650 35777 -25638
rect 34977 -25862 35777 -25850
rect 34977 -25896 34989 -25862
rect 35765 -25896 35777 -25862
rect 34977 -25908 35777 -25896
rect 34977 -26120 35777 -26108
rect 34977 -26154 34989 -26120
rect 35765 -26154 35777 -26120
rect 34977 -26166 35777 -26154
rect 34977 -26378 35777 -26366
rect 34977 -26412 34989 -26378
rect 35765 -26412 35777 -26378
rect 34977 -26424 35777 -26412
rect 34977 -26636 35777 -26624
rect 34977 -26670 34989 -26636
rect 35765 -26670 35777 -26636
rect 34977 -26682 35777 -26670
rect 34977 -26894 35777 -26882
rect 34977 -26928 34989 -26894
rect 35765 -26928 35777 -26894
rect 34977 -26940 35777 -26928
rect 36317 -24830 37117 -24818
rect 36317 -24864 36329 -24830
rect 37105 -24864 37117 -24830
rect 36317 -24876 37117 -24864
rect 36317 -25088 37117 -25076
rect 36317 -25122 36329 -25088
rect 37105 -25122 37117 -25088
rect 36317 -25134 37117 -25122
rect 36317 -25346 37117 -25334
rect 36317 -25380 36329 -25346
rect 37105 -25380 37117 -25346
rect 36317 -25392 37117 -25380
rect 36317 -25604 37117 -25592
rect 36317 -25638 36329 -25604
rect 37105 -25638 37117 -25604
rect 36317 -25650 37117 -25638
rect 36317 -25862 37117 -25850
rect 36317 -25896 36329 -25862
rect 37105 -25896 37117 -25862
rect 36317 -25908 37117 -25896
rect 36317 -26120 37117 -26108
rect 36317 -26154 36329 -26120
rect 37105 -26154 37117 -26120
rect 36317 -26166 37117 -26154
rect 36317 -26378 37117 -26366
rect 36317 -26412 36329 -26378
rect 37105 -26412 37117 -26378
rect 36317 -26424 37117 -26412
rect 36317 -26636 37117 -26624
rect 36317 -26670 36329 -26636
rect 37105 -26670 37117 -26636
rect 36317 -26682 37117 -26670
rect 36317 -26894 37117 -26882
rect 36317 -26928 36329 -26894
rect 37105 -26928 37117 -26894
rect 36317 -26940 37117 -26928
rect 31800 -28533 31858 -28521
rect 31800 -28909 31812 -28533
rect 31846 -28909 31858 -28533
rect 31800 -28921 31858 -28909
rect 31958 -28533 32016 -28521
rect 31958 -28909 31970 -28533
rect 32004 -28909 32016 -28533
rect 31958 -28921 32016 -28909
rect 32240 -28533 32298 -28521
rect 32240 -28909 32252 -28533
rect 32286 -28909 32298 -28533
rect 32240 -28921 32298 -28909
rect 32398 -28533 32456 -28521
rect 32398 -28909 32410 -28533
rect 32444 -28909 32456 -28533
rect 32398 -28921 32456 -28909
rect 32680 -28533 32738 -28521
rect 32680 -28909 32692 -28533
rect 32726 -28909 32738 -28533
rect 32680 -28921 32738 -28909
rect 32838 -28533 32896 -28521
rect 32838 -28909 32850 -28533
rect 32884 -28909 32896 -28533
rect 32838 -28921 32896 -28909
rect 33094 -28833 33152 -28821
rect 33094 -28909 33106 -28833
rect 33140 -28909 33152 -28833
rect 33094 -28921 33152 -28909
rect 33552 -28833 33610 -28821
rect 33552 -28909 33564 -28833
rect 33598 -28909 33610 -28833
rect 33552 -28921 33610 -28909
rect 34000 -28533 34058 -28521
rect 34000 -28909 34012 -28533
rect 34046 -28909 34058 -28533
rect 34000 -28921 34058 -28909
rect 34158 -28533 34216 -28521
rect 34158 -28909 34170 -28533
rect 34204 -28909 34216 -28533
rect 34158 -28921 34216 -28909
rect 34440 -28533 34498 -28521
rect 34440 -28909 34452 -28533
rect 34486 -28909 34498 -28533
rect 34440 -28921 34498 -28909
rect 34598 -28533 34656 -28521
rect 34598 -28909 34610 -28533
rect 34644 -28909 34656 -28533
rect 34598 -28921 34656 -28909
rect 34880 -28533 34938 -28521
rect 34880 -28909 34892 -28533
rect 34926 -28909 34938 -28533
rect 34880 -28921 34938 -28909
rect 35038 -28533 35096 -28521
rect 35038 -28909 35050 -28533
rect 35084 -28909 35096 -28533
rect 35038 -28921 35096 -28909
rect 35294 -28833 35352 -28821
rect 35294 -28909 35306 -28833
rect 35340 -28909 35352 -28833
rect 35294 -28921 35352 -28909
rect 35752 -28833 35810 -28821
rect 35752 -28909 35764 -28833
rect 35798 -28909 35810 -28833
rect 35752 -28921 35810 -28909
rect 36200 -28533 36258 -28521
rect 36200 -28909 36212 -28533
rect 36246 -28909 36258 -28533
rect 36200 -28921 36258 -28909
rect 36358 -28533 36416 -28521
rect 36358 -28909 36370 -28533
rect 36404 -28909 36416 -28533
rect 36358 -28921 36416 -28909
rect 36640 -28533 36698 -28521
rect 36640 -28909 36652 -28533
rect 36686 -28909 36698 -28533
rect 36640 -28921 36698 -28909
rect 36798 -28533 36856 -28521
rect 36798 -28909 36810 -28533
rect 36844 -28909 36856 -28533
rect 36798 -28921 36856 -28909
rect 37080 -28533 37138 -28521
rect 37080 -28909 37092 -28533
rect 37126 -28909 37138 -28533
rect 37080 -28921 37138 -28909
rect 37238 -28533 37296 -28521
rect 37238 -28909 37250 -28533
rect 37284 -28909 37296 -28533
rect 37238 -28921 37296 -28909
rect 37494 -28833 37552 -28821
rect 37494 -28909 37506 -28833
rect 37540 -28909 37552 -28833
rect 37494 -28921 37552 -28909
rect 37952 -28833 38010 -28821
rect 37952 -28909 37964 -28833
rect 37998 -28909 38010 -28833
rect 37952 -28921 38010 -28909
rect 31812 -31115 31870 -31103
rect 31812 -31191 31824 -31115
rect 31858 -31191 31870 -31115
rect 31812 -31203 31870 -31191
rect 32270 -31115 32328 -31103
rect 32270 -31191 32282 -31115
rect 32316 -31191 32328 -31115
rect 32270 -31203 32328 -31191
rect 32526 -31115 32584 -31103
rect 32526 -31491 32538 -31115
rect 32572 -31491 32584 -31115
rect 32526 -31503 32584 -31491
rect 32684 -31115 32742 -31103
rect 32684 -31491 32696 -31115
rect 32730 -31491 32742 -31115
rect 32684 -31503 32742 -31491
rect 32966 -31115 33024 -31103
rect 32966 -31491 32978 -31115
rect 33012 -31491 33024 -31115
rect 32966 -31503 33024 -31491
rect 33124 -31115 33182 -31103
rect 33124 -31491 33136 -31115
rect 33170 -31491 33182 -31115
rect 33124 -31503 33182 -31491
rect 33406 -31115 33464 -31103
rect 33406 -31491 33418 -31115
rect 33452 -31491 33464 -31115
rect 33406 -31503 33464 -31491
rect 33564 -31115 33622 -31103
rect 33564 -31491 33576 -31115
rect 33610 -31491 33622 -31115
rect 33564 -31503 33622 -31491
rect 34012 -31115 34070 -31103
rect 34012 -31191 34024 -31115
rect 34058 -31191 34070 -31115
rect 34012 -31203 34070 -31191
rect 34470 -31115 34528 -31103
rect 34470 -31191 34482 -31115
rect 34516 -31191 34528 -31115
rect 34470 -31203 34528 -31191
rect 34726 -31115 34784 -31103
rect 34726 -31491 34738 -31115
rect 34772 -31491 34784 -31115
rect 34726 -31503 34784 -31491
rect 34884 -31115 34942 -31103
rect 34884 -31491 34896 -31115
rect 34930 -31491 34942 -31115
rect 34884 -31503 34942 -31491
rect 35166 -31115 35224 -31103
rect 35166 -31491 35178 -31115
rect 35212 -31491 35224 -31115
rect 35166 -31503 35224 -31491
rect 35324 -31115 35382 -31103
rect 35324 -31491 35336 -31115
rect 35370 -31491 35382 -31115
rect 35324 -31503 35382 -31491
rect 35606 -31115 35664 -31103
rect 35606 -31491 35618 -31115
rect 35652 -31491 35664 -31115
rect 35606 -31503 35664 -31491
rect 35764 -31115 35822 -31103
rect 35764 -31491 35776 -31115
rect 35810 -31491 35822 -31115
rect 35764 -31503 35822 -31491
rect 36212 -31115 36270 -31103
rect 36212 -31191 36224 -31115
rect 36258 -31191 36270 -31115
rect 36212 -31203 36270 -31191
rect 36670 -31115 36728 -31103
rect 36670 -31191 36682 -31115
rect 36716 -31191 36728 -31115
rect 36670 -31203 36728 -31191
rect 36926 -31115 36984 -31103
rect 36926 -31491 36938 -31115
rect 36972 -31491 36984 -31115
rect 36926 -31503 36984 -31491
rect 37084 -31115 37142 -31103
rect 37084 -31491 37096 -31115
rect 37130 -31491 37142 -31115
rect 37084 -31503 37142 -31491
rect 37366 -31115 37424 -31103
rect 37366 -31491 37378 -31115
rect 37412 -31491 37424 -31115
rect 37366 -31503 37424 -31491
rect 37524 -31115 37582 -31103
rect 37524 -31491 37536 -31115
rect 37570 -31491 37582 -31115
rect 37524 -31503 37582 -31491
rect 37806 -31115 37864 -31103
rect 37806 -31491 37818 -31115
rect 37852 -31491 37864 -31115
rect 37806 -31503 37864 -31491
rect 37964 -31115 38022 -31103
rect 37964 -31491 37976 -31115
rect 38010 -31491 38022 -31115
rect 37964 -31503 38022 -31491
<< ndiffc >>
rect 34590 7142 34624 7318
rect 34678 7142 34712 7318
rect 35010 7142 35044 7318
rect 35098 7142 35132 7318
rect 35430 7142 35464 7318
rect 35518 7142 35552 7318
<< pdiffc >>
rect 32910 8071 32944 8847
rect 33168 8071 33202 8847
rect 33426 8071 33460 8847
rect 33750 8071 33784 8847
rect 34008 8071 34042 8847
rect 34266 8071 34300 8847
rect 34590 8251 34624 8627
rect 34678 8251 34712 8627
rect 35010 8251 35044 8627
rect 35098 8251 35132 8627
rect 35430 8251 35464 8627
rect 35518 8251 35552 8627
<< mvndiffc >>
rect 271 11741 1847 11775
rect 271 11383 1847 11417
rect 2471 11741 4047 11775
rect 2471 11383 4047 11417
rect 4671 11741 6247 11775
rect 4671 11383 6247 11417
rect 6871 11741 8447 11775
rect 6871 11383 8447 11417
rect 9071 11741 10647 11775
rect 9071 11383 10647 11417
rect 11271 11741 12847 11775
rect 11271 11383 12847 11417
rect 13471 11741 15047 11775
rect 13471 11383 15047 11417
rect 15671 11741 17247 11775
rect 15671 11383 17247 11417
rect 17871 11741 19447 11775
rect 17871 11383 19447 11417
rect 20071 11741 21647 11775
rect 20071 11383 21647 11417
rect 271 10941 1847 10975
rect 271 10583 1847 10617
rect 2470 10940 4046 10974
rect 2470 10582 4046 10616
rect 4670 10940 6246 10974
rect 4670 10582 6246 10616
rect 6870 10940 8446 10974
rect 6870 10582 8446 10616
rect 9070 10940 10646 10974
rect 9070 10582 10646 10616
rect 11270 10940 12846 10974
rect 11270 10582 12846 10616
rect 13470 10940 15046 10974
rect 13470 10582 15046 10616
rect 15670 10940 17246 10974
rect 15670 10582 17246 10616
rect 17870 10940 19446 10974
rect 17870 10582 19446 10616
rect 20071 10941 21647 10975
rect 20071 10583 21647 10617
rect 271 10141 1847 10175
rect 271 9783 1847 9817
rect 2470 10140 4046 10174
rect 2470 9782 4046 9816
rect 4670 10140 6246 10174
rect 4670 9782 6246 9816
rect 6870 10140 8446 10174
rect 6870 9782 8446 9816
rect 9070 10140 10646 10174
rect 9070 9782 10646 9816
rect 11270 10140 12846 10174
rect 11270 9782 12846 9816
rect 13470 10140 15046 10174
rect 13470 9782 15046 9816
rect 15670 10140 17246 10174
rect 15670 9782 17246 9816
rect 17870 10140 19446 10174
rect 17870 9782 19446 9816
rect 20071 10141 21647 10175
rect 20071 9783 21647 9817
rect 271 9341 1847 9375
rect 271 8983 1847 9017
rect 2470 9340 4046 9374
rect 2470 8982 4046 9016
rect 4670 9340 6246 9374
rect 4670 8982 6246 9016
rect 6870 9340 8446 9374
rect 6870 8982 8446 9016
rect 9070 9340 10646 9374
rect 9070 8982 10646 9016
rect 11270 9340 12846 9374
rect 11270 8982 12846 9016
rect 13470 9340 15046 9374
rect 13470 8982 15046 9016
rect 15670 9340 17246 9374
rect 15670 8982 17246 9016
rect 17870 9340 19446 9374
rect 17870 8982 19446 9016
rect 20071 9341 21647 9375
rect 20071 8983 21647 9017
rect 271 8541 1847 8575
rect 271 8183 1847 8217
rect 2470 8540 4046 8574
rect 2470 8182 4046 8216
rect 4670 8540 6246 8574
rect 4670 8182 6246 8216
rect 6870 8540 8446 8574
rect 6870 8182 8446 8216
rect 9070 8540 10646 8574
rect 9070 8182 10646 8216
rect 11270 8540 12846 8574
rect 11270 8182 12846 8216
rect 13470 8540 15046 8574
rect 13470 8182 15046 8216
rect 15670 8540 17246 8574
rect 15670 8182 17246 8216
rect 17870 8540 19446 8574
rect 17870 8182 19446 8216
rect 20071 8541 21647 8575
rect 20071 8183 21647 8217
rect 271 7741 1847 7775
rect 271 7383 1847 7417
rect 2470 7740 4046 7774
rect 2470 7382 4046 7416
rect 4670 7740 6246 7774
rect 4670 7382 6246 7416
rect 6870 7740 8446 7774
rect 6870 7382 8446 7416
rect 9070 7740 10646 7774
rect 9070 7382 10646 7416
rect 11270 7740 12846 7774
rect 11270 7382 12846 7416
rect 13470 7740 15046 7774
rect 13470 7382 15046 7416
rect 15670 7740 17246 7774
rect 15670 7382 17246 7416
rect 17870 7740 19446 7774
rect 17870 7382 19446 7416
rect 20071 7741 21647 7775
rect 20071 7383 21647 7417
rect 271 6941 1847 6975
rect 271 6583 1847 6617
rect 2470 6940 4046 6974
rect 2470 6582 4046 6616
rect 4670 6940 6246 6974
rect 4670 6582 6246 6616
rect 6870 6940 8446 6974
rect 6870 6582 8446 6616
rect 9070 6940 10646 6974
rect 9070 6582 10646 6616
rect 11270 6940 12846 6974
rect 11270 6582 12846 6616
rect 13470 6940 15046 6974
rect 13470 6582 15046 6616
rect 15670 6940 17246 6974
rect 15670 6582 17246 6616
rect 17870 6940 19446 6974
rect 17870 6582 19446 6616
rect 20071 6941 21647 6975
rect 20071 6583 21647 6617
rect 271 6141 1847 6175
rect 271 5783 1847 5817
rect 2470 6140 4046 6174
rect 2470 5782 4046 5816
rect 4670 6140 6246 6174
rect 4670 5782 6246 5816
rect 6870 6140 8446 6174
rect 6870 5782 8446 5816
rect 9070 6140 10646 6174
rect 9070 5782 10646 5816
rect 11270 6140 12846 6174
rect 11270 5782 12846 5816
rect 13470 6140 15046 6174
rect 13470 5782 15046 5816
rect 15670 6140 17246 6174
rect 15670 5782 17246 5816
rect 17870 6140 19446 6174
rect 17870 5782 19446 5816
rect 20071 6141 21647 6175
rect 20071 5783 21647 5817
rect 271 5341 1847 5375
rect 271 4983 1847 5017
rect 2470 5340 4046 5374
rect 2470 4982 4046 5016
rect 4670 5340 6246 5374
rect 4670 4982 6246 5016
rect 6870 5340 8446 5374
rect 6870 4982 8446 5016
rect 9070 5340 10646 5374
rect 9070 4982 10646 5016
rect 11270 5340 12846 5374
rect 11270 4982 12846 5016
rect 13470 5340 15046 5374
rect 13470 4982 15046 5016
rect 15670 5340 17246 5374
rect 15670 4982 17246 5016
rect 17870 5340 19446 5374
rect 17870 4982 19446 5016
rect 20071 5341 21647 5375
rect 20071 4983 21647 5017
rect 271 4541 1847 4575
rect 271 4183 1847 4217
rect 2471 4541 4047 4575
rect 2471 4183 4047 4217
rect 4671 4541 6247 4575
rect 4671 4183 6247 4217
rect 6871 4541 8447 4575
rect 6871 4183 8447 4217
rect 9072 4542 10648 4576
rect 9072 4184 10648 4218
rect 11272 4542 12848 4576
rect 11272 4184 12848 4218
rect 13471 4541 15047 4575
rect 13471 4183 15047 4217
rect 15671 4541 17247 4575
rect 15671 4183 17247 4217
rect 17871 4541 19447 4575
rect 17871 4183 19447 4217
rect 20071 4541 21647 4575
rect 20071 4183 21647 4217
rect 30102 11539 30136 11715
rect 30260 11539 30294 11715
rect 30418 11539 30452 11715
rect 30576 11539 30610 11715
rect 30857 11539 30891 11715
rect 31015 11539 31049 11715
rect 31297 11539 31331 11715
rect 31455 11539 31489 11715
rect 31737 11539 31771 11715
rect 31895 11539 31929 11715
rect 32302 11539 32336 11715
rect 32460 11539 32494 11715
rect 32618 11539 32652 11715
rect 32776 11539 32810 11715
rect 33057 11539 33091 11715
rect 33215 11539 33249 11715
rect 33497 11539 33531 11715
rect 33655 11539 33689 11715
rect 33937 11539 33971 11715
rect 34095 11539 34129 11715
rect 34502 11539 34536 11715
rect 34660 11539 34694 11715
rect 34818 11539 34852 11715
rect 34976 11539 35010 11715
rect 35257 11539 35291 11715
rect 35415 11539 35449 11715
rect 35697 11539 35731 11715
rect 35855 11539 35889 11715
rect 36137 11539 36171 11715
rect 36295 11539 36329 11715
rect 33472 7050 33506 7426
rect 33630 7050 33664 7426
rect 33788 7050 33822 7426
rect 33946 7050 33980 7426
rect 34104 7050 34138 7426
rect 29770 6200 30546 6234
rect 29770 5942 30546 5976
rect 31110 6200 31886 6234
rect 31110 5942 31886 5976
rect 29922 5420 29956 5496
rect 30380 5420 30414 5496
rect 31232 5420 31266 5496
rect 31690 5420 31724 5496
rect 29770 4940 30546 4974
rect 29770 4682 30546 4716
rect 31110 4940 31886 4974
rect 31110 4682 31886 4716
rect 17102 2528 17136 3304
rect 17260 2528 17294 3304
rect 17418 2528 17452 3304
rect 17576 2528 17610 3304
rect 17734 2528 17768 3304
rect 32722 3570 32756 3946
rect 32880 3570 32914 3946
rect 33038 3570 33072 3946
rect 33196 3570 33230 3946
rect 33354 3570 33388 3946
rect 33512 3570 33546 3946
rect 33670 3570 33704 3946
rect 33828 3570 33862 3946
rect 33986 3570 34020 3946
rect 34912 3570 34946 3946
rect 35070 3570 35104 3946
rect 35228 3570 35262 3946
rect 35386 3570 35420 3946
rect 36460 5966 36836 6000
rect 36460 5708 36836 5742
rect 36460 5450 36836 5484
rect 36460 5192 36836 5226
rect 36460 4934 36836 4968
rect 36460 4676 36836 4710
rect 36460 4418 36836 4452
rect 36460 4160 36836 4194
rect 36460 3902 36836 3936
rect 37246 5966 37622 6000
rect 37246 5708 37622 5742
rect 37246 5450 37622 5484
rect 37246 5192 37622 5226
rect 37246 4934 37622 4968
rect 37246 4676 37622 4710
rect 37246 4418 37622 4452
rect 37246 4160 37622 4194
rect 37246 3902 37622 3936
rect 32392 2640 32426 3016
rect 32550 2640 32584 3016
rect 32708 2640 32742 3016
rect 33992 2640 34026 3016
rect 34150 2640 34184 3016
rect 34308 2640 34342 3016
rect 35592 2640 35626 3016
rect 35750 2640 35784 3016
rect 35908 2640 35942 3016
rect 71 2061 447 2095
rect 689 2061 1065 2095
rect 71 1203 447 1237
rect 689 1203 1065 1237
rect 71 915 447 949
rect 689 915 1065 949
rect 71 657 447 691
rect 689 657 1065 691
rect 1671 2061 2047 2095
rect 2289 2061 2665 2095
rect 1671 1203 2047 1237
rect 2289 1203 2665 1237
rect 1671 915 2047 949
rect 2289 915 2665 949
rect 1671 657 2047 691
rect 2289 657 2665 691
rect 3271 2061 3647 2095
rect 3889 2061 4265 2095
rect 3271 1203 3647 1237
rect 3889 1203 4265 1237
rect 3271 915 3647 949
rect 3889 915 4265 949
rect 3271 657 3647 691
rect 3889 657 4265 691
rect 4871 2061 5247 2095
rect 5489 2061 5865 2095
rect 4871 1203 5247 1237
rect 5489 1203 5865 1237
rect 4871 915 5247 949
rect 5489 915 5865 949
rect 4871 657 5247 691
rect 5489 657 5865 691
rect 6471 2061 6847 2095
rect 7089 2061 7465 2095
rect 6471 1203 6847 1237
rect 7089 1203 7465 1237
rect 6471 915 6847 949
rect 7089 915 7465 949
rect 6471 657 6847 691
rect 7089 657 7465 691
rect 8071 2061 8447 2095
rect 8689 2061 9065 2095
rect 8071 1203 8447 1237
rect 8689 1203 9065 1237
rect 8071 915 8447 949
rect 8689 915 9065 949
rect 8071 657 8447 691
rect 8689 657 9065 691
rect 9671 2061 10047 2095
rect 10289 2061 10665 2095
rect 9671 1203 10047 1237
rect 10289 1203 10665 1237
rect 9671 915 10047 949
rect 10289 915 10665 949
rect 9671 657 10047 691
rect 10289 657 10665 691
rect 11271 2061 11647 2095
rect 11889 2061 12265 2095
rect 11271 1203 11647 1237
rect 11889 1203 12265 1237
rect 11271 915 11647 949
rect 11889 915 12265 949
rect 11271 657 11647 691
rect 11889 657 12265 691
rect 12871 2061 13247 2095
rect 13489 2061 13865 2095
rect 12871 1203 13247 1237
rect 13489 1203 13865 1237
rect 12871 915 13247 949
rect 13489 915 13865 949
rect 12871 657 13247 691
rect 13489 657 13865 691
rect 14471 2061 14847 2095
rect 15089 2061 15465 2095
rect 14471 1203 14847 1237
rect 15089 1203 15465 1237
rect 14471 915 14847 949
rect 15089 915 15465 949
rect 14471 657 14847 691
rect 15089 657 15465 691
rect 16071 2061 16447 2095
rect 16689 2061 17065 2095
rect 16071 1203 16447 1237
rect 16689 1203 17065 1237
rect 16071 915 16447 949
rect 16689 915 17065 949
rect 16071 657 16447 691
rect 16689 657 17065 691
rect 17671 2061 18047 2095
rect 18289 2061 18665 2095
rect 17671 1203 18047 1237
rect 18289 1203 18665 1237
rect 17671 915 18047 949
rect 18289 915 18665 949
rect 17671 657 18047 691
rect 18289 657 18665 691
rect 19271 2061 19647 2095
rect 19889 2061 20265 2095
rect 19271 1203 19647 1237
rect 19889 1203 20265 1237
rect 19271 915 19647 949
rect 19889 915 20265 949
rect 19271 657 19647 691
rect 19889 657 20265 691
rect 20871 2061 21247 2095
rect 21489 2061 21865 2095
rect 20871 1203 21247 1237
rect 21489 1203 21865 1237
rect 20871 915 21247 949
rect 21489 915 21865 949
rect 20871 657 21247 691
rect 21489 657 21865 691
rect 22471 2061 22847 2095
rect 23089 2061 23465 2095
rect 22471 1203 22847 1237
rect 23089 1203 23465 1237
rect 22471 915 22847 949
rect 23089 915 23465 949
rect 22471 657 22847 691
rect 23089 657 23465 691
rect 24071 2061 24447 2095
rect 24689 2061 25065 2095
rect 24071 1203 24447 1237
rect 24689 1203 25065 1237
rect 24071 915 24447 949
rect 24689 915 25065 949
rect 24071 657 24447 691
rect 24689 657 25065 691
rect 25671 2061 26047 2095
rect 26289 2061 26665 2095
rect 25671 1203 26047 1237
rect 26289 1203 26665 1237
rect 25671 915 26047 949
rect 26289 915 26665 949
rect 25671 657 26047 691
rect 26289 657 26665 691
rect 27271 2061 27647 2095
rect 27889 2061 28265 2095
rect 27271 1203 27647 1237
rect 27889 1203 28265 1237
rect 27271 915 27647 949
rect 27889 915 28265 949
rect 27271 657 27647 691
rect 27889 657 28265 691
rect 28871 2061 29247 2095
rect 29489 2061 29865 2095
rect 28871 1203 29247 1237
rect 29489 1203 29865 1237
rect 28871 915 29247 949
rect 29489 915 29865 949
rect 28871 657 29247 691
rect 29489 657 29865 691
rect 30471 2061 30847 2095
rect 31089 2061 31465 2095
rect 30471 1203 30847 1237
rect 31089 1203 31465 1237
rect 30471 915 30847 949
rect 31089 915 31465 949
rect 30471 657 30847 691
rect 31089 657 31465 691
rect 32071 2061 32447 2095
rect 32689 2061 33065 2095
rect 32071 1203 32447 1237
rect 32689 1203 33065 1237
rect 32071 915 32447 949
rect 32689 915 33065 949
rect 32071 657 32447 691
rect 32689 657 33065 691
rect 33671 2061 34047 2095
rect 34289 2061 34665 2095
rect 33671 1203 34047 1237
rect 34289 1203 34665 1237
rect 33671 915 34047 949
rect 34289 915 34665 949
rect 33671 657 34047 691
rect 34289 657 34665 691
rect 35271 2061 35647 2095
rect 35889 2061 36265 2095
rect 35271 1203 35647 1237
rect 35889 1203 36265 1237
rect 35271 915 35647 949
rect 35889 915 36265 949
rect 35271 657 35647 691
rect 35889 657 36265 691
rect 36871 2061 37247 2095
rect 37489 2061 37865 2095
rect 36871 1203 37247 1237
rect 37489 1203 37865 1237
rect 36871 915 37247 949
rect 37489 915 37865 949
rect 36871 657 37247 691
rect 37489 657 37865 691
rect 71 261 447 295
rect 689 261 1065 295
rect 71 -597 447 -563
rect 689 -597 1065 -563
rect 71 -885 447 -851
rect 689 -885 1065 -851
rect 71 -1143 447 -1109
rect 689 -1143 1065 -1109
rect 1671 261 2047 295
rect 2289 261 2665 295
rect 1671 -597 2047 -563
rect 2289 -597 2665 -563
rect 1671 -885 2047 -851
rect 2289 -885 2665 -851
rect 1671 -1143 2047 -1109
rect 2289 -1143 2665 -1109
rect 3271 261 3647 295
rect 3889 261 4265 295
rect 3271 -597 3647 -563
rect 3889 -597 4265 -563
rect 3271 -885 3647 -851
rect 3889 -885 4265 -851
rect 3271 -1143 3647 -1109
rect 3889 -1143 4265 -1109
rect 4871 261 5247 295
rect 5489 261 5865 295
rect 4871 -597 5247 -563
rect 5489 -597 5865 -563
rect 4871 -885 5247 -851
rect 5489 -885 5865 -851
rect 4871 -1143 5247 -1109
rect 5489 -1143 5865 -1109
rect 6471 261 6847 295
rect 7089 261 7465 295
rect 6471 -597 6847 -563
rect 7089 -597 7465 -563
rect 6471 -885 6847 -851
rect 7089 -885 7465 -851
rect 6471 -1143 6847 -1109
rect 7089 -1143 7465 -1109
rect 8071 261 8447 295
rect 8689 261 9065 295
rect 8071 -597 8447 -563
rect 8689 -597 9065 -563
rect 8071 -885 8447 -851
rect 8689 -885 9065 -851
rect 8071 -1143 8447 -1109
rect 8689 -1143 9065 -1109
rect 9671 261 10047 295
rect 10289 261 10665 295
rect 9671 -597 10047 -563
rect 10289 -597 10665 -563
rect 9671 -885 10047 -851
rect 10289 -885 10665 -851
rect 9671 -1143 10047 -1109
rect 10289 -1143 10665 -1109
rect 11271 261 11647 295
rect 11889 261 12265 295
rect 11271 -597 11647 -563
rect 11889 -597 12265 -563
rect 11271 -885 11647 -851
rect 11889 -885 12265 -851
rect 11271 -1143 11647 -1109
rect 11889 -1143 12265 -1109
rect 12871 261 13247 295
rect 13489 261 13865 295
rect 12871 -597 13247 -563
rect 13489 -597 13865 -563
rect 12871 -885 13247 -851
rect 13489 -885 13865 -851
rect 12871 -1143 13247 -1109
rect 13489 -1143 13865 -1109
rect 14471 261 14847 295
rect 15089 261 15465 295
rect 14471 -597 14847 -563
rect 15089 -597 15465 -563
rect 14471 -885 14847 -851
rect 15089 -885 15465 -851
rect 14471 -1143 14847 -1109
rect 15089 -1143 15465 -1109
rect 16071 261 16447 295
rect 16689 261 17065 295
rect 16071 -597 16447 -563
rect 16689 -597 17065 -563
rect 16071 -885 16447 -851
rect 16689 -885 17065 -851
rect 16071 -1143 16447 -1109
rect 16689 -1143 17065 -1109
rect 17671 261 18047 295
rect 18289 261 18665 295
rect 17671 -597 18047 -563
rect 18289 -597 18665 -563
rect 17671 -885 18047 -851
rect 18289 -885 18665 -851
rect 17671 -1143 18047 -1109
rect 18289 -1143 18665 -1109
rect 19271 261 19647 295
rect 19889 261 20265 295
rect 19271 -597 19647 -563
rect 19889 -597 20265 -563
rect 19271 -885 19647 -851
rect 19889 -885 20265 -851
rect 19271 -1143 19647 -1109
rect 19889 -1143 20265 -1109
rect 20871 261 21247 295
rect 21489 261 21865 295
rect 20871 -597 21247 -563
rect 21489 -597 21865 -563
rect 20871 -885 21247 -851
rect 21489 -885 21865 -851
rect 20871 -1143 21247 -1109
rect 21489 -1143 21865 -1109
rect 22471 261 22847 295
rect 23089 261 23465 295
rect 22471 -597 22847 -563
rect 23089 -597 23465 -563
rect 22471 -885 22847 -851
rect 23089 -885 23465 -851
rect 22471 -1143 22847 -1109
rect 23089 -1143 23465 -1109
rect 24071 261 24447 295
rect 24689 261 25065 295
rect 24071 -597 24447 -563
rect 24689 -597 25065 -563
rect 24071 -885 24447 -851
rect 24689 -885 25065 -851
rect 24071 -1143 24447 -1109
rect 24689 -1143 25065 -1109
rect 25671 261 26047 295
rect 26289 261 26665 295
rect 25671 -597 26047 -563
rect 26289 -597 26665 -563
rect 25671 -885 26047 -851
rect 26289 -885 26665 -851
rect 25671 -1143 26047 -1109
rect 26289 -1143 26665 -1109
rect 27271 261 27647 295
rect 27889 261 28265 295
rect 27271 -597 27647 -563
rect 27889 -597 28265 -563
rect 27271 -885 27647 -851
rect 27889 -885 28265 -851
rect 27271 -1143 27647 -1109
rect 27889 -1143 28265 -1109
rect 28871 261 29247 295
rect 29489 261 29865 295
rect 28871 -597 29247 -563
rect 29489 -597 29865 -563
rect 28871 -885 29247 -851
rect 29489 -885 29865 -851
rect 28871 -1143 29247 -1109
rect 29489 -1143 29865 -1109
rect 30471 261 30847 295
rect 31089 261 31465 295
rect 30471 -597 30847 -563
rect 31089 -597 31465 -563
rect 30471 -885 30847 -851
rect 31089 -885 31465 -851
rect 30471 -1143 30847 -1109
rect 31089 -1143 31465 -1109
rect 32071 261 32447 295
rect 32689 261 33065 295
rect 32071 -597 32447 -563
rect 32689 -597 33065 -563
rect 32071 -885 32447 -851
rect 32689 -885 33065 -851
rect 32071 -1143 32447 -1109
rect 32689 -1143 33065 -1109
rect 33671 261 34047 295
rect 34289 261 34665 295
rect 33671 -597 34047 -563
rect 34289 -597 34665 -563
rect 33671 -885 34047 -851
rect 34289 -885 34665 -851
rect 33671 -1143 34047 -1109
rect 34289 -1143 34665 -1109
rect 35271 261 35647 295
rect 35889 261 36265 295
rect 35271 -597 35647 -563
rect 35889 -597 36265 -563
rect 35271 -885 35647 -851
rect 35889 -885 36265 -851
rect 35271 -1143 35647 -1109
rect 35889 -1143 36265 -1109
rect 36871 261 37247 295
rect 37489 261 37865 295
rect 36871 -597 37247 -563
rect 37489 -597 37865 -563
rect 36871 -885 37247 -851
rect 37489 -885 37865 -851
rect 36871 -1143 37247 -1109
rect 37489 -1143 37865 -1109
rect 71 -1539 447 -1505
rect 689 -1539 1065 -1505
rect 71 -2397 447 -2363
rect 689 -2397 1065 -2363
rect 71 -2685 447 -2651
rect 689 -2685 1065 -2651
rect 71 -2943 447 -2909
rect 689 -2943 1065 -2909
rect 1671 -1539 2047 -1505
rect 2289 -1539 2665 -1505
rect 1671 -2397 2047 -2363
rect 2289 -2397 2665 -2363
rect 1671 -2685 2047 -2651
rect 2289 -2685 2665 -2651
rect 1671 -2943 2047 -2909
rect 2289 -2943 2665 -2909
rect 3271 -1539 3647 -1505
rect 3889 -1539 4265 -1505
rect 3271 -2397 3647 -2363
rect 3889 -2397 4265 -2363
rect 3271 -2685 3647 -2651
rect 3889 -2685 4265 -2651
rect 3271 -2943 3647 -2909
rect 3889 -2943 4265 -2909
rect 4871 -1539 5247 -1505
rect 5489 -1539 5865 -1505
rect 4871 -2397 5247 -2363
rect 5489 -2397 5865 -2363
rect 4871 -2685 5247 -2651
rect 5489 -2685 5865 -2651
rect 4871 -2943 5247 -2909
rect 5489 -2943 5865 -2909
rect 6471 -1539 6847 -1505
rect 7089 -1539 7465 -1505
rect 6471 -2397 6847 -2363
rect 7089 -2397 7465 -2363
rect 6471 -2685 6847 -2651
rect 7089 -2685 7465 -2651
rect 6471 -2943 6847 -2909
rect 7089 -2943 7465 -2909
rect 8071 -1539 8447 -1505
rect 8689 -1539 9065 -1505
rect 8071 -2397 8447 -2363
rect 8689 -2397 9065 -2363
rect 8071 -2685 8447 -2651
rect 8689 -2685 9065 -2651
rect 8071 -2943 8447 -2909
rect 8689 -2943 9065 -2909
rect 9671 -1539 10047 -1505
rect 10289 -1539 10665 -1505
rect 9671 -2397 10047 -2363
rect 10289 -2397 10665 -2363
rect 9671 -2685 10047 -2651
rect 10289 -2685 10665 -2651
rect 9671 -2943 10047 -2909
rect 10289 -2943 10665 -2909
rect 11271 -1539 11647 -1505
rect 11889 -1539 12265 -1505
rect 11271 -2397 11647 -2363
rect 11889 -2397 12265 -2363
rect 11271 -2685 11647 -2651
rect 11889 -2685 12265 -2651
rect 11271 -2943 11647 -2909
rect 11889 -2943 12265 -2909
rect 12871 -1539 13247 -1505
rect 13489 -1539 13865 -1505
rect 12871 -2397 13247 -2363
rect 13489 -2397 13865 -2363
rect 12871 -2685 13247 -2651
rect 13489 -2685 13865 -2651
rect 12871 -2943 13247 -2909
rect 13489 -2943 13865 -2909
rect 14471 -1539 14847 -1505
rect 15089 -1539 15465 -1505
rect 14471 -2397 14847 -2363
rect 15089 -2397 15465 -2363
rect 14471 -2685 14847 -2651
rect 15089 -2685 15465 -2651
rect 14471 -2943 14847 -2909
rect 15089 -2943 15465 -2909
rect 16071 -1539 16447 -1505
rect 16689 -1539 17065 -1505
rect 16071 -2397 16447 -2363
rect 16689 -2397 17065 -2363
rect 16071 -2685 16447 -2651
rect 16689 -2685 17065 -2651
rect 16071 -2943 16447 -2909
rect 16689 -2943 17065 -2909
rect 17671 -1539 18047 -1505
rect 18289 -1539 18665 -1505
rect 17671 -2397 18047 -2363
rect 18289 -2397 18665 -2363
rect 17671 -2685 18047 -2651
rect 18289 -2685 18665 -2651
rect 17671 -2943 18047 -2909
rect 18289 -2943 18665 -2909
rect 19271 -1539 19647 -1505
rect 19889 -1539 20265 -1505
rect 19271 -2397 19647 -2363
rect 19889 -2397 20265 -2363
rect 19271 -2685 19647 -2651
rect 19889 -2685 20265 -2651
rect 19271 -2943 19647 -2909
rect 19889 -2943 20265 -2909
rect 20871 -1539 21247 -1505
rect 21489 -1539 21865 -1505
rect 20871 -2397 21247 -2363
rect 21489 -2397 21865 -2363
rect 20871 -2685 21247 -2651
rect 21489 -2685 21865 -2651
rect 20871 -2943 21247 -2909
rect 21489 -2943 21865 -2909
rect 22471 -1539 22847 -1505
rect 23089 -1539 23465 -1505
rect 22471 -2397 22847 -2363
rect 23089 -2397 23465 -2363
rect 22471 -2685 22847 -2651
rect 23089 -2685 23465 -2651
rect 22471 -2943 22847 -2909
rect 23089 -2943 23465 -2909
rect 24071 -1539 24447 -1505
rect 24689 -1539 25065 -1505
rect 24071 -2397 24447 -2363
rect 24689 -2397 25065 -2363
rect 24071 -2685 24447 -2651
rect 24689 -2685 25065 -2651
rect 24071 -2943 24447 -2909
rect 24689 -2943 25065 -2909
rect 25671 -1539 26047 -1505
rect 26289 -1539 26665 -1505
rect 25671 -2397 26047 -2363
rect 26289 -2397 26665 -2363
rect 25671 -2685 26047 -2651
rect 26289 -2685 26665 -2651
rect 25671 -2943 26047 -2909
rect 26289 -2943 26665 -2909
rect 27271 -1539 27647 -1505
rect 27889 -1539 28265 -1505
rect 27271 -2397 27647 -2363
rect 27889 -2397 28265 -2363
rect 27271 -2685 27647 -2651
rect 27889 -2685 28265 -2651
rect 27271 -2943 27647 -2909
rect 27889 -2943 28265 -2909
rect 28871 -1539 29247 -1505
rect 29489 -1539 29865 -1505
rect 28871 -2397 29247 -2363
rect 29489 -2397 29865 -2363
rect 28871 -2685 29247 -2651
rect 29489 -2685 29865 -2651
rect 28871 -2943 29247 -2909
rect 29489 -2943 29865 -2909
rect 30471 -1539 30847 -1505
rect 31089 -1539 31465 -1505
rect 30471 -2397 30847 -2363
rect 31089 -2397 31465 -2363
rect 30471 -2685 30847 -2651
rect 31089 -2685 31465 -2651
rect 30471 -2943 30847 -2909
rect 31089 -2943 31465 -2909
rect 32071 -1539 32447 -1505
rect 32689 -1539 33065 -1505
rect 32071 -2397 32447 -2363
rect 32689 -2397 33065 -2363
rect 32071 -2685 32447 -2651
rect 32689 -2685 33065 -2651
rect 32071 -2943 32447 -2909
rect 32689 -2943 33065 -2909
rect 33671 -1539 34047 -1505
rect 34289 -1539 34665 -1505
rect 33671 -2397 34047 -2363
rect 34289 -2397 34665 -2363
rect 33671 -2685 34047 -2651
rect 34289 -2685 34665 -2651
rect 33671 -2943 34047 -2909
rect 34289 -2943 34665 -2909
rect 35271 -1539 35647 -1505
rect 35889 -1539 36265 -1505
rect 35271 -2397 35647 -2363
rect 35889 -2397 36265 -2363
rect 35271 -2685 35647 -2651
rect 35889 -2685 36265 -2651
rect 35271 -2943 35647 -2909
rect 35889 -2943 36265 -2909
rect 36871 -1539 37247 -1505
rect 37489 -1539 37865 -1505
rect 36871 -2397 37247 -2363
rect 37489 -2397 37865 -2363
rect 36871 -2685 37247 -2651
rect 37489 -2685 37865 -2651
rect 36871 -2943 37247 -2909
rect 37489 -2943 37865 -2909
rect 71 -3339 447 -3305
rect 689 -3339 1065 -3305
rect 71 -4197 447 -4163
rect 689 -4197 1065 -4163
rect 71 -4485 447 -4451
rect 689 -4485 1065 -4451
rect 71 -4743 447 -4709
rect 689 -4743 1065 -4709
rect 1671 -3339 2047 -3305
rect 2289 -3339 2665 -3305
rect 1671 -4197 2047 -4163
rect 2289 -4197 2665 -4163
rect 1671 -4485 2047 -4451
rect 2289 -4485 2665 -4451
rect 1671 -4743 2047 -4709
rect 2289 -4743 2665 -4709
rect 3271 -3339 3647 -3305
rect 3889 -3339 4265 -3305
rect 3271 -4197 3647 -4163
rect 3889 -4197 4265 -4163
rect 3271 -4485 3647 -4451
rect 3889 -4485 4265 -4451
rect 3271 -4743 3647 -4709
rect 3889 -4743 4265 -4709
rect 4871 -3339 5247 -3305
rect 5489 -3339 5865 -3305
rect 4871 -4197 5247 -4163
rect 5489 -4197 5865 -4163
rect 4871 -4485 5247 -4451
rect 5489 -4485 5865 -4451
rect 4871 -4743 5247 -4709
rect 5489 -4743 5865 -4709
rect 6471 -3339 6847 -3305
rect 7089 -3339 7465 -3305
rect 6471 -4197 6847 -4163
rect 7089 -4197 7465 -4163
rect 6471 -4485 6847 -4451
rect 7089 -4485 7465 -4451
rect 6471 -4743 6847 -4709
rect 7089 -4743 7465 -4709
rect 8071 -3339 8447 -3305
rect 8689 -3339 9065 -3305
rect 8071 -4197 8447 -4163
rect 8689 -4197 9065 -4163
rect 8071 -4485 8447 -4451
rect 8689 -4485 9065 -4451
rect 8071 -4743 8447 -4709
rect 8689 -4743 9065 -4709
rect 9671 -3339 10047 -3305
rect 10289 -3339 10665 -3305
rect 9671 -4197 10047 -4163
rect 10289 -4197 10665 -4163
rect 9671 -4485 10047 -4451
rect 10289 -4485 10665 -4451
rect 9671 -4743 10047 -4709
rect 10289 -4743 10665 -4709
rect 11271 -3339 11647 -3305
rect 11889 -3339 12265 -3305
rect 11271 -4197 11647 -4163
rect 11889 -4197 12265 -4163
rect 11271 -4485 11647 -4451
rect 11889 -4485 12265 -4451
rect 11271 -4743 11647 -4709
rect 11889 -4743 12265 -4709
rect 12871 -3339 13247 -3305
rect 13489 -3339 13865 -3305
rect 12871 -4197 13247 -4163
rect 13489 -4197 13865 -4163
rect 12871 -4485 13247 -4451
rect 13489 -4485 13865 -4451
rect 12871 -4743 13247 -4709
rect 13489 -4743 13865 -4709
rect 14471 -3339 14847 -3305
rect 15089 -3339 15465 -3305
rect 14471 -4197 14847 -4163
rect 15089 -4197 15465 -4163
rect 14471 -4485 14847 -4451
rect 15089 -4485 15465 -4451
rect 14471 -4743 14847 -4709
rect 15089 -4743 15465 -4709
rect 16071 -3339 16447 -3305
rect 16689 -3339 17065 -3305
rect 16071 -4197 16447 -4163
rect 16689 -4197 17065 -4163
rect 16071 -4485 16447 -4451
rect 16689 -4485 17065 -4451
rect 16071 -4743 16447 -4709
rect 16689 -4743 17065 -4709
rect 17671 -3339 18047 -3305
rect 18289 -3339 18665 -3305
rect 17671 -4197 18047 -4163
rect 18289 -4197 18665 -4163
rect 17671 -4485 18047 -4451
rect 18289 -4485 18665 -4451
rect 17671 -4743 18047 -4709
rect 18289 -4743 18665 -4709
rect 19271 -3339 19647 -3305
rect 19889 -3339 20265 -3305
rect 19271 -4197 19647 -4163
rect 19889 -4197 20265 -4163
rect 19271 -4485 19647 -4451
rect 19889 -4485 20265 -4451
rect 19271 -4743 19647 -4709
rect 19889 -4743 20265 -4709
rect 20871 -3339 21247 -3305
rect 21489 -3339 21865 -3305
rect 20871 -4197 21247 -4163
rect 21489 -4197 21865 -4163
rect 20871 -4485 21247 -4451
rect 21489 -4485 21865 -4451
rect 20871 -4743 21247 -4709
rect 21489 -4743 21865 -4709
rect 22471 -3339 22847 -3305
rect 23089 -3339 23465 -3305
rect 22471 -4197 22847 -4163
rect 23089 -4197 23465 -4163
rect 22471 -4485 22847 -4451
rect 23089 -4485 23465 -4451
rect 22471 -4743 22847 -4709
rect 23089 -4743 23465 -4709
rect 24071 -3339 24447 -3305
rect 24689 -3339 25065 -3305
rect 24071 -4197 24447 -4163
rect 24689 -4197 25065 -4163
rect 24071 -4485 24447 -4451
rect 24689 -4485 25065 -4451
rect 24071 -4743 24447 -4709
rect 24689 -4743 25065 -4709
rect 25671 -3339 26047 -3305
rect 26289 -3339 26665 -3305
rect 25671 -4197 26047 -4163
rect 26289 -4197 26665 -4163
rect 25671 -4485 26047 -4451
rect 26289 -4485 26665 -4451
rect 25671 -4743 26047 -4709
rect 26289 -4743 26665 -4709
rect 27271 -3339 27647 -3305
rect 27889 -3339 28265 -3305
rect 27271 -4197 27647 -4163
rect 27889 -4197 28265 -4163
rect 27271 -4485 27647 -4451
rect 27889 -4485 28265 -4451
rect 27271 -4743 27647 -4709
rect 27889 -4743 28265 -4709
rect 28871 -3339 29247 -3305
rect 29489 -3339 29865 -3305
rect 28871 -4197 29247 -4163
rect 29489 -4197 29865 -4163
rect 28871 -4485 29247 -4451
rect 29489 -4485 29865 -4451
rect 28871 -4743 29247 -4709
rect 29489 -4743 29865 -4709
rect 30471 -3339 30847 -3305
rect 31089 -3339 31465 -3305
rect 30471 -4197 30847 -4163
rect 31089 -4197 31465 -4163
rect 30471 -4485 30847 -4451
rect 31089 -4485 31465 -4451
rect 30471 -4743 30847 -4709
rect 31089 -4743 31465 -4709
rect 32071 -3339 32447 -3305
rect 32689 -3339 33065 -3305
rect 32071 -4197 32447 -4163
rect 32689 -4197 33065 -4163
rect 32071 -4485 32447 -4451
rect 32689 -4485 33065 -4451
rect 32071 -4743 32447 -4709
rect 32689 -4743 33065 -4709
rect 33671 -3339 34047 -3305
rect 34289 -3339 34665 -3305
rect 33671 -4197 34047 -4163
rect 34289 -4197 34665 -4163
rect 33671 -4485 34047 -4451
rect 34289 -4485 34665 -4451
rect 33671 -4743 34047 -4709
rect 34289 -4743 34665 -4709
rect 35271 -3339 35647 -3305
rect 35889 -3339 36265 -3305
rect 35271 -4197 35647 -4163
rect 35889 -4197 36265 -4163
rect 35271 -4485 35647 -4451
rect 35889 -4485 36265 -4451
rect 35271 -4743 35647 -4709
rect 35889 -4743 36265 -4709
rect 36871 -3339 37247 -3305
rect 37489 -3339 37865 -3305
rect 36871 -4197 37247 -4163
rect 37489 -4197 37865 -4163
rect 36871 -4485 37247 -4451
rect 37489 -4485 37865 -4451
rect 36871 -4743 37247 -4709
rect 37489 -4743 37865 -4709
rect 27922 -25100 27956 -24724
rect 28780 -25100 28814 -24724
rect 27948 -25576 28724 -25542
rect 27948 -25734 28724 -25700
rect 27948 -25892 28724 -25858
rect 27948 -26050 28724 -26016
rect 27948 -26208 28724 -26174
rect 27948 -26616 28724 -26582
rect 27948 -26774 28724 -26740
rect 27948 -26932 28724 -26898
rect 27948 -27090 28724 -27056
rect 27948 -27248 28724 -27214
rect 27948 -27656 28724 -27622
rect 27948 -27814 28724 -27780
rect 27948 -27972 28724 -27938
rect 27948 -28130 28724 -28096
rect 27948 -28288 28724 -28254
rect 27948 -28696 28724 -28662
rect 27948 -28854 28724 -28820
rect 27948 -29012 28724 -28978
rect 27948 -29170 28724 -29136
rect 27948 -29328 28724 -29294
rect 27948 -29736 28724 -29702
rect 27948 -29894 28724 -29860
rect 27948 -30052 28724 -30018
rect 27948 -30210 28724 -30176
rect 27948 -30368 28724 -30334
rect 31813 -29729 31847 -29553
rect 31971 -29729 32005 -29553
rect 32253 -29729 32287 -29553
rect 32411 -29729 32445 -29553
rect 32693 -29729 32727 -29553
rect 32851 -29729 32885 -29553
rect 33132 -29729 33166 -29553
rect 33290 -29729 33324 -29553
rect 33448 -29729 33482 -29553
rect 33606 -29729 33640 -29553
rect 34013 -29729 34047 -29553
rect 34171 -29729 34205 -29553
rect 34453 -29729 34487 -29553
rect 34611 -29729 34645 -29553
rect 34893 -29729 34927 -29553
rect 35051 -29729 35085 -29553
rect 35332 -29729 35366 -29553
rect 35490 -29729 35524 -29553
rect 35648 -29729 35682 -29553
rect 35806 -29729 35840 -29553
rect 36213 -29729 36247 -29553
rect 36371 -29729 36405 -29553
rect 36653 -29729 36687 -29553
rect 36811 -29729 36845 -29553
rect 37093 -29729 37127 -29553
rect 37251 -29729 37285 -29553
rect 37532 -29729 37566 -29553
rect 37690 -29729 37724 -29553
rect 37848 -29729 37882 -29553
rect 38006 -29729 38040 -29553
rect 27948 -30776 28724 -30742
rect 27948 -30934 28724 -30900
rect 27948 -31092 28724 -31058
rect 27948 -31250 28724 -31216
rect 27948 -31408 28724 -31374
rect 31782 -30471 31816 -30295
rect 31940 -30471 31974 -30295
rect 32098 -30471 32132 -30295
rect 32256 -30471 32290 -30295
rect 32537 -30471 32571 -30295
rect 32695 -30471 32729 -30295
rect 32977 -30471 33011 -30295
rect 33135 -30471 33169 -30295
rect 33417 -30471 33451 -30295
rect 33575 -30471 33609 -30295
rect 33982 -30471 34016 -30295
rect 34140 -30471 34174 -30295
rect 34298 -30471 34332 -30295
rect 34456 -30471 34490 -30295
rect 34737 -30471 34771 -30295
rect 34895 -30471 34929 -30295
rect 35177 -30471 35211 -30295
rect 35335 -30471 35369 -30295
rect 35617 -30471 35651 -30295
rect 35775 -30471 35809 -30295
rect 36182 -30471 36216 -30295
rect 36340 -30471 36374 -30295
rect 36498 -30471 36532 -30295
rect 36656 -30471 36690 -30295
rect 36937 -30471 36971 -30295
rect 37095 -30471 37129 -30295
rect 37377 -30471 37411 -30295
rect 37535 -30471 37569 -30295
rect 37817 -30471 37851 -30295
rect 37975 -30471 38009 -30295
<< mvpdiffc >>
rect 27938 11424 28714 11458
rect 27938 11266 28714 11300
rect 27938 11108 28714 11142
rect 27938 10950 28714 10984
rect 27938 10792 28714 10826
rect 30144 10819 30178 10895
rect 30602 10819 30636 10895
rect 27938 10384 28714 10418
rect 27938 10226 28714 10260
rect 27938 10068 28714 10102
rect 27938 9910 28714 9944
rect 27938 9752 28714 9786
rect 30858 10519 30892 10895
rect 31016 10519 31050 10895
rect 31298 10519 31332 10895
rect 31456 10519 31490 10895
rect 31738 10519 31772 10895
rect 31896 10519 31930 10895
rect 32344 10819 32378 10895
rect 32802 10819 32836 10895
rect 33058 10519 33092 10895
rect 33216 10519 33250 10895
rect 33498 10519 33532 10895
rect 33656 10519 33690 10895
rect 33938 10519 33972 10895
rect 34096 10519 34130 10895
rect 34544 10819 34578 10895
rect 35002 10819 35036 10895
rect 35258 10519 35292 10895
rect 35416 10519 35450 10895
rect 35698 10519 35732 10895
rect 35856 10519 35890 10895
rect 36138 10519 36172 10895
rect 36296 10519 36330 10895
rect 27938 9344 28714 9378
rect 27938 9186 28714 9220
rect 27938 9028 28714 9062
rect 27938 8870 28714 8904
rect 27938 8712 28714 8746
rect 29732 9209 29766 9585
rect 30590 9209 30624 9585
rect 31448 9209 31482 9585
rect 27938 8304 28714 8338
rect 27938 8146 28714 8180
rect 27938 7988 28714 8022
rect 27938 7830 28714 7864
rect 27938 7672 28714 7706
rect 27938 7264 28714 7298
rect 27938 7106 28714 7140
rect 27938 6948 28714 6982
rect 27938 6790 28714 6824
rect 27938 6632 28714 6666
rect 29732 8205 29766 8581
rect 30590 8205 30624 8581
rect 31448 8205 31482 8581
rect 29732 7569 29766 7945
rect 30590 7569 30624 7945
rect 31448 7569 31482 7945
rect 29769 7030 30545 7064
rect 29769 6772 30545 6806
rect 31109 7030 31885 7064
rect 31109 6772 31885 6806
rect 27938 6224 28714 6258
rect 27938 6066 28714 6100
rect 27938 5908 28714 5942
rect 27938 5750 28714 5784
rect 27938 5592 28714 5626
rect 27912 4369 27946 5145
rect 28770 4369 28804 5145
rect 69 -8204 445 -8170
rect 705 -8204 1081 -8170
rect 69 -8462 445 -8428
rect 705 -8462 1081 -8428
rect 69 -8730 445 -8696
rect 705 -8730 1081 -8696
rect 69 -9588 445 -9554
rect 705 -9588 1081 -9554
rect 1669 -8204 2045 -8170
rect 2305 -8204 2681 -8170
rect 1669 -8462 2045 -8428
rect 2305 -8462 2681 -8428
rect 1669 -8730 2045 -8696
rect 2305 -8730 2681 -8696
rect 1669 -9588 2045 -9554
rect 2305 -9588 2681 -9554
rect 3269 -8204 3645 -8170
rect 3905 -8204 4281 -8170
rect 3269 -8462 3645 -8428
rect 3905 -8462 4281 -8428
rect 3269 -8730 3645 -8696
rect 3905 -8730 4281 -8696
rect 3269 -9588 3645 -9554
rect 3905 -9588 4281 -9554
rect 4869 -8204 5245 -8170
rect 5505 -8204 5881 -8170
rect 4869 -8462 5245 -8428
rect 5505 -8462 5881 -8428
rect 4869 -8730 5245 -8696
rect 5505 -8730 5881 -8696
rect 4869 -9588 5245 -9554
rect 5505 -9588 5881 -9554
rect 6469 -8204 6845 -8170
rect 7105 -8204 7481 -8170
rect 6469 -8462 6845 -8428
rect 7105 -8462 7481 -8428
rect 6469 -8730 6845 -8696
rect 7105 -8730 7481 -8696
rect 6469 -9588 6845 -9554
rect 7105 -9588 7481 -9554
rect 8069 -8204 8445 -8170
rect 8705 -8204 9081 -8170
rect 8069 -8462 8445 -8428
rect 8705 -8462 9081 -8428
rect 8069 -8730 8445 -8696
rect 8705 -8730 9081 -8696
rect 8069 -9588 8445 -9554
rect 8705 -9588 9081 -9554
rect 9669 -8204 10045 -8170
rect 10305 -8204 10681 -8170
rect 9669 -8462 10045 -8428
rect 10305 -8462 10681 -8428
rect 9669 -8730 10045 -8696
rect 10305 -8730 10681 -8696
rect 9669 -9588 10045 -9554
rect 10305 -9588 10681 -9554
rect 11269 -8204 11645 -8170
rect 11905 -8204 12281 -8170
rect 11269 -8462 11645 -8428
rect 11905 -8462 12281 -8428
rect 11269 -8730 11645 -8696
rect 11905 -8730 12281 -8696
rect 11269 -9588 11645 -9554
rect 11905 -9588 12281 -9554
rect 12869 -8204 13245 -8170
rect 13505 -8204 13881 -8170
rect 12869 -8462 13245 -8428
rect 13505 -8462 13881 -8428
rect 12869 -8730 13245 -8696
rect 13505 -8730 13881 -8696
rect 12869 -9588 13245 -9554
rect 13505 -9588 13881 -9554
rect 14469 -8204 14845 -8170
rect 15105 -8204 15481 -8170
rect 14469 -8462 14845 -8428
rect 15105 -8462 15481 -8428
rect 14469 -8730 14845 -8696
rect 15105 -8730 15481 -8696
rect 14469 -9588 14845 -9554
rect 15105 -9588 15481 -9554
rect 16069 -8204 16445 -8170
rect 16705 -8204 17081 -8170
rect 16069 -8462 16445 -8428
rect 16705 -8462 17081 -8428
rect 16069 -8730 16445 -8696
rect 16705 -8730 17081 -8696
rect 16069 -9588 16445 -9554
rect 16705 -9588 17081 -9554
rect 17669 -8204 18045 -8170
rect 18305 -8204 18681 -8170
rect 17669 -8462 18045 -8428
rect 18305 -8462 18681 -8428
rect 17669 -8730 18045 -8696
rect 18305 -8730 18681 -8696
rect 17669 -9588 18045 -9554
rect 18305 -9588 18681 -9554
rect 19269 -8204 19645 -8170
rect 19905 -8204 20281 -8170
rect 19269 -8462 19645 -8428
rect 19905 -8462 20281 -8428
rect 19269 -8730 19645 -8696
rect 19905 -8730 20281 -8696
rect 19269 -9588 19645 -9554
rect 19905 -9588 20281 -9554
rect 20869 -8204 21245 -8170
rect 21505 -8204 21881 -8170
rect 20869 -8462 21245 -8428
rect 21505 -8462 21881 -8428
rect 20869 -8730 21245 -8696
rect 21505 -8730 21881 -8696
rect 20869 -9588 21245 -9554
rect 21505 -9588 21881 -9554
rect 22469 -8204 22845 -8170
rect 23105 -8204 23481 -8170
rect 22469 -8462 22845 -8428
rect 23105 -8462 23481 -8428
rect 22469 -8730 22845 -8696
rect 23105 -8730 23481 -8696
rect 22469 -9588 22845 -9554
rect 23105 -9588 23481 -9554
rect 24069 -8204 24445 -8170
rect 24705 -8204 25081 -8170
rect 24069 -8462 24445 -8428
rect 24705 -8462 25081 -8428
rect 24069 -8730 24445 -8696
rect 24705 -8730 25081 -8696
rect 24069 -9588 24445 -9554
rect 24705 -9588 25081 -9554
rect 25669 -8204 26045 -8170
rect 26305 -8204 26681 -8170
rect 25669 -8462 26045 -8428
rect 26305 -8462 26681 -8428
rect 25669 -8730 26045 -8696
rect 26305 -8730 26681 -8696
rect 25669 -9588 26045 -9554
rect 26305 -9588 26681 -9554
rect 27269 -8204 27645 -8170
rect 27905 -8204 28281 -8170
rect 27269 -8462 27645 -8428
rect 27905 -8462 28281 -8428
rect 27269 -8730 27645 -8696
rect 27905 -8730 28281 -8696
rect 27269 -9588 27645 -9554
rect 27905 -9588 28281 -9554
rect 28869 -8204 29245 -8170
rect 29505 -8204 29881 -8170
rect 28869 -8462 29245 -8428
rect 29505 -8462 29881 -8428
rect 28869 -8730 29245 -8696
rect 29505 -8730 29881 -8696
rect 28869 -9588 29245 -9554
rect 29505 -9588 29881 -9554
rect 30469 -8204 30845 -8170
rect 31105 -8204 31481 -8170
rect 30469 -8462 30845 -8428
rect 31105 -8462 31481 -8428
rect 30469 -8730 30845 -8696
rect 31105 -8730 31481 -8696
rect 30469 -9588 30845 -9554
rect 31105 -9588 31481 -9554
rect 32069 -8204 32445 -8170
rect 32705 -8204 33081 -8170
rect 32069 -8462 32445 -8428
rect 32705 -8462 33081 -8428
rect 32069 -8730 32445 -8696
rect 32705 -8730 33081 -8696
rect 32069 -9588 32445 -9554
rect 32705 -9588 33081 -9554
rect 33669 -8204 34045 -8170
rect 34305 -8204 34681 -8170
rect 33669 -8462 34045 -8428
rect 34305 -8462 34681 -8428
rect 33669 -8730 34045 -8696
rect 34305 -8730 34681 -8696
rect 33669 -9588 34045 -9554
rect 34305 -9588 34681 -9554
rect 35269 -8204 35645 -8170
rect 35905 -8204 36281 -8170
rect 35269 -8462 35645 -8428
rect 35905 -8462 36281 -8428
rect 35269 -8730 35645 -8696
rect 35905 -8730 36281 -8696
rect 35269 -9588 35645 -9554
rect 35905 -9588 36281 -9554
rect 36869 -8204 37245 -8170
rect 37505 -8204 37881 -8170
rect 36869 -8462 37245 -8428
rect 37505 -8462 37881 -8428
rect 36869 -8730 37245 -8696
rect 37505 -8730 37881 -8696
rect 36869 -9588 37245 -9554
rect 37505 -9588 37881 -9554
rect 69 -10004 445 -9970
rect 705 -10004 1081 -9970
rect 69 -10262 445 -10228
rect 705 -10262 1081 -10228
rect 69 -10530 445 -10496
rect 705 -10530 1081 -10496
rect 69 -11388 445 -11354
rect 705 -11388 1081 -11354
rect 1669 -10004 2045 -9970
rect 2305 -10004 2681 -9970
rect 1669 -10262 2045 -10228
rect 2305 -10262 2681 -10228
rect 1669 -10530 2045 -10496
rect 2305 -10530 2681 -10496
rect 1669 -11388 2045 -11354
rect 2305 -11388 2681 -11354
rect 3269 -10004 3645 -9970
rect 3905 -10004 4281 -9970
rect 3269 -10262 3645 -10228
rect 3905 -10262 4281 -10228
rect 3269 -10530 3645 -10496
rect 3905 -10530 4281 -10496
rect 3269 -11388 3645 -11354
rect 3905 -11388 4281 -11354
rect 4869 -10004 5245 -9970
rect 5505 -10004 5881 -9970
rect 4869 -10262 5245 -10228
rect 5505 -10262 5881 -10228
rect 4869 -10530 5245 -10496
rect 5505 -10530 5881 -10496
rect 4869 -11388 5245 -11354
rect 5505 -11388 5881 -11354
rect 6469 -10004 6845 -9970
rect 7105 -10004 7481 -9970
rect 6469 -10262 6845 -10228
rect 7105 -10262 7481 -10228
rect 6469 -10530 6845 -10496
rect 7105 -10530 7481 -10496
rect 6469 -11388 6845 -11354
rect 7105 -11388 7481 -11354
rect 8069 -10004 8445 -9970
rect 8705 -10004 9081 -9970
rect 8069 -10262 8445 -10228
rect 8705 -10262 9081 -10228
rect 8069 -10530 8445 -10496
rect 8705 -10530 9081 -10496
rect 8069 -11388 8445 -11354
rect 8705 -11388 9081 -11354
rect 9669 -10004 10045 -9970
rect 10305 -10004 10681 -9970
rect 9669 -10262 10045 -10228
rect 10305 -10262 10681 -10228
rect 9669 -10530 10045 -10496
rect 10305 -10530 10681 -10496
rect 9669 -11388 10045 -11354
rect 10305 -11388 10681 -11354
rect 11269 -10004 11645 -9970
rect 11905 -10004 12281 -9970
rect 11269 -10262 11645 -10228
rect 11905 -10262 12281 -10228
rect 11269 -10530 11645 -10496
rect 11905 -10530 12281 -10496
rect 11269 -11388 11645 -11354
rect 11905 -11388 12281 -11354
rect 12869 -10004 13245 -9970
rect 13505 -10004 13881 -9970
rect 12869 -10262 13245 -10228
rect 13505 -10262 13881 -10228
rect 12869 -10530 13245 -10496
rect 13505 -10530 13881 -10496
rect 12869 -11388 13245 -11354
rect 13505 -11388 13881 -11354
rect 14469 -10004 14845 -9970
rect 15105 -10004 15481 -9970
rect 14469 -10262 14845 -10228
rect 15105 -10262 15481 -10228
rect 14469 -10530 14845 -10496
rect 15105 -10530 15481 -10496
rect 14469 -11388 14845 -11354
rect 15105 -11388 15481 -11354
rect 16069 -10004 16445 -9970
rect 16705 -10004 17081 -9970
rect 16069 -10262 16445 -10228
rect 16705 -10262 17081 -10228
rect 16069 -10530 16445 -10496
rect 16705 -10530 17081 -10496
rect 16069 -11388 16445 -11354
rect 16705 -11388 17081 -11354
rect 17669 -10004 18045 -9970
rect 18305 -10004 18681 -9970
rect 17669 -10262 18045 -10228
rect 18305 -10262 18681 -10228
rect 17669 -10530 18045 -10496
rect 18305 -10530 18681 -10496
rect 17669 -11388 18045 -11354
rect 18305 -11388 18681 -11354
rect 19269 -10004 19645 -9970
rect 19905 -10004 20281 -9970
rect 19269 -10262 19645 -10228
rect 19905 -10262 20281 -10228
rect 19269 -10530 19645 -10496
rect 19905 -10530 20281 -10496
rect 19269 -11388 19645 -11354
rect 19905 -11388 20281 -11354
rect 20869 -10004 21245 -9970
rect 21505 -10004 21881 -9970
rect 20869 -10262 21245 -10228
rect 21505 -10262 21881 -10228
rect 20869 -10530 21245 -10496
rect 21505 -10530 21881 -10496
rect 20869 -11388 21245 -11354
rect 21505 -11388 21881 -11354
rect 22469 -10004 22845 -9970
rect 23105 -10004 23481 -9970
rect 22469 -10262 22845 -10228
rect 23105 -10262 23481 -10228
rect 22469 -10530 22845 -10496
rect 23105 -10530 23481 -10496
rect 22469 -11388 22845 -11354
rect 23105 -11388 23481 -11354
rect 24069 -10004 24445 -9970
rect 24705 -10004 25081 -9970
rect 24069 -10262 24445 -10228
rect 24705 -10262 25081 -10228
rect 24069 -10530 24445 -10496
rect 24705 -10530 25081 -10496
rect 24069 -11388 24445 -11354
rect 24705 -11388 25081 -11354
rect 25669 -10004 26045 -9970
rect 26305 -10004 26681 -9970
rect 25669 -10262 26045 -10228
rect 26305 -10262 26681 -10228
rect 25669 -10530 26045 -10496
rect 26305 -10530 26681 -10496
rect 25669 -11388 26045 -11354
rect 26305 -11388 26681 -11354
rect 27269 -10004 27645 -9970
rect 27905 -10004 28281 -9970
rect 27269 -10262 27645 -10228
rect 27905 -10262 28281 -10228
rect 27269 -10530 27645 -10496
rect 27905 -10530 28281 -10496
rect 27269 -11388 27645 -11354
rect 27905 -11388 28281 -11354
rect 28869 -10004 29245 -9970
rect 29505 -10004 29881 -9970
rect 28869 -10262 29245 -10228
rect 29505 -10262 29881 -10228
rect 28869 -10530 29245 -10496
rect 29505 -10530 29881 -10496
rect 28869 -11388 29245 -11354
rect 29505 -11388 29881 -11354
rect 30469 -10004 30845 -9970
rect 31105 -10004 31481 -9970
rect 30469 -10262 30845 -10228
rect 31105 -10262 31481 -10228
rect 30469 -10530 30845 -10496
rect 31105 -10530 31481 -10496
rect 30469 -11388 30845 -11354
rect 31105 -11388 31481 -11354
rect 32069 -10004 32445 -9970
rect 32705 -10004 33081 -9970
rect 32069 -10262 32445 -10228
rect 32705 -10262 33081 -10228
rect 32069 -10530 32445 -10496
rect 32705 -10530 33081 -10496
rect 32069 -11388 32445 -11354
rect 32705 -11388 33081 -11354
rect 33669 -10004 34045 -9970
rect 34305 -10004 34681 -9970
rect 33669 -10262 34045 -10228
rect 34305 -10262 34681 -10228
rect 33669 -10530 34045 -10496
rect 34305 -10530 34681 -10496
rect 33669 -11388 34045 -11354
rect 34305 -11388 34681 -11354
rect 35269 -10004 35645 -9970
rect 35905 -10004 36281 -9970
rect 35269 -10262 35645 -10228
rect 35905 -10262 36281 -10228
rect 35269 -10530 35645 -10496
rect 35905 -10530 36281 -10496
rect 35269 -11388 35645 -11354
rect 35905 -11388 36281 -11354
rect 36869 -10004 37245 -9970
rect 37505 -10004 37881 -9970
rect 36869 -10262 37245 -10228
rect 37505 -10262 37881 -10228
rect 36869 -10530 37245 -10496
rect 37505 -10530 37881 -10496
rect 36869 -11388 37245 -11354
rect 37505 -11388 37881 -11354
rect 69 -11804 445 -11770
rect 705 -11804 1081 -11770
rect 69 -12062 445 -12028
rect 705 -12062 1081 -12028
rect 69 -12330 445 -12296
rect 705 -12330 1081 -12296
rect 69 -13188 445 -13154
rect 705 -13188 1081 -13154
rect 1669 -11804 2045 -11770
rect 2305 -11804 2681 -11770
rect 1669 -12062 2045 -12028
rect 2305 -12062 2681 -12028
rect 1669 -12330 2045 -12296
rect 2305 -12330 2681 -12296
rect 1669 -13188 2045 -13154
rect 2305 -13188 2681 -13154
rect 3269 -11804 3645 -11770
rect 3905 -11804 4281 -11770
rect 3269 -12062 3645 -12028
rect 3905 -12062 4281 -12028
rect 3269 -12330 3645 -12296
rect 3905 -12330 4281 -12296
rect 3269 -13188 3645 -13154
rect 3905 -13188 4281 -13154
rect 4869 -11804 5245 -11770
rect 5505 -11804 5881 -11770
rect 4869 -12062 5245 -12028
rect 5505 -12062 5881 -12028
rect 4869 -12330 5245 -12296
rect 5505 -12330 5881 -12296
rect 4869 -13188 5245 -13154
rect 5505 -13188 5881 -13154
rect 6469 -11804 6845 -11770
rect 7105 -11804 7481 -11770
rect 6469 -12062 6845 -12028
rect 7105 -12062 7481 -12028
rect 6469 -12330 6845 -12296
rect 7105 -12330 7481 -12296
rect 6469 -13188 6845 -13154
rect 7105 -13188 7481 -13154
rect 8069 -11804 8445 -11770
rect 8705 -11804 9081 -11770
rect 8069 -12062 8445 -12028
rect 8705 -12062 9081 -12028
rect 8069 -12330 8445 -12296
rect 8705 -12330 9081 -12296
rect 8069 -13188 8445 -13154
rect 8705 -13188 9081 -13154
rect 9669 -11804 10045 -11770
rect 10305 -11804 10681 -11770
rect 9669 -12062 10045 -12028
rect 10305 -12062 10681 -12028
rect 9669 -12330 10045 -12296
rect 10305 -12330 10681 -12296
rect 9669 -13188 10045 -13154
rect 10305 -13188 10681 -13154
rect 11269 -11804 11645 -11770
rect 11905 -11804 12281 -11770
rect 11269 -12062 11645 -12028
rect 11905 -12062 12281 -12028
rect 11269 -12330 11645 -12296
rect 11905 -12330 12281 -12296
rect 11269 -13188 11645 -13154
rect 11905 -13188 12281 -13154
rect 12869 -11804 13245 -11770
rect 13505 -11804 13881 -11770
rect 12869 -12062 13245 -12028
rect 13505 -12062 13881 -12028
rect 12869 -12330 13245 -12296
rect 13505 -12330 13881 -12296
rect 12869 -13188 13245 -13154
rect 13505 -13188 13881 -13154
rect 14469 -11804 14845 -11770
rect 15105 -11804 15481 -11770
rect 14469 -12062 14845 -12028
rect 15105 -12062 15481 -12028
rect 14469 -12330 14845 -12296
rect 15105 -12330 15481 -12296
rect 14469 -13188 14845 -13154
rect 15105 -13188 15481 -13154
rect 16069 -11804 16445 -11770
rect 16705 -11804 17081 -11770
rect 16069 -12062 16445 -12028
rect 16705 -12062 17081 -12028
rect 16069 -12330 16445 -12296
rect 16705 -12330 17081 -12296
rect 16069 -13188 16445 -13154
rect 16705 -13188 17081 -13154
rect 17669 -11804 18045 -11770
rect 18305 -11804 18681 -11770
rect 17669 -12062 18045 -12028
rect 18305 -12062 18681 -12028
rect 17669 -12330 18045 -12296
rect 18305 -12330 18681 -12296
rect 17669 -13188 18045 -13154
rect 18305 -13188 18681 -13154
rect 19269 -11804 19645 -11770
rect 19905 -11804 20281 -11770
rect 19269 -12062 19645 -12028
rect 19905 -12062 20281 -12028
rect 19269 -12330 19645 -12296
rect 19905 -12330 20281 -12296
rect 19269 -13188 19645 -13154
rect 19905 -13188 20281 -13154
rect 20869 -11804 21245 -11770
rect 21505 -11804 21881 -11770
rect 20869 -12062 21245 -12028
rect 21505 -12062 21881 -12028
rect 20869 -12330 21245 -12296
rect 21505 -12330 21881 -12296
rect 20869 -13188 21245 -13154
rect 21505 -13188 21881 -13154
rect 22469 -11804 22845 -11770
rect 23105 -11804 23481 -11770
rect 22469 -12062 22845 -12028
rect 23105 -12062 23481 -12028
rect 22469 -12330 22845 -12296
rect 23105 -12330 23481 -12296
rect 22469 -13188 22845 -13154
rect 23105 -13188 23481 -13154
rect 24069 -11804 24445 -11770
rect 24705 -11804 25081 -11770
rect 24069 -12062 24445 -12028
rect 24705 -12062 25081 -12028
rect 24069 -12330 24445 -12296
rect 24705 -12330 25081 -12296
rect 24069 -13188 24445 -13154
rect 24705 -13188 25081 -13154
rect 25669 -11804 26045 -11770
rect 26305 -11804 26681 -11770
rect 25669 -12062 26045 -12028
rect 26305 -12062 26681 -12028
rect 25669 -12330 26045 -12296
rect 26305 -12330 26681 -12296
rect 25669 -13188 26045 -13154
rect 26305 -13188 26681 -13154
rect 27269 -11804 27645 -11770
rect 27905 -11804 28281 -11770
rect 27269 -12062 27645 -12028
rect 27905 -12062 28281 -12028
rect 27269 -12330 27645 -12296
rect 27905 -12330 28281 -12296
rect 27269 -13188 27645 -13154
rect 27905 -13188 28281 -13154
rect 28869 -11804 29245 -11770
rect 29505 -11804 29881 -11770
rect 28869 -12062 29245 -12028
rect 29505 -12062 29881 -12028
rect 28869 -12330 29245 -12296
rect 29505 -12330 29881 -12296
rect 28869 -13188 29245 -13154
rect 29505 -13188 29881 -13154
rect 30469 -11804 30845 -11770
rect 31105 -11804 31481 -11770
rect 30469 -12062 30845 -12028
rect 31105 -12062 31481 -12028
rect 30469 -12330 30845 -12296
rect 31105 -12330 31481 -12296
rect 30469 -13188 30845 -13154
rect 31105 -13188 31481 -13154
rect 32069 -11804 32445 -11770
rect 32705 -11804 33081 -11770
rect 32069 -12062 32445 -12028
rect 32705 -12062 33081 -12028
rect 32069 -12330 32445 -12296
rect 32705 -12330 33081 -12296
rect 32069 -13188 32445 -13154
rect 32705 -13188 33081 -13154
rect 33669 -11804 34045 -11770
rect 34305 -11804 34681 -11770
rect 33669 -12062 34045 -12028
rect 34305 -12062 34681 -12028
rect 33669 -12330 34045 -12296
rect 34305 -12330 34681 -12296
rect 33669 -13188 34045 -13154
rect 34305 -13188 34681 -13154
rect 35269 -11804 35645 -11770
rect 35905 -11804 36281 -11770
rect 35269 -12062 35645 -12028
rect 35905 -12062 36281 -12028
rect 35269 -12330 35645 -12296
rect 35905 -12330 36281 -12296
rect 35269 -13188 35645 -13154
rect 35905 -13188 36281 -13154
rect 36869 -11804 37245 -11770
rect 37505 -11804 37881 -11770
rect 36869 -12062 37245 -12028
rect 37505 -12062 37881 -12028
rect 36869 -12330 37245 -12296
rect 37505 -12330 37881 -12296
rect 36869 -13188 37245 -13154
rect 37505 -13188 37881 -13154
rect 69 -13604 445 -13570
rect 705 -13604 1081 -13570
rect 69 -13862 445 -13828
rect 705 -13862 1081 -13828
rect 69 -14130 445 -14096
rect 705 -14130 1081 -14096
rect 69 -14988 445 -14954
rect 705 -14988 1081 -14954
rect 1669 -13604 2045 -13570
rect 2305 -13604 2681 -13570
rect 1669 -13862 2045 -13828
rect 2305 -13862 2681 -13828
rect 1669 -14130 2045 -14096
rect 2305 -14130 2681 -14096
rect 1669 -14988 2045 -14954
rect 2305 -14988 2681 -14954
rect 3269 -13604 3645 -13570
rect 3905 -13604 4281 -13570
rect 3269 -13862 3645 -13828
rect 3905 -13862 4281 -13828
rect 3269 -14130 3645 -14096
rect 3905 -14130 4281 -14096
rect 3269 -14988 3645 -14954
rect 3905 -14988 4281 -14954
rect 4869 -13604 5245 -13570
rect 5505 -13604 5881 -13570
rect 4869 -13862 5245 -13828
rect 5505 -13862 5881 -13828
rect 4869 -14130 5245 -14096
rect 5505 -14130 5881 -14096
rect 4869 -14988 5245 -14954
rect 5505 -14988 5881 -14954
rect 6469 -13604 6845 -13570
rect 7105 -13604 7481 -13570
rect 6469 -13862 6845 -13828
rect 7105 -13862 7481 -13828
rect 6469 -14130 6845 -14096
rect 7105 -14130 7481 -14096
rect 6469 -14988 6845 -14954
rect 7105 -14988 7481 -14954
rect 8069 -13604 8445 -13570
rect 8705 -13604 9081 -13570
rect 8069 -13862 8445 -13828
rect 8705 -13862 9081 -13828
rect 8069 -14130 8445 -14096
rect 8705 -14130 9081 -14096
rect 8069 -14988 8445 -14954
rect 8705 -14988 9081 -14954
rect 9669 -13604 10045 -13570
rect 10305 -13604 10681 -13570
rect 9669 -13862 10045 -13828
rect 10305 -13862 10681 -13828
rect 9669 -14130 10045 -14096
rect 10305 -14130 10681 -14096
rect 9669 -14988 10045 -14954
rect 10305 -14988 10681 -14954
rect 11269 -13604 11645 -13570
rect 11905 -13604 12281 -13570
rect 11269 -13862 11645 -13828
rect 11905 -13862 12281 -13828
rect 11269 -14130 11645 -14096
rect 11905 -14130 12281 -14096
rect 11269 -14988 11645 -14954
rect 11905 -14988 12281 -14954
rect 12869 -13604 13245 -13570
rect 13505 -13604 13881 -13570
rect 12869 -13862 13245 -13828
rect 13505 -13862 13881 -13828
rect 12869 -14130 13245 -14096
rect 13505 -14130 13881 -14096
rect 12869 -14988 13245 -14954
rect 13505 -14988 13881 -14954
rect 14469 -13604 14845 -13570
rect 15105 -13604 15481 -13570
rect 14469 -13862 14845 -13828
rect 15105 -13862 15481 -13828
rect 14469 -14130 14845 -14096
rect 15105 -14130 15481 -14096
rect 14469 -14988 14845 -14954
rect 15105 -14988 15481 -14954
rect 16069 -13604 16445 -13570
rect 16705 -13604 17081 -13570
rect 16069 -13862 16445 -13828
rect 16705 -13862 17081 -13828
rect 16069 -14130 16445 -14096
rect 16705 -14130 17081 -14096
rect 16069 -14988 16445 -14954
rect 16705 -14988 17081 -14954
rect 17669 -13604 18045 -13570
rect 18305 -13604 18681 -13570
rect 17669 -13862 18045 -13828
rect 18305 -13862 18681 -13828
rect 17669 -14130 18045 -14096
rect 18305 -14130 18681 -14096
rect 17669 -14988 18045 -14954
rect 18305 -14988 18681 -14954
rect 19269 -13604 19645 -13570
rect 19905 -13604 20281 -13570
rect 19269 -13862 19645 -13828
rect 19905 -13862 20281 -13828
rect 19269 -14130 19645 -14096
rect 19905 -14130 20281 -14096
rect 19269 -14988 19645 -14954
rect 19905 -14988 20281 -14954
rect 20869 -13604 21245 -13570
rect 21505 -13604 21881 -13570
rect 20869 -13862 21245 -13828
rect 21505 -13862 21881 -13828
rect 20869 -14130 21245 -14096
rect 21505 -14130 21881 -14096
rect 20869 -14988 21245 -14954
rect 21505 -14988 21881 -14954
rect 22469 -13604 22845 -13570
rect 23105 -13604 23481 -13570
rect 22469 -13862 22845 -13828
rect 23105 -13862 23481 -13828
rect 22469 -14130 22845 -14096
rect 23105 -14130 23481 -14096
rect 22469 -14988 22845 -14954
rect 23105 -14988 23481 -14954
rect 24069 -13604 24445 -13570
rect 24705 -13604 25081 -13570
rect 24069 -13862 24445 -13828
rect 24705 -13862 25081 -13828
rect 24069 -14130 24445 -14096
rect 24705 -14130 25081 -14096
rect 24069 -14988 24445 -14954
rect 24705 -14988 25081 -14954
rect 25669 -13604 26045 -13570
rect 26305 -13604 26681 -13570
rect 25669 -13862 26045 -13828
rect 26305 -13862 26681 -13828
rect 25669 -14130 26045 -14096
rect 26305 -14130 26681 -14096
rect 25669 -14988 26045 -14954
rect 26305 -14988 26681 -14954
rect 27269 -13604 27645 -13570
rect 27905 -13604 28281 -13570
rect 27269 -13862 27645 -13828
rect 27905 -13862 28281 -13828
rect 27269 -14130 27645 -14096
rect 27905 -14130 28281 -14096
rect 27269 -14988 27645 -14954
rect 27905 -14988 28281 -14954
rect 28869 -13604 29245 -13570
rect 29505 -13604 29881 -13570
rect 28869 -13862 29245 -13828
rect 29505 -13862 29881 -13828
rect 28869 -14130 29245 -14096
rect 29505 -14130 29881 -14096
rect 28869 -14988 29245 -14954
rect 29505 -14988 29881 -14954
rect 30469 -13604 30845 -13570
rect 31105 -13604 31481 -13570
rect 30469 -13862 30845 -13828
rect 31105 -13862 31481 -13828
rect 30469 -14130 30845 -14096
rect 31105 -14130 31481 -14096
rect 30469 -14988 30845 -14954
rect 31105 -14988 31481 -14954
rect 32069 -13604 32445 -13570
rect 32705 -13604 33081 -13570
rect 32069 -13862 32445 -13828
rect 32705 -13862 33081 -13828
rect 32069 -14130 32445 -14096
rect 32705 -14130 33081 -14096
rect 32069 -14988 32445 -14954
rect 32705 -14988 33081 -14954
rect 33669 -13604 34045 -13570
rect 34305 -13604 34681 -13570
rect 33669 -13862 34045 -13828
rect 34305 -13862 34681 -13828
rect 33669 -14130 34045 -14096
rect 34305 -14130 34681 -14096
rect 33669 -14988 34045 -14954
rect 34305 -14988 34681 -14954
rect 35269 -13604 35645 -13570
rect 35905 -13604 36281 -13570
rect 35269 -13862 35645 -13828
rect 35905 -13862 36281 -13828
rect 35269 -14130 35645 -14096
rect 35905 -14130 36281 -14096
rect 35269 -14988 35645 -14954
rect 35905 -14988 36281 -14954
rect 36869 -13604 37245 -13570
rect 37505 -13604 37881 -13570
rect 36869 -13862 37245 -13828
rect 37505 -13862 37881 -13828
rect 36869 -14130 37245 -14096
rect 37505 -14130 37881 -14096
rect 36869 -14988 37245 -14954
rect 37505 -14988 37881 -14954
rect 69 -15404 445 -15370
rect 705 -15404 1081 -15370
rect 69 -15662 445 -15628
rect 705 -15662 1081 -15628
rect 69 -15930 445 -15896
rect 705 -15930 1081 -15896
rect 69 -16788 445 -16754
rect 705 -16788 1081 -16754
rect 1669 -15404 2045 -15370
rect 2305 -15404 2681 -15370
rect 1669 -15662 2045 -15628
rect 2305 -15662 2681 -15628
rect 1669 -15930 2045 -15896
rect 2305 -15930 2681 -15896
rect 1669 -16788 2045 -16754
rect 2305 -16788 2681 -16754
rect 3269 -15404 3645 -15370
rect 3905 -15404 4281 -15370
rect 3269 -15662 3645 -15628
rect 3905 -15662 4281 -15628
rect 3269 -15930 3645 -15896
rect 3905 -15930 4281 -15896
rect 3269 -16788 3645 -16754
rect 3905 -16788 4281 -16754
rect 4869 -15404 5245 -15370
rect 5505 -15404 5881 -15370
rect 4869 -15662 5245 -15628
rect 5505 -15662 5881 -15628
rect 4869 -15930 5245 -15896
rect 5505 -15930 5881 -15896
rect 4869 -16788 5245 -16754
rect 5505 -16788 5881 -16754
rect 6469 -15404 6845 -15370
rect 7105 -15404 7481 -15370
rect 6469 -15662 6845 -15628
rect 7105 -15662 7481 -15628
rect 6469 -15930 6845 -15896
rect 7105 -15930 7481 -15896
rect 6469 -16788 6845 -16754
rect 7105 -16788 7481 -16754
rect 8069 -15404 8445 -15370
rect 8705 -15404 9081 -15370
rect 8069 -15662 8445 -15628
rect 8705 -15662 9081 -15628
rect 8069 -15930 8445 -15896
rect 8705 -15930 9081 -15896
rect 8069 -16788 8445 -16754
rect 8705 -16788 9081 -16754
rect 9669 -15404 10045 -15370
rect 10305 -15404 10681 -15370
rect 9669 -15662 10045 -15628
rect 10305 -15662 10681 -15628
rect 9669 -15930 10045 -15896
rect 10305 -15930 10681 -15896
rect 9669 -16788 10045 -16754
rect 10305 -16788 10681 -16754
rect 11269 -15404 11645 -15370
rect 11905 -15404 12281 -15370
rect 11269 -15662 11645 -15628
rect 11905 -15662 12281 -15628
rect 11269 -15930 11645 -15896
rect 11905 -15930 12281 -15896
rect 11269 -16788 11645 -16754
rect 11905 -16788 12281 -16754
rect 12869 -15404 13245 -15370
rect 13505 -15404 13881 -15370
rect 12869 -15662 13245 -15628
rect 13505 -15662 13881 -15628
rect 12869 -15930 13245 -15896
rect 13505 -15930 13881 -15896
rect 12869 -16788 13245 -16754
rect 13505 -16788 13881 -16754
rect 14469 -15404 14845 -15370
rect 15105 -15404 15481 -15370
rect 14469 -15662 14845 -15628
rect 15105 -15662 15481 -15628
rect 14469 -15930 14845 -15896
rect 15105 -15930 15481 -15896
rect 14469 -16788 14845 -16754
rect 15105 -16788 15481 -16754
rect 16069 -15404 16445 -15370
rect 16705 -15404 17081 -15370
rect 16069 -15662 16445 -15628
rect 16705 -15662 17081 -15628
rect 16069 -15930 16445 -15896
rect 16705 -15930 17081 -15896
rect 16069 -16788 16445 -16754
rect 16705 -16788 17081 -16754
rect 17669 -15404 18045 -15370
rect 18305 -15404 18681 -15370
rect 17669 -15662 18045 -15628
rect 18305 -15662 18681 -15628
rect 17669 -15930 18045 -15896
rect 18305 -15930 18681 -15896
rect 17669 -16788 18045 -16754
rect 18305 -16788 18681 -16754
rect 19269 -15404 19645 -15370
rect 19905 -15404 20281 -15370
rect 19269 -15662 19645 -15628
rect 19905 -15662 20281 -15628
rect 19269 -15930 19645 -15896
rect 19905 -15930 20281 -15896
rect 19269 -16788 19645 -16754
rect 19905 -16788 20281 -16754
rect 20869 -15404 21245 -15370
rect 21505 -15404 21881 -15370
rect 20869 -15662 21245 -15628
rect 21505 -15662 21881 -15628
rect 20869 -15930 21245 -15896
rect 21505 -15930 21881 -15896
rect 20869 -16788 21245 -16754
rect 21505 -16788 21881 -16754
rect 22469 -15404 22845 -15370
rect 23105 -15404 23481 -15370
rect 22469 -15662 22845 -15628
rect 23105 -15662 23481 -15628
rect 22469 -15930 22845 -15896
rect 23105 -15930 23481 -15896
rect 22469 -16788 22845 -16754
rect 23105 -16788 23481 -16754
rect 24069 -15404 24445 -15370
rect 24705 -15404 25081 -15370
rect 24069 -15662 24445 -15628
rect 24705 -15662 25081 -15628
rect 24069 -15930 24445 -15896
rect 24705 -15930 25081 -15896
rect 24069 -16788 24445 -16754
rect 24705 -16788 25081 -16754
rect 25669 -15404 26045 -15370
rect 26305 -15404 26681 -15370
rect 25669 -15662 26045 -15628
rect 26305 -15662 26681 -15628
rect 25669 -15930 26045 -15896
rect 26305 -15930 26681 -15896
rect 25669 -16788 26045 -16754
rect 26305 -16788 26681 -16754
rect 27269 -15404 27645 -15370
rect 27905 -15404 28281 -15370
rect 27269 -15662 27645 -15628
rect 27905 -15662 28281 -15628
rect 27269 -15930 27645 -15896
rect 27905 -15930 28281 -15896
rect 27269 -16788 27645 -16754
rect 27905 -16788 28281 -16754
rect 28869 -15404 29245 -15370
rect 29505 -15404 29881 -15370
rect 28869 -15662 29245 -15628
rect 29505 -15662 29881 -15628
rect 28869 -15930 29245 -15896
rect 29505 -15930 29881 -15896
rect 28869 -16788 29245 -16754
rect 29505 -16788 29881 -16754
rect 30469 -15404 30845 -15370
rect 31105 -15404 31481 -15370
rect 30469 -15662 30845 -15628
rect 31105 -15662 31481 -15628
rect 30469 -15930 30845 -15896
rect 31105 -15930 31481 -15896
rect 30469 -16788 30845 -16754
rect 31105 -16788 31481 -16754
rect 32069 -15404 32445 -15370
rect 32705 -15404 33081 -15370
rect 32069 -15662 32445 -15628
rect 32705 -15662 33081 -15628
rect 32069 -15930 32445 -15896
rect 32705 -15930 33081 -15896
rect 32069 -16788 32445 -16754
rect 32705 -16788 33081 -16754
rect 33669 -15404 34045 -15370
rect 34305 -15404 34681 -15370
rect 33669 -15662 34045 -15628
rect 34305 -15662 34681 -15628
rect 33669 -15930 34045 -15896
rect 34305 -15930 34681 -15896
rect 33669 -16788 34045 -16754
rect 34305 -16788 34681 -16754
rect 35269 -15404 35645 -15370
rect 35905 -15404 36281 -15370
rect 35269 -15662 35645 -15628
rect 35905 -15662 36281 -15628
rect 35269 -15930 35645 -15896
rect 35905 -15930 36281 -15896
rect 35269 -16788 35645 -16754
rect 35905 -16788 36281 -16754
rect 36869 -15404 37245 -15370
rect 37505 -15404 37881 -15370
rect 36869 -15662 37245 -15628
rect 37505 -15662 37881 -15628
rect 36869 -15930 37245 -15896
rect 37505 -15930 37881 -15896
rect 36869 -16788 37245 -16754
rect 37505 -16788 37881 -16754
rect 69 -17204 445 -17170
rect 705 -17204 1081 -17170
rect 69 -17462 445 -17428
rect 705 -17462 1081 -17428
rect 69 -17730 445 -17696
rect 705 -17730 1081 -17696
rect 69 -18588 445 -18554
rect 705 -18588 1081 -18554
rect 1669 -17204 2045 -17170
rect 2305 -17204 2681 -17170
rect 1669 -17462 2045 -17428
rect 2305 -17462 2681 -17428
rect 1669 -17730 2045 -17696
rect 2305 -17730 2681 -17696
rect 1669 -18588 2045 -18554
rect 2305 -18588 2681 -18554
rect 3269 -17204 3645 -17170
rect 3905 -17204 4281 -17170
rect 3269 -17462 3645 -17428
rect 3905 -17462 4281 -17428
rect 3269 -17730 3645 -17696
rect 3905 -17730 4281 -17696
rect 3269 -18588 3645 -18554
rect 3905 -18588 4281 -18554
rect 4869 -17204 5245 -17170
rect 5505 -17204 5881 -17170
rect 4869 -17462 5245 -17428
rect 5505 -17462 5881 -17428
rect 4869 -17730 5245 -17696
rect 5505 -17730 5881 -17696
rect 4869 -18588 5245 -18554
rect 5505 -18588 5881 -18554
rect 6469 -17204 6845 -17170
rect 7105 -17204 7481 -17170
rect 6469 -17462 6845 -17428
rect 7105 -17462 7481 -17428
rect 6469 -17730 6845 -17696
rect 7105 -17730 7481 -17696
rect 6469 -18588 6845 -18554
rect 7105 -18588 7481 -18554
rect 8069 -17204 8445 -17170
rect 8705 -17204 9081 -17170
rect 8069 -17462 8445 -17428
rect 8705 -17462 9081 -17428
rect 8069 -17730 8445 -17696
rect 8705 -17730 9081 -17696
rect 8069 -18588 8445 -18554
rect 8705 -18588 9081 -18554
rect 9669 -17204 10045 -17170
rect 10305 -17204 10681 -17170
rect 9669 -17462 10045 -17428
rect 10305 -17462 10681 -17428
rect 9669 -17730 10045 -17696
rect 10305 -17730 10681 -17696
rect 9669 -18588 10045 -18554
rect 10305 -18588 10681 -18554
rect 11269 -17204 11645 -17170
rect 11905 -17204 12281 -17170
rect 11269 -17462 11645 -17428
rect 11905 -17462 12281 -17428
rect 11269 -17730 11645 -17696
rect 11905 -17730 12281 -17696
rect 11269 -18588 11645 -18554
rect 11905 -18588 12281 -18554
rect 12869 -17204 13245 -17170
rect 13505 -17204 13881 -17170
rect 12869 -17462 13245 -17428
rect 13505 -17462 13881 -17428
rect 12869 -17730 13245 -17696
rect 13505 -17730 13881 -17696
rect 12869 -18588 13245 -18554
rect 13505 -18588 13881 -18554
rect 14469 -17204 14845 -17170
rect 15105 -17204 15481 -17170
rect 14469 -17462 14845 -17428
rect 15105 -17462 15481 -17428
rect 14469 -17730 14845 -17696
rect 15105 -17730 15481 -17696
rect 14469 -18588 14845 -18554
rect 15105 -18588 15481 -18554
rect 16069 -17204 16445 -17170
rect 16705 -17204 17081 -17170
rect 16069 -17462 16445 -17428
rect 16705 -17462 17081 -17428
rect 16069 -17730 16445 -17696
rect 16705 -17730 17081 -17696
rect 16069 -18588 16445 -18554
rect 16705 -18588 17081 -18554
rect 17669 -17204 18045 -17170
rect 18305 -17204 18681 -17170
rect 17669 -17462 18045 -17428
rect 18305 -17462 18681 -17428
rect 17669 -17730 18045 -17696
rect 18305 -17730 18681 -17696
rect 17669 -18588 18045 -18554
rect 18305 -18588 18681 -18554
rect 19269 -17204 19645 -17170
rect 19905 -17204 20281 -17170
rect 19269 -17462 19645 -17428
rect 19905 -17462 20281 -17428
rect 19269 -17730 19645 -17696
rect 19905 -17730 20281 -17696
rect 19269 -18588 19645 -18554
rect 19905 -18588 20281 -18554
rect 20869 -17204 21245 -17170
rect 21505 -17204 21881 -17170
rect 20869 -17462 21245 -17428
rect 21505 -17462 21881 -17428
rect 20869 -17730 21245 -17696
rect 21505 -17730 21881 -17696
rect 20869 -18588 21245 -18554
rect 21505 -18588 21881 -18554
rect 22469 -17204 22845 -17170
rect 23105 -17204 23481 -17170
rect 22469 -17462 22845 -17428
rect 23105 -17462 23481 -17428
rect 22469 -17730 22845 -17696
rect 23105 -17730 23481 -17696
rect 22469 -18588 22845 -18554
rect 23105 -18588 23481 -18554
rect 24069 -17204 24445 -17170
rect 24705 -17204 25081 -17170
rect 24069 -17462 24445 -17428
rect 24705 -17462 25081 -17428
rect 24069 -17730 24445 -17696
rect 24705 -17730 25081 -17696
rect 24069 -18588 24445 -18554
rect 24705 -18588 25081 -18554
rect 25669 -17204 26045 -17170
rect 26305 -17204 26681 -17170
rect 25669 -17462 26045 -17428
rect 26305 -17462 26681 -17428
rect 25669 -17730 26045 -17696
rect 26305 -17730 26681 -17696
rect 25669 -18588 26045 -18554
rect 26305 -18588 26681 -18554
rect 27269 -17204 27645 -17170
rect 27905 -17204 28281 -17170
rect 27269 -17462 27645 -17428
rect 27905 -17462 28281 -17428
rect 27269 -17730 27645 -17696
rect 27905 -17730 28281 -17696
rect 27269 -18588 27645 -18554
rect 27905 -18588 28281 -18554
rect 28869 -17204 29245 -17170
rect 29505 -17204 29881 -17170
rect 28869 -17462 29245 -17428
rect 29505 -17462 29881 -17428
rect 28869 -17730 29245 -17696
rect 29505 -17730 29881 -17696
rect 28869 -18588 29245 -18554
rect 29505 -18588 29881 -18554
rect 30469 -17204 30845 -17170
rect 31105 -17204 31481 -17170
rect 30469 -17462 30845 -17428
rect 31105 -17462 31481 -17428
rect 30469 -17730 30845 -17696
rect 31105 -17730 31481 -17696
rect 30469 -18588 30845 -18554
rect 31105 -18588 31481 -18554
rect 32069 -17204 32445 -17170
rect 32705 -17204 33081 -17170
rect 32069 -17462 32445 -17428
rect 32705 -17462 33081 -17428
rect 32069 -17730 32445 -17696
rect 32705 -17730 33081 -17696
rect 32069 -18588 32445 -18554
rect 32705 -18588 33081 -18554
rect 33669 -17204 34045 -17170
rect 34305 -17204 34681 -17170
rect 33669 -17462 34045 -17428
rect 34305 -17462 34681 -17428
rect 33669 -17730 34045 -17696
rect 34305 -17730 34681 -17696
rect 33669 -18588 34045 -18554
rect 34305 -18588 34681 -18554
rect 35269 -17204 35645 -17170
rect 35905 -17204 36281 -17170
rect 35269 -17462 35645 -17428
rect 35905 -17462 36281 -17428
rect 35269 -17730 35645 -17696
rect 35905 -17730 36281 -17696
rect 35269 -18588 35645 -18554
rect 35905 -18588 36281 -18554
rect 36869 -17204 37245 -17170
rect 37505 -17204 37881 -17170
rect 36869 -17462 37245 -17428
rect 37505 -17462 37881 -17428
rect 36869 -17730 37245 -17696
rect 37505 -17730 37881 -17696
rect 36869 -18588 37245 -18554
rect 37505 -18588 37881 -18554
rect 69 -19004 445 -18970
rect 705 -19004 1081 -18970
rect 69 -19262 445 -19228
rect 705 -19262 1081 -19228
rect 69 -19530 445 -19496
rect 705 -19530 1081 -19496
rect 69 -20388 445 -20354
rect 705 -20388 1081 -20354
rect 1669 -19004 2045 -18970
rect 2305 -19004 2681 -18970
rect 1669 -19262 2045 -19228
rect 2305 -19262 2681 -19228
rect 1669 -19530 2045 -19496
rect 2305 -19530 2681 -19496
rect 1669 -20388 2045 -20354
rect 2305 -20388 2681 -20354
rect 3269 -19004 3645 -18970
rect 3905 -19004 4281 -18970
rect 3269 -19262 3645 -19228
rect 3905 -19262 4281 -19228
rect 3269 -19530 3645 -19496
rect 3905 -19530 4281 -19496
rect 3269 -20388 3645 -20354
rect 3905 -20388 4281 -20354
rect 4869 -19004 5245 -18970
rect 5505 -19004 5881 -18970
rect 4869 -19262 5245 -19228
rect 5505 -19262 5881 -19228
rect 4869 -19530 5245 -19496
rect 5505 -19530 5881 -19496
rect 4869 -20388 5245 -20354
rect 5505 -20388 5881 -20354
rect 6469 -19004 6845 -18970
rect 7105 -19004 7481 -18970
rect 6469 -19262 6845 -19228
rect 7105 -19262 7481 -19228
rect 6469 -19530 6845 -19496
rect 7105 -19530 7481 -19496
rect 6469 -20388 6845 -20354
rect 7105 -20388 7481 -20354
rect 8069 -19004 8445 -18970
rect 8705 -19004 9081 -18970
rect 8069 -19262 8445 -19228
rect 8705 -19262 9081 -19228
rect 8069 -19530 8445 -19496
rect 8705 -19530 9081 -19496
rect 8069 -20388 8445 -20354
rect 8705 -20388 9081 -20354
rect 9669 -19004 10045 -18970
rect 10305 -19004 10681 -18970
rect 9669 -19262 10045 -19228
rect 10305 -19262 10681 -19228
rect 9669 -19530 10045 -19496
rect 10305 -19530 10681 -19496
rect 9669 -20388 10045 -20354
rect 10305 -20388 10681 -20354
rect 11269 -19004 11645 -18970
rect 11905 -19004 12281 -18970
rect 11269 -19262 11645 -19228
rect 11905 -19262 12281 -19228
rect 11269 -19530 11645 -19496
rect 11905 -19530 12281 -19496
rect 11269 -20388 11645 -20354
rect 11905 -20388 12281 -20354
rect 12869 -19004 13245 -18970
rect 13505 -19004 13881 -18970
rect 12869 -19262 13245 -19228
rect 13505 -19262 13881 -19228
rect 12869 -19530 13245 -19496
rect 13505 -19530 13881 -19496
rect 12869 -20388 13245 -20354
rect 13505 -20388 13881 -20354
rect 14469 -19004 14845 -18970
rect 15105 -19004 15481 -18970
rect 14469 -19262 14845 -19228
rect 15105 -19262 15481 -19228
rect 14469 -19530 14845 -19496
rect 15105 -19530 15481 -19496
rect 14469 -20388 14845 -20354
rect 15105 -20388 15481 -20354
rect 16069 -19004 16445 -18970
rect 16705 -19004 17081 -18970
rect 16069 -19262 16445 -19228
rect 16705 -19262 17081 -19228
rect 16069 -19530 16445 -19496
rect 16705 -19530 17081 -19496
rect 16069 -20388 16445 -20354
rect 16705 -20388 17081 -20354
rect 17669 -19004 18045 -18970
rect 18305 -19004 18681 -18970
rect 17669 -19262 18045 -19228
rect 18305 -19262 18681 -19228
rect 17669 -19530 18045 -19496
rect 18305 -19530 18681 -19496
rect 17669 -20388 18045 -20354
rect 18305 -20388 18681 -20354
rect 19269 -19004 19645 -18970
rect 19905 -19004 20281 -18970
rect 19269 -19262 19645 -19228
rect 19905 -19262 20281 -19228
rect 19269 -19530 19645 -19496
rect 19905 -19530 20281 -19496
rect 19269 -20388 19645 -20354
rect 19905 -20388 20281 -20354
rect 20869 -19004 21245 -18970
rect 21505 -19004 21881 -18970
rect 20869 -19262 21245 -19228
rect 21505 -19262 21881 -19228
rect 20869 -19530 21245 -19496
rect 21505 -19530 21881 -19496
rect 20869 -20388 21245 -20354
rect 21505 -20388 21881 -20354
rect 22469 -19004 22845 -18970
rect 23105 -19004 23481 -18970
rect 22469 -19262 22845 -19228
rect 23105 -19262 23481 -19228
rect 22469 -19530 22845 -19496
rect 23105 -19530 23481 -19496
rect 22469 -20388 22845 -20354
rect 23105 -20388 23481 -20354
rect 24069 -19004 24445 -18970
rect 24705 -19004 25081 -18970
rect 24069 -19262 24445 -19228
rect 24705 -19262 25081 -19228
rect 24069 -19530 24445 -19496
rect 24705 -19530 25081 -19496
rect 24069 -20388 24445 -20354
rect 24705 -20388 25081 -20354
rect 25669 -19004 26045 -18970
rect 26305 -19004 26681 -18970
rect 25669 -19262 26045 -19228
rect 26305 -19262 26681 -19228
rect 25669 -19530 26045 -19496
rect 26305 -19530 26681 -19496
rect 25669 -20388 26045 -20354
rect 26305 -20388 26681 -20354
rect 27269 -19004 27645 -18970
rect 27905 -19004 28281 -18970
rect 27269 -19262 27645 -19228
rect 27905 -19262 28281 -19228
rect 27269 -19530 27645 -19496
rect 27905 -19530 28281 -19496
rect 27269 -20388 27645 -20354
rect 27905 -20388 28281 -20354
rect 28869 -19004 29245 -18970
rect 29505 -19004 29881 -18970
rect 28869 -19262 29245 -19228
rect 29505 -19262 29881 -19228
rect 28869 -19530 29245 -19496
rect 29505 -19530 29881 -19496
rect 28869 -20388 29245 -20354
rect 29505 -20388 29881 -20354
rect 30469 -19004 30845 -18970
rect 31105 -19004 31481 -18970
rect 30469 -19262 30845 -19228
rect 31105 -19262 31481 -19228
rect 30469 -19530 30845 -19496
rect 31105 -19530 31481 -19496
rect 30469 -20388 30845 -20354
rect 31105 -20388 31481 -20354
rect 32069 -19004 32445 -18970
rect 32705 -19004 33081 -18970
rect 32069 -19262 32445 -19228
rect 32705 -19262 33081 -19228
rect 32069 -19530 32445 -19496
rect 32705 -19530 33081 -19496
rect 32069 -20388 32445 -20354
rect 32705 -20388 33081 -20354
rect 33669 -19004 34045 -18970
rect 34305 -19004 34681 -18970
rect 33669 -19262 34045 -19228
rect 34305 -19262 34681 -19228
rect 33669 -19530 34045 -19496
rect 34305 -19530 34681 -19496
rect 33669 -20388 34045 -20354
rect 34305 -20388 34681 -20354
rect 35269 -19004 35645 -18970
rect 35905 -19004 36281 -18970
rect 35269 -19262 35645 -19228
rect 35905 -19262 36281 -19228
rect 35269 -19530 35645 -19496
rect 35905 -19530 36281 -19496
rect 35269 -20388 35645 -20354
rect 35905 -20388 36281 -20354
rect 36869 -19004 37245 -18970
rect 37505 -19004 37881 -18970
rect 36869 -19262 37245 -19228
rect 37505 -19262 37881 -19228
rect 36869 -19530 37245 -19496
rect 37505 -19530 37881 -19496
rect 36869 -20388 37245 -20354
rect 37505 -20388 37881 -20354
rect 69 -20804 445 -20770
rect 705 -20804 1081 -20770
rect 69 -21062 445 -21028
rect 705 -21062 1081 -21028
rect 69 -21330 445 -21296
rect 705 -21330 1081 -21296
rect 69 -22188 445 -22154
rect 705 -22188 1081 -22154
rect 1669 -20804 2045 -20770
rect 2305 -20804 2681 -20770
rect 1669 -21062 2045 -21028
rect 2305 -21062 2681 -21028
rect 1669 -21330 2045 -21296
rect 2305 -21330 2681 -21296
rect 1669 -22188 2045 -22154
rect 2305 -22188 2681 -22154
rect 3269 -20804 3645 -20770
rect 3905 -20804 4281 -20770
rect 3269 -21062 3645 -21028
rect 3905 -21062 4281 -21028
rect 3269 -21330 3645 -21296
rect 3905 -21330 4281 -21296
rect 3269 -22188 3645 -22154
rect 3905 -22188 4281 -22154
rect 4869 -20804 5245 -20770
rect 5505 -20804 5881 -20770
rect 4869 -21062 5245 -21028
rect 5505 -21062 5881 -21028
rect 4869 -21330 5245 -21296
rect 5505 -21330 5881 -21296
rect 4869 -22188 5245 -22154
rect 5505 -22188 5881 -22154
rect 6469 -20804 6845 -20770
rect 7105 -20804 7481 -20770
rect 6469 -21062 6845 -21028
rect 7105 -21062 7481 -21028
rect 6469 -21330 6845 -21296
rect 7105 -21330 7481 -21296
rect 6469 -22188 6845 -22154
rect 7105 -22188 7481 -22154
rect 8069 -20804 8445 -20770
rect 8705 -20804 9081 -20770
rect 8069 -21062 8445 -21028
rect 8705 -21062 9081 -21028
rect 8069 -21330 8445 -21296
rect 8705 -21330 9081 -21296
rect 8069 -22188 8445 -22154
rect 8705 -22188 9081 -22154
rect 9669 -20804 10045 -20770
rect 10305 -20804 10681 -20770
rect 9669 -21062 10045 -21028
rect 10305 -21062 10681 -21028
rect 9669 -21330 10045 -21296
rect 10305 -21330 10681 -21296
rect 9669 -22188 10045 -22154
rect 10305 -22188 10681 -22154
rect 11269 -20804 11645 -20770
rect 11905 -20804 12281 -20770
rect 11269 -21062 11645 -21028
rect 11905 -21062 12281 -21028
rect 11269 -21330 11645 -21296
rect 11905 -21330 12281 -21296
rect 11269 -22188 11645 -22154
rect 11905 -22188 12281 -22154
rect 12869 -20804 13245 -20770
rect 13505 -20804 13881 -20770
rect 12869 -21062 13245 -21028
rect 13505 -21062 13881 -21028
rect 12869 -21330 13245 -21296
rect 13505 -21330 13881 -21296
rect 12869 -22188 13245 -22154
rect 13505 -22188 13881 -22154
rect 14469 -20804 14845 -20770
rect 15105 -20804 15481 -20770
rect 14469 -21062 14845 -21028
rect 15105 -21062 15481 -21028
rect 14469 -21330 14845 -21296
rect 15105 -21330 15481 -21296
rect 14469 -22188 14845 -22154
rect 15105 -22188 15481 -22154
rect 16069 -20804 16445 -20770
rect 16705 -20804 17081 -20770
rect 16069 -21062 16445 -21028
rect 16705 -21062 17081 -21028
rect 16069 -21330 16445 -21296
rect 16705 -21330 17081 -21296
rect 16069 -22188 16445 -22154
rect 16705 -22188 17081 -22154
rect 17669 -20804 18045 -20770
rect 18305 -20804 18681 -20770
rect 17669 -21062 18045 -21028
rect 18305 -21062 18681 -21028
rect 17669 -21330 18045 -21296
rect 18305 -21330 18681 -21296
rect 17669 -22188 18045 -22154
rect 18305 -22188 18681 -22154
rect 19269 -20804 19645 -20770
rect 19905 -20804 20281 -20770
rect 19269 -21062 19645 -21028
rect 19905 -21062 20281 -21028
rect 19269 -21330 19645 -21296
rect 19905 -21330 20281 -21296
rect 19269 -22188 19645 -22154
rect 19905 -22188 20281 -22154
rect 20869 -20804 21245 -20770
rect 21505 -20804 21881 -20770
rect 20869 -21062 21245 -21028
rect 21505 -21062 21881 -21028
rect 20869 -21330 21245 -21296
rect 21505 -21330 21881 -21296
rect 20869 -22188 21245 -22154
rect 21505 -22188 21881 -22154
rect 22469 -20804 22845 -20770
rect 23105 -20804 23481 -20770
rect 22469 -21062 22845 -21028
rect 23105 -21062 23481 -21028
rect 22469 -21330 22845 -21296
rect 23105 -21330 23481 -21296
rect 22469 -22188 22845 -22154
rect 23105 -22188 23481 -22154
rect 24069 -20804 24445 -20770
rect 24705 -20804 25081 -20770
rect 24069 -21062 24445 -21028
rect 24705 -21062 25081 -21028
rect 24069 -21330 24445 -21296
rect 24705 -21330 25081 -21296
rect 24069 -22188 24445 -22154
rect 24705 -22188 25081 -22154
rect 25669 -20804 26045 -20770
rect 26305 -20804 26681 -20770
rect 25669 -21062 26045 -21028
rect 26305 -21062 26681 -21028
rect 25669 -21330 26045 -21296
rect 26305 -21330 26681 -21296
rect 25669 -22188 26045 -22154
rect 26305 -22188 26681 -22154
rect 27269 -20804 27645 -20770
rect 27905 -20804 28281 -20770
rect 27269 -21062 27645 -21028
rect 27905 -21062 28281 -21028
rect 27269 -21330 27645 -21296
rect 27905 -21330 28281 -21296
rect 27269 -22188 27645 -22154
rect 27905 -22188 28281 -22154
rect 28869 -20804 29245 -20770
rect 29505 -20804 29881 -20770
rect 28869 -21062 29245 -21028
rect 29505 -21062 29881 -21028
rect 28869 -21330 29245 -21296
rect 29505 -21330 29881 -21296
rect 28869 -22188 29245 -22154
rect 29505 -22188 29881 -22154
rect 30469 -20804 30845 -20770
rect 31105 -20804 31481 -20770
rect 30469 -21062 30845 -21028
rect 31105 -21062 31481 -21028
rect 30469 -21330 30845 -21296
rect 31105 -21330 31481 -21296
rect 30469 -22188 30845 -22154
rect 31105 -22188 31481 -22154
rect 32069 -20804 32445 -20770
rect 32705 -20804 33081 -20770
rect 32069 -21062 32445 -21028
rect 32705 -21062 33081 -21028
rect 32069 -21330 32445 -21296
rect 32705 -21330 33081 -21296
rect 32069 -22188 32445 -22154
rect 32705 -22188 33081 -22154
rect 33669 -20804 34045 -20770
rect 34305 -20804 34681 -20770
rect 33669 -21062 34045 -21028
rect 34305 -21062 34681 -21028
rect 33669 -21330 34045 -21296
rect 34305 -21330 34681 -21296
rect 33669 -22188 34045 -22154
rect 34305 -22188 34681 -22154
rect 35269 -20804 35645 -20770
rect 35905 -20804 36281 -20770
rect 35269 -21062 35645 -21028
rect 35905 -21062 36281 -21028
rect 35269 -21330 35645 -21296
rect 35905 -21330 36281 -21296
rect 35269 -22188 35645 -22154
rect 35905 -22188 36281 -22154
rect 36869 -20804 37245 -20770
rect 37505 -20804 37881 -20770
rect 36869 -21062 37245 -21028
rect 37505 -21062 37881 -21028
rect 36869 -21330 37245 -21296
rect 37505 -21330 37881 -21296
rect 36869 -22188 37245 -22154
rect 37505 -22188 37881 -22154
rect 28352 -23460 28386 -22684
rect 28510 -23460 28544 -22684
rect 28668 -23460 28702 -22684
rect 28826 -23460 28860 -22684
rect 28984 -23460 29018 -22684
rect 32632 -23011 32666 -22635
rect 32790 -23011 32824 -22635
rect 32948 -23011 32982 -22635
rect 33106 -23011 33140 -22635
rect 33264 -23011 33298 -22635
rect 34002 -23031 34036 -22655
rect 34160 -23031 34194 -22655
rect 34318 -23031 34352 -22655
rect 279 -24340 1855 -24306
rect 279 -24698 1855 -24664
rect 2479 -24340 4055 -24306
rect 2479 -24698 4055 -24664
rect 4679 -24340 6255 -24306
rect 4679 -24698 6255 -24664
rect 6879 -24340 8455 -24306
rect 6879 -24698 8455 -24664
rect 9079 -24340 10655 -24306
rect 9079 -24698 10655 -24664
rect 11279 -24340 12855 -24306
rect 11279 -24698 12855 -24664
rect 13479 -24340 15055 -24306
rect 13479 -24698 15055 -24664
rect 15679 -24340 17255 -24306
rect 15679 -24698 17255 -24664
rect 17879 -24340 19455 -24306
rect 17879 -24698 19455 -24664
rect 20079 -24340 21655 -24306
rect 20079 -24698 21655 -24664
rect 33170 -24153 33204 -23777
rect 33328 -24153 33362 -23777
rect 33486 -24153 33520 -23777
rect 33644 -24153 33678 -23777
rect 33802 -24153 33836 -23777
rect 33960 -24153 33994 -23777
rect 34118 -24153 34152 -23777
rect 34542 -24151 34576 -23775
rect 34700 -24151 34734 -23775
rect 34858 -24151 34892 -23775
rect 35016 -24151 35050 -23775
rect 35174 -24151 35208 -23775
rect 35332 -24151 35366 -23775
rect 35490 -24151 35524 -23775
rect 35648 -24151 35682 -23775
rect 35806 -24151 35840 -23775
rect 35964 -24151 35998 -23775
rect 36122 -24151 36156 -23775
rect 36280 -24151 36314 -23775
rect 36438 -24151 36472 -23775
rect 36596 -24151 36630 -23775
rect 36754 -24151 36788 -23775
rect 36912 -24151 36946 -23775
rect 37070 -24151 37104 -23775
rect 279 -25140 1855 -25106
rect 279 -25498 1855 -25464
rect 2479 -25140 4055 -25106
rect 2479 -25498 4055 -25464
rect 4679 -25140 6255 -25106
rect 4679 -25498 6255 -25464
rect 6879 -25140 8455 -25106
rect 6879 -25498 8455 -25464
rect 9079 -25140 10655 -25106
rect 9079 -25498 10655 -25464
rect 11279 -25140 12855 -25106
rect 11279 -25498 12855 -25464
rect 13479 -25140 15055 -25106
rect 13479 -25498 15055 -25464
rect 15679 -25140 17255 -25106
rect 15679 -25498 17255 -25464
rect 17879 -25140 19455 -25106
rect 17879 -25498 19455 -25464
rect 20079 -25140 21655 -25106
rect 20079 -25498 21655 -25464
rect 279 -25940 1855 -25906
rect 279 -26298 1855 -26264
rect 2479 -25940 4055 -25906
rect 2479 -26298 4055 -26264
rect 4679 -25940 6255 -25906
rect 4679 -26298 6255 -26264
rect 6879 -25940 8455 -25906
rect 6879 -26298 8455 -26264
rect 9079 -25940 10655 -25906
rect 9079 -26298 10655 -26264
rect 11279 -25940 12855 -25906
rect 11279 -26298 12855 -26264
rect 13479 -25940 15055 -25906
rect 13479 -26298 15055 -26264
rect 15679 -25940 17255 -25906
rect 15679 -26298 17255 -26264
rect 17879 -25940 19455 -25906
rect 17879 -26298 19455 -26264
rect 20079 -25940 21655 -25906
rect 20079 -26298 21655 -26264
rect 279 -26740 1855 -26706
rect 279 -27098 1855 -27064
rect 2479 -26740 4055 -26706
rect 2479 -27098 4055 -27064
rect 4679 -26740 6255 -26706
rect 4679 -27098 6255 -27064
rect 6879 -26740 8455 -26706
rect 6879 -27098 8455 -27064
rect 9079 -26740 10655 -26706
rect 9079 -27098 10655 -27064
rect 11279 -26740 12855 -26706
rect 11279 -27098 12855 -27064
rect 13479 -26740 15055 -26706
rect 13479 -27098 15055 -27064
rect 15679 -26740 17255 -26706
rect 15679 -27098 17255 -27064
rect 17879 -26740 19455 -26706
rect 17879 -27098 19455 -27064
rect 20079 -26740 21655 -26706
rect 20079 -27098 21655 -27064
rect 279 -27540 1855 -27506
rect 279 -27898 1855 -27864
rect 2479 -27540 4055 -27506
rect 2479 -27898 4055 -27864
rect 4679 -27540 6255 -27506
rect 4679 -27898 6255 -27864
rect 6879 -27540 8455 -27506
rect 6879 -27898 8455 -27864
rect 9079 -27540 10655 -27506
rect 9079 -27898 10655 -27864
rect 11279 -27540 12855 -27506
rect 11279 -27898 12855 -27864
rect 13479 -27540 15055 -27506
rect 13479 -27898 15055 -27864
rect 15679 -27540 17255 -27506
rect 15679 -27898 17255 -27864
rect 17879 -27540 19455 -27506
rect 17879 -27898 19455 -27864
rect 20079 -27540 21655 -27506
rect 20079 -27898 21655 -27864
rect 279 -28340 1855 -28306
rect 279 -28698 1855 -28664
rect 2479 -28340 4055 -28306
rect 2479 -28698 4055 -28664
rect 4679 -28340 6255 -28306
rect 4679 -28698 6255 -28664
rect 6879 -28340 8455 -28306
rect 6879 -28698 8455 -28664
rect 9079 -28340 10655 -28306
rect 9079 -28698 10655 -28664
rect 11279 -28340 12855 -28306
rect 11279 -28698 12855 -28664
rect 13479 -28340 15055 -28306
rect 13479 -28698 15055 -28664
rect 15679 -28340 17255 -28306
rect 15679 -28698 17255 -28664
rect 17879 -28340 19455 -28306
rect 17879 -28698 19455 -28664
rect 20079 -28340 21655 -28306
rect 20079 -28698 21655 -28664
rect 279 -29140 1855 -29106
rect 279 -29498 1855 -29464
rect 2479 -29140 4055 -29106
rect 2479 -29498 4055 -29464
rect 4679 -29140 6255 -29106
rect 4679 -29498 6255 -29464
rect 6879 -29140 8455 -29106
rect 6879 -29498 8455 -29464
rect 9079 -29140 10655 -29106
rect 9079 -29498 10655 -29464
rect 11279 -29140 12855 -29106
rect 11279 -29498 12855 -29464
rect 13479 -29140 15055 -29106
rect 13479 -29498 15055 -29464
rect 15679 -29140 17255 -29106
rect 15679 -29498 17255 -29464
rect 17879 -29140 19455 -29106
rect 17879 -29498 19455 -29464
rect 20079 -29140 21655 -29106
rect 20079 -29498 21655 -29464
rect 279 -29940 1855 -29906
rect 279 -30298 1855 -30264
rect 2479 -29940 4055 -29906
rect 2479 -30298 4055 -30264
rect 4679 -29940 6255 -29906
rect 4679 -30298 6255 -30264
rect 6879 -29940 8455 -29906
rect 6879 -30298 8455 -30264
rect 9079 -29940 10655 -29906
rect 9079 -30298 10655 -30264
rect 11279 -29940 12855 -29906
rect 11279 -30298 12855 -30264
rect 13479 -29940 15055 -29906
rect 13479 -30298 15055 -30264
rect 15679 -29940 17255 -29906
rect 15679 -30298 17255 -30264
rect 17879 -29940 19455 -29906
rect 17879 -30298 19455 -30264
rect 20079 -29940 21655 -29906
rect 20079 -30298 21655 -30264
rect 279 -30740 1855 -30706
rect 279 -31098 1855 -31064
rect 2479 -30740 4055 -30706
rect 2479 -31098 4055 -31064
rect 4679 -30740 6255 -30706
rect 4679 -31098 6255 -31064
rect 6879 -30740 8455 -30706
rect 6879 -31098 8455 -31064
rect 9079 -30740 10655 -30706
rect 9079 -31098 10655 -31064
rect 11279 -30740 12855 -30706
rect 11279 -31098 12855 -31064
rect 13479 -30740 15055 -30706
rect 13479 -31098 15055 -31064
rect 15679 -30740 17255 -30706
rect 15679 -31098 17255 -31064
rect 17879 -30740 19455 -30706
rect 17879 -31098 19455 -31064
rect 20079 -30740 21655 -30706
rect 20079 -31098 21655 -31064
rect 279 -31540 1855 -31506
rect 279 -31898 1855 -31864
rect 2479 -31540 4055 -31506
rect 2479 -31898 4055 -31864
rect 4679 -31540 6255 -31506
rect 4679 -31898 6255 -31864
rect 6879 -31540 8455 -31506
rect 6879 -31898 8455 -31864
rect 9079 -31540 10655 -31506
rect 9079 -31898 10655 -31864
rect 11279 -31540 12855 -31506
rect 11279 -31898 12855 -31864
rect 13479 -31540 15055 -31506
rect 13479 -31898 15055 -31864
rect 15679 -31540 17255 -31506
rect 15679 -31898 17255 -31864
rect 17879 -31540 19455 -31506
rect 17879 -31898 19455 -31864
rect 20079 -31540 21655 -31506
rect 20079 -31898 21655 -31864
rect 34989 -24864 35765 -24830
rect 34989 -25122 35765 -25088
rect 34989 -25380 35765 -25346
rect 34989 -25638 35765 -25604
rect 34989 -25896 35765 -25862
rect 34989 -26154 35765 -26120
rect 34989 -26412 35765 -26378
rect 34989 -26670 35765 -26636
rect 34989 -26928 35765 -26894
rect 36329 -24864 37105 -24830
rect 36329 -25122 37105 -25088
rect 36329 -25380 37105 -25346
rect 36329 -25638 37105 -25604
rect 36329 -25896 37105 -25862
rect 36329 -26154 37105 -26120
rect 36329 -26412 37105 -26378
rect 36329 -26670 37105 -26636
rect 36329 -26928 37105 -26894
rect 31812 -28909 31846 -28533
rect 31970 -28909 32004 -28533
rect 32252 -28909 32286 -28533
rect 32410 -28909 32444 -28533
rect 32692 -28909 32726 -28533
rect 32850 -28909 32884 -28533
rect 33106 -28909 33140 -28833
rect 33564 -28909 33598 -28833
rect 34012 -28909 34046 -28533
rect 34170 -28909 34204 -28533
rect 34452 -28909 34486 -28533
rect 34610 -28909 34644 -28533
rect 34892 -28909 34926 -28533
rect 35050 -28909 35084 -28533
rect 35306 -28909 35340 -28833
rect 35764 -28909 35798 -28833
rect 36212 -28909 36246 -28533
rect 36370 -28909 36404 -28533
rect 36652 -28909 36686 -28533
rect 36810 -28909 36844 -28533
rect 37092 -28909 37126 -28533
rect 37250 -28909 37284 -28533
rect 37506 -28909 37540 -28833
rect 37964 -28909 37998 -28833
rect 31824 -31191 31858 -31115
rect 32282 -31191 32316 -31115
rect 32538 -31491 32572 -31115
rect 32696 -31491 32730 -31115
rect 32978 -31491 33012 -31115
rect 33136 -31491 33170 -31115
rect 33418 -31491 33452 -31115
rect 33576 -31491 33610 -31115
rect 34024 -31191 34058 -31115
rect 34482 -31191 34516 -31115
rect 34738 -31491 34772 -31115
rect 34896 -31491 34930 -31115
rect 35178 -31491 35212 -31115
rect 35336 -31491 35370 -31115
rect 35618 -31491 35652 -31115
rect 35776 -31491 35810 -31115
rect 36224 -31191 36258 -31115
rect 36682 -31191 36716 -31115
rect 36938 -31491 36972 -31115
rect 37096 -31491 37130 -31115
rect 37378 -31491 37412 -31115
rect 37536 -31491 37570 -31115
rect 37818 -31491 37852 -31115
rect 37976 -31491 38010 -31115
<< psubdiff >>
rect 22236 11910 22332 11944
rect 26966 11910 27062 11944
rect 22236 11848 22270 11910
rect 27028 11848 27062 11910
rect 22236 4470 22270 4532
rect 34476 7470 34572 7504
rect 34730 7470 34826 7504
rect 34476 7408 34510 7470
rect 34792 7408 34826 7470
rect 34476 6990 34510 7052
rect 34792 6990 34826 7052
rect 34476 6956 34572 6990
rect 34730 6956 34826 6990
rect 34896 7470 34992 7504
rect 35150 7470 35246 7504
rect 34896 7408 34930 7470
rect 35212 7408 35246 7470
rect 34896 6990 34930 7052
rect 35212 6990 35246 7052
rect 34896 6956 34992 6990
rect 35150 6956 35246 6990
rect 35316 7470 35412 7504
rect 35570 7470 35666 7504
rect 35316 7408 35350 7470
rect 35632 7408 35666 7470
rect 35316 6990 35350 7052
rect 35632 6990 35666 7052
rect 35316 6956 35412 6990
rect 35570 6956 35666 6990
rect 27028 4470 27062 4532
rect 22236 4436 22332 4470
rect 26966 4436 27062 4470
<< nsubdiff >>
rect 32796 9008 32892 9042
rect 33478 9008 33574 9042
rect 32796 8946 32830 9008
rect 33540 8946 33574 9008
rect 32796 7910 32830 7972
rect 33540 7910 33574 7972
rect 32796 7876 32892 7910
rect 33478 7876 33574 7910
rect 33636 9008 33732 9042
rect 34318 9008 34414 9042
rect 33636 8946 33670 9008
rect 34380 8946 34414 9008
rect 33636 7910 33670 7972
rect 34476 8788 34572 8822
rect 34730 8788 34826 8822
rect 34476 8726 34510 8788
rect 34792 8726 34826 8788
rect 34476 8090 34510 8152
rect 34792 8090 34826 8152
rect 34476 8056 34572 8090
rect 34730 8056 34826 8090
rect 34896 8788 34992 8822
rect 35150 8788 35246 8822
rect 34896 8726 34930 8788
rect 35212 8726 35246 8788
rect 34896 8090 34930 8152
rect 35212 8090 35246 8152
rect 34896 8056 34992 8090
rect 35150 8056 35246 8090
rect 35316 8788 35412 8822
rect 35570 8788 35666 8822
rect 35316 8726 35350 8788
rect 35632 8726 35666 8788
rect 35316 8090 35350 8152
rect 35632 8090 35666 8152
rect 35316 8056 35412 8090
rect 35570 8056 35666 8090
rect 34380 7910 34414 7972
rect 33636 7876 33732 7910
rect 34318 7876 34414 7910
<< mvpsubdiff >>
rect 37 11909 2081 11921
rect 37 11875 145 11909
rect 1973 11875 2081 11909
rect 37 11863 2081 11875
rect 37 11813 95 11863
rect 37 11345 49 11813
rect 83 11345 95 11813
rect 2023 11813 2081 11863
rect 37 11295 95 11345
rect 2023 11345 2035 11813
rect 2069 11345 2081 11813
rect 2023 11295 2081 11345
rect 37 11283 2081 11295
rect 37 11249 145 11283
rect 1973 11249 2081 11283
rect 37 11237 2081 11249
rect 2237 11909 4281 11921
rect 2237 11875 2345 11909
rect 4173 11875 4281 11909
rect 2237 11863 4281 11875
rect 2237 11813 2295 11863
rect 2237 11345 2249 11813
rect 2283 11345 2295 11813
rect 4223 11813 4281 11863
rect 2237 11295 2295 11345
rect 4223 11345 4235 11813
rect 4269 11345 4281 11813
rect 4223 11295 4281 11345
rect 2237 11283 4281 11295
rect 2237 11249 2345 11283
rect 4173 11249 4281 11283
rect 2237 11237 4281 11249
rect 4437 11909 6481 11921
rect 4437 11875 4545 11909
rect 6373 11875 6481 11909
rect 4437 11863 6481 11875
rect 4437 11813 4495 11863
rect 4437 11345 4449 11813
rect 4483 11345 4495 11813
rect 6423 11813 6481 11863
rect 4437 11295 4495 11345
rect 6423 11345 6435 11813
rect 6469 11345 6481 11813
rect 6423 11295 6481 11345
rect 4437 11283 6481 11295
rect 4437 11249 4545 11283
rect 6373 11249 6481 11283
rect 4437 11237 6481 11249
rect 6637 11909 8681 11921
rect 6637 11875 6745 11909
rect 8573 11875 8681 11909
rect 6637 11863 8681 11875
rect 6637 11813 6695 11863
rect 6637 11345 6649 11813
rect 6683 11345 6695 11813
rect 8623 11813 8681 11863
rect 6637 11295 6695 11345
rect 8623 11345 8635 11813
rect 8669 11345 8681 11813
rect 8623 11295 8681 11345
rect 6637 11283 8681 11295
rect 6637 11249 6745 11283
rect 8573 11249 8681 11283
rect 6637 11237 8681 11249
rect 8837 11909 10881 11921
rect 8837 11875 8945 11909
rect 10773 11875 10881 11909
rect 8837 11863 10881 11875
rect 8837 11813 8895 11863
rect 8837 11345 8849 11813
rect 8883 11345 8895 11813
rect 10823 11813 10881 11863
rect 8837 11295 8895 11345
rect 10823 11345 10835 11813
rect 10869 11345 10881 11813
rect 10823 11295 10881 11345
rect 8837 11283 10881 11295
rect 8837 11249 8945 11283
rect 10773 11249 10881 11283
rect 8837 11237 10881 11249
rect 11037 11909 13081 11921
rect 11037 11875 11145 11909
rect 12973 11875 13081 11909
rect 11037 11863 13081 11875
rect 11037 11813 11095 11863
rect 11037 11345 11049 11813
rect 11083 11345 11095 11813
rect 13023 11813 13081 11863
rect 11037 11295 11095 11345
rect 13023 11345 13035 11813
rect 13069 11345 13081 11813
rect 13023 11295 13081 11345
rect 11037 11283 13081 11295
rect 11037 11249 11145 11283
rect 12973 11249 13081 11283
rect 11037 11237 13081 11249
rect 13237 11909 15281 11921
rect 13237 11875 13345 11909
rect 15173 11875 15281 11909
rect 13237 11863 15281 11875
rect 13237 11813 13295 11863
rect 13237 11345 13249 11813
rect 13283 11345 13295 11813
rect 15223 11813 15281 11863
rect 13237 11295 13295 11345
rect 15223 11345 15235 11813
rect 15269 11345 15281 11813
rect 15223 11295 15281 11345
rect 13237 11283 15281 11295
rect 13237 11249 13345 11283
rect 15173 11249 15281 11283
rect 13237 11237 15281 11249
rect 15437 11909 17481 11921
rect 15437 11875 15545 11909
rect 17373 11875 17481 11909
rect 15437 11863 17481 11875
rect 15437 11813 15495 11863
rect 15437 11345 15449 11813
rect 15483 11345 15495 11813
rect 17423 11813 17481 11863
rect 15437 11295 15495 11345
rect 17423 11345 17435 11813
rect 17469 11345 17481 11813
rect 17423 11295 17481 11345
rect 15437 11283 17481 11295
rect 15437 11249 15545 11283
rect 17373 11249 17481 11283
rect 15437 11237 17481 11249
rect 17637 11909 19681 11921
rect 17637 11875 17745 11909
rect 19573 11875 19681 11909
rect 17637 11863 19681 11875
rect 17637 11813 17695 11863
rect 17637 11345 17649 11813
rect 17683 11345 17695 11813
rect 19623 11813 19681 11863
rect 17637 11295 17695 11345
rect 19623 11345 19635 11813
rect 19669 11345 19681 11813
rect 19623 11295 19681 11345
rect 17637 11283 19681 11295
rect 17637 11249 17745 11283
rect 19573 11249 19681 11283
rect 17637 11237 19681 11249
rect 19837 11909 21881 11921
rect 19837 11875 19945 11909
rect 21773 11875 21881 11909
rect 19837 11863 21881 11875
rect 19837 11813 19895 11863
rect 19837 11345 19849 11813
rect 19883 11345 19895 11813
rect 21823 11813 21881 11863
rect 19837 11295 19895 11345
rect 21823 11345 21835 11813
rect 21869 11345 21881 11813
rect 21823 11295 21881 11345
rect 19837 11283 21881 11295
rect 19837 11249 19945 11283
rect 21773 11249 21881 11283
rect 19837 11237 21881 11249
rect 37 11109 2081 11121
rect 37 11075 145 11109
rect 1973 11075 2081 11109
rect 37 11063 2081 11075
rect 37 11013 95 11063
rect 37 10545 49 11013
rect 83 10545 95 11013
rect 2023 11013 2081 11063
rect 37 10495 95 10545
rect 2023 10545 2035 11013
rect 2069 10545 2081 11013
rect 2023 10495 2081 10545
rect 37 10483 2081 10495
rect 37 10449 145 10483
rect 1973 10449 2081 10483
rect 37 10437 2081 10449
rect 2236 11108 4280 11120
rect 2236 11074 2344 11108
rect 4172 11074 4280 11108
rect 2236 11062 4280 11074
rect 2236 11012 2294 11062
rect 2236 10544 2248 11012
rect 2282 10544 2294 11012
rect 4222 11012 4280 11062
rect 2236 10494 2294 10544
rect 4222 10544 4234 11012
rect 4268 10544 4280 11012
rect 4222 10494 4280 10544
rect 2236 10482 4280 10494
rect 2236 10448 2344 10482
rect 4172 10448 4280 10482
rect 2236 10436 4280 10448
rect 4436 11108 6480 11120
rect 4436 11074 4544 11108
rect 6372 11074 6480 11108
rect 4436 11062 6480 11074
rect 4436 11012 4494 11062
rect 4436 10544 4448 11012
rect 4482 10544 4494 11012
rect 6422 11012 6480 11062
rect 4436 10494 4494 10544
rect 6422 10544 6434 11012
rect 6468 10544 6480 11012
rect 6422 10494 6480 10544
rect 4436 10482 6480 10494
rect 4436 10448 4544 10482
rect 6372 10448 6480 10482
rect 4436 10436 6480 10448
rect 6636 11108 8680 11120
rect 6636 11074 6744 11108
rect 8572 11074 8680 11108
rect 6636 11062 8680 11074
rect 6636 11012 6694 11062
rect 6636 10544 6648 11012
rect 6682 10544 6694 11012
rect 8622 11012 8680 11062
rect 6636 10494 6694 10544
rect 8622 10544 8634 11012
rect 8668 10544 8680 11012
rect 8622 10494 8680 10544
rect 6636 10482 8680 10494
rect 6636 10448 6744 10482
rect 8572 10448 8680 10482
rect 6636 10436 8680 10448
rect 8836 11108 10880 11120
rect 8836 11074 8944 11108
rect 10772 11074 10880 11108
rect 8836 11062 10880 11074
rect 8836 11012 8894 11062
rect 8836 10544 8848 11012
rect 8882 10544 8894 11012
rect 10822 11012 10880 11062
rect 8836 10494 8894 10544
rect 10822 10544 10834 11012
rect 10868 10544 10880 11012
rect 10822 10494 10880 10544
rect 8836 10482 10880 10494
rect 8836 10448 8944 10482
rect 10772 10448 10880 10482
rect 8836 10436 10880 10448
rect 11036 11108 13080 11120
rect 11036 11074 11144 11108
rect 12972 11074 13080 11108
rect 11036 11062 13080 11074
rect 11036 11012 11094 11062
rect 11036 10544 11048 11012
rect 11082 10544 11094 11012
rect 13022 11012 13080 11062
rect 11036 10494 11094 10544
rect 13022 10544 13034 11012
rect 13068 10544 13080 11012
rect 13022 10494 13080 10544
rect 11036 10482 13080 10494
rect 11036 10448 11144 10482
rect 12972 10448 13080 10482
rect 11036 10436 13080 10448
rect 13236 11108 15280 11120
rect 13236 11074 13344 11108
rect 15172 11074 15280 11108
rect 13236 11062 15280 11074
rect 13236 11012 13294 11062
rect 13236 10544 13248 11012
rect 13282 10544 13294 11012
rect 15222 11012 15280 11062
rect 13236 10494 13294 10544
rect 15222 10544 15234 11012
rect 15268 10544 15280 11012
rect 15222 10494 15280 10544
rect 13236 10482 15280 10494
rect 13236 10448 13344 10482
rect 15172 10448 15280 10482
rect 13236 10436 15280 10448
rect 15436 11108 17480 11120
rect 15436 11074 15544 11108
rect 17372 11074 17480 11108
rect 15436 11062 17480 11074
rect 15436 11012 15494 11062
rect 15436 10544 15448 11012
rect 15482 10544 15494 11012
rect 17422 11012 17480 11062
rect 15436 10494 15494 10544
rect 17422 10544 17434 11012
rect 17468 10544 17480 11012
rect 17422 10494 17480 10544
rect 15436 10482 17480 10494
rect 15436 10448 15544 10482
rect 17372 10448 17480 10482
rect 15436 10436 17480 10448
rect 17636 11108 19680 11120
rect 17636 11074 17744 11108
rect 19572 11074 19680 11108
rect 17636 11062 19680 11074
rect 17636 11012 17694 11062
rect 17636 10544 17648 11012
rect 17682 10544 17694 11012
rect 19622 11012 19680 11062
rect 17636 10494 17694 10544
rect 19622 10544 19634 11012
rect 19668 10544 19680 11012
rect 19622 10494 19680 10544
rect 17636 10482 19680 10494
rect 17636 10448 17744 10482
rect 19572 10448 19680 10482
rect 17636 10436 19680 10448
rect 19837 11109 21881 11121
rect 19837 11075 19945 11109
rect 21773 11075 21881 11109
rect 19837 11063 21881 11075
rect 19837 11013 19895 11063
rect 19837 10545 19849 11013
rect 19883 10545 19895 11013
rect 21823 11013 21881 11063
rect 19837 10495 19895 10545
rect 21823 10545 21835 11013
rect 21869 10545 21881 11013
rect 21823 10495 21881 10545
rect 19837 10483 21881 10495
rect 19837 10449 19945 10483
rect 21773 10449 21881 10483
rect 19837 10437 21881 10449
rect 37 10309 2081 10321
rect 37 10275 145 10309
rect 1973 10275 2081 10309
rect 37 10263 2081 10275
rect 37 10213 95 10263
rect 37 9745 49 10213
rect 83 9745 95 10213
rect 2023 10213 2081 10263
rect 37 9695 95 9745
rect 2023 9745 2035 10213
rect 2069 9745 2081 10213
rect 2023 9695 2081 9745
rect 37 9683 2081 9695
rect 37 9649 145 9683
rect 1973 9649 2081 9683
rect 37 9637 2081 9649
rect 2236 10308 4280 10320
rect 2236 10274 2344 10308
rect 4172 10274 4280 10308
rect 2236 10262 4280 10274
rect 2236 10212 2294 10262
rect 2236 9744 2248 10212
rect 2282 9744 2294 10212
rect 4222 10212 4280 10262
rect 2236 9694 2294 9744
rect 4222 9744 4234 10212
rect 4268 9744 4280 10212
rect 4222 9694 4280 9744
rect 2236 9682 4280 9694
rect 2236 9648 2344 9682
rect 4172 9648 4280 9682
rect 2236 9636 4280 9648
rect 4436 10308 6480 10320
rect 4436 10274 4544 10308
rect 6372 10274 6480 10308
rect 4436 10262 6480 10274
rect 4436 10212 4494 10262
rect 4436 9744 4448 10212
rect 4482 9744 4494 10212
rect 6422 10212 6480 10262
rect 4436 9694 4494 9744
rect 6422 9744 6434 10212
rect 6468 9744 6480 10212
rect 6422 9694 6480 9744
rect 4436 9682 6480 9694
rect 4436 9648 4544 9682
rect 6372 9648 6480 9682
rect 4436 9636 6480 9648
rect 6636 10308 8680 10320
rect 6636 10274 6744 10308
rect 8572 10274 8680 10308
rect 6636 10262 8680 10274
rect 6636 10212 6694 10262
rect 6636 9744 6648 10212
rect 6682 9744 6694 10212
rect 8622 10212 8680 10262
rect 6636 9694 6694 9744
rect 8622 9744 8634 10212
rect 8668 9744 8680 10212
rect 8622 9694 8680 9744
rect 6636 9682 8680 9694
rect 6636 9648 6744 9682
rect 8572 9648 8680 9682
rect 6636 9636 8680 9648
rect 8836 10308 10880 10320
rect 8836 10274 8944 10308
rect 10772 10274 10880 10308
rect 8836 10262 10880 10274
rect 8836 10212 8894 10262
rect 8836 9744 8848 10212
rect 8882 9744 8894 10212
rect 10822 10212 10880 10262
rect 8836 9694 8894 9744
rect 10822 9744 10834 10212
rect 10868 9744 10880 10212
rect 10822 9694 10880 9744
rect 8836 9682 10880 9694
rect 8836 9648 8944 9682
rect 10772 9648 10880 9682
rect 8836 9636 10880 9648
rect 11036 10308 13080 10320
rect 11036 10274 11144 10308
rect 12972 10274 13080 10308
rect 11036 10262 13080 10274
rect 11036 10212 11094 10262
rect 11036 9744 11048 10212
rect 11082 9744 11094 10212
rect 13022 10212 13080 10262
rect 11036 9694 11094 9744
rect 13022 9744 13034 10212
rect 13068 9744 13080 10212
rect 13022 9694 13080 9744
rect 11036 9682 13080 9694
rect 11036 9648 11144 9682
rect 12972 9648 13080 9682
rect 11036 9636 13080 9648
rect 13236 10308 15280 10320
rect 13236 10274 13344 10308
rect 15172 10274 15280 10308
rect 13236 10262 15280 10274
rect 13236 10212 13294 10262
rect 13236 9744 13248 10212
rect 13282 9744 13294 10212
rect 15222 10212 15280 10262
rect 13236 9694 13294 9744
rect 15222 9744 15234 10212
rect 15268 9744 15280 10212
rect 15222 9694 15280 9744
rect 13236 9682 15280 9694
rect 13236 9648 13344 9682
rect 15172 9648 15280 9682
rect 13236 9636 15280 9648
rect 15436 10308 17480 10320
rect 15436 10274 15544 10308
rect 17372 10274 17480 10308
rect 15436 10262 17480 10274
rect 15436 10212 15494 10262
rect 15436 9744 15448 10212
rect 15482 9744 15494 10212
rect 17422 10212 17480 10262
rect 15436 9694 15494 9744
rect 17422 9744 17434 10212
rect 17468 9744 17480 10212
rect 17422 9694 17480 9744
rect 15436 9682 17480 9694
rect 15436 9648 15544 9682
rect 17372 9648 17480 9682
rect 15436 9636 17480 9648
rect 17636 10308 19680 10320
rect 17636 10274 17744 10308
rect 19572 10274 19680 10308
rect 17636 10262 19680 10274
rect 17636 10212 17694 10262
rect 17636 9744 17648 10212
rect 17682 9744 17694 10212
rect 19622 10212 19680 10262
rect 17636 9694 17694 9744
rect 19622 9744 19634 10212
rect 19668 9744 19680 10212
rect 19622 9694 19680 9744
rect 17636 9682 19680 9694
rect 17636 9648 17744 9682
rect 19572 9648 19680 9682
rect 17636 9636 19680 9648
rect 19837 10309 21881 10321
rect 19837 10275 19945 10309
rect 21773 10275 21881 10309
rect 19837 10263 21881 10275
rect 19837 10213 19895 10263
rect 19837 9745 19849 10213
rect 19883 9745 19895 10213
rect 21823 10213 21881 10263
rect 19837 9695 19895 9745
rect 21823 9745 21835 10213
rect 21869 9745 21881 10213
rect 21823 9695 21881 9745
rect 19837 9683 21881 9695
rect 19837 9649 19945 9683
rect 21773 9649 21881 9683
rect 19837 9637 21881 9649
rect 37 9509 2081 9521
rect 37 9475 145 9509
rect 1973 9475 2081 9509
rect 37 9463 2081 9475
rect 37 9413 95 9463
rect 37 8945 49 9413
rect 83 8945 95 9413
rect 2023 9413 2081 9463
rect 37 8895 95 8945
rect 2023 8945 2035 9413
rect 2069 8945 2081 9413
rect 2023 8895 2081 8945
rect 37 8883 2081 8895
rect 37 8849 145 8883
rect 1973 8849 2081 8883
rect 37 8837 2081 8849
rect 2236 9508 4280 9520
rect 2236 9474 2344 9508
rect 4172 9474 4280 9508
rect 2236 9462 4280 9474
rect 2236 9412 2294 9462
rect 2236 8944 2248 9412
rect 2282 8944 2294 9412
rect 4222 9412 4280 9462
rect 2236 8894 2294 8944
rect 4222 8944 4234 9412
rect 4268 8944 4280 9412
rect 4222 8894 4280 8944
rect 2236 8882 4280 8894
rect 2236 8848 2344 8882
rect 4172 8848 4280 8882
rect 2236 8836 4280 8848
rect 4436 9508 6480 9520
rect 4436 9474 4544 9508
rect 6372 9474 6480 9508
rect 4436 9462 6480 9474
rect 4436 9412 4494 9462
rect 4436 8944 4448 9412
rect 4482 8944 4494 9412
rect 6422 9412 6480 9462
rect 4436 8894 4494 8944
rect 6422 8944 6434 9412
rect 6468 8944 6480 9412
rect 6422 8894 6480 8944
rect 4436 8882 6480 8894
rect 4436 8848 4544 8882
rect 6372 8848 6480 8882
rect 4436 8836 6480 8848
rect 6636 9508 8680 9520
rect 6636 9474 6744 9508
rect 8572 9474 8680 9508
rect 6636 9462 8680 9474
rect 6636 9412 6694 9462
rect 6636 8944 6648 9412
rect 6682 8944 6694 9412
rect 8622 9412 8680 9462
rect 6636 8894 6694 8944
rect 8622 8944 8634 9412
rect 8668 8944 8680 9412
rect 8622 8894 8680 8944
rect 6636 8882 8680 8894
rect 6636 8848 6744 8882
rect 8572 8848 8680 8882
rect 6636 8836 8680 8848
rect 8836 9508 10880 9520
rect 8836 9474 8944 9508
rect 10772 9474 10880 9508
rect 8836 9462 10880 9474
rect 8836 9412 8894 9462
rect 8836 8944 8848 9412
rect 8882 8944 8894 9412
rect 10822 9412 10880 9462
rect 8836 8894 8894 8944
rect 10822 8944 10834 9412
rect 10868 8944 10880 9412
rect 10822 8894 10880 8944
rect 8836 8882 10880 8894
rect 8836 8848 8944 8882
rect 10772 8848 10880 8882
rect 8836 8836 10880 8848
rect 11036 9508 13080 9520
rect 11036 9474 11144 9508
rect 12972 9474 13080 9508
rect 11036 9462 13080 9474
rect 11036 9412 11094 9462
rect 11036 8944 11048 9412
rect 11082 8944 11094 9412
rect 13022 9412 13080 9462
rect 11036 8894 11094 8944
rect 13022 8944 13034 9412
rect 13068 8944 13080 9412
rect 13022 8894 13080 8944
rect 11036 8882 13080 8894
rect 11036 8848 11144 8882
rect 12972 8848 13080 8882
rect 11036 8836 13080 8848
rect 13236 9508 15280 9520
rect 13236 9474 13344 9508
rect 15172 9474 15280 9508
rect 13236 9462 15280 9474
rect 13236 9412 13294 9462
rect 13236 8944 13248 9412
rect 13282 8944 13294 9412
rect 15222 9412 15280 9462
rect 13236 8894 13294 8944
rect 15222 8944 15234 9412
rect 15268 8944 15280 9412
rect 15222 8894 15280 8944
rect 13236 8882 15280 8894
rect 13236 8848 13344 8882
rect 15172 8848 15280 8882
rect 13236 8836 15280 8848
rect 15436 9508 17480 9520
rect 15436 9474 15544 9508
rect 17372 9474 17480 9508
rect 15436 9462 17480 9474
rect 15436 9412 15494 9462
rect 15436 8944 15448 9412
rect 15482 8944 15494 9412
rect 17422 9412 17480 9462
rect 15436 8894 15494 8944
rect 17422 8944 17434 9412
rect 17468 8944 17480 9412
rect 17422 8894 17480 8944
rect 15436 8882 17480 8894
rect 15436 8848 15544 8882
rect 17372 8848 17480 8882
rect 15436 8836 17480 8848
rect 17636 9508 19680 9520
rect 17636 9474 17744 9508
rect 19572 9474 19680 9508
rect 17636 9462 19680 9474
rect 17636 9412 17694 9462
rect 17636 8944 17648 9412
rect 17682 8944 17694 9412
rect 19622 9412 19680 9462
rect 17636 8894 17694 8944
rect 19622 8944 19634 9412
rect 19668 8944 19680 9412
rect 19622 8894 19680 8944
rect 17636 8882 19680 8894
rect 17636 8848 17744 8882
rect 19572 8848 19680 8882
rect 17636 8836 19680 8848
rect 19837 9509 21881 9521
rect 19837 9475 19945 9509
rect 21773 9475 21881 9509
rect 19837 9463 21881 9475
rect 19837 9413 19895 9463
rect 19837 8945 19849 9413
rect 19883 8945 19895 9413
rect 21823 9413 21881 9463
rect 19837 8895 19895 8945
rect 21823 8945 21835 9413
rect 21869 8945 21881 9413
rect 21823 8895 21881 8945
rect 19837 8883 21881 8895
rect 19837 8849 19945 8883
rect 21773 8849 21881 8883
rect 19837 8837 21881 8849
rect 37 8709 2081 8721
rect 37 8675 145 8709
rect 1973 8675 2081 8709
rect 37 8663 2081 8675
rect 37 8613 95 8663
rect 37 8145 49 8613
rect 83 8145 95 8613
rect 2023 8613 2081 8663
rect 37 8095 95 8145
rect 2023 8145 2035 8613
rect 2069 8145 2081 8613
rect 2023 8095 2081 8145
rect 37 8083 2081 8095
rect 37 8049 145 8083
rect 1973 8049 2081 8083
rect 37 8037 2081 8049
rect 2236 8708 4280 8720
rect 2236 8674 2344 8708
rect 4172 8674 4280 8708
rect 2236 8662 4280 8674
rect 2236 8612 2294 8662
rect 2236 8144 2248 8612
rect 2282 8144 2294 8612
rect 4222 8612 4280 8662
rect 2236 8094 2294 8144
rect 4222 8144 4234 8612
rect 4268 8144 4280 8612
rect 4222 8094 4280 8144
rect 2236 8082 4280 8094
rect 2236 8048 2344 8082
rect 4172 8048 4280 8082
rect 2236 8036 4280 8048
rect 4436 8708 6480 8720
rect 4436 8674 4544 8708
rect 6372 8674 6480 8708
rect 4436 8662 6480 8674
rect 4436 8612 4494 8662
rect 4436 8144 4448 8612
rect 4482 8144 4494 8612
rect 6422 8612 6480 8662
rect 4436 8094 4494 8144
rect 6422 8144 6434 8612
rect 6468 8144 6480 8612
rect 6422 8094 6480 8144
rect 4436 8082 6480 8094
rect 4436 8048 4544 8082
rect 6372 8048 6480 8082
rect 4436 8036 6480 8048
rect 6636 8708 8680 8720
rect 6636 8674 6744 8708
rect 8572 8674 8680 8708
rect 6636 8662 8680 8674
rect 6636 8612 6694 8662
rect 6636 8144 6648 8612
rect 6682 8144 6694 8612
rect 8622 8612 8680 8662
rect 6636 8094 6694 8144
rect 8622 8144 8634 8612
rect 8668 8144 8680 8612
rect 8622 8094 8680 8144
rect 6636 8082 8680 8094
rect 6636 8048 6744 8082
rect 8572 8048 8680 8082
rect 6636 8036 8680 8048
rect 8836 8708 10880 8720
rect 8836 8674 8944 8708
rect 10772 8674 10880 8708
rect 8836 8662 10880 8674
rect 8836 8612 8894 8662
rect 8836 8144 8848 8612
rect 8882 8144 8894 8612
rect 10822 8612 10880 8662
rect 8836 8094 8894 8144
rect 10822 8144 10834 8612
rect 10868 8144 10880 8612
rect 10822 8094 10880 8144
rect 8836 8082 10880 8094
rect 8836 8048 8944 8082
rect 10772 8048 10880 8082
rect 8836 8036 10880 8048
rect 11036 8708 13080 8720
rect 11036 8674 11144 8708
rect 12972 8674 13080 8708
rect 11036 8662 13080 8674
rect 11036 8612 11094 8662
rect 11036 8144 11048 8612
rect 11082 8144 11094 8612
rect 13022 8612 13080 8662
rect 11036 8094 11094 8144
rect 13022 8144 13034 8612
rect 13068 8144 13080 8612
rect 13022 8094 13080 8144
rect 11036 8082 13080 8094
rect 11036 8048 11144 8082
rect 12972 8048 13080 8082
rect 11036 8036 13080 8048
rect 13236 8708 15280 8720
rect 13236 8674 13344 8708
rect 15172 8674 15280 8708
rect 13236 8662 15280 8674
rect 13236 8612 13294 8662
rect 13236 8144 13248 8612
rect 13282 8144 13294 8612
rect 15222 8612 15280 8662
rect 13236 8094 13294 8144
rect 15222 8144 15234 8612
rect 15268 8144 15280 8612
rect 15222 8094 15280 8144
rect 13236 8082 15280 8094
rect 13236 8048 13344 8082
rect 15172 8048 15280 8082
rect 13236 8036 15280 8048
rect 15436 8708 17480 8720
rect 15436 8674 15544 8708
rect 17372 8674 17480 8708
rect 15436 8662 17480 8674
rect 15436 8612 15494 8662
rect 15436 8144 15448 8612
rect 15482 8144 15494 8612
rect 17422 8612 17480 8662
rect 15436 8094 15494 8144
rect 17422 8144 17434 8612
rect 17468 8144 17480 8612
rect 17422 8094 17480 8144
rect 15436 8082 17480 8094
rect 15436 8048 15544 8082
rect 17372 8048 17480 8082
rect 15436 8036 17480 8048
rect 17636 8708 19680 8720
rect 17636 8674 17744 8708
rect 19572 8674 19680 8708
rect 17636 8662 19680 8674
rect 17636 8612 17694 8662
rect 17636 8144 17648 8612
rect 17682 8144 17694 8612
rect 19622 8612 19680 8662
rect 17636 8094 17694 8144
rect 19622 8144 19634 8612
rect 19668 8144 19680 8612
rect 19622 8094 19680 8144
rect 17636 8082 19680 8094
rect 17636 8048 17744 8082
rect 19572 8048 19680 8082
rect 17636 8036 19680 8048
rect 19837 8709 21881 8721
rect 19837 8675 19945 8709
rect 21773 8675 21881 8709
rect 19837 8663 21881 8675
rect 19837 8613 19895 8663
rect 19837 8145 19849 8613
rect 19883 8145 19895 8613
rect 21823 8613 21881 8663
rect 19837 8095 19895 8145
rect 21823 8145 21835 8613
rect 21869 8145 21881 8613
rect 21823 8095 21881 8145
rect 19837 8083 21881 8095
rect 19837 8049 19945 8083
rect 21773 8049 21881 8083
rect 19837 8037 21881 8049
rect 37 7909 2081 7921
rect 37 7875 145 7909
rect 1973 7875 2081 7909
rect 37 7863 2081 7875
rect 37 7813 95 7863
rect 37 7345 49 7813
rect 83 7345 95 7813
rect 2023 7813 2081 7863
rect 37 7295 95 7345
rect 2023 7345 2035 7813
rect 2069 7345 2081 7813
rect 2023 7295 2081 7345
rect 37 7283 2081 7295
rect 37 7249 145 7283
rect 1973 7249 2081 7283
rect 37 7237 2081 7249
rect 2236 7908 4280 7920
rect 2236 7874 2344 7908
rect 4172 7874 4280 7908
rect 2236 7862 4280 7874
rect 2236 7812 2294 7862
rect 2236 7344 2248 7812
rect 2282 7344 2294 7812
rect 4222 7812 4280 7862
rect 2236 7294 2294 7344
rect 4222 7344 4234 7812
rect 4268 7344 4280 7812
rect 4222 7294 4280 7344
rect 2236 7282 4280 7294
rect 2236 7248 2344 7282
rect 4172 7248 4280 7282
rect 2236 7236 4280 7248
rect 4436 7908 6480 7920
rect 4436 7874 4544 7908
rect 6372 7874 6480 7908
rect 4436 7862 6480 7874
rect 4436 7812 4494 7862
rect 4436 7344 4448 7812
rect 4482 7344 4494 7812
rect 6422 7812 6480 7862
rect 4436 7294 4494 7344
rect 6422 7344 6434 7812
rect 6468 7344 6480 7812
rect 6422 7294 6480 7344
rect 4436 7282 6480 7294
rect 4436 7248 4544 7282
rect 6372 7248 6480 7282
rect 4436 7236 6480 7248
rect 6636 7908 8680 7920
rect 6636 7874 6744 7908
rect 8572 7874 8680 7908
rect 6636 7862 8680 7874
rect 6636 7812 6694 7862
rect 6636 7344 6648 7812
rect 6682 7344 6694 7812
rect 8622 7812 8680 7862
rect 6636 7294 6694 7344
rect 8622 7344 8634 7812
rect 8668 7344 8680 7812
rect 8622 7294 8680 7344
rect 6636 7282 8680 7294
rect 6636 7248 6744 7282
rect 8572 7248 8680 7282
rect 6636 7236 8680 7248
rect 8836 7908 10880 7920
rect 8836 7874 8944 7908
rect 10772 7874 10880 7908
rect 8836 7862 10880 7874
rect 8836 7812 8894 7862
rect 8836 7344 8848 7812
rect 8882 7344 8894 7812
rect 10822 7812 10880 7862
rect 8836 7294 8894 7344
rect 10822 7344 10834 7812
rect 10868 7344 10880 7812
rect 10822 7294 10880 7344
rect 8836 7282 10880 7294
rect 8836 7248 8944 7282
rect 10772 7248 10880 7282
rect 8836 7236 10880 7248
rect 11036 7908 13080 7920
rect 11036 7874 11144 7908
rect 12972 7874 13080 7908
rect 11036 7862 13080 7874
rect 11036 7812 11094 7862
rect 11036 7344 11048 7812
rect 11082 7344 11094 7812
rect 13022 7812 13080 7862
rect 11036 7294 11094 7344
rect 13022 7344 13034 7812
rect 13068 7344 13080 7812
rect 13022 7294 13080 7344
rect 11036 7282 13080 7294
rect 11036 7248 11144 7282
rect 12972 7248 13080 7282
rect 11036 7236 13080 7248
rect 13236 7908 15280 7920
rect 13236 7874 13344 7908
rect 15172 7874 15280 7908
rect 13236 7862 15280 7874
rect 13236 7812 13294 7862
rect 13236 7344 13248 7812
rect 13282 7344 13294 7812
rect 15222 7812 15280 7862
rect 13236 7294 13294 7344
rect 15222 7344 15234 7812
rect 15268 7344 15280 7812
rect 15222 7294 15280 7344
rect 13236 7282 15280 7294
rect 13236 7248 13344 7282
rect 15172 7248 15280 7282
rect 13236 7236 15280 7248
rect 15436 7908 17480 7920
rect 15436 7874 15544 7908
rect 17372 7874 17480 7908
rect 15436 7862 17480 7874
rect 15436 7812 15494 7862
rect 15436 7344 15448 7812
rect 15482 7344 15494 7812
rect 17422 7812 17480 7862
rect 15436 7294 15494 7344
rect 17422 7344 17434 7812
rect 17468 7344 17480 7812
rect 17422 7294 17480 7344
rect 15436 7282 17480 7294
rect 15436 7248 15544 7282
rect 17372 7248 17480 7282
rect 15436 7236 17480 7248
rect 17636 7908 19680 7920
rect 17636 7874 17744 7908
rect 19572 7874 19680 7908
rect 17636 7862 19680 7874
rect 17636 7812 17694 7862
rect 17636 7344 17648 7812
rect 17682 7344 17694 7812
rect 19622 7812 19680 7862
rect 17636 7294 17694 7344
rect 19622 7344 19634 7812
rect 19668 7344 19680 7812
rect 19622 7294 19680 7344
rect 17636 7282 19680 7294
rect 17636 7248 17744 7282
rect 19572 7248 19680 7282
rect 17636 7236 19680 7248
rect 19837 7909 21881 7921
rect 19837 7875 19945 7909
rect 21773 7875 21881 7909
rect 19837 7863 21881 7875
rect 19837 7813 19895 7863
rect 19837 7345 19849 7813
rect 19883 7345 19895 7813
rect 21823 7813 21881 7863
rect 19837 7295 19895 7345
rect 21823 7345 21835 7813
rect 21869 7345 21881 7813
rect 21823 7295 21881 7345
rect 19837 7283 21881 7295
rect 19837 7249 19945 7283
rect 21773 7249 21881 7283
rect 19837 7237 21881 7249
rect 37 7109 2081 7121
rect 37 7075 145 7109
rect 1973 7075 2081 7109
rect 37 7063 2081 7075
rect 37 7013 95 7063
rect 37 6545 49 7013
rect 83 6545 95 7013
rect 2023 7013 2081 7063
rect 37 6495 95 6545
rect 2023 6545 2035 7013
rect 2069 6545 2081 7013
rect 2023 6495 2081 6545
rect 37 6483 2081 6495
rect 37 6449 145 6483
rect 1973 6449 2081 6483
rect 37 6437 2081 6449
rect 2236 7108 4280 7120
rect 2236 7074 2344 7108
rect 4172 7074 4280 7108
rect 2236 7062 4280 7074
rect 2236 7012 2294 7062
rect 2236 6544 2248 7012
rect 2282 6544 2294 7012
rect 4222 7012 4280 7062
rect 2236 6494 2294 6544
rect 4222 6544 4234 7012
rect 4268 6544 4280 7012
rect 4222 6494 4280 6544
rect 2236 6482 4280 6494
rect 2236 6448 2344 6482
rect 4172 6448 4280 6482
rect 2236 6436 4280 6448
rect 4436 7108 6480 7120
rect 4436 7074 4544 7108
rect 6372 7074 6480 7108
rect 4436 7062 6480 7074
rect 4436 7012 4494 7062
rect 4436 6544 4448 7012
rect 4482 6544 4494 7012
rect 6422 7012 6480 7062
rect 4436 6494 4494 6544
rect 6422 6544 6434 7012
rect 6468 6544 6480 7012
rect 6422 6494 6480 6544
rect 4436 6482 6480 6494
rect 4436 6448 4544 6482
rect 6372 6448 6480 6482
rect 4436 6436 6480 6448
rect 6636 7108 8680 7120
rect 6636 7074 6744 7108
rect 8572 7074 8680 7108
rect 6636 7062 8680 7074
rect 6636 7012 6694 7062
rect 6636 6544 6648 7012
rect 6682 6544 6694 7012
rect 8622 7012 8680 7062
rect 6636 6494 6694 6544
rect 8622 6544 8634 7012
rect 8668 6544 8680 7012
rect 8622 6494 8680 6544
rect 6636 6482 8680 6494
rect 6636 6448 6744 6482
rect 8572 6448 8680 6482
rect 6636 6436 8680 6448
rect 8836 7108 10880 7120
rect 8836 7074 8944 7108
rect 10772 7074 10880 7108
rect 8836 7062 10880 7074
rect 8836 7012 8894 7062
rect 8836 6544 8848 7012
rect 8882 6544 8894 7012
rect 10822 7012 10880 7062
rect 8836 6494 8894 6544
rect 10822 6544 10834 7012
rect 10868 6544 10880 7012
rect 10822 6494 10880 6544
rect 8836 6482 10880 6494
rect 8836 6448 8944 6482
rect 10772 6448 10880 6482
rect 8836 6436 10880 6448
rect 11036 7108 13080 7120
rect 11036 7074 11144 7108
rect 12972 7074 13080 7108
rect 11036 7062 13080 7074
rect 11036 7012 11094 7062
rect 11036 6544 11048 7012
rect 11082 6544 11094 7012
rect 13022 7012 13080 7062
rect 11036 6494 11094 6544
rect 13022 6544 13034 7012
rect 13068 6544 13080 7012
rect 13022 6494 13080 6544
rect 11036 6482 13080 6494
rect 11036 6448 11144 6482
rect 12972 6448 13080 6482
rect 11036 6436 13080 6448
rect 13236 7108 15280 7120
rect 13236 7074 13344 7108
rect 15172 7074 15280 7108
rect 13236 7062 15280 7074
rect 13236 7012 13294 7062
rect 13236 6544 13248 7012
rect 13282 6544 13294 7012
rect 15222 7012 15280 7062
rect 13236 6494 13294 6544
rect 15222 6544 15234 7012
rect 15268 6544 15280 7012
rect 15222 6494 15280 6544
rect 13236 6482 15280 6494
rect 13236 6448 13344 6482
rect 15172 6448 15280 6482
rect 13236 6436 15280 6448
rect 15436 7108 17480 7120
rect 15436 7074 15544 7108
rect 17372 7074 17480 7108
rect 15436 7062 17480 7074
rect 15436 7012 15494 7062
rect 15436 6544 15448 7012
rect 15482 6544 15494 7012
rect 17422 7012 17480 7062
rect 15436 6494 15494 6544
rect 17422 6544 17434 7012
rect 17468 6544 17480 7012
rect 17422 6494 17480 6544
rect 15436 6482 17480 6494
rect 15436 6448 15544 6482
rect 17372 6448 17480 6482
rect 15436 6436 17480 6448
rect 17636 7108 19680 7120
rect 17636 7074 17744 7108
rect 19572 7074 19680 7108
rect 17636 7062 19680 7074
rect 17636 7012 17694 7062
rect 17636 6544 17648 7012
rect 17682 6544 17694 7012
rect 19622 7012 19680 7062
rect 17636 6494 17694 6544
rect 19622 6544 19634 7012
rect 19668 6544 19680 7012
rect 19622 6494 19680 6544
rect 17636 6482 19680 6494
rect 17636 6448 17744 6482
rect 19572 6448 19680 6482
rect 17636 6436 19680 6448
rect 19837 7109 21881 7121
rect 19837 7075 19945 7109
rect 21773 7075 21881 7109
rect 19837 7063 21881 7075
rect 19837 7013 19895 7063
rect 19837 6545 19849 7013
rect 19883 6545 19895 7013
rect 21823 7013 21881 7063
rect 19837 6495 19895 6545
rect 21823 6545 21835 7013
rect 21869 6545 21881 7013
rect 21823 6495 21881 6545
rect 19837 6483 21881 6495
rect 19837 6449 19945 6483
rect 21773 6449 21881 6483
rect 19837 6437 21881 6449
rect 37 6309 2081 6321
rect 37 6275 145 6309
rect 1973 6275 2081 6309
rect 37 6263 2081 6275
rect 37 6213 95 6263
rect 37 5745 49 6213
rect 83 5745 95 6213
rect 2023 6213 2081 6263
rect 37 5695 95 5745
rect 2023 5745 2035 6213
rect 2069 5745 2081 6213
rect 2023 5695 2081 5745
rect 37 5683 2081 5695
rect 37 5649 145 5683
rect 1973 5649 2081 5683
rect 37 5637 2081 5649
rect 2236 6308 4280 6320
rect 2236 6274 2344 6308
rect 4172 6274 4280 6308
rect 2236 6262 4280 6274
rect 2236 6212 2294 6262
rect 2236 5744 2248 6212
rect 2282 5744 2294 6212
rect 4222 6212 4280 6262
rect 2236 5694 2294 5744
rect 4222 5744 4234 6212
rect 4268 5744 4280 6212
rect 4222 5694 4280 5744
rect 2236 5682 4280 5694
rect 2236 5648 2344 5682
rect 4172 5648 4280 5682
rect 2236 5636 4280 5648
rect 4436 6308 6480 6320
rect 4436 6274 4544 6308
rect 6372 6274 6480 6308
rect 4436 6262 6480 6274
rect 4436 6212 4494 6262
rect 4436 5744 4448 6212
rect 4482 5744 4494 6212
rect 6422 6212 6480 6262
rect 4436 5694 4494 5744
rect 6422 5744 6434 6212
rect 6468 5744 6480 6212
rect 6422 5694 6480 5744
rect 4436 5682 6480 5694
rect 4436 5648 4544 5682
rect 6372 5648 6480 5682
rect 4436 5636 6480 5648
rect 6636 6308 8680 6320
rect 6636 6274 6744 6308
rect 8572 6274 8680 6308
rect 6636 6262 8680 6274
rect 6636 6212 6694 6262
rect 6636 5744 6648 6212
rect 6682 5744 6694 6212
rect 8622 6212 8680 6262
rect 6636 5694 6694 5744
rect 8622 5744 8634 6212
rect 8668 5744 8680 6212
rect 8622 5694 8680 5744
rect 6636 5682 8680 5694
rect 6636 5648 6744 5682
rect 8572 5648 8680 5682
rect 6636 5636 8680 5648
rect 8836 6308 10880 6320
rect 8836 6274 8944 6308
rect 10772 6274 10880 6308
rect 8836 6262 10880 6274
rect 8836 6212 8894 6262
rect 8836 5744 8848 6212
rect 8882 5744 8894 6212
rect 10822 6212 10880 6262
rect 8836 5694 8894 5744
rect 10822 5744 10834 6212
rect 10868 5744 10880 6212
rect 10822 5694 10880 5744
rect 8836 5682 10880 5694
rect 8836 5648 8944 5682
rect 10772 5648 10880 5682
rect 8836 5636 10880 5648
rect 11036 6308 13080 6320
rect 11036 6274 11144 6308
rect 12972 6274 13080 6308
rect 11036 6262 13080 6274
rect 11036 6212 11094 6262
rect 11036 5744 11048 6212
rect 11082 5744 11094 6212
rect 13022 6212 13080 6262
rect 11036 5694 11094 5744
rect 13022 5744 13034 6212
rect 13068 5744 13080 6212
rect 13022 5694 13080 5744
rect 11036 5682 13080 5694
rect 11036 5648 11144 5682
rect 12972 5648 13080 5682
rect 11036 5636 13080 5648
rect 13236 6308 15280 6320
rect 13236 6274 13344 6308
rect 15172 6274 15280 6308
rect 13236 6262 15280 6274
rect 13236 6212 13294 6262
rect 13236 5744 13248 6212
rect 13282 5744 13294 6212
rect 15222 6212 15280 6262
rect 13236 5694 13294 5744
rect 15222 5744 15234 6212
rect 15268 5744 15280 6212
rect 15222 5694 15280 5744
rect 13236 5682 15280 5694
rect 13236 5648 13344 5682
rect 15172 5648 15280 5682
rect 13236 5636 15280 5648
rect 15436 6308 17480 6320
rect 15436 6274 15544 6308
rect 17372 6274 17480 6308
rect 15436 6262 17480 6274
rect 15436 6212 15494 6262
rect 15436 5744 15448 6212
rect 15482 5744 15494 6212
rect 17422 6212 17480 6262
rect 15436 5694 15494 5744
rect 17422 5744 17434 6212
rect 17468 5744 17480 6212
rect 17422 5694 17480 5744
rect 15436 5682 17480 5694
rect 15436 5648 15544 5682
rect 17372 5648 17480 5682
rect 15436 5636 17480 5648
rect 17636 6308 19680 6320
rect 17636 6274 17744 6308
rect 19572 6274 19680 6308
rect 17636 6262 19680 6274
rect 17636 6212 17694 6262
rect 17636 5744 17648 6212
rect 17682 5744 17694 6212
rect 19622 6212 19680 6262
rect 17636 5694 17694 5744
rect 19622 5744 19634 6212
rect 19668 5744 19680 6212
rect 19622 5694 19680 5744
rect 17636 5682 19680 5694
rect 17636 5648 17744 5682
rect 19572 5648 19680 5682
rect 17636 5636 19680 5648
rect 19837 6309 21881 6321
rect 19837 6275 19945 6309
rect 21773 6275 21881 6309
rect 19837 6263 21881 6275
rect 19837 6213 19895 6263
rect 19837 5745 19849 6213
rect 19883 5745 19895 6213
rect 21823 6213 21881 6263
rect 19837 5695 19895 5745
rect 21823 5745 21835 6213
rect 21869 5745 21881 6213
rect 21823 5695 21881 5745
rect 19837 5683 21881 5695
rect 19837 5649 19945 5683
rect 21773 5649 21881 5683
rect 19837 5637 21881 5649
rect 37 5509 2081 5521
rect 37 5475 145 5509
rect 1973 5475 2081 5509
rect 37 5463 2081 5475
rect 37 5413 95 5463
rect 37 4945 49 5413
rect 83 4945 95 5413
rect 2023 5413 2081 5463
rect 37 4895 95 4945
rect 2023 4945 2035 5413
rect 2069 4945 2081 5413
rect 2023 4895 2081 4945
rect 37 4883 2081 4895
rect 37 4849 145 4883
rect 1973 4849 2081 4883
rect 37 4837 2081 4849
rect 2236 5508 4280 5520
rect 2236 5474 2344 5508
rect 4172 5474 4280 5508
rect 2236 5462 4280 5474
rect 2236 5412 2294 5462
rect 2236 4944 2248 5412
rect 2282 4944 2294 5412
rect 4222 5412 4280 5462
rect 2236 4894 2294 4944
rect 4222 4944 4234 5412
rect 4268 4944 4280 5412
rect 4222 4894 4280 4944
rect 2236 4882 4280 4894
rect 2236 4848 2344 4882
rect 4172 4848 4280 4882
rect 2236 4836 4280 4848
rect 4436 5508 6480 5520
rect 4436 5474 4544 5508
rect 6372 5474 6480 5508
rect 4436 5462 6480 5474
rect 4436 5412 4494 5462
rect 4436 4944 4448 5412
rect 4482 4944 4494 5412
rect 6422 5412 6480 5462
rect 4436 4894 4494 4944
rect 6422 4944 6434 5412
rect 6468 4944 6480 5412
rect 6422 4894 6480 4944
rect 4436 4882 6480 4894
rect 4436 4848 4544 4882
rect 6372 4848 6480 4882
rect 4436 4836 6480 4848
rect 6636 5508 8680 5520
rect 6636 5474 6744 5508
rect 8572 5474 8680 5508
rect 6636 5462 8680 5474
rect 6636 5412 6694 5462
rect 6636 4944 6648 5412
rect 6682 4944 6694 5412
rect 8622 5412 8680 5462
rect 6636 4894 6694 4944
rect 8622 4944 8634 5412
rect 8668 4944 8680 5412
rect 8622 4894 8680 4944
rect 6636 4882 8680 4894
rect 6636 4848 6744 4882
rect 8572 4848 8680 4882
rect 6636 4836 8680 4848
rect 8836 5508 10880 5520
rect 8836 5474 8944 5508
rect 10772 5474 10880 5508
rect 8836 5462 10880 5474
rect 8836 5412 8894 5462
rect 8836 4944 8848 5412
rect 8882 4944 8894 5412
rect 10822 5412 10880 5462
rect 8836 4894 8894 4944
rect 10822 4944 10834 5412
rect 10868 4944 10880 5412
rect 10822 4894 10880 4944
rect 8836 4882 10880 4894
rect 8836 4848 8944 4882
rect 10772 4848 10880 4882
rect 8836 4836 10880 4848
rect 11036 5508 13080 5520
rect 11036 5474 11144 5508
rect 12972 5474 13080 5508
rect 11036 5462 13080 5474
rect 11036 5412 11094 5462
rect 11036 4944 11048 5412
rect 11082 4944 11094 5412
rect 13022 5412 13080 5462
rect 11036 4894 11094 4944
rect 13022 4944 13034 5412
rect 13068 4944 13080 5412
rect 13022 4894 13080 4944
rect 11036 4882 13080 4894
rect 11036 4848 11144 4882
rect 12972 4848 13080 4882
rect 11036 4836 13080 4848
rect 13236 5508 15280 5520
rect 13236 5474 13344 5508
rect 15172 5474 15280 5508
rect 13236 5462 15280 5474
rect 13236 5412 13294 5462
rect 13236 4944 13248 5412
rect 13282 4944 13294 5412
rect 15222 5412 15280 5462
rect 13236 4894 13294 4944
rect 15222 4944 15234 5412
rect 15268 4944 15280 5412
rect 15222 4894 15280 4944
rect 13236 4882 15280 4894
rect 13236 4848 13344 4882
rect 15172 4848 15280 4882
rect 13236 4836 15280 4848
rect 15436 5508 17480 5520
rect 15436 5474 15544 5508
rect 17372 5474 17480 5508
rect 15436 5462 17480 5474
rect 15436 5412 15494 5462
rect 15436 4944 15448 5412
rect 15482 4944 15494 5412
rect 17422 5412 17480 5462
rect 15436 4894 15494 4944
rect 17422 4944 17434 5412
rect 17468 4944 17480 5412
rect 17422 4894 17480 4944
rect 15436 4882 17480 4894
rect 15436 4848 15544 4882
rect 17372 4848 17480 4882
rect 15436 4836 17480 4848
rect 17636 5508 19680 5520
rect 17636 5474 17744 5508
rect 19572 5474 19680 5508
rect 17636 5462 19680 5474
rect 17636 5412 17694 5462
rect 17636 4944 17648 5412
rect 17682 4944 17694 5412
rect 19622 5412 19680 5462
rect 17636 4894 17694 4944
rect 19622 4944 19634 5412
rect 19668 4944 19680 5412
rect 19622 4894 19680 4944
rect 17636 4882 19680 4894
rect 17636 4848 17744 4882
rect 19572 4848 19680 4882
rect 17636 4836 19680 4848
rect 19837 5509 21881 5521
rect 19837 5475 19945 5509
rect 21773 5475 21881 5509
rect 19837 5463 21881 5475
rect 19837 5413 19895 5463
rect 19837 4945 19849 5413
rect 19883 4945 19895 5413
rect 21823 5413 21881 5463
rect 19837 4895 19895 4945
rect 21823 4945 21835 5413
rect 21869 4945 21881 5413
rect 21823 4895 21881 4945
rect 19837 4883 21881 4895
rect 19837 4849 19945 4883
rect 21773 4849 21881 4883
rect 19837 4837 21881 4849
rect 37 4709 2081 4721
rect 37 4675 145 4709
rect 1973 4675 2081 4709
rect 37 4663 2081 4675
rect 37 4613 95 4663
rect 37 4145 49 4613
rect 83 4145 95 4613
rect 2023 4613 2081 4663
rect 37 4095 95 4145
rect 2023 4145 2035 4613
rect 2069 4145 2081 4613
rect 2023 4095 2081 4145
rect 37 4083 2081 4095
rect 37 4049 145 4083
rect 1973 4049 2081 4083
rect 37 4037 2081 4049
rect 2237 4709 4281 4721
rect 2237 4675 2345 4709
rect 4173 4675 4281 4709
rect 2237 4663 4281 4675
rect 2237 4613 2295 4663
rect 2237 4145 2249 4613
rect 2283 4145 2295 4613
rect 4223 4613 4281 4663
rect 2237 4095 2295 4145
rect 4223 4145 4235 4613
rect 4269 4145 4281 4613
rect 4223 4095 4281 4145
rect 2237 4083 4281 4095
rect 2237 4049 2345 4083
rect 4173 4049 4281 4083
rect 2237 4037 4281 4049
rect 4437 4709 6481 4721
rect 4437 4675 4545 4709
rect 6373 4675 6481 4709
rect 4437 4663 6481 4675
rect 4437 4613 4495 4663
rect 4437 4145 4449 4613
rect 4483 4145 4495 4613
rect 6423 4613 6481 4663
rect 4437 4095 4495 4145
rect 6423 4145 6435 4613
rect 6469 4145 6481 4613
rect 6423 4095 6481 4145
rect 4437 4083 6481 4095
rect 4437 4049 4545 4083
rect 6373 4049 6481 4083
rect 4437 4037 6481 4049
rect 6637 4709 8681 4721
rect 6637 4675 6745 4709
rect 8573 4675 8681 4709
rect 6637 4663 8681 4675
rect 6637 4613 6695 4663
rect 6637 4145 6649 4613
rect 6683 4145 6695 4613
rect 8623 4613 8681 4663
rect 6637 4095 6695 4145
rect 8623 4145 8635 4613
rect 8669 4145 8681 4613
rect 8623 4095 8681 4145
rect 6637 4083 8681 4095
rect 6637 4049 6745 4083
rect 8573 4049 8681 4083
rect 6637 4037 8681 4049
rect 8838 4710 10882 4722
rect 8838 4676 8946 4710
rect 10774 4676 10882 4710
rect 8838 4664 10882 4676
rect 8838 4614 8896 4664
rect 8838 4146 8850 4614
rect 8884 4146 8896 4614
rect 10824 4614 10882 4664
rect 8838 4096 8896 4146
rect 10824 4146 10836 4614
rect 10870 4146 10882 4614
rect 10824 4096 10882 4146
rect 8838 4084 10882 4096
rect 8838 4050 8946 4084
rect 10774 4050 10882 4084
rect 8838 4038 10882 4050
rect 11038 4710 13082 4722
rect 11038 4676 11146 4710
rect 12974 4676 13082 4710
rect 11038 4664 13082 4676
rect 11038 4614 11096 4664
rect 11038 4146 11050 4614
rect 11084 4146 11096 4614
rect 13024 4614 13082 4664
rect 11038 4096 11096 4146
rect 13024 4146 13036 4614
rect 13070 4146 13082 4614
rect 13024 4096 13082 4146
rect 11038 4084 13082 4096
rect 11038 4050 11146 4084
rect 12974 4050 13082 4084
rect 11038 4038 13082 4050
rect 13237 4709 15281 4721
rect 13237 4675 13345 4709
rect 15173 4675 15281 4709
rect 13237 4663 15281 4675
rect 13237 4613 13295 4663
rect 13237 4145 13249 4613
rect 13283 4145 13295 4613
rect 15223 4613 15281 4663
rect 13237 4095 13295 4145
rect 15223 4145 15235 4613
rect 15269 4145 15281 4613
rect 15223 4095 15281 4145
rect 13237 4083 15281 4095
rect 13237 4049 13345 4083
rect 15173 4049 15281 4083
rect 13237 4037 15281 4049
rect 15437 4709 17481 4721
rect 15437 4675 15545 4709
rect 17373 4675 17481 4709
rect 15437 4663 17481 4675
rect 15437 4613 15495 4663
rect 15437 4145 15449 4613
rect 15483 4145 15495 4613
rect 17423 4613 17481 4663
rect 15437 4095 15495 4145
rect 17423 4145 17435 4613
rect 17469 4145 17481 4613
rect 17423 4095 17481 4145
rect 15437 4083 17481 4095
rect 15437 4049 15545 4083
rect 17373 4049 17481 4083
rect 15437 4037 17481 4049
rect 17637 4709 19681 4721
rect 17637 4675 17745 4709
rect 19573 4675 19681 4709
rect 17637 4663 19681 4675
rect 17637 4613 17695 4663
rect 17637 4145 17649 4613
rect 17683 4145 17695 4613
rect 19623 4613 19681 4663
rect 17637 4095 17695 4145
rect 19623 4145 19635 4613
rect 19669 4145 19681 4613
rect 19623 4095 19681 4145
rect 17637 4083 19681 4095
rect 17637 4049 17745 4083
rect 19573 4049 19681 4083
rect 17637 4037 19681 4049
rect 19837 4709 21881 4721
rect 19837 4675 19945 4709
rect 21773 4675 21881 4709
rect 19837 4663 21881 4675
rect 19837 4613 19895 4663
rect 19837 4145 19849 4613
rect 19883 4145 19895 4613
rect 21823 4613 21881 4663
rect 19837 4095 19895 4145
rect 21823 4145 21835 4613
rect 21869 4145 21881 4613
rect 29956 11937 32075 11949
rect 29956 11903 30064 11937
rect 30648 11903 30819 11937
rect 31087 11903 31259 11937
rect 31527 11903 31699 11937
rect 31967 11903 32075 11937
rect 29956 11891 32075 11903
rect 29956 11841 30014 11891
rect 29956 11413 29968 11841
rect 30002 11413 30014 11841
rect 30698 11841 30769 11891
rect 29956 11363 30014 11413
rect 30698 11413 30710 11841
rect 30744 11413 30769 11841
rect 30698 11363 30769 11413
rect 31137 11363 31209 11891
rect 31577 11841 31649 11891
rect 31577 11413 31603 11841
rect 31637 11413 31649 11841
rect 32017 11841 32075 11891
rect 31577 11363 31649 11413
rect 32017 11413 32029 11841
rect 32063 11413 32075 11841
rect 32017 11363 32075 11413
rect 29956 11351 32075 11363
rect 29956 11317 30064 11351
rect 30648 11317 30819 11351
rect 31087 11317 31259 11351
rect 31527 11317 31699 11351
rect 31967 11317 32075 11351
rect 29956 11305 32075 11317
rect 32156 11937 34275 11949
rect 32156 11903 32264 11937
rect 32848 11903 33019 11937
rect 33287 11903 33459 11937
rect 33727 11903 33899 11937
rect 34167 11903 34275 11937
rect 32156 11891 34275 11903
rect 32156 11841 32214 11891
rect 32156 11413 32168 11841
rect 32202 11413 32214 11841
rect 32898 11841 32969 11891
rect 32156 11363 32214 11413
rect 32898 11413 32910 11841
rect 32944 11413 32969 11841
rect 32898 11363 32969 11413
rect 33337 11363 33409 11891
rect 33777 11841 33849 11891
rect 33777 11413 33803 11841
rect 33837 11413 33849 11841
rect 34217 11841 34275 11891
rect 33777 11363 33849 11413
rect 34217 11413 34229 11841
rect 34263 11413 34275 11841
rect 34217 11363 34275 11413
rect 32156 11351 34275 11363
rect 32156 11317 32264 11351
rect 32848 11317 33019 11351
rect 33287 11317 33459 11351
rect 33727 11317 33899 11351
rect 34167 11317 34275 11351
rect 32156 11305 34275 11317
rect 34356 11937 36475 11949
rect 34356 11903 34464 11937
rect 35048 11903 35219 11937
rect 35487 11903 35659 11937
rect 35927 11903 36099 11937
rect 36367 11903 36475 11937
rect 34356 11891 36475 11903
rect 34356 11841 34414 11891
rect 34356 11413 34368 11841
rect 34402 11413 34414 11841
rect 35098 11841 35169 11891
rect 34356 11363 34414 11413
rect 35098 11413 35110 11841
rect 35144 11413 35169 11841
rect 35098 11363 35169 11413
rect 35537 11363 35609 11891
rect 35977 11841 36049 11891
rect 35977 11413 36003 11841
rect 36037 11413 36049 11841
rect 36417 11841 36475 11891
rect 35977 11363 36049 11413
rect 36417 11413 36429 11841
rect 36463 11413 36475 11841
rect 36417 11363 36475 11413
rect 34356 11351 36475 11363
rect 34356 11317 34464 11351
rect 35048 11317 35219 11351
rect 35487 11317 35659 11351
rect 35927 11317 36099 11351
rect 36367 11317 36475 11351
rect 34356 11305 36475 11317
rect 33326 7648 34284 7660
rect 33326 7614 33434 7648
rect 34176 7614 34284 7648
rect 33326 7602 34284 7614
rect 33326 7552 33384 7602
rect 33326 6924 33338 7552
rect 33372 6924 33384 7552
rect 34226 7552 34284 7602
rect 33326 6874 33384 6924
rect 34226 6924 34238 7552
rect 34272 6924 34284 7552
rect 34226 6874 34284 6924
rect 33326 6862 34284 6874
rect 33326 6828 33434 6862
rect 34176 6828 34284 6862
rect 33326 6816 34284 6828
rect 29536 6368 30780 6380
rect 29536 6334 29644 6368
rect 30672 6334 30780 6368
rect 29536 6322 30780 6334
rect 29536 6272 29594 6322
rect 29536 5904 29548 6272
rect 29582 5904 29594 6272
rect 30722 6272 30780 6322
rect 29536 5854 29594 5904
rect 30722 5904 30734 6272
rect 30768 5904 30780 6272
rect 30722 5854 30780 5904
rect 29536 5842 30780 5854
rect 29536 5808 29644 5842
rect 30672 5808 30780 5842
rect 29536 5796 30780 5808
rect 30876 6368 32120 6380
rect 30876 6334 30984 6368
rect 32012 6334 32120 6368
rect 30876 6322 32120 6334
rect 30876 6272 30934 6322
rect 30876 5904 30888 6272
rect 30922 5904 30934 6272
rect 32062 6272 32120 6322
rect 30876 5854 30934 5904
rect 32062 5904 32074 6272
rect 32108 5904 32120 6272
rect 32062 5854 32120 5904
rect 30876 5842 32120 5854
rect 30876 5808 30984 5842
rect 32012 5808 32120 5842
rect 30876 5796 32120 5808
rect 36226 6134 37856 6146
rect 36226 6100 36334 6134
rect 36962 6100 37120 6134
rect 37748 6100 37856 6134
rect 36226 6088 37856 6100
rect 36226 6038 36284 6088
rect 29776 5718 30560 5730
rect 29776 5684 29884 5718
rect 30452 5684 30560 5718
rect 29776 5672 30560 5684
rect 29776 5622 29834 5672
rect 21823 4095 21881 4145
rect 29776 5294 29788 5622
rect 29822 5294 29834 5622
rect 30502 5622 30560 5672
rect 29776 5244 29834 5294
rect 30502 5294 30514 5622
rect 30548 5294 30560 5622
rect 30502 5244 30560 5294
rect 29776 5232 30560 5244
rect 29776 5198 29884 5232
rect 30452 5198 30560 5232
rect 29776 5186 30560 5198
rect 31086 5718 31870 5730
rect 31086 5684 31194 5718
rect 31762 5684 31870 5718
rect 31086 5672 31870 5684
rect 31086 5622 31144 5672
rect 31086 5294 31098 5622
rect 31132 5294 31144 5622
rect 31812 5622 31870 5672
rect 31086 5244 31144 5294
rect 31812 5294 31824 5622
rect 31858 5294 31870 5622
rect 31812 5244 31870 5294
rect 31086 5232 31870 5244
rect 31086 5198 31194 5232
rect 31762 5198 31870 5232
rect 31086 5186 31870 5198
rect 29536 5108 30780 5120
rect 29536 5074 29644 5108
rect 30672 5074 30780 5108
rect 29536 5062 30780 5074
rect 29536 5012 29594 5062
rect 29536 4644 29548 5012
rect 29582 4644 29594 5012
rect 30722 5012 30780 5062
rect 29536 4594 29594 4644
rect 30722 4644 30734 5012
rect 30768 4644 30780 5012
rect 30722 4594 30780 4644
rect 29536 4582 30780 4594
rect 29536 4548 29644 4582
rect 30672 4548 30780 4582
rect 29536 4536 30780 4548
rect 30876 5108 32120 5120
rect 30876 5074 30984 5108
rect 32012 5074 32120 5108
rect 30876 5062 32120 5074
rect 30876 5012 30934 5062
rect 30876 4644 30888 5012
rect 30922 4644 30934 5012
rect 32062 5012 32120 5062
rect 30876 4594 30934 4644
rect 32062 4644 32074 5012
rect 32108 4644 32120 5012
rect 32062 4594 32120 4644
rect 30876 4582 32120 4594
rect 30876 4548 30984 4582
rect 32012 4548 32120 4582
rect 30876 4536 32120 4548
rect 32576 4168 34166 4180
rect 32576 4134 32684 4168
rect 34058 4134 34166 4168
rect 19837 4083 21881 4095
rect 19837 4049 19945 4083
rect 21773 4049 21881 4083
rect 19837 4037 21881 4049
rect 32576 4122 34166 4134
rect 32576 4072 32634 4122
rect 16956 3526 17914 3538
rect 16956 3492 17064 3526
rect 17806 3492 17914 3526
rect 16956 3480 17914 3492
rect 16956 3430 17014 3480
rect 16956 2464 16968 3430
rect 17002 2464 17014 3430
rect 17856 3430 17914 3480
rect 16956 2414 17014 2464
rect 17856 2464 17868 3430
rect 17902 2464 17914 3430
rect 32576 3444 32588 4072
rect 32622 3444 32634 4072
rect 34108 4072 34166 4122
rect 32576 3394 32634 3444
rect 34108 3444 34120 4072
rect 34154 3444 34166 4072
rect 34108 3394 34166 3444
rect 32576 3382 34166 3394
rect 32576 3348 32684 3382
rect 34058 3348 34166 3382
rect 32576 3336 34166 3348
rect 34766 4168 35566 4180
rect 34766 4134 34874 4168
rect 35458 4134 35566 4168
rect 34766 4122 35566 4134
rect 34766 4072 34824 4122
rect 34766 3444 34778 4072
rect 34812 3444 34824 4072
rect 35508 4072 35566 4122
rect 34766 3394 34824 3444
rect 35508 3444 35520 4072
rect 35554 3444 35566 4072
rect 36226 3864 36238 6038
rect 36272 3864 36284 6038
rect 37012 6038 37070 6088
rect 36226 3814 36284 3864
rect 37012 3864 37024 6038
rect 37058 3864 37070 6038
rect 37798 6038 37856 6088
rect 37012 3814 37070 3864
rect 37798 3864 37810 6038
rect 37844 3864 37856 6038
rect 37798 3814 37856 3864
rect 36226 3802 37856 3814
rect 36226 3768 36334 3802
rect 36962 3768 37120 3802
rect 37748 3768 37856 3802
rect 36226 3756 37856 3768
rect 35508 3394 35566 3444
rect 34766 3382 35566 3394
rect 34766 3348 34874 3382
rect 35458 3348 35566 3382
rect 34766 3336 35566 3348
rect 17856 2414 17914 2464
rect 16956 2402 17914 2414
rect 32246 3238 32888 3250
rect 32246 3204 32354 3238
rect 32780 3204 32888 3238
rect 32246 3192 32888 3204
rect 32246 3142 32304 3192
rect 32246 2514 32258 3142
rect 32292 2514 32304 3142
rect 32830 3142 32888 3192
rect 32246 2464 32304 2514
rect 32830 2514 32842 3142
rect 32876 2514 32888 3142
rect 32830 2464 32888 2514
rect 32246 2452 32888 2464
rect 32246 2418 32354 2452
rect 32780 2418 32888 2452
rect 32246 2406 32888 2418
rect 33846 3238 34488 3250
rect 33846 3204 33954 3238
rect 34380 3204 34488 3238
rect 33846 3192 34488 3204
rect 33846 3142 33904 3192
rect 33846 2514 33858 3142
rect 33892 2514 33904 3142
rect 34430 3142 34488 3192
rect 33846 2464 33904 2514
rect 34430 2514 34442 3142
rect 34476 2514 34488 3142
rect 34430 2464 34488 2514
rect 33846 2452 34488 2464
rect 33846 2418 33954 2452
rect 34380 2418 34488 2452
rect 33846 2406 34488 2418
rect 35446 3238 36088 3250
rect 35446 3204 35554 3238
rect 35980 3204 36088 3238
rect 35446 3192 36088 3204
rect 35446 3142 35504 3192
rect 35446 2514 35458 3142
rect 35492 2514 35504 3142
rect 36030 3142 36088 3192
rect 35446 2464 35504 2514
rect 36030 2514 36042 3142
rect 36076 2514 36088 3142
rect 36030 2464 36088 2514
rect 35446 2452 36088 2464
rect 35446 2418 35554 2452
rect 35980 2418 36088 2452
rect 35446 2406 36088 2418
rect 16956 2368 17064 2402
rect 17806 2368 17914 2402
rect 16956 2356 17914 2368
rect -163 2229 1299 2241
rect -163 2195 -55 2229
rect 1191 2195 1299 2229
rect -163 2183 1299 2195
rect -163 2133 -105 2183
rect -163 1165 -151 2133
rect -117 1165 -105 2133
rect 1241 2133 1299 2183
rect -163 1115 -105 1165
rect 1241 1165 1253 2133
rect 1287 1165 1299 2133
rect 1241 1115 1299 1165
rect -163 1103 1299 1115
rect -163 1069 -55 1103
rect 1191 1069 1299 1103
rect -163 1037 1299 1069
rect -163 987 -105 1037
rect -163 619 -151 987
rect -117 619 -105 987
rect 1241 987 1299 1037
rect -163 569 -105 619
rect 1241 619 1253 987
rect 1287 619 1299 987
rect 1241 569 1299 619
rect -163 511 1299 569
rect 1437 2229 2899 2241
rect 1437 2195 1545 2229
rect 2791 2195 2899 2229
rect 1437 2183 2899 2195
rect 1437 2133 1495 2183
rect 1437 1165 1449 2133
rect 1483 1165 1495 2133
rect 2841 2133 2899 2183
rect 1437 1115 1495 1165
rect 2841 1165 2853 2133
rect 2887 1165 2899 2133
rect 2841 1115 2899 1165
rect 1437 1103 2899 1115
rect 1437 1069 1545 1103
rect 2791 1069 2899 1103
rect 1437 1037 2899 1069
rect 1437 987 1495 1037
rect 1437 619 1449 987
rect 1483 619 1495 987
rect 2841 987 2899 1037
rect 1437 569 1495 619
rect 2841 619 2853 987
rect 2887 619 2899 987
rect 2841 569 2899 619
rect 1437 511 2899 569
rect 3037 2229 4499 2241
rect 3037 2195 3145 2229
rect 4391 2195 4499 2229
rect 3037 2183 4499 2195
rect 3037 2133 3095 2183
rect 3037 1165 3049 2133
rect 3083 1165 3095 2133
rect 4441 2133 4499 2183
rect 3037 1115 3095 1165
rect 4441 1165 4453 2133
rect 4487 1165 4499 2133
rect 4441 1115 4499 1165
rect 3037 1103 4499 1115
rect 3037 1069 3145 1103
rect 4391 1069 4499 1103
rect 3037 1037 4499 1069
rect 3037 987 3095 1037
rect 3037 619 3049 987
rect 3083 619 3095 987
rect 4441 987 4499 1037
rect 3037 569 3095 619
rect 4441 619 4453 987
rect 4487 619 4499 987
rect 4441 569 4499 619
rect 3037 511 4499 569
rect 4637 2229 6099 2241
rect 4637 2195 4745 2229
rect 5991 2195 6099 2229
rect 4637 2183 6099 2195
rect 4637 2133 4695 2183
rect 4637 1165 4649 2133
rect 4683 1165 4695 2133
rect 6041 2133 6099 2183
rect 4637 1115 4695 1165
rect 6041 1165 6053 2133
rect 6087 1165 6099 2133
rect 6041 1115 6099 1165
rect 4637 1103 6099 1115
rect 4637 1069 4745 1103
rect 5991 1069 6099 1103
rect 4637 1037 6099 1069
rect 4637 987 4695 1037
rect 4637 619 4649 987
rect 4683 619 4695 987
rect 6041 987 6099 1037
rect 4637 569 4695 619
rect 6041 619 6053 987
rect 6087 619 6099 987
rect 6041 569 6099 619
rect 4637 511 6099 569
rect 6237 2229 7699 2241
rect 6237 2195 6345 2229
rect 7591 2195 7699 2229
rect 6237 2183 7699 2195
rect 6237 2133 6295 2183
rect 6237 1165 6249 2133
rect 6283 1165 6295 2133
rect 7641 2133 7699 2183
rect 6237 1115 6295 1165
rect 7641 1165 7653 2133
rect 7687 1165 7699 2133
rect 7641 1115 7699 1165
rect 6237 1103 7699 1115
rect 6237 1069 6345 1103
rect 7591 1069 7699 1103
rect 6237 1037 7699 1069
rect 6237 987 6295 1037
rect 6237 619 6249 987
rect 6283 619 6295 987
rect 7641 987 7699 1037
rect 6237 569 6295 619
rect 7641 619 7653 987
rect 7687 619 7699 987
rect 7641 569 7699 619
rect 6237 511 7699 569
rect 7837 2229 9299 2241
rect 7837 2195 7945 2229
rect 9191 2195 9299 2229
rect 7837 2183 9299 2195
rect 7837 2133 7895 2183
rect 7837 1165 7849 2133
rect 7883 1165 7895 2133
rect 9241 2133 9299 2183
rect 7837 1115 7895 1165
rect 9241 1165 9253 2133
rect 9287 1165 9299 2133
rect 9241 1115 9299 1165
rect 7837 1103 9299 1115
rect 7837 1069 7945 1103
rect 9191 1069 9299 1103
rect 7837 1037 9299 1069
rect 7837 987 7895 1037
rect 7837 619 7849 987
rect 7883 619 7895 987
rect 9241 987 9299 1037
rect 7837 569 7895 619
rect 9241 619 9253 987
rect 9287 619 9299 987
rect 9241 569 9299 619
rect 7837 511 9299 569
rect 9437 2229 10899 2241
rect 9437 2195 9545 2229
rect 10791 2195 10899 2229
rect 9437 2183 10899 2195
rect 9437 2133 9495 2183
rect 9437 1165 9449 2133
rect 9483 1165 9495 2133
rect 10841 2133 10899 2183
rect 9437 1115 9495 1165
rect 10841 1165 10853 2133
rect 10887 1165 10899 2133
rect 10841 1115 10899 1165
rect 9437 1103 10899 1115
rect 9437 1069 9545 1103
rect 10791 1069 10899 1103
rect 9437 1037 10899 1069
rect 9437 987 9495 1037
rect 9437 619 9449 987
rect 9483 619 9495 987
rect 10841 987 10899 1037
rect 9437 569 9495 619
rect 10841 619 10853 987
rect 10887 619 10899 987
rect 10841 569 10899 619
rect 9437 511 10899 569
rect 11037 2229 12499 2241
rect 11037 2195 11145 2229
rect 12391 2195 12499 2229
rect 11037 2183 12499 2195
rect 11037 2133 11095 2183
rect 11037 1165 11049 2133
rect 11083 1165 11095 2133
rect 12441 2133 12499 2183
rect 11037 1115 11095 1165
rect 12441 1165 12453 2133
rect 12487 1165 12499 2133
rect 12441 1115 12499 1165
rect 11037 1103 12499 1115
rect 11037 1069 11145 1103
rect 12391 1069 12499 1103
rect 11037 1037 12499 1069
rect 11037 987 11095 1037
rect 11037 619 11049 987
rect 11083 619 11095 987
rect 12441 987 12499 1037
rect 11037 569 11095 619
rect 12441 619 12453 987
rect 12487 619 12499 987
rect 12441 569 12499 619
rect 11037 511 12499 569
rect 12637 2229 14099 2241
rect 12637 2195 12745 2229
rect 13991 2195 14099 2229
rect 12637 2183 14099 2195
rect 12637 2133 12695 2183
rect 12637 1165 12649 2133
rect 12683 1165 12695 2133
rect 14041 2133 14099 2183
rect 12637 1115 12695 1165
rect 14041 1165 14053 2133
rect 14087 1165 14099 2133
rect 14041 1115 14099 1165
rect 12637 1103 14099 1115
rect 12637 1069 12745 1103
rect 13991 1069 14099 1103
rect 12637 1037 14099 1069
rect 12637 987 12695 1037
rect 12637 619 12649 987
rect 12683 619 12695 987
rect 14041 987 14099 1037
rect 12637 569 12695 619
rect 14041 619 14053 987
rect 14087 619 14099 987
rect 14041 569 14099 619
rect 12637 511 14099 569
rect 14237 2229 15699 2241
rect 14237 2195 14345 2229
rect 15591 2195 15699 2229
rect 14237 2183 15699 2195
rect 14237 2133 14295 2183
rect 14237 1165 14249 2133
rect 14283 1165 14295 2133
rect 15641 2133 15699 2183
rect 14237 1115 14295 1165
rect 15641 1165 15653 2133
rect 15687 1165 15699 2133
rect 15641 1115 15699 1165
rect 14237 1103 15699 1115
rect 14237 1069 14345 1103
rect 15591 1069 15699 1103
rect 14237 1037 15699 1069
rect 14237 987 14295 1037
rect 14237 619 14249 987
rect 14283 619 14295 987
rect 15641 987 15699 1037
rect 14237 569 14295 619
rect 15641 619 15653 987
rect 15687 619 15699 987
rect 15641 569 15699 619
rect 14237 511 15699 569
rect 15837 2229 17299 2241
rect 15837 2195 15945 2229
rect 17191 2195 17299 2229
rect 15837 2183 17299 2195
rect 15837 2133 15895 2183
rect 15837 1165 15849 2133
rect 15883 1165 15895 2133
rect 17241 2133 17299 2183
rect 15837 1115 15895 1165
rect 17241 1165 17253 2133
rect 17287 1165 17299 2133
rect 17241 1115 17299 1165
rect 15837 1103 17299 1115
rect 15837 1069 15945 1103
rect 17191 1069 17299 1103
rect 15837 1037 17299 1069
rect 15837 987 15895 1037
rect 15837 619 15849 987
rect 15883 619 15895 987
rect 17241 987 17299 1037
rect 15837 569 15895 619
rect 17241 619 17253 987
rect 17287 619 17299 987
rect 17241 569 17299 619
rect 15837 511 17299 569
rect 17437 2229 18899 2241
rect 17437 2195 17545 2229
rect 18791 2195 18899 2229
rect 17437 2183 18899 2195
rect 17437 2133 17495 2183
rect 17437 1165 17449 2133
rect 17483 1165 17495 2133
rect 18841 2133 18899 2183
rect 17437 1115 17495 1165
rect 18841 1165 18853 2133
rect 18887 1165 18899 2133
rect 18841 1115 18899 1165
rect 17437 1103 18899 1115
rect 17437 1069 17545 1103
rect 18791 1069 18899 1103
rect 17437 1037 18899 1069
rect 17437 987 17495 1037
rect 17437 619 17449 987
rect 17483 619 17495 987
rect 18841 987 18899 1037
rect 17437 569 17495 619
rect 18841 619 18853 987
rect 18887 619 18899 987
rect 18841 569 18899 619
rect 17437 511 18899 569
rect 19037 2229 20499 2241
rect 19037 2195 19145 2229
rect 20391 2195 20499 2229
rect 19037 2183 20499 2195
rect 19037 2133 19095 2183
rect 19037 1165 19049 2133
rect 19083 1165 19095 2133
rect 20441 2133 20499 2183
rect 19037 1115 19095 1165
rect 20441 1165 20453 2133
rect 20487 1165 20499 2133
rect 20441 1115 20499 1165
rect 19037 1103 20499 1115
rect 19037 1069 19145 1103
rect 20391 1069 20499 1103
rect 19037 1037 20499 1069
rect 19037 987 19095 1037
rect 19037 619 19049 987
rect 19083 619 19095 987
rect 20441 987 20499 1037
rect 19037 569 19095 619
rect 20441 619 20453 987
rect 20487 619 20499 987
rect 20441 569 20499 619
rect 19037 511 20499 569
rect 20637 2229 22099 2241
rect 20637 2195 20745 2229
rect 21991 2195 22099 2229
rect 20637 2183 22099 2195
rect 20637 2133 20695 2183
rect 20637 1165 20649 2133
rect 20683 1165 20695 2133
rect 22041 2133 22099 2183
rect 20637 1115 20695 1165
rect 22041 1165 22053 2133
rect 22087 1165 22099 2133
rect 22041 1115 22099 1165
rect 20637 1103 22099 1115
rect 20637 1069 20745 1103
rect 21991 1069 22099 1103
rect 20637 1037 22099 1069
rect 20637 987 20695 1037
rect 20637 619 20649 987
rect 20683 619 20695 987
rect 22041 987 22099 1037
rect 20637 569 20695 619
rect 22041 619 22053 987
rect 22087 619 22099 987
rect 22041 569 22099 619
rect 20637 511 22099 569
rect 22237 2229 23699 2241
rect 22237 2195 22345 2229
rect 23591 2195 23699 2229
rect 22237 2183 23699 2195
rect 22237 2133 22295 2183
rect 22237 1165 22249 2133
rect 22283 1165 22295 2133
rect 23641 2133 23699 2183
rect 22237 1115 22295 1165
rect 23641 1165 23653 2133
rect 23687 1165 23699 2133
rect 23641 1115 23699 1165
rect 22237 1103 23699 1115
rect 22237 1069 22345 1103
rect 23591 1069 23699 1103
rect 22237 1037 23699 1069
rect 22237 987 22295 1037
rect 22237 619 22249 987
rect 22283 619 22295 987
rect 23641 987 23699 1037
rect 22237 569 22295 619
rect 23641 619 23653 987
rect 23687 619 23699 987
rect 23641 569 23699 619
rect 22237 511 23699 569
rect 23837 2229 25299 2241
rect 23837 2195 23945 2229
rect 25191 2195 25299 2229
rect 23837 2183 25299 2195
rect 23837 2133 23895 2183
rect 23837 1165 23849 2133
rect 23883 1165 23895 2133
rect 25241 2133 25299 2183
rect 23837 1115 23895 1165
rect 25241 1165 25253 2133
rect 25287 1165 25299 2133
rect 25241 1115 25299 1165
rect 23837 1103 25299 1115
rect 23837 1069 23945 1103
rect 25191 1069 25299 1103
rect 23837 1037 25299 1069
rect 23837 987 23895 1037
rect 23837 619 23849 987
rect 23883 619 23895 987
rect 25241 987 25299 1037
rect 23837 569 23895 619
rect 25241 619 25253 987
rect 25287 619 25299 987
rect 25241 569 25299 619
rect 23837 511 25299 569
rect 25437 2229 26899 2241
rect 25437 2195 25545 2229
rect 26791 2195 26899 2229
rect 25437 2183 26899 2195
rect 25437 2133 25495 2183
rect 25437 1165 25449 2133
rect 25483 1165 25495 2133
rect 26841 2133 26899 2183
rect 25437 1115 25495 1165
rect 26841 1165 26853 2133
rect 26887 1165 26899 2133
rect 26841 1115 26899 1165
rect 25437 1103 26899 1115
rect 25437 1069 25545 1103
rect 26791 1069 26899 1103
rect 25437 1037 26899 1069
rect 25437 987 25495 1037
rect 25437 619 25449 987
rect 25483 619 25495 987
rect 26841 987 26899 1037
rect 25437 569 25495 619
rect 26841 619 26853 987
rect 26887 619 26899 987
rect 26841 569 26899 619
rect 25437 511 26899 569
rect 27037 2229 28499 2241
rect 27037 2195 27145 2229
rect 28391 2195 28499 2229
rect 27037 2183 28499 2195
rect 27037 2133 27095 2183
rect 27037 1165 27049 2133
rect 27083 1165 27095 2133
rect 28441 2133 28499 2183
rect 27037 1115 27095 1165
rect 28441 1165 28453 2133
rect 28487 1165 28499 2133
rect 28441 1115 28499 1165
rect 27037 1103 28499 1115
rect 27037 1069 27145 1103
rect 28391 1069 28499 1103
rect 27037 1037 28499 1069
rect 27037 987 27095 1037
rect 27037 619 27049 987
rect 27083 619 27095 987
rect 28441 987 28499 1037
rect 27037 569 27095 619
rect 28441 619 28453 987
rect 28487 619 28499 987
rect 28441 569 28499 619
rect 27037 511 28499 569
rect 28637 2229 30099 2241
rect 28637 2195 28745 2229
rect 29991 2195 30099 2229
rect 28637 2183 30099 2195
rect 28637 2133 28695 2183
rect 28637 1165 28649 2133
rect 28683 1165 28695 2133
rect 30041 2133 30099 2183
rect 28637 1115 28695 1165
rect 30041 1165 30053 2133
rect 30087 1165 30099 2133
rect 30041 1115 30099 1165
rect 28637 1103 30099 1115
rect 28637 1069 28745 1103
rect 29991 1069 30099 1103
rect 28637 1037 30099 1069
rect 28637 987 28695 1037
rect 28637 619 28649 987
rect 28683 619 28695 987
rect 30041 987 30099 1037
rect 28637 569 28695 619
rect 30041 619 30053 987
rect 30087 619 30099 987
rect 30041 569 30099 619
rect 28637 511 30099 569
rect 30237 2229 31699 2241
rect 30237 2195 30345 2229
rect 31591 2195 31699 2229
rect 30237 2183 31699 2195
rect 30237 2133 30295 2183
rect 30237 1165 30249 2133
rect 30283 1165 30295 2133
rect 31641 2133 31699 2183
rect 30237 1115 30295 1165
rect 31641 1165 31653 2133
rect 31687 1165 31699 2133
rect 31641 1115 31699 1165
rect 30237 1103 31699 1115
rect 30237 1069 30345 1103
rect 31591 1069 31699 1103
rect 30237 1037 31699 1069
rect 30237 987 30295 1037
rect 30237 619 30249 987
rect 30283 619 30295 987
rect 31641 987 31699 1037
rect 30237 569 30295 619
rect 31641 619 31653 987
rect 31687 619 31699 987
rect 31641 569 31699 619
rect 30237 511 31699 569
rect 31837 2229 33299 2241
rect 31837 2195 31945 2229
rect 33191 2195 33299 2229
rect 31837 2183 33299 2195
rect 31837 2133 31895 2183
rect 31837 1165 31849 2133
rect 31883 1165 31895 2133
rect 33241 2133 33299 2183
rect 31837 1115 31895 1165
rect 33241 1165 33253 2133
rect 33287 1165 33299 2133
rect 33241 1115 33299 1165
rect 31837 1103 33299 1115
rect 31837 1069 31945 1103
rect 33191 1069 33299 1103
rect 31837 1037 33299 1069
rect 31837 987 31895 1037
rect 31837 619 31849 987
rect 31883 619 31895 987
rect 33241 987 33299 1037
rect 31837 569 31895 619
rect 33241 619 33253 987
rect 33287 619 33299 987
rect 33241 569 33299 619
rect 31837 511 33299 569
rect 33437 2229 34899 2241
rect 33437 2195 33545 2229
rect 34791 2195 34899 2229
rect 33437 2183 34899 2195
rect 33437 2133 33495 2183
rect 33437 1165 33449 2133
rect 33483 1165 33495 2133
rect 34841 2133 34899 2183
rect 33437 1115 33495 1165
rect 34841 1165 34853 2133
rect 34887 1165 34899 2133
rect 34841 1115 34899 1165
rect 33437 1103 34899 1115
rect 33437 1069 33545 1103
rect 34791 1069 34899 1103
rect 33437 1037 34899 1069
rect 33437 987 33495 1037
rect 33437 619 33449 987
rect 33483 619 33495 987
rect 34841 987 34899 1037
rect 33437 569 33495 619
rect 34841 619 34853 987
rect 34887 619 34899 987
rect 34841 569 34899 619
rect 33437 511 34899 569
rect 35037 2229 36499 2241
rect 35037 2195 35145 2229
rect 36391 2195 36499 2229
rect 35037 2183 36499 2195
rect 35037 2133 35095 2183
rect 35037 1165 35049 2133
rect 35083 1165 35095 2133
rect 36441 2133 36499 2183
rect 35037 1115 35095 1165
rect 36441 1165 36453 2133
rect 36487 1165 36499 2133
rect 36441 1115 36499 1165
rect 35037 1103 36499 1115
rect 35037 1069 35145 1103
rect 36391 1069 36499 1103
rect 35037 1037 36499 1069
rect 35037 987 35095 1037
rect 35037 619 35049 987
rect 35083 619 35095 987
rect 36441 987 36499 1037
rect 35037 569 35095 619
rect 36441 619 36453 987
rect 36487 619 36499 987
rect 36441 569 36499 619
rect 35037 511 36499 569
rect 36637 2229 38099 2241
rect 36637 2195 36745 2229
rect 37991 2195 38099 2229
rect 36637 2183 38099 2195
rect 36637 2133 36695 2183
rect 36637 1165 36649 2133
rect 36683 1165 36695 2133
rect 38041 2133 38099 2183
rect 36637 1115 36695 1165
rect 38041 1165 38053 2133
rect 38087 1165 38099 2133
rect 38041 1115 38099 1165
rect 36637 1103 38099 1115
rect 36637 1069 36745 1103
rect 37991 1069 38099 1103
rect 36637 1037 38099 1069
rect 36637 987 36695 1037
rect 36637 619 36649 987
rect 36683 619 36695 987
rect 38041 987 38099 1037
rect 36637 569 36695 619
rect 38041 619 38053 987
rect 38087 619 38099 987
rect 38041 569 38099 619
rect 36637 511 38099 569
rect -163 429 1299 441
rect -163 395 -55 429
rect 1191 395 1299 429
rect -163 383 1299 395
rect -163 333 -105 383
rect -163 -635 -151 333
rect -117 -635 -105 333
rect 1241 333 1299 383
rect -163 -685 -105 -635
rect 1241 -635 1253 333
rect 1287 -635 1299 333
rect 1241 -685 1299 -635
rect -163 -697 1299 -685
rect -163 -731 -55 -697
rect 1191 -731 1299 -697
rect -163 -763 1299 -731
rect -163 -813 -105 -763
rect -163 -1181 -151 -813
rect -117 -1181 -105 -813
rect 1241 -813 1299 -763
rect -163 -1231 -105 -1181
rect 1241 -1181 1253 -813
rect 1287 -1181 1299 -813
rect 1241 -1231 1299 -1181
rect -163 -1289 1299 -1231
rect 1437 429 2899 441
rect 1437 395 1545 429
rect 2791 395 2899 429
rect 1437 383 2899 395
rect 1437 333 1495 383
rect 1437 -635 1449 333
rect 1483 -635 1495 333
rect 2841 333 2899 383
rect 1437 -685 1495 -635
rect 2841 -635 2853 333
rect 2887 -635 2899 333
rect 2841 -685 2899 -635
rect 1437 -697 2899 -685
rect 1437 -731 1545 -697
rect 2791 -731 2899 -697
rect 1437 -763 2899 -731
rect 1437 -813 1495 -763
rect 1437 -1181 1449 -813
rect 1483 -1181 1495 -813
rect 2841 -813 2899 -763
rect 1437 -1231 1495 -1181
rect 2841 -1181 2853 -813
rect 2887 -1181 2899 -813
rect 2841 -1231 2899 -1181
rect 1437 -1289 2899 -1231
rect 3037 429 4499 441
rect 3037 395 3145 429
rect 4391 395 4499 429
rect 3037 383 4499 395
rect 3037 333 3095 383
rect 3037 -635 3049 333
rect 3083 -635 3095 333
rect 4441 333 4499 383
rect 3037 -685 3095 -635
rect 4441 -635 4453 333
rect 4487 -635 4499 333
rect 4441 -685 4499 -635
rect 3037 -697 4499 -685
rect 3037 -731 3145 -697
rect 4391 -731 4499 -697
rect 3037 -763 4499 -731
rect 3037 -813 3095 -763
rect 3037 -1181 3049 -813
rect 3083 -1181 3095 -813
rect 4441 -813 4499 -763
rect 3037 -1231 3095 -1181
rect 4441 -1181 4453 -813
rect 4487 -1181 4499 -813
rect 4441 -1231 4499 -1181
rect 3037 -1289 4499 -1231
rect 4637 429 6099 441
rect 4637 395 4745 429
rect 5991 395 6099 429
rect 4637 383 6099 395
rect 4637 333 4695 383
rect 4637 -635 4649 333
rect 4683 -635 4695 333
rect 6041 333 6099 383
rect 4637 -685 4695 -635
rect 6041 -635 6053 333
rect 6087 -635 6099 333
rect 6041 -685 6099 -635
rect 4637 -697 6099 -685
rect 4637 -731 4745 -697
rect 5991 -731 6099 -697
rect 4637 -763 6099 -731
rect 4637 -813 4695 -763
rect 4637 -1181 4649 -813
rect 4683 -1181 4695 -813
rect 6041 -813 6099 -763
rect 4637 -1231 4695 -1181
rect 6041 -1181 6053 -813
rect 6087 -1181 6099 -813
rect 6041 -1231 6099 -1181
rect 4637 -1289 6099 -1231
rect 6237 429 7699 441
rect 6237 395 6345 429
rect 7591 395 7699 429
rect 6237 383 7699 395
rect 6237 333 6295 383
rect 6237 -635 6249 333
rect 6283 -635 6295 333
rect 7641 333 7699 383
rect 6237 -685 6295 -635
rect 7641 -635 7653 333
rect 7687 -635 7699 333
rect 7641 -685 7699 -635
rect 6237 -697 7699 -685
rect 6237 -731 6345 -697
rect 7591 -731 7699 -697
rect 6237 -763 7699 -731
rect 6237 -813 6295 -763
rect 6237 -1181 6249 -813
rect 6283 -1181 6295 -813
rect 7641 -813 7699 -763
rect 6237 -1231 6295 -1181
rect 7641 -1181 7653 -813
rect 7687 -1181 7699 -813
rect 7641 -1231 7699 -1181
rect 6237 -1289 7699 -1231
rect 7837 429 9299 441
rect 7837 395 7945 429
rect 9191 395 9299 429
rect 7837 383 9299 395
rect 7837 333 7895 383
rect 7837 -635 7849 333
rect 7883 -635 7895 333
rect 9241 333 9299 383
rect 7837 -685 7895 -635
rect 9241 -635 9253 333
rect 9287 -635 9299 333
rect 9241 -685 9299 -635
rect 7837 -697 9299 -685
rect 7837 -731 7945 -697
rect 9191 -731 9299 -697
rect 7837 -763 9299 -731
rect 7837 -813 7895 -763
rect 7837 -1181 7849 -813
rect 7883 -1181 7895 -813
rect 9241 -813 9299 -763
rect 7837 -1231 7895 -1181
rect 9241 -1181 9253 -813
rect 9287 -1181 9299 -813
rect 9241 -1231 9299 -1181
rect 7837 -1289 9299 -1231
rect 9437 429 10899 441
rect 9437 395 9545 429
rect 10791 395 10899 429
rect 9437 383 10899 395
rect 9437 333 9495 383
rect 9437 -635 9449 333
rect 9483 -635 9495 333
rect 10841 333 10899 383
rect 9437 -685 9495 -635
rect 10841 -635 10853 333
rect 10887 -635 10899 333
rect 10841 -685 10899 -635
rect 9437 -697 10899 -685
rect 9437 -731 9545 -697
rect 10791 -731 10899 -697
rect 9437 -763 10899 -731
rect 9437 -813 9495 -763
rect 9437 -1181 9449 -813
rect 9483 -1181 9495 -813
rect 10841 -813 10899 -763
rect 9437 -1231 9495 -1181
rect 10841 -1181 10853 -813
rect 10887 -1181 10899 -813
rect 10841 -1231 10899 -1181
rect 9437 -1289 10899 -1231
rect 11037 429 12499 441
rect 11037 395 11145 429
rect 12391 395 12499 429
rect 11037 383 12499 395
rect 11037 333 11095 383
rect 11037 -635 11049 333
rect 11083 -635 11095 333
rect 12441 333 12499 383
rect 11037 -685 11095 -635
rect 12441 -635 12453 333
rect 12487 -635 12499 333
rect 12441 -685 12499 -635
rect 11037 -697 12499 -685
rect 11037 -731 11145 -697
rect 12391 -731 12499 -697
rect 11037 -763 12499 -731
rect 11037 -813 11095 -763
rect 11037 -1181 11049 -813
rect 11083 -1181 11095 -813
rect 12441 -813 12499 -763
rect 11037 -1231 11095 -1181
rect 12441 -1181 12453 -813
rect 12487 -1181 12499 -813
rect 12441 -1231 12499 -1181
rect 11037 -1289 12499 -1231
rect 12637 429 14099 441
rect 12637 395 12745 429
rect 13991 395 14099 429
rect 12637 383 14099 395
rect 12637 333 12695 383
rect 12637 -635 12649 333
rect 12683 -635 12695 333
rect 14041 333 14099 383
rect 12637 -685 12695 -635
rect 14041 -635 14053 333
rect 14087 -635 14099 333
rect 14041 -685 14099 -635
rect 12637 -697 14099 -685
rect 12637 -731 12745 -697
rect 13991 -731 14099 -697
rect 12637 -763 14099 -731
rect 12637 -813 12695 -763
rect 12637 -1181 12649 -813
rect 12683 -1181 12695 -813
rect 14041 -813 14099 -763
rect 12637 -1231 12695 -1181
rect 14041 -1181 14053 -813
rect 14087 -1181 14099 -813
rect 14041 -1231 14099 -1181
rect 12637 -1289 14099 -1231
rect 14237 429 15699 441
rect 14237 395 14345 429
rect 15591 395 15699 429
rect 14237 383 15699 395
rect 14237 333 14295 383
rect 14237 -635 14249 333
rect 14283 -635 14295 333
rect 15641 333 15699 383
rect 14237 -685 14295 -635
rect 15641 -635 15653 333
rect 15687 -635 15699 333
rect 15641 -685 15699 -635
rect 14237 -697 15699 -685
rect 14237 -731 14345 -697
rect 15591 -731 15699 -697
rect 14237 -763 15699 -731
rect 14237 -813 14295 -763
rect 14237 -1181 14249 -813
rect 14283 -1181 14295 -813
rect 15641 -813 15699 -763
rect 14237 -1231 14295 -1181
rect 15641 -1181 15653 -813
rect 15687 -1181 15699 -813
rect 15641 -1231 15699 -1181
rect 14237 -1289 15699 -1231
rect 15837 429 17299 441
rect 15837 395 15945 429
rect 17191 395 17299 429
rect 15837 383 17299 395
rect 15837 333 15895 383
rect 15837 -635 15849 333
rect 15883 -635 15895 333
rect 17241 333 17299 383
rect 15837 -685 15895 -635
rect 17241 -635 17253 333
rect 17287 -635 17299 333
rect 17241 -685 17299 -635
rect 15837 -697 17299 -685
rect 15837 -731 15945 -697
rect 17191 -731 17299 -697
rect 15837 -763 17299 -731
rect 15837 -813 15895 -763
rect 15837 -1181 15849 -813
rect 15883 -1181 15895 -813
rect 17241 -813 17299 -763
rect 15837 -1231 15895 -1181
rect 17241 -1181 17253 -813
rect 17287 -1181 17299 -813
rect 17241 -1231 17299 -1181
rect 15837 -1289 17299 -1231
rect 17437 429 18899 441
rect 17437 395 17545 429
rect 18791 395 18899 429
rect 17437 383 18899 395
rect 17437 333 17495 383
rect 17437 -635 17449 333
rect 17483 -635 17495 333
rect 18841 333 18899 383
rect 17437 -685 17495 -635
rect 18841 -635 18853 333
rect 18887 -635 18899 333
rect 18841 -685 18899 -635
rect 17437 -697 18899 -685
rect 17437 -731 17545 -697
rect 18791 -731 18899 -697
rect 17437 -763 18899 -731
rect 17437 -813 17495 -763
rect 17437 -1181 17449 -813
rect 17483 -1181 17495 -813
rect 18841 -813 18899 -763
rect 17437 -1231 17495 -1181
rect 18841 -1181 18853 -813
rect 18887 -1181 18899 -813
rect 18841 -1231 18899 -1181
rect 17437 -1289 18899 -1231
rect 19037 429 20499 441
rect 19037 395 19145 429
rect 20391 395 20499 429
rect 19037 383 20499 395
rect 19037 333 19095 383
rect 19037 -635 19049 333
rect 19083 -635 19095 333
rect 20441 333 20499 383
rect 19037 -685 19095 -635
rect 20441 -635 20453 333
rect 20487 -635 20499 333
rect 20441 -685 20499 -635
rect 19037 -697 20499 -685
rect 19037 -731 19145 -697
rect 20391 -731 20499 -697
rect 19037 -763 20499 -731
rect 19037 -813 19095 -763
rect 19037 -1181 19049 -813
rect 19083 -1181 19095 -813
rect 20441 -813 20499 -763
rect 19037 -1231 19095 -1181
rect 20441 -1181 20453 -813
rect 20487 -1181 20499 -813
rect 20441 -1231 20499 -1181
rect 19037 -1289 20499 -1231
rect 20637 429 22099 441
rect 20637 395 20745 429
rect 21991 395 22099 429
rect 20637 383 22099 395
rect 20637 333 20695 383
rect 20637 -635 20649 333
rect 20683 -635 20695 333
rect 22041 333 22099 383
rect 20637 -685 20695 -635
rect 22041 -635 22053 333
rect 22087 -635 22099 333
rect 22041 -685 22099 -635
rect 20637 -697 22099 -685
rect 20637 -731 20745 -697
rect 21991 -731 22099 -697
rect 20637 -763 22099 -731
rect 20637 -813 20695 -763
rect 20637 -1181 20649 -813
rect 20683 -1181 20695 -813
rect 22041 -813 22099 -763
rect 20637 -1231 20695 -1181
rect 22041 -1181 22053 -813
rect 22087 -1181 22099 -813
rect 22041 -1231 22099 -1181
rect 20637 -1289 22099 -1231
rect 22237 429 23699 441
rect 22237 395 22345 429
rect 23591 395 23699 429
rect 22237 383 23699 395
rect 22237 333 22295 383
rect 22237 -635 22249 333
rect 22283 -635 22295 333
rect 23641 333 23699 383
rect 22237 -685 22295 -635
rect 23641 -635 23653 333
rect 23687 -635 23699 333
rect 23641 -685 23699 -635
rect 22237 -697 23699 -685
rect 22237 -731 22345 -697
rect 23591 -731 23699 -697
rect 22237 -763 23699 -731
rect 22237 -813 22295 -763
rect 22237 -1181 22249 -813
rect 22283 -1181 22295 -813
rect 23641 -813 23699 -763
rect 22237 -1231 22295 -1181
rect 23641 -1181 23653 -813
rect 23687 -1181 23699 -813
rect 23641 -1231 23699 -1181
rect 22237 -1289 23699 -1231
rect 23837 429 25299 441
rect 23837 395 23945 429
rect 25191 395 25299 429
rect 23837 383 25299 395
rect 23837 333 23895 383
rect 23837 -635 23849 333
rect 23883 -635 23895 333
rect 25241 333 25299 383
rect 23837 -685 23895 -635
rect 25241 -635 25253 333
rect 25287 -635 25299 333
rect 25241 -685 25299 -635
rect 23837 -697 25299 -685
rect 23837 -731 23945 -697
rect 25191 -731 25299 -697
rect 23837 -763 25299 -731
rect 23837 -813 23895 -763
rect 23837 -1181 23849 -813
rect 23883 -1181 23895 -813
rect 25241 -813 25299 -763
rect 23837 -1231 23895 -1181
rect 25241 -1181 25253 -813
rect 25287 -1181 25299 -813
rect 25241 -1231 25299 -1181
rect 23837 -1289 25299 -1231
rect 25437 429 26899 441
rect 25437 395 25545 429
rect 26791 395 26899 429
rect 25437 383 26899 395
rect 25437 333 25495 383
rect 25437 -635 25449 333
rect 25483 -635 25495 333
rect 26841 333 26899 383
rect 25437 -685 25495 -635
rect 26841 -635 26853 333
rect 26887 -635 26899 333
rect 26841 -685 26899 -635
rect 25437 -697 26899 -685
rect 25437 -731 25545 -697
rect 26791 -731 26899 -697
rect 25437 -763 26899 -731
rect 25437 -813 25495 -763
rect 25437 -1181 25449 -813
rect 25483 -1181 25495 -813
rect 26841 -813 26899 -763
rect 25437 -1231 25495 -1181
rect 26841 -1181 26853 -813
rect 26887 -1181 26899 -813
rect 26841 -1231 26899 -1181
rect 25437 -1289 26899 -1231
rect 27037 429 28499 441
rect 27037 395 27145 429
rect 28391 395 28499 429
rect 27037 383 28499 395
rect 27037 333 27095 383
rect 27037 -635 27049 333
rect 27083 -635 27095 333
rect 28441 333 28499 383
rect 27037 -685 27095 -635
rect 28441 -635 28453 333
rect 28487 -635 28499 333
rect 28441 -685 28499 -635
rect 27037 -697 28499 -685
rect 27037 -731 27145 -697
rect 28391 -731 28499 -697
rect 27037 -763 28499 -731
rect 27037 -813 27095 -763
rect 27037 -1181 27049 -813
rect 27083 -1181 27095 -813
rect 28441 -813 28499 -763
rect 27037 -1231 27095 -1181
rect 28441 -1181 28453 -813
rect 28487 -1181 28499 -813
rect 28441 -1231 28499 -1181
rect 27037 -1289 28499 -1231
rect 28637 429 30099 441
rect 28637 395 28745 429
rect 29991 395 30099 429
rect 28637 383 30099 395
rect 28637 333 28695 383
rect 28637 -635 28649 333
rect 28683 -635 28695 333
rect 30041 333 30099 383
rect 28637 -685 28695 -635
rect 30041 -635 30053 333
rect 30087 -635 30099 333
rect 30041 -685 30099 -635
rect 28637 -697 30099 -685
rect 28637 -731 28745 -697
rect 29991 -731 30099 -697
rect 28637 -763 30099 -731
rect 28637 -813 28695 -763
rect 28637 -1181 28649 -813
rect 28683 -1181 28695 -813
rect 30041 -813 30099 -763
rect 28637 -1231 28695 -1181
rect 30041 -1181 30053 -813
rect 30087 -1181 30099 -813
rect 30041 -1231 30099 -1181
rect 28637 -1289 30099 -1231
rect 30237 429 31699 441
rect 30237 395 30345 429
rect 31591 395 31699 429
rect 30237 383 31699 395
rect 30237 333 30295 383
rect 30237 -635 30249 333
rect 30283 -635 30295 333
rect 31641 333 31699 383
rect 30237 -685 30295 -635
rect 31641 -635 31653 333
rect 31687 -635 31699 333
rect 31641 -685 31699 -635
rect 30237 -697 31699 -685
rect 30237 -731 30345 -697
rect 31591 -731 31699 -697
rect 30237 -763 31699 -731
rect 30237 -813 30295 -763
rect 30237 -1181 30249 -813
rect 30283 -1181 30295 -813
rect 31641 -813 31699 -763
rect 30237 -1231 30295 -1181
rect 31641 -1181 31653 -813
rect 31687 -1181 31699 -813
rect 31641 -1231 31699 -1181
rect 30237 -1289 31699 -1231
rect 31837 429 33299 441
rect 31837 395 31945 429
rect 33191 395 33299 429
rect 31837 383 33299 395
rect 31837 333 31895 383
rect 31837 -635 31849 333
rect 31883 -635 31895 333
rect 33241 333 33299 383
rect 31837 -685 31895 -635
rect 33241 -635 33253 333
rect 33287 -635 33299 333
rect 33241 -685 33299 -635
rect 31837 -697 33299 -685
rect 31837 -731 31945 -697
rect 33191 -731 33299 -697
rect 31837 -763 33299 -731
rect 31837 -813 31895 -763
rect 31837 -1181 31849 -813
rect 31883 -1181 31895 -813
rect 33241 -813 33299 -763
rect 31837 -1231 31895 -1181
rect 33241 -1181 33253 -813
rect 33287 -1181 33299 -813
rect 33241 -1231 33299 -1181
rect 31837 -1289 33299 -1231
rect 33437 429 34899 441
rect 33437 395 33545 429
rect 34791 395 34899 429
rect 33437 383 34899 395
rect 33437 333 33495 383
rect 33437 -635 33449 333
rect 33483 -635 33495 333
rect 34841 333 34899 383
rect 33437 -685 33495 -635
rect 34841 -635 34853 333
rect 34887 -635 34899 333
rect 34841 -685 34899 -635
rect 33437 -697 34899 -685
rect 33437 -731 33545 -697
rect 34791 -731 34899 -697
rect 33437 -763 34899 -731
rect 33437 -813 33495 -763
rect 33437 -1181 33449 -813
rect 33483 -1181 33495 -813
rect 34841 -813 34899 -763
rect 33437 -1231 33495 -1181
rect 34841 -1181 34853 -813
rect 34887 -1181 34899 -813
rect 34841 -1231 34899 -1181
rect 33437 -1289 34899 -1231
rect 35037 429 36499 441
rect 35037 395 35145 429
rect 36391 395 36499 429
rect 35037 383 36499 395
rect 35037 333 35095 383
rect 35037 -635 35049 333
rect 35083 -635 35095 333
rect 36441 333 36499 383
rect 35037 -685 35095 -635
rect 36441 -635 36453 333
rect 36487 -635 36499 333
rect 36441 -685 36499 -635
rect 35037 -697 36499 -685
rect 35037 -731 35145 -697
rect 36391 -731 36499 -697
rect 35037 -763 36499 -731
rect 35037 -813 35095 -763
rect 35037 -1181 35049 -813
rect 35083 -1181 35095 -813
rect 36441 -813 36499 -763
rect 35037 -1231 35095 -1181
rect 36441 -1181 36453 -813
rect 36487 -1181 36499 -813
rect 36441 -1231 36499 -1181
rect 35037 -1289 36499 -1231
rect 36637 429 38099 441
rect 36637 395 36745 429
rect 37991 395 38099 429
rect 36637 383 38099 395
rect 36637 333 36695 383
rect 36637 -635 36649 333
rect 36683 -635 36695 333
rect 38041 333 38099 383
rect 36637 -685 36695 -635
rect 38041 -635 38053 333
rect 38087 -635 38099 333
rect 38041 -685 38099 -635
rect 36637 -697 38099 -685
rect 36637 -731 36745 -697
rect 37991 -731 38099 -697
rect 36637 -763 38099 -731
rect 36637 -813 36695 -763
rect 36637 -1181 36649 -813
rect 36683 -1181 36695 -813
rect 38041 -813 38099 -763
rect 36637 -1231 36695 -1181
rect 38041 -1181 38053 -813
rect 38087 -1181 38099 -813
rect 38041 -1231 38099 -1181
rect 36637 -1289 38099 -1231
rect -163 -1371 1299 -1359
rect -163 -1405 -55 -1371
rect 1191 -1405 1299 -1371
rect -163 -1417 1299 -1405
rect -163 -1467 -105 -1417
rect -163 -2435 -151 -1467
rect -117 -2435 -105 -1467
rect 1241 -1467 1299 -1417
rect -163 -2485 -105 -2435
rect 1241 -2435 1253 -1467
rect 1287 -2435 1299 -1467
rect 1241 -2485 1299 -2435
rect -163 -2497 1299 -2485
rect -163 -2531 -55 -2497
rect 1191 -2531 1299 -2497
rect -163 -2563 1299 -2531
rect -163 -2613 -105 -2563
rect -163 -2981 -151 -2613
rect -117 -2981 -105 -2613
rect 1241 -2613 1299 -2563
rect -163 -3031 -105 -2981
rect 1241 -2981 1253 -2613
rect 1287 -2981 1299 -2613
rect 1241 -3031 1299 -2981
rect -163 -3089 1299 -3031
rect 1437 -1371 2899 -1359
rect 1437 -1405 1545 -1371
rect 2791 -1405 2899 -1371
rect 1437 -1417 2899 -1405
rect 1437 -1467 1495 -1417
rect 1437 -2435 1449 -1467
rect 1483 -2435 1495 -1467
rect 2841 -1467 2899 -1417
rect 1437 -2485 1495 -2435
rect 2841 -2435 2853 -1467
rect 2887 -2435 2899 -1467
rect 2841 -2485 2899 -2435
rect 1437 -2497 2899 -2485
rect 1437 -2531 1545 -2497
rect 2791 -2531 2899 -2497
rect 1437 -2563 2899 -2531
rect 1437 -2613 1495 -2563
rect 1437 -2981 1449 -2613
rect 1483 -2981 1495 -2613
rect 2841 -2613 2899 -2563
rect 1437 -3031 1495 -2981
rect 2841 -2981 2853 -2613
rect 2887 -2981 2899 -2613
rect 2841 -3031 2899 -2981
rect 1437 -3089 2899 -3031
rect 3037 -1371 4499 -1359
rect 3037 -1405 3145 -1371
rect 4391 -1405 4499 -1371
rect 3037 -1417 4499 -1405
rect 3037 -1467 3095 -1417
rect 3037 -2435 3049 -1467
rect 3083 -2435 3095 -1467
rect 4441 -1467 4499 -1417
rect 3037 -2485 3095 -2435
rect 4441 -2435 4453 -1467
rect 4487 -2435 4499 -1467
rect 4441 -2485 4499 -2435
rect 3037 -2497 4499 -2485
rect 3037 -2531 3145 -2497
rect 4391 -2531 4499 -2497
rect 3037 -2563 4499 -2531
rect 3037 -2613 3095 -2563
rect 3037 -2981 3049 -2613
rect 3083 -2981 3095 -2613
rect 4441 -2613 4499 -2563
rect 3037 -3031 3095 -2981
rect 4441 -2981 4453 -2613
rect 4487 -2981 4499 -2613
rect 4441 -3031 4499 -2981
rect 3037 -3089 4499 -3031
rect 4637 -1371 6099 -1359
rect 4637 -1405 4745 -1371
rect 5991 -1405 6099 -1371
rect 4637 -1417 6099 -1405
rect 4637 -1467 4695 -1417
rect 4637 -2435 4649 -1467
rect 4683 -2435 4695 -1467
rect 6041 -1467 6099 -1417
rect 4637 -2485 4695 -2435
rect 6041 -2435 6053 -1467
rect 6087 -2435 6099 -1467
rect 6041 -2485 6099 -2435
rect 4637 -2497 6099 -2485
rect 4637 -2531 4745 -2497
rect 5991 -2531 6099 -2497
rect 4637 -2563 6099 -2531
rect 4637 -2613 4695 -2563
rect 4637 -2981 4649 -2613
rect 4683 -2981 4695 -2613
rect 6041 -2613 6099 -2563
rect 4637 -3031 4695 -2981
rect 6041 -2981 6053 -2613
rect 6087 -2981 6099 -2613
rect 6041 -3031 6099 -2981
rect 4637 -3089 6099 -3031
rect 6237 -1371 7699 -1359
rect 6237 -1405 6345 -1371
rect 7591 -1405 7699 -1371
rect 6237 -1417 7699 -1405
rect 6237 -1467 6295 -1417
rect 6237 -2435 6249 -1467
rect 6283 -2435 6295 -1467
rect 7641 -1467 7699 -1417
rect 6237 -2485 6295 -2435
rect 7641 -2435 7653 -1467
rect 7687 -2435 7699 -1467
rect 7641 -2485 7699 -2435
rect 6237 -2497 7699 -2485
rect 6237 -2531 6345 -2497
rect 7591 -2531 7699 -2497
rect 6237 -2563 7699 -2531
rect 6237 -2613 6295 -2563
rect 6237 -2981 6249 -2613
rect 6283 -2981 6295 -2613
rect 7641 -2613 7699 -2563
rect 6237 -3031 6295 -2981
rect 7641 -2981 7653 -2613
rect 7687 -2981 7699 -2613
rect 7641 -3031 7699 -2981
rect 6237 -3089 7699 -3031
rect 7837 -1371 9299 -1359
rect 7837 -1405 7945 -1371
rect 9191 -1405 9299 -1371
rect 7837 -1417 9299 -1405
rect 7837 -1467 7895 -1417
rect 7837 -2435 7849 -1467
rect 7883 -2435 7895 -1467
rect 9241 -1467 9299 -1417
rect 7837 -2485 7895 -2435
rect 9241 -2435 9253 -1467
rect 9287 -2435 9299 -1467
rect 9241 -2485 9299 -2435
rect 7837 -2497 9299 -2485
rect 7837 -2531 7945 -2497
rect 9191 -2531 9299 -2497
rect 7837 -2563 9299 -2531
rect 7837 -2613 7895 -2563
rect 7837 -2981 7849 -2613
rect 7883 -2981 7895 -2613
rect 9241 -2613 9299 -2563
rect 7837 -3031 7895 -2981
rect 9241 -2981 9253 -2613
rect 9287 -2981 9299 -2613
rect 9241 -3031 9299 -2981
rect 7837 -3089 9299 -3031
rect 9437 -1371 10899 -1359
rect 9437 -1405 9545 -1371
rect 10791 -1405 10899 -1371
rect 9437 -1417 10899 -1405
rect 9437 -1467 9495 -1417
rect 9437 -2435 9449 -1467
rect 9483 -2435 9495 -1467
rect 10841 -1467 10899 -1417
rect 9437 -2485 9495 -2435
rect 10841 -2435 10853 -1467
rect 10887 -2435 10899 -1467
rect 10841 -2485 10899 -2435
rect 9437 -2497 10899 -2485
rect 9437 -2531 9545 -2497
rect 10791 -2531 10899 -2497
rect 9437 -2563 10899 -2531
rect 9437 -2613 9495 -2563
rect 9437 -2981 9449 -2613
rect 9483 -2981 9495 -2613
rect 10841 -2613 10899 -2563
rect 9437 -3031 9495 -2981
rect 10841 -2981 10853 -2613
rect 10887 -2981 10899 -2613
rect 10841 -3031 10899 -2981
rect 9437 -3089 10899 -3031
rect 11037 -1371 12499 -1359
rect 11037 -1405 11145 -1371
rect 12391 -1405 12499 -1371
rect 11037 -1417 12499 -1405
rect 11037 -1467 11095 -1417
rect 11037 -2435 11049 -1467
rect 11083 -2435 11095 -1467
rect 12441 -1467 12499 -1417
rect 11037 -2485 11095 -2435
rect 12441 -2435 12453 -1467
rect 12487 -2435 12499 -1467
rect 12441 -2485 12499 -2435
rect 11037 -2497 12499 -2485
rect 11037 -2531 11145 -2497
rect 12391 -2531 12499 -2497
rect 11037 -2563 12499 -2531
rect 11037 -2613 11095 -2563
rect 11037 -2981 11049 -2613
rect 11083 -2981 11095 -2613
rect 12441 -2613 12499 -2563
rect 11037 -3031 11095 -2981
rect 12441 -2981 12453 -2613
rect 12487 -2981 12499 -2613
rect 12441 -3031 12499 -2981
rect 11037 -3089 12499 -3031
rect 12637 -1371 14099 -1359
rect 12637 -1405 12745 -1371
rect 13991 -1405 14099 -1371
rect 12637 -1417 14099 -1405
rect 12637 -1467 12695 -1417
rect 12637 -2435 12649 -1467
rect 12683 -2435 12695 -1467
rect 14041 -1467 14099 -1417
rect 12637 -2485 12695 -2435
rect 14041 -2435 14053 -1467
rect 14087 -2435 14099 -1467
rect 14041 -2485 14099 -2435
rect 12637 -2497 14099 -2485
rect 12637 -2531 12745 -2497
rect 13991 -2531 14099 -2497
rect 12637 -2563 14099 -2531
rect 12637 -2613 12695 -2563
rect 12637 -2981 12649 -2613
rect 12683 -2981 12695 -2613
rect 14041 -2613 14099 -2563
rect 12637 -3031 12695 -2981
rect 14041 -2981 14053 -2613
rect 14087 -2981 14099 -2613
rect 14041 -3031 14099 -2981
rect 12637 -3089 14099 -3031
rect 14237 -1371 15699 -1359
rect 14237 -1405 14345 -1371
rect 15591 -1405 15699 -1371
rect 14237 -1417 15699 -1405
rect 14237 -1467 14295 -1417
rect 14237 -2435 14249 -1467
rect 14283 -2435 14295 -1467
rect 15641 -1467 15699 -1417
rect 14237 -2485 14295 -2435
rect 15641 -2435 15653 -1467
rect 15687 -2435 15699 -1467
rect 15641 -2485 15699 -2435
rect 14237 -2497 15699 -2485
rect 14237 -2531 14345 -2497
rect 15591 -2531 15699 -2497
rect 14237 -2563 15699 -2531
rect 14237 -2613 14295 -2563
rect 14237 -2981 14249 -2613
rect 14283 -2981 14295 -2613
rect 15641 -2613 15699 -2563
rect 14237 -3031 14295 -2981
rect 15641 -2981 15653 -2613
rect 15687 -2981 15699 -2613
rect 15641 -3031 15699 -2981
rect 14237 -3089 15699 -3031
rect 15837 -1371 17299 -1359
rect 15837 -1405 15945 -1371
rect 17191 -1405 17299 -1371
rect 15837 -1417 17299 -1405
rect 15837 -1467 15895 -1417
rect 15837 -2435 15849 -1467
rect 15883 -2435 15895 -1467
rect 17241 -1467 17299 -1417
rect 15837 -2485 15895 -2435
rect 17241 -2435 17253 -1467
rect 17287 -2435 17299 -1467
rect 17241 -2485 17299 -2435
rect 15837 -2497 17299 -2485
rect 15837 -2531 15945 -2497
rect 17191 -2531 17299 -2497
rect 15837 -2563 17299 -2531
rect 15837 -2613 15895 -2563
rect 15837 -2981 15849 -2613
rect 15883 -2981 15895 -2613
rect 17241 -2613 17299 -2563
rect 15837 -3031 15895 -2981
rect 17241 -2981 17253 -2613
rect 17287 -2981 17299 -2613
rect 17241 -3031 17299 -2981
rect 15837 -3089 17299 -3031
rect 17437 -1371 18899 -1359
rect 17437 -1405 17545 -1371
rect 18791 -1405 18899 -1371
rect 17437 -1417 18899 -1405
rect 17437 -1467 17495 -1417
rect 17437 -2435 17449 -1467
rect 17483 -2435 17495 -1467
rect 18841 -1467 18899 -1417
rect 17437 -2485 17495 -2435
rect 18841 -2435 18853 -1467
rect 18887 -2435 18899 -1467
rect 18841 -2485 18899 -2435
rect 17437 -2497 18899 -2485
rect 17437 -2531 17545 -2497
rect 18791 -2531 18899 -2497
rect 17437 -2563 18899 -2531
rect 17437 -2613 17495 -2563
rect 17437 -2981 17449 -2613
rect 17483 -2981 17495 -2613
rect 18841 -2613 18899 -2563
rect 17437 -3031 17495 -2981
rect 18841 -2981 18853 -2613
rect 18887 -2981 18899 -2613
rect 18841 -3031 18899 -2981
rect 17437 -3089 18899 -3031
rect 19037 -1371 20499 -1359
rect 19037 -1405 19145 -1371
rect 20391 -1405 20499 -1371
rect 19037 -1417 20499 -1405
rect 19037 -1467 19095 -1417
rect 19037 -2435 19049 -1467
rect 19083 -2435 19095 -1467
rect 20441 -1467 20499 -1417
rect 19037 -2485 19095 -2435
rect 20441 -2435 20453 -1467
rect 20487 -2435 20499 -1467
rect 20441 -2485 20499 -2435
rect 19037 -2497 20499 -2485
rect 19037 -2531 19145 -2497
rect 20391 -2531 20499 -2497
rect 19037 -2563 20499 -2531
rect 19037 -2613 19095 -2563
rect 19037 -2981 19049 -2613
rect 19083 -2981 19095 -2613
rect 20441 -2613 20499 -2563
rect 19037 -3031 19095 -2981
rect 20441 -2981 20453 -2613
rect 20487 -2981 20499 -2613
rect 20441 -3031 20499 -2981
rect 19037 -3089 20499 -3031
rect 20637 -1371 22099 -1359
rect 20637 -1405 20745 -1371
rect 21991 -1405 22099 -1371
rect 20637 -1417 22099 -1405
rect 20637 -1467 20695 -1417
rect 20637 -2435 20649 -1467
rect 20683 -2435 20695 -1467
rect 22041 -1467 22099 -1417
rect 20637 -2485 20695 -2435
rect 22041 -2435 22053 -1467
rect 22087 -2435 22099 -1467
rect 22041 -2485 22099 -2435
rect 20637 -2497 22099 -2485
rect 20637 -2531 20745 -2497
rect 21991 -2531 22099 -2497
rect 20637 -2563 22099 -2531
rect 20637 -2613 20695 -2563
rect 20637 -2981 20649 -2613
rect 20683 -2981 20695 -2613
rect 22041 -2613 22099 -2563
rect 20637 -3031 20695 -2981
rect 22041 -2981 22053 -2613
rect 22087 -2981 22099 -2613
rect 22041 -3031 22099 -2981
rect 20637 -3089 22099 -3031
rect 22237 -1371 23699 -1359
rect 22237 -1405 22345 -1371
rect 23591 -1405 23699 -1371
rect 22237 -1417 23699 -1405
rect 22237 -1467 22295 -1417
rect 22237 -2435 22249 -1467
rect 22283 -2435 22295 -1467
rect 23641 -1467 23699 -1417
rect 22237 -2485 22295 -2435
rect 23641 -2435 23653 -1467
rect 23687 -2435 23699 -1467
rect 23641 -2485 23699 -2435
rect 22237 -2497 23699 -2485
rect 22237 -2531 22345 -2497
rect 23591 -2531 23699 -2497
rect 22237 -2563 23699 -2531
rect 22237 -2613 22295 -2563
rect 22237 -2981 22249 -2613
rect 22283 -2981 22295 -2613
rect 23641 -2613 23699 -2563
rect 22237 -3031 22295 -2981
rect 23641 -2981 23653 -2613
rect 23687 -2981 23699 -2613
rect 23641 -3031 23699 -2981
rect 22237 -3089 23699 -3031
rect 23837 -1371 25299 -1359
rect 23837 -1405 23945 -1371
rect 25191 -1405 25299 -1371
rect 23837 -1417 25299 -1405
rect 23837 -1467 23895 -1417
rect 23837 -2435 23849 -1467
rect 23883 -2435 23895 -1467
rect 25241 -1467 25299 -1417
rect 23837 -2485 23895 -2435
rect 25241 -2435 25253 -1467
rect 25287 -2435 25299 -1467
rect 25241 -2485 25299 -2435
rect 23837 -2497 25299 -2485
rect 23837 -2531 23945 -2497
rect 25191 -2531 25299 -2497
rect 23837 -2563 25299 -2531
rect 23837 -2613 23895 -2563
rect 23837 -2981 23849 -2613
rect 23883 -2981 23895 -2613
rect 25241 -2613 25299 -2563
rect 23837 -3031 23895 -2981
rect 25241 -2981 25253 -2613
rect 25287 -2981 25299 -2613
rect 25241 -3031 25299 -2981
rect 23837 -3089 25299 -3031
rect 25437 -1371 26899 -1359
rect 25437 -1405 25545 -1371
rect 26791 -1405 26899 -1371
rect 25437 -1417 26899 -1405
rect 25437 -1467 25495 -1417
rect 25437 -2435 25449 -1467
rect 25483 -2435 25495 -1467
rect 26841 -1467 26899 -1417
rect 25437 -2485 25495 -2435
rect 26841 -2435 26853 -1467
rect 26887 -2435 26899 -1467
rect 26841 -2485 26899 -2435
rect 25437 -2497 26899 -2485
rect 25437 -2531 25545 -2497
rect 26791 -2531 26899 -2497
rect 25437 -2563 26899 -2531
rect 25437 -2613 25495 -2563
rect 25437 -2981 25449 -2613
rect 25483 -2981 25495 -2613
rect 26841 -2613 26899 -2563
rect 25437 -3031 25495 -2981
rect 26841 -2981 26853 -2613
rect 26887 -2981 26899 -2613
rect 26841 -3031 26899 -2981
rect 25437 -3089 26899 -3031
rect 27037 -1371 28499 -1359
rect 27037 -1405 27145 -1371
rect 28391 -1405 28499 -1371
rect 27037 -1417 28499 -1405
rect 27037 -1467 27095 -1417
rect 27037 -2435 27049 -1467
rect 27083 -2435 27095 -1467
rect 28441 -1467 28499 -1417
rect 27037 -2485 27095 -2435
rect 28441 -2435 28453 -1467
rect 28487 -2435 28499 -1467
rect 28441 -2485 28499 -2435
rect 27037 -2497 28499 -2485
rect 27037 -2531 27145 -2497
rect 28391 -2531 28499 -2497
rect 27037 -2563 28499 -2531
rect 27037 -2613 27095 -2563
rect 27037 -2981 27049 -2613
rect 27083 -2981 27095 -2613
rect 28441 -2613 28499 -2563
rect 27037 -3031 27095 -2981
rect 28441 -2981 28453 -2613
rect 28487 -2981 28499 -2613
rect 28441 -3031 28499 -2981
rect 27037 -3089 28499 -3031
rect 28637 -1371 30099 -1359
rect 28637 -1405 28745 -1371
rect 29991 -1405 30099 -1371
rect 28637 -1417 30099 -1405
rect 28637 -1467 28695 -1417
rect 28637 -2435 28649 -1467
rect 28683 -2435 28695 -1467
rect 30041 -1467 30099 -1417
rect 28637 -2485 28695 -2435
rect 30041 -2435 30053 -1467
rect 30087 -2435 30099 -1467
rect 30041 -2485 30099 -2435
rect 28637 -2497 30099 -2485
rect 28637 -2531 28745 -2497
rect 29991 -2531 30099 -2497
rect 28637 -2563 30099 -2531
rect 28637 -2613 28695 -2563
rect 28637 -2981 28649 -2613
rect 28683 -2981 28695 -2613
rect 30041 -2613 30099 -2563
rect 28637 -3031 28695 -2981
rect 30041 -2981 30053 -2613
rect 30087 -2981 30099 -2613
rect 30041 -3031 30099 -2981
rect 28637 -3089 30099 -3031
rect 30237 -1371 31699 -1359
rect 30237 -1405 30345 -1371
rect 31591 -1405 31699 -1371
rect 30237 -1417 31699 -1405
rect 30237 -1467 30295 -1417
rect 30237 -2435 30249 -1467
rect 30283 -2435 30295 -1467
rect 31641 -1467 31699 -1417
rect 30237 -2485 30295 -2435
rect 31641 -2435 31653 -1467
rect 31687 -2435 31699 -1467
rect 31641 -2485 31699 -2435
rect 30237 -2497 31699 -2485
rect 30237 -2531 30345 -2497
rect 31591 -2531 31699 -2497
rect 30237 -2563 31699 -2531
rect 30237 -2613 30295 -2563
rect 30237 -2981 30249 -2613
rect 30283 -2981 30295 -2613
rect 31641 -2613 31699 -2563
rect 30237 -3031 30295 -2981
rect 31641 -2981 31653 -2613
rect 31687 -2981 31699 -2613
rect 31641 -3031 31699 -2981
rect 30237 -3089 31699 -3031
rect 31837 -1371 33299 -1359
rect 31837 -1405 31945 -1371
rect 33191 -1405 33299 -1371
rect 31837 -1417 33299 -1405
rect 31837 -1467 31895 -1417
rect 31837 -2435 31849 -1467
rect 31883 -2435 31895 -1467
rect 33241 -1467 33299 -1417
rect 31837 -2485 31895 -2435
rect 33241 -2435 33253 -1467
rect 33287 -2435 33299 -1467
rect 33241 -2485 33299 -2435
rect 31837 -2497 33299 -2485
rect 31837 -2531 31945 -2497
rect 33191 -2531 33299 -2497
rect 31837 -2563 33299 -2531
rect 31837 -2613 31895 -2563
rect 31837 -2981 31849 -2613
rect 31883 -2981 31895 -2613
rect 33241 -2613 33299 -2563
rect 31837 -3031 31895 -2981
rect 33241 -2981 33253 -2613
rect 33287 -2981 33299 -2613
rect 33241 -3031 33299 -2981
rect 31837 -3089 33299 -3031
rect 33437 -1371 34899 -1359
rect 33437 -1405 33545 -1371
rect 34791 -1405 34899 -1371
rect 33437 -1417 34899 -1405
rect 33437 -1467 33495 -1417
rect 33437 -2435 33449 -1467
rect 33483 -2435 33495 -1467
rect 34841 -1467 34899 -1417
rect 33437 -2485 33495 -2435
rect 34841 -2435 34853 -1467
rect 34887 -2435 34899 -1467
rect 34841 -2485 34899 -2435
rect 33437 -2497 34899 -2485
rect 33437 -2531 33545 -2497
rect 34791 -2531 34899 -2497
rect 33437 -2563 34899 -2531
rect 33437 -2613 33495 -2563
rect 33437 -2981 33449 -2613
rect 33483 -2981 33495 -2613
rect 34841 -2613 34899 -2563
rect 33437 -3031 33495 -2981
rect 34841 -2981 34853 -2613
rect 34887 -2981 34899 -2613
rect 34841 -3031 34899 -2981
rect 33437 -3089 34899 -3031
rect 35037 -1371 36499 -1359
rect 35037 -1405 35145 -1371
rect 36391 -1405 36499 -1371
rect 35037 -1417 36499 -1405
rect 35037 -1467 35095 -1417
rect 35037 -2435 35049 -1467
rect 35083 -2435 35095 -1467
rect 36441 -1467 36499 -1417
rect 35037 -2485 35095 -2435
rect 36441 -2435 36453 -1467
rect 36487 -2435 36499 -1467
rect 36441 -2485 36499 -2435
rect 35037 -2497 36499 -2485
rect 35037 -2531 35145 -2497
rect 36391 -2531 36499 -2497
rect 35037 -2563 36499 -2531
rect 35037 -2613 35095 -2563
rect 35037 -2981 35049 -2613
rect 35083 -2981 35095 -2613
rect 36441 -2613 36499 -2563
rect 35037 -3031 35095 -2981
rect 36441 -2981 36453 -2613
rect 36487 -2981 36499 -2613
rect 36441 -3031 36499 -2981
rect 35037 -3089 36499 -3031
rect 36637 -1371 38099 -1359
rect 36637 -1405 36745 -1371
rect 37991 -1405 38099 -1371
rect 36637 -1417 38099 -1405
rect 36637 -1467 36695 -1417
rect 36637 -2435 36649 -1467
rect 36683 -2435 36695 -1467
rect 38041 -1467 38099 -1417
rect 36637 -2485 36695 -2435
rect 38041 -2435 38053 -1467
rect 38087 -2435 38099 -1467
rect 38041 -2485 38099 -2435
rect 36637 -2497 38099 -2485
rect 36637 -2531 36745 -2497
rect 37991 -2531 38099 -2497
rect 36637 -2563 38099 -2531
rect 36637 -2613 36695 -2563
rect 36637 -2981 36649 -2613
rect 36683 -2981 36695 -2613
rect 38041 -2613 38099 -2563
rect 36637 -3031 36695 -2981
rect 38041 -2981 38053 -2613
rect 38087 -2981 38099 -2613
rect 38041 -3031 38099 -2981
rect 36637 -3089 38099 -3031
rect -163 -3171 1299 -3159
rect -163 -3205 -55 -3171
rect 1191 -3205 1299 -3171
rect -163 -3217 1299 -3205
rect -163 -3267 -105 -3217
rect -163 -4235 -151 -3267
rect -117 -4235 -105 -3267
rect 1241 -3267 1299 -3217
rect -163 -4285 -105 -4235
rect 1241 -4235 1253 -3267
rect 1287 -4235 1299 -3267
rect 1241 -4285 1299 -4235
rect -163 -4297 1299 -4285
rect -163 -4331 -55 -4297
rect 1191 -4331 1299 -4297
rect -163 -4363 1299 -4331
rect -163 -4413 -105 -4363
rect -163 -4781 -151 -4413
rect -117 -4781 -105 -4413
rect 1241 -4413 1299 -4363
rect -163 -4831 -105 -4781
rect 1241 -4781 1253 -4413
rect 1287 -4781 1299 -4413
rect 1241 -4831 1299 -4781
rect -163 -4889 1299 -4831
rect 1437 -3171 2899 -3159
rect 1437 -3205 1545 -3171
rect 2791 -3205 2899 -3171
rect 1437 -3217 2899 -3205
rect 1437 -3267 1495 -3217
rect 1437 -4235 1449 -3267
rect 1483 -4235 1495 -3267
rect 2841 -3267 2899 -3217
rect 1437 -4285 1495 -4235
rect 2841 -4235 2853 -3267
rect 2887 -4235 2899 -3267
rect 2841 -4285 2899 -4235
rect 1437 -4297 2899 -4285
rect 1437 -4331 1545 -4297
rect 2791 -4331 2899 -4297
rect 1437 -4363 2899 -4331
rect 1437 -4413 1495 -4363
rect 1437 -4781 1449 -4413
rect 1483 -4781 1495 -4413
rect 2841 -4413 2899 -4363
rect 1437 -4831 1495 -4781
rect 2841 -4781 2853 -4413
rect 2887 -4781 2899 -4413
rect 2841 -4831 2899 -4781
rect 1437 -4889 2899 -4831
rect 3037 -3171 4499 -3159
rect 3037 -3205 3145 -3171
rect 4391 -3205 4499 -3171
rect 3037 -3217 4499 -3205
rect 3037 -3267 3095 -3217
rect 3037 -4235 3049 -3267
rect 3083 -4235 3095 -3267
rect 4441 -3267 4499 -3217
rect 3037 -4285 3095 -4235
rect 4441 -4235 4453 -3267
rect 4487 -4235 4499 -3267
rect 4441 -4285 4499 -4235
rect 3037 -4297 4499 -4285
rect 3037 -4331 3145 -4297
rect 4391 -4331 4499 -4297
rect 3037 -4363 4499 -4331
rect 3037 -4413 3095 -4363
rect 3037 -4781 3049 -4413
rect 3083 -4781 3095 -4413
rect 4441 -4413 4499 -4363
rect 3037 -4831 3095 -4781
rect 4441 -4781 4453 -4413
rect 4487 -4781 4499 -4413
rect 4441 -4831 4499 -4781
rect 3037 -4889 4499 -4831
rect 4637 -3171 6099 -3159
rect 4637 -3205 4745 -3171
rect 5991 -3205 6099 -3171
rect 4637 -3217 6099 -3205
rect 4637 -3267 4695 -3217
rect 4637 -4235 4649 -3267
rect 4683 -4235 4695 -3267
rect 6041 -3267 6099 -3217
rect 4637 -4285 4695 -4235
rect 6041 -4235 6053 -3267
rect 6087 -4235 6099 -3267
rect 6041 -4285 6099 -4235
rect 4637 -4297 6099 -4285
rect 4637 -4331 4745 -4297
rect 5991 -4331 6099 -4297
rect 4637 -4363 6099 -4331
rect 4637 -4413 4695 -4363
rect 4637 -4781 4649 -4413
rect 4683 -4781 4695 -4413
rect 6041 -4413 6099 -4363
rect 4637 -4831 4695 -4781
rect 6041 -4781 6053 -4413
rect 6087 -4781 6099 -4413
rect 6041 -4831 6099 -4781
rect 4637 -4889 6099 -4831
rect 6237 -3171 7699 -3159
rect 6237 -3205 6345 -3171
rect 7591 -3205 7699 -3171
rect 6237 -3217 7699 -3205
rect 6237 -3267 6295 -3217
rect 6237 -4235 6249 -3267
rect 6283 -4235 6295 -3267
rect 7641 -3267 7699 -3217
rect 6237 -4285 6295 -4235
rect 7641 -4235 7653 -3267
rect 7687 -4235 7699 -3267
rect 7641 -4285 7699 -4235
rect 6237 -4297 7699 -4285
rect 6237 -4331 6345 -4297
rect 7591 -4331 7699 -4297
rect 6237 -4363 7699 -4331
rect 6237 -4413 6295 -4363
rect 6237 -4781 6249 -4413
rect 6283 -4781 6295 -4413
rect 7641 -4413 7699 -4363
rect 6237 -4831 6295 -4781
rect 7641 -4781 7653 -4413
rect 7687 -4781 7699 -4413
rect 7641 -4831 7699 -4781
rect 6237 -4889 7699 -4831
rect 7837 -3171 9299 -3159
rect 7837 -3205 7945 -3171
rect 9191 -3205 9299 -3171
rect 7837 -3217 9299 -3205
rect 7837 -3267 7895 -3217
rect 7837 -4235 7849 -3267
rect 7883 -4235 7895 -3267
rect 9241 -3267 9299 -3217
rect 7837 -4285 7895 -4235
rect 9241 -4235 9253 -3267
rect 9287 -4235 9299 -3267
rect 9241 -4285 9299 -4235
rect 7837 -4297 9299 -4285
rect 7837 -4331 7945 -4297
rect 9191 -4331 9299 -4297
rect 7837 -4363 9299 -4331
rect 7837 -4413 7895 -4363
rect 7837 -4781 7849 -4413
rect 7883 -4781 7895 -4413
rect 9241 -4413 9299 -4363
rect 7837 -4831 7895 -4781
rect 9241 -4781 9253 -4413
rect 9287 -4781 9299 -4413
rect 9241 -4831 9299 -4781
rect 7837 -4889 9299 -4831
rect 9437 -3171 10899 -3159
rect 9437 -3205 9545 -3171
rect 10791 -3205 10899 -3171
rect 9437 -3217 10899 -3205
rect 9437 -3267 9495 -3217
rect 9437 -4235 9449 -3267
rect 9483 -4235 9495 -3267
rect 10841 -3267 10899 -3217
rect 9437 -4285 9495 -4235
rect 10841 -4235 10853 -3267
rect 10887 -4235 10899 -3267
rect 10841 -4285 10899 -4235
rect 9437 -4297 10899 -4285
rect 9437 -4331 9545 -4297
rect 10791 -4331 10899 -4297
rect 9437 -4363 10899 -4331
rect 9437 -4413 9495 -4363
rect 9437 -4781 9449 -4413
rect 9483 -4781 9495 -4413
rect 10841 -4413 10899 -4363
rect 9437 -4831 9495 -4781
rect 10841 -4781 10853 -4413
rect 10887 -4781 10899 -4413
rect 10841 -4831 10899 -4781
rect 9437 -4889 10899 -4831
rect 11037 -3171 12499 -3159
rect 11037 -3205 11145 -3171
rect 12391 -3205 12499 -3171
rect 11037 -3217 12499 -3205
rect 11037 -3267 11095 -3217
rect 11037 -4235 11049 -3267
rect 11083 -4235 11095 -3267
rect 12441 -3267 12499 -3217
rect 11037 -4285 11095 -4235
rect 12441 -4235 12453 -3267
rect 12487 -4235 12499 -3267
rect 12441 -4285 12499 -4235
rect 11037 -4297 12499 -4285
rect 11037 -4331 11145 -4297
rect 12391 -4331 12499 -4297
rect 11037 -4363 12499 -4331
rect 11037 -4413 11095 -4363
rect 11037 -4781 11049 -4413
rect 11083 -4781 11095 -4413
rect 12441 -4413 12499 -4363
rect 11037 -4831 11095 -4781
rect 12441 -4781 12453 -4413
rect 12487 -4781 12499 -4413
rect 12441 -4831 12499 -4781
rect 11037 -4889 12499 -4831
rect 12637 -3171 14099 -3159
rect 12637 -3205 12745 -3171
rect 13991 -3205 14099 -3171
rect 12637 -3217 14099 -3205
rect 12637 -3267 12695 -3217
rect 12637 -4235 12649 -3267
rect 12683 -4235 12695 -3267
rect 14041 -3267 14099 -3217
rect 12637 -4285 12695 -4235
rect 14041 -4235 14053 -3267
rect 14087 -4235 14099 -3267
rect 14041 -4285 14099 -4235
rect 12637 -4297 14099 -4285
rect 12637 -4331 12745 -4297
rect 13991 -4331 14099 -4297
rect 12637 -4363 14099 -4331
rect 12637 -4413 12695 -4363
rect 12637 -4781 12649 -4413
rect 12683 -4781 12695 -4413
rect 14041 -4413 14099 -4363
rect 12637 -4831 12695 -4781
rect 14041 -4781 14053 -4413
rect 14087 -4781 14099 -4413
rect 14041 -4831 14099 -4781
rect 12637 -4889 14099 -4831
rect 14237 -3171 15699 -3159
rect 14237 -3205 14345 -3171
rect 15591 -3205 15699 -3171
rect 14237 -3217 15699 -3205
rect 14237 -3267 14295 -3217
rect 14237 -4235 14249 -3267
rect 14283 -4235 14295 -3267
rect 15641 -3267 15699 -3217
rect 14237 -4285 14295 -4235
rect 15641 -4235 15653 -3267
rect 15687 -4235 15699 -3267
rect 15641 -4285 15699 -4235
rect 14237 -4297 15699 -4285
rect 14237 -4331 14345 -4297
rect 15591 -4331 15699 -4297
rect 14237 -4363 15699 -4331
rect 14237 -4413 14295 -4363
rect 14237 -4781 14249 -4413
rect 14283 -4781 14295 -4413
rect 15641 -4413 15699 -4363
rect 14237 -4831 14295 -4781
rect 15641 -4781 15653 -4413
rect 15687 -4781 15699 -4413
rect 15641 -4831 15699 -4781
rect 14237 -4889 15699 -4831
rect 15837 -3171 17299 -3159
rect 15837 -3205 15945 -3171
rect 17191 -3205 17299 -3171
rect 15837 -3217 17299 -3205
rect 15837 -3267 15895 -3217
rect 15837 -4235 15849 -3267
rect 15883 -4235 15895 -3267
rect 17241 -3267 17299 -3217
rect 15837 -4285 15895 -4235
rect 17241 -4235 17253 -3267
rect 17287 -4235 17299 -3267
rect 17241 -4285 17299 -4235
rect 15837 -4297 17299 -4285
rect 15837 -4331 15945 -4297
rect 17191 -4331 17299 -4297
rect 15837 -4363 17299 -4331
rect 15837 -4413 15895 -4363
rect 15837 -4781 15849 -4413
rect 15883 -4781 15895 -4413
rect 17241 -4413 17299 -4363
rect 15837 -4831 15895 -4781
rect 17241 -4781 17253 -4413
rect 17287 -4781 17299 -4413
rect 17241 -4831 17299 -4781
rect 15837 -4889 17299 -4831
rect 17437 -3171 18899 -3159
rect 17437 -3205 17545 -3171
rect 18791 -3205 18899 -3171
rect 17437 -3217 18899 -3205
rect 17437 -3267 17495 -3217
rect 17437 -4235 17449 -3267
rect 17483 -4235 17495 -3267
rect 18841 -3267 18899 -3217
rect 17437 -4285 17495 -4235
rect 18841 -4235 18853 -3267
rect 18887 -4235 18899 -3267
rect 18841 -4285 18899 -4235
rect 17437 -4297 18899 -4285
rect 17437 -4331 17545 -4297
rect 18791 -4331 18899 -4297
rect 17437 -4363 18899 -4331
rect 17437 -4413 17495 -4363
rect 17437 -4781 17449 -4413
rect 17483 -4781 17495 -4413
rect 18841 -4413 18899 -4363
rect 17437 -4831 17495 -4781
rect 18841 -4781 18853 -4413
rect 18887 -4781 18899 -4413
rect 18841 -4831 18899 -4781
rect 17437 -4889 18899 -4831
rect 19037 -3171 20499 -3159
rect 19037 -3205 19145 -3171
rect 20391 -3205 20499 -3171
rect 19037 -3217 20499 -3205
rect 19037 -3267 19095 -3217
rect 19037 -4235 19049 -3267
rect 19083 -4235 19095 -3267
rect 20441 -3267 20499 -3217
rect 19037 -4285 19095 -4235
rect 20441 -4235 20453 -3267
rect 20487 -4235 20499 -3267
rect 20441 -4285 20499 -4235
rect 19037 -4297 20499 -4285
rect 19037 -4331 19145 -4297
rect 20391 -4331 20499 -4297
rect 19037 -4363 20499 -4331
rect 19037 -4413 19095 -4363
rect 19037 -4781 19049 -4413
rect 19083 -4781 19095 -4413
rect 20441 -4413 20499 -4363
rect 19037 -4831 19095 -4781
rect 20441 -4781 20453 -4413
rect 20487 -4781 20499 -4413
rect 20441 -4831 20499 -4781
rect 19037 -4889 20499 -4831
rect 20637 -3171 22099 -3159
rect 20637 -3205 20745 -3171
rect 21991 -3205 22099 -3171
rect 20637 -3217 22099 -3205
rect 20637 -3267 20695 -3217
rect 20637 -4235 20649 -3267
rect 20683 -4235 20695 -3267
rect 22041 -3267 22099 -3217
rect 20637 -4285 20695 -4235
rect 22041 -4235 22053 -3267
rect 22087 -4235 22099 -3267
rect 22041 -4285 22099 -4235
rect 20637 -4297 22099 -4285
rect 20637 -4331 20745 -4297
rect 21991 -4331 22099 -4297
rect 20637 -4363 22099 -4331
rect 20637 -4413 20695 -4363
rect 20637 -4781 20649 -4413
rect 20683 -4781 20695 -4413
rect 22041 -4413 22099 -4363
rect 20637 -4831 20695 -4781
rect 22041 -4781 22053 -4413
rect 22087 -4781 22099 -4413
rect 22041 -4831 22099 -4781
rect 20637 -4889 22099 -4831
rect 22237 -3171 23699 -3159
rect 22237 -3205 22345 -3171
rect 23591 -3205 23699 -3171
rect 22237 -3217 23699 -3205
rect 22237 -3267 22295 -3217
rect 22237 -4235 22249 -3267
rect 22283 -4235 22295 -3267
rect 23641 -3267 23699 -3217
rect 22237 -4285 22295 -4235
rect 23641 -4235 23653 -3267
rect 23687 -4235 23699 -3267
rect 23641 -4285 23699 -4235
rect 22237 -4297 23699 -4285
rect 22237 -4331 22345 -4297
rect 23591 -4331 23699 -4297
rect 22237 -4363 23699 -4331
rect 22237 -4413 22295 -4363
rect 22237 -4781 22249 -4413
rect 22283 -4781 22295 -4413
rect 23641 -4413 23699 -4363
rect 22237 -4831 22295 -4781
rect 23641 -4781 23653 -4413
rect 23687 -4781 23699 -4413
rect 23641 -4831 23699 -4781
rect 22237 -4889 23699 -4831
rect 23837 -3171 25299 -3159
rect 23837 -3205 23945 -3171
rect 25191 -3205 25299 -3171
rect 23837 -3217 25299 -3205
rect 23837 -3267 23895 -3217
rect 23837 -4235 23849 -3267
rect 23883 -4235 23895 -3267
rect 25241 -3267 25299 -3217
rect 23837 -4285 23895 -4235
rect 25241 -4235 25253 -3267
rect 25287 -4235 25299 -3267
rect 25241 -4285 25299 -4235
rect 23837 -4297 25299 -4285
rect 23837 -4331 23945 -4297
rect 25191 -4331 25299 -4297
rect 23837 -4363 25299 -4331
rect 23837 -4413 23895 -4363
rect 23837 -4781 23849 -4413
rect 23883 -4781 23895 -4413
rect 25241 -4413 25299 -4363
rect 23837 -4831 23895 -4781
rect 25241 -4781 25253 -4413
rect 25287 -4781 25299 -4413
rect 25241 -4831 25299 -4781
rect 23837 -4889 25299 -4831
rect 25437 -3171 26899 -3159
rect 25437 -3205 25545 -3171
rect 26791 -3205 26899 -3171
rect 25437 -3217 26899 -3205
rect 25437 -3267 25495 -3217
rect 25437 -4235 25449 -3267
rect 25483 -4235 25495 -3267
rect 26841 -3267 26899 -3217
rect 25437 -4285 25495 -4235
rect 26841 -4235 26853 -3267
rect 26887 -4235 26899 -3267
rect 26841 -4285 26899 -4235
rect 25437 -4297 26899 -4285
rect 25437 -4331 25545 -4297
rect 26791 -4331 26899 -4297
rect 25437 -4363 26899 -4331
rect 25437 -4413 25495 -4363
rect 25437 -4781 25449 -4413
rect 25483 -4781 25495 -4413
rect 26841 -4413 26899 -4363
rect 25437 -4831 25495 -4781
rect 26841 -4781 26853 -4413
rect 26887 -4781 26899 -4413
rect 26841 -4831 26899 -4781
rect 25437 -4889 26899 -4831
rect 27037 -3171 28499 -3159
rect 27037 -3205 27145 -3171
rect 28391 -3205 28499 -3171
rect 27037 -3217 28499 -3205
rect 27037 -3267 27095 -3217
rect 27037 -4235 27049 -3267
rect 27083 -4235 27095 -3267
rect 28441 -3267 28499 -3217
rect 27037 -4285 27095 -4235
rect 28441 -4235 28453 -3267
rect 28487 -4235 28499 -3267
rect 28441 -4285 28499 -4235
rect 27037 -4297 28499 -4285
rect 27037 -4331 27145 -4297
rect 28391 -4331 28499 -4297
rect 27037 -4363 28499 -4331
rect 27037 -4413 27095 -4363
rect 27037 -4781 27049 -4413
rect 27083 -4781 27095 -4413
rect 28441 -4413 28499 -4363
rect 27037 -4831 27095 -4781
rect 28441 -4781 28453 -4413
rect 28487 -4781 28499 -4413
rect 28441 -4831 28499 -4781
rect 27037 -4889 28499 -4831
rect 28637 -3171 30099 -3159
rect 28637 -3205 28745 -3171
rect 29991 -3205 30099 -3171
rect 28637 -3217 30099 -3205
rect 28637 -3267 28695 -3217
rect 28637 -4235 28649 -3267
rect 28683 -4235 28695 -3267
rect 30041 -3267 30099 -3217
rect 28637 -4285 28695 -4235
rect 30041 -4235 30053 -3267
rect 30087 -4235 30099 -3267
rect 30041 -4285 30099 -4235
rect 28637 -4297 30099 -4285
rect 28637 -4331 28745 -4297
rect 29991 -4331 30099 -4297
rect 28637 -4363 30099 -4331
rect 28637 -4413 28695 -4363
rect 28637 -4781 28649 -4413
rect 28683 -4781 28695 -4413
rect 30041 -4413 30099 -4363
rect 28637 -4831 28695 -4781
rect 30041 -4781 30053 -4413
rect 30087 -4781 30099 -4413
rect 30041 -4831 30099 -4781
rect 28637 -4889 30099 -4831
rect 30237 -3171 31699 -3159
rect 30237 -3205 30345 -3171
rect 31591 -3205 31699 -3171
rect 30237 -3217 31699 -3205
rect 30237 -3267 30295 -3217
rect 30237 -4235 30249 -3267
rect 30283 -4235 30295 -3267
rect 31641 -3267 31699 -3217
rect 30237 -4285 30295 -4235
rect 31641 -4235 31653 -3267
rect 31687 -4235 31699 -3267
rect 31641 -4285 31699 -4235
rect 30237 -4297 31699 -4285
rect 30237 -4331 30345 -4297
rect 31591 -4331 31699 -4297
rect 30237 -4363 31699 -4331
rect 30237 -4413 30295 -4363
rect 30237 -4781 30249 -4413
rect 30283 -4781 30295 -4413
rect 31641 -4413 31699 -4363
rect 30237 -4831 30295 -4781
rect 31641 -4781 31653 -4413
rect 31687 -4781 31699 -4413
rect 31641 -4831 31699 -4781
rect 30237 -4889 31699 -4831
rect 31837 -3171 33299 -3159
rect 31837 -3205 31945 -3171
rect 33191 -3205 33299 -3171
rect 31837 -3217 33299 -3205
rect 31837 -3267 31895 -3217
rect 31837 -4235 31849 -3267
rect 31883 -4235 31895 -3267
rect 33241 -3267 33299 -3217
rect 31837 -4285 31895 -4235
rect 33241 -4235 33253 -3267
rect 33287 -4235 33299 -3267
rect 33241 -4285 33299 -4235
rect 31837 -4297 33299 -4285
rect 31837 -4331 31945 -4297
rect 33191 -4331 33299 -4297
rect 31837 -4363 33299 -4331
rect 31837 -4413 31895 -4363
rect 31837 -4781 31849 -4413
rect 31883 -4781 31895 -4413
rect 33241 -4413 33299 -4363
rect 31837 -4831 31895 -4781
rect 33241 -4781 33253 -4413
rect 33287 -4781 33299 -4413
rect 33241 -4831 33299 -4781
rect 31837 -4889 33299 -4831
rect 33437 -3171 34899 -3159
rect 33437 -3205 33545 -3171
rect 34791 -3205 34899 -3171
rect 33437 -3217 34899 -3205
rect 33437 -3267 33495 -3217
rect 33437 -4235 33449 -3267
rect 33483 -4235 33495 -3267
rect 34841 -3267 34899 -3217
rect 33437 -4285 33495 -4235
rect 34841 -4235 34853 -3267
rect 34887 -4235 34899 -3267
rect 34841 -4285 34899 -4235
rect 33437 -4297 34899 -4285
rect 33437 -4331 33545 -4297
rect 34791 -4331 34899 -4297
rect 33437 -4363 34899 -4331
rect 33437 -4413 33495 -4363
rect 33437 -4781 33449 -4413
rect 33483 -4781 33495 -4413
rect 34841 -4413 34899 -4363
rect 33437 -4831 33495 -4781
rect 34841 -4781 34853 -4413
rect 34887 -4781 34899 -4413
rect 34841 -4831 34899 -4781
rect 33437 -4889 34899 -4831
rect 35037 -3171 36499 -3159
rect 35037 -3205 35145 -3171
rect 36391 -3205 36499 -3171
rect 35037 -3217 36499 -3205
rect 35037 -3267 35095 -3217
rect 35037 -4235 35049 -3267
rect 35083 -4235 35095 -3267
rect 36441 -3267 36499 -3217
rect 35037 -4285 35095 -4235
rect 36441 -4235 36453 -3267
rect 36487 -4235 36499 -3267
rect 36441 -4285 36499 -4235
rect 35037 -4297 36499 -4285
rect 35037 -4331 35145 -4297
rect 36391 -4331 36499 -4297
rect 35037 -4363 36499 -4331
rect 35037 -4413 35095 -4363
rect 35037 -4781 35049 -4413
rect 35083 -4781 35095 -4413
rect 36441 -4413 36499 -4363
rect 35037 -4831 35095 -4781
rect 36441 -4781 36453 -4413
rect 36487 -4781 36499 -4413
rect 36441 -4831 36499 -4781
rect 35037 -4889 36499 -4831
rect 36637 -3171 38099 -3159
rect 36637 -3205 36745 -3171
rect 37991 -3205 38099 -3171
rect 36637 -3217 38099 -3205
rect 36637 -3267 36695 -3217
rect 36637 -4235 36649 -3267
rect 36683 -4235 36695 -3267
rect 38041 -3267 38099 -3217
rect 36637 -4285 36695 -4235
rect 38041 -4235 38053 -3267
rect 38087 -4235 38099 -3267
rect 38041 -4285 38099 -4235
rect 36637 -4297 38099 -4285
rect 36637 -4331 36745 -4297
rect 37991 -4331 38099 -4297
rect 36637 -4363 38099 -4331
rect 36637 -4413 36695 -4363
rect 36637 -4781 36649 -4413
rect 36683 -4781 36695 -4413
rect 38041 -4413 38099 -4363
rect 36637 -4831 36695 -4781
rect 38041 -4781 38053 -4413
rect 38087 -4781 38099 -4413
rect 38041 -4831 38099 -4781
rect 36637 -4889 38099 -4831
rect 27776 -24502 28960 -24490
rect 27776 -24536 27884 -24502
rect 28852 -24536 28960 -24502
rect 27776 -24548 28960 -24536
rect 27776 -24598 27834 -24548
rect 27776 -25226 27788 -24598
rect 27822 -25226 27834 -24598
rect 28902 -24598 28960 -24548
rect 27776 -25276 27834 -25226
rect 28902 -25226 28914 -24598
rect 28948 -25226 28960 -24598
rect 28902 -25276 28960 -25226
rect 27776 -25288 28960 -25276
rect 27776 -25322 27884 -25288
rect 28852 -25322 28960 -25288
rect 27776 -25334 28960 -25322
rect 27776 -25408 28958 -25396
rect 27776 -25442 27884 -25408
rect 28850 -25442 28958 -25408
rect 27776 -25454 28958 -25442
rect 27776 -25504 27834 -25454
rect 27776 -26246 27788 -25504
rect 27822 -26246 27834 -25504
rect 28900 -25504 28958 -25454
rect 27776 -26296 27834 -26246
rect 28900 -26246 28912 -25504
rect 28946 -26246 28958 -25504
rect 28900 -26296 28958 -26246
rect 27776 -26308 28958 -26296
rect 27776 -26342 27884 -26308
rect 28850 -26342 28958 -26308
rect 27776 -26354 28958 -26342
rect 27776 -26448 28958 -26436
rect 27776 -26482 27884 -26448
rect 28850 -26482 28958 -26448
rect 27776 -26494 28958 -26482
rect 27776 -26544 27834 -26494
rect 27776 -27286 27788 -26544
rect 27822 -27286 27834 -26544
rect 28900 -26544 28958 -26494
rect 27776 -27336 27834 -27286
rect 28900 -27286 28912 -26544
rect 28946 -27286 28958 -26544
rect 28900 -27336 28958 -27286
rect 27776 -27348 28958 -27336
rect 27776 -27382 27884 -27348
rect 28850 -27382 28958 -27348
rect 27776 -27394 28958 -27382
rect 27776 -27488 28958 -27476
rect 27776 -27522 27884 -27488
rect 28850 -27522 28958 -27488
rect 27776 -27534 28958 -27522
rect 27776 -27584 27834 -27534
rect 27776 -28326 27788 -27584
rect 27822 -28326 27834 -27584
rect 28900 -27584 28958 -27534
rect 27776 -28376 27834 -28326
rect 28900 -28326 28912 -27584
rect 28946 -28326 28958 -27584
rect 28900 -28376 28958 -28326
rect 27776 -28388 28958 -28376
rect 27776 -28422 27884 -28388
rect 28850 -28422 28958 -28388
rect 27776 -28434 28958 -28422
rect 27776 -28528 28958 -28516
rect 27776 -28562 27884 -28528
rect 28850 -28562 28958 -28528
rect 27776 -28574 28958 -28562
rect 27776 -28624 27834 -28574
rect 27776 -29366 27788 -28624
rect 27822 -29366 27834 -28624
rect 28900 -28624 28958 -28574
rect 27776 -29416 27834 -29366
rect 28900 -29366 28912 -28624
rect 28946 -29366 28958 -28624
rect 28900 -29416 28958 -29366
rect 27776 -29428 28958 -29416
rect 27776 -29462 27884 -29428
rect 28850 -29462 28958 -29428
rect 27776 -29474 28958 -29462
rect 31667 -29331 33786 -29319
rect 31667 -29365 31775 -29331
rect 32043 -29365 32215 -29331
rect 32483 -29365 32655 -29331
rect 32923 -29365 33094 -29331
rect 33678 -29365 33786 -29331
rect 31667 -29377 33786 -29365
rect 31667 -29427 31725 -29377
rect 27776 -29568 28958 -29556
rect 27776 -29602 27884 -29568
rect 28850 -29602 28958 -29568
rect 27776 -29614 28958 -29602
rect 27776 -29664 27834 -29614
rect 27776 -30406 27788 -29664
rect 27822 -30406 27834 -29664
rect 28900 -29664 28958 -29614
rect 27776 -30456 27834 -30406
rect 28900 -30406 28912 -29664
rect 28946 -30406 28958 -29664
rect 31667 -29855 31679 -29427
rect 31713 -29855 31725 -29427
rect 32093 -29427 32165 -29377
rect 31667 -29905 31725 -29855
rect 32093 -29855 32105 -29427
rect 32139 -29855 32165 -29427
rect 32093 -29905 32165 -29855
rect 32533 -29905 32605 -29377
rect 32973 -29427 33044 -29377
rect 32973 -29855 32998 -29427
rect 33032 -29855 33044 -29427
rect 33728 -29427 33786 -29377
rect 32973 -29905 33044 -29855
rect 33728 -29855 33740 -29427
rect 33774 -29855 33786 -29427
rect 33728 -29905 33786 -29855
rect 31667 -29917 33786 -29905
rect 31667 -29951 31775 -29917
rect 32043 -29951 32215 -29917
rect 32483 -29951 32655 -29917
rect 32923 -29951 33094 -29917
rect 33678 -29951 33786 -29917
rect 31667 -29963 33786 -29951
rect 33867 -29331 35986 -29319
rect 33867 -29365 33975 -29331
rect 34243 -29365 34415 -29331
rect 34683 -29365 34855 -29331
rect 35123 -29365 35294 -29331
rect 35878 -29365 35986 -29331
rect 33867 -29377 35986 -29365
rect 33867 -29427 33925 -29377
rect 33867 -29855 33879 -29427
rect 33913 -29855 33925 -29427
rect 34293 -29427 34365 -29377
rect 33867 -29905 33925 -29855
rect 34293 -29855 34305 -29427
rect 34339 -29855 34365 -29427
rect 34293 -29905 34365 -29855
rect 34733 -29905 34805 -29377
rect 35173 -29427 35244 -29377
rect 35173 -29855 35198 -29427
rect 35232 -29855 35244 -29427
rect 35928 -29427 35986 -29377
rect 35173 -29905 35244 -29855
rect 35928 -29855 35940 -29427
rect 35974 -29855 35986 -29427
rect 35928 -29905 35986 -29855
rect 33867 -29917 35986 -29905
rect 33867 -29951 33975 -29917
rect 34243 -29951 34415 -29917
rect 34683 -29951 34855 -29917
rect 35123 -29951 35294 -29917
rect 35878 -29951 35986 -29917
rect 33867 -29963 35986 -29951
rect 36067 -29331 38186 -29319
rect 36067 -29365 36175 -29331
rect 36443 -29365 36615 -29331
rect 36883 -29365 37055 -29331
rect 37323 -29365 37494 -29331
rect 38078 -29365 38186 -29331
rect 36067 -29377 38186 -29365
rect 36067 -29427 36125 -29377
rect 36067 -29855 36079 -29427
rect 36113 -29855 36125 -29427
rect 36493 -29427 36565 -29377
rect 36067 -29905 36125 -29855
rect 36493 -29855 36505 -29427
rect 36539 -29855 36565 -29427
rect 36493 -29905 36565 -29855
rect 36933 -29905 37005 -29377
rect 37373 -29427 37444 -29377
rect 37373 -29855 37398 -29427
rect 37432 -29855 37444 -29427
rect 38128 -29427 38186 -29377
rect 37373 -29905 37444 -29855
rect 38128 -29855 38140 -29427
rect 38174 -29855 38186 -29427
rect 38128 -29905 38186 -29855
rect 36067 -29917 38186 -29905
rect 36067 -29951 36175 -29917
rect 36443 -29951 36615 -29917
rect 36883 -29951 37055 -29917
rect 37323 -29951 37494 -29917
rect 38078 -29951 38186 -29917
rect 36067 -29963 38186 -29951
rect 28900 -30456 28958 -30406
rect 27776 -30468 28958 -30456
rect 27776 -30502 27884 -30468
rect 28850 -30502 28958 -30468
rect 27776 -30514 28958 -30502
rect 31636 -30073 33755 -30061
rect 31636 -30107 31744 -30073
rect 32328 -30107 32499 -30073
rect 32767 -30107 32939 -30073
rect 33207 -30107 33379 -30073
rect 33647 -30107 33755 -30073
rect 31636 -30119 33755 -30107
rect 31636 -30169 31694 -30119
rect 27776 -30608 28958 -30596
rect 27776 -30642 27884 -30608
rect 28850 -30642 28958 -30608
rect 27776 -30654 28958 -30642
rect 27776 -30704 27834 -30654
rect 27776 -31446 27788 -30704
rect 27822 -31446 27834 -30704
rect 28900 -30704 28958 -30654
rect 27776 -31496 27834 -31446
rect 28900 -31446 28912 -30704
rect 28946 -31446 28958 -30704
rect 31636 -30597 31648 -30169
rect 31682 -30597 31694 -30169
rect 32378 -30169 32449 -30119
rect 31636 -30647 31694 -30597
rect 32378 -30597 32390 -30169
rect 32424 -30597 32449 -30169
rect 32378 -30647 32449 -30597
rect 32817 -30647 32889 -30119
rect 33257 -30169 33329 -30119
rect 33257 -30597 33283 -30169
rect 33317 -30597 33329 -30169
rect 33697 -30169 33755 -30119
rect 33257 -30647 33329 -30597
rect 33697 -30597 33709 -30169
rect 33743 -30597 33755 -30169
rect 33697 -30647 33755 -30597
rect 31636 -30659 33755 -30647
rect 31636 -30693 31744 -30659
rect 32328 -30693 32499 -30659
rect 32767 -30693 32939 -30659
rect 33207 -30693 33379 -30659
rect 33647 -30693 33755 -30659
rect 31636 -30705 33755 -30693
rect 33836 -30073 35955 -30061
rect 33836 -30107 33944 -30073
rect 34528 -30107 34699 -30073
rect 34967 -30107 35139 -30073
rect 35407 -30107 35579 -30073
rect 35847 -30107 35955 -30073
rect 33836 -30119 35955 -30107
rect 33836 -30169 33894 -30119
rect 33836 -30597 33848 -30169
rect 33882 -30597 33894 -30169
rect 34578 -30169 34649 -30119
rect 33836 -30647 33894 -30597
rect 34578 -30597 34590 -30169
rect 34624 -30597 34649 -30169
rect 34578 -30647 34649 -30597
rect 35017 -30647 35089 -30119
rect 35457 -30169 35529 -30119
rect 35457 -30597 35483 -30169
rect 35517 -30597 35529 -30169
rect 35897 -30169 35955 -30119
rect 35457 -30647 35529 -30597
rect 35897 -30597 35909 -30169
rect 35943 -30597 35955 -30169
rect 35897 -30647 35955 -30597
rect 33836 -30659 35955 -30647
rect 33836 -30693 33944 -30659
rect 34528 -30693 34699 -30659
rect 34967 -30693 35139 -30659
rect 35407 -30693 35579 -30659
rect 35847 -30693 35955 -30659
rect 33836 -30705 35955 -30693
rect 36036 -30073 38155 -30061
rect 36036 -30107 36144 -30073
rect 36728 -30107 36899 -30073
rect 37167 -30107 37339 -30073
rect 37607 -30107 37779 -30073
rect 38047 -30107 38155 -30073
rect 36036 -30119 38155 -30107
rect 36036 -30169 36094 -30119
rect 36036 -30597 36048 -30169
rect 36082 -30597 36094 -30169
rect 36778 -30169 36849 -30119
rect 36036 -30647 36094 -30597
rect 36778 -30597 36790 -30169
rect 36824 -30597 36849 -30169
rect 36778 -30647 36849 -30597
rect 37217 -30647 37289 -30119
rect 37657 -30169 37729 -30119
rect 37657 -30597 37683 -30169
rect 37717 -30597 37729 -30169
rect 38097 -30169 38155 -30119
rect 37657 -30647 37729 -30597
rect 38097 -30597 38109 -30169
rect 38143 -30597 38155 -30169
rect 38097 -30647 38155 -30597
rect 36036 -30659 38155 -30647
rect 36036 -30693 36144 -30659
rect 36728 -30693 36899 -30659
rect 37167 -30693 37339 -30659
rect 37607 -30693 37779 -30659
rect 38047 -30693 38155 -30659
rect 36036 -30705 38155 -30693
rect 28900 -31496 28958 -31446
rect 27776 -31508 28958 -31496
rect 27776 -31542 27884 -31508
rect 28850 -31542 28958 -31508
rect 27776 -31554 28958 -31542
<< mvnsubdiff >>
rect 27766 11592 28958 11604
rect 27766 11558 27874 11592
rect 28850 11558 28958 11592
rect 27766 11546 28958 11558
rect 27766 11496 27824 11546
rect 27766 10754 27778 11496
rect 27812 10754 27824 11496
rect 28900 11496 28958 11546
rect 27766 10704 27824 10754
rect 28900 10754 28912 11496
rect 28946 10754 28958 11496
rect 28900 10704 28958 10754
rect 27766 10692 28958 10704
rect 27766 10658 27874 10692
rect 28850 10658 28958 10692
rect 27766 10646 28958 10658
rect 29998 11126 32076 11138
rect 29998 11092 30106 11126
rect 30674 11092 30820 11126
rect 31088 11092 31260 11126
rect 31528 11092 31700 11126
rect 31968 11092 32076 11126
rect 29998 11080 32076 11092
rect 29998 11030 30056 11080
rect 29998 10684 30010 11030
rect 30044 10684 30056 11030
rect 30712 11030 30782 11080
rect 29998 10634 30056 10684
rect 30712 10684 30736 11030
rect 30770 10684 30782 11030
rect 30712 10634 30782 10684
rect 29998 10622 30782 10634
rect 29998 10588 30106 10622
rect 30674 10588 30782 10622
rect 29998 10576 30782 10588
rect 27766 10552 28958 10564
rect 27766 10518 27874 10552
rect 28850 10518 28958 10552
rect 27766 10506 28958 10518
rect 27766 10456 27824 10506
rect 27766 9714 27778 10456
rect 27812 9714 27824 10456
rect 28900 10456 28958 10506
rect 27766 9664 27824 9714
rect 28900 9714 28912 10456
rect 28946 9714 28958 10456
rect 30712 10334 30770 10576
rect 31138 10334 31210 11080
rect 31578 11030 31650 11080
rect 31578 10384 31604 11030
rect 31638 10384 31650 11030
rect 32018 11030 32076 11080
rect 31578 10334 31650 10384
rect 32018 10384 32030 11030
rect 32064 10384 32076 11030
rect 32198 11126 34276 11138
rect 32198 11092 32306 11126
rect 32874 11092 33020 11126
rect 33288 11092 33460 11126
rect 33728 11092 33900 11126
rect 34168 11092 34276 11126
rect 32198 11080 34276 11092
rect 32198 11030 32256 11080
rect 32198 10684 32210 11030
rect 32244 10684 32256 11030
rect 32912 11030 32982 11080
rect 32198 10634 32256 10684
rect 32912 10684 32936 11030
rect 32970 10684 32982 11030
rect 32912 10634 32982 10684
rect 32198 10622 32982 10634
rect 32198 10588 32306 10622
rect 32874 10588 32982 10622
rect 32198 10576 32982 10588
rect 32018 10334 32076 10384
rect 30712 10322 32076 10334
rect 30712 10288 30820 10322
rect 31088 10288 31260 10322
rect 31528 10288 31700 10322
rect 31968 10288 32076 10322
rect 30712 10276 32076 10288
rect 32912 10334 32970 10576
rect 33338 10334 33410 11080
rect 33778 11030 33850 11080
rect 33778 10384 33804 11030
rect 33838 10384 33850 11030
rect 34218 11030 34276 11080
rect 33778 10334 33850 10384
rect 34218 10384 34230 11030
rect 34264 10384 34276 11030
rect 34398 11126 36476 11138
rect 34398 11092 34506 11126
rect 35074 11092 35220 11126
rect 35488 11092 35660 11126
rect 35928 11092 36100 11126
rect 36368 11092 36476 11126
rect 34398 11080 36476 11092
rect 34398 11030 34456 11080
rect 34398 10684 34410 11030
rect 34444 10684 34456 11030
rect 35112 11030 35182 11080
rect 34398 10634 34456 10684
rect 35112 10684 35136 11030
rect 35170 10684 35182 11030
rect 35112 10634 35182 10684
rect 34398 10622 35182 10634
rect 34398 10588 34506 10622
rect 35074 10588 35182 10622
rect 34398 10576 35182 10588
rect 34218 10334 34276 10384
rect 32912 10322 34276 10334
rect 32912 10288 33020 10322
rect 33288 10288 33460 10322
rect 33728 10288 33900 10322
rect 34168 10288 34276 10322
rect 32912 10276 34276 10288
rect 35112 10334 35170 10576
rect 35538 10334 35610 11080
rect 35978 11030 36050 11080
rect 35978 10384 36004 11030
rect 36038 10384 36050 11030
rect 36418 11030 36476 11080
rect 35978 10334 36050 10384
rect 36418 10384 36430 11030
rect 36464 10384 36476 11030
rect 36418 10334 36476 10384
rect 35112 10322 36476 10334
rect 35112 10288 35220 10322
rect 35488 10288 35660 10322
rect 35928 10288 36100 10322
rect 36368 10288 36476 10322
rect 35112 10276 36476 10288
rect 28900 9664 28958 9714
rect 27766 9652 28958 9664
rect 27766 9618 27874 9652
rect 28850 9618 28958 9652
rect 27766 9606 28958 9618
rect 29586 9816 31628 9828
rect 29586 9782 29694 9816
rect 31520 9782 31628 9816
rect 29586 9770 31628 9782
rect 29586 9720 29644 9770
rect 27766 9512 28958 9524
rect 27766 9478 27874 9512
rect 28850 9478 28958 9512
rect 27766 9466 28958 9478
rect 27766 9416 27824 9466
rect 27766 8674 27778 9416
rect 27812 8674 27824 9416
rect 28900 9416 28958 9466
rect 27766 8624 27824 8674
rect 28900 8674 28912 9416
rect 28946 8674 28958 9416
rect 29586 9074 29598 9720
rect 29632 9074 29644 9720
rect 31570 9720 31628 9770
rect 29586 9024 29644 9074
rect 31570 9074 31582 9720
rect 31616 9074 31628 9720
rect 31570 9024 31628 9074
rect 29586 9012 31628 9024
rect 29586 8978 29694 9012
rect 31520 8978 31628 9012
rect 29586 8966 31628 8978
rect 28900 8624 28958 8674
rect 27766 8612 28958 8624
rect 27766 8578 27874 8612
rect 28850 8578 28958 8612
rect 27766 8566 28958 8578
rect 29586 8812 31628 8824
rect 29586 8778 29694 8812
rect 31520 8778 31628 8812
rect 29586 8766 31628 8778
rect 29586 8716 29644 8766
rect 27766 8472 28958 8484
rect 27766 8438 27874 8472
rect 28850 8438 28958 8472
rect 27766 8426 28958 8438
rect 27766 8376 27824 8426
rect 27766 7634 27778 8376
rect 27812 7634 27824 8376
rect 28900 8376 28958 8426
rect 27766 7584 27824 7634
rect 28900 7634 28912 8376
rect 28946 7634 28958 8376
rect 28900 7584 28958 7634
rect 27766 7572 28958 7584
rect 27766 7538 27874 7572
rect 28850 7538 28958 7572
rect 27766 7526 28958 7538
rect 27766 7432 28958 7444
rect 27766 7398 27874 7432
rect 28850 7398 28958 7432
rect 27766 7386 28958 7398
rect 27766 7336 27824 7386
rect 27766 6594 27778 7336
rect 27812 6594 27824 7336
rect 28900 7336 28958 7386
rect 27766 6544 27824 6594
rect 28900 6594 28912 7336
rect 28946 6594 28958 7336
rect 29586 7434 29598 8716
rect 29632 7434 29644 8716
rect 31570 8716 31628 8766
rect 29586 7384 29644 7434
rect 31570 7434 31582 8716
rect 31616 7434 31628 8716
rect 31570 7384 31628 7434
rect 29586 7372 31628 7384
rect 29586 7338 29694 7372
rect 31520 7338 31628 7372
rect 29586 7326 31628 7338
rect 29526 7152 30788 7210
rect 29526 7102 29584 7152
rect 29526 6734 29538 7102
rect 29572 6734 29584 7102
rect 30730 7102 30788 7152
rect 29526 6684 29584 6734
rect 30730 6734 30742 7102
rect 30776 6734 30788 7102
rect 30730 6684 30788 6734
rect 29526 6626 30788 6684
rect 30866 7152 32128 7210
rect 30866 7102 30924 7152
rect 30866 6734 30878 7102
rect 30912 6734 30924 7102
rect 32070 7102 32128 7152
rect 30866 6684 30924 6734
rect 32070 6734 32082 7102
rect 32116 6734 32128 7102
rect 32070 6684 32128 6734
rect 30866 6626 32128 6684
rect 28900 6544 28958 6594
rect 27766 6532 28958 6544
rect 27766 6498 27874 6532
rect 28850 6498 28958 6532
rect 27766 6486 28958 6498
rect 27766 6392 28958 6404
rect 27766 6358 27874 6392
rect 28850 6358 28958 6392
rect 27766 6346 28958 6358
rect 27766 6296 27824 6346
rect 27766 5554 27778 6296
rect 27812 5554 27824 6296
rect 28900 6296 28958 6346
rect 27766 5504 27824 5554
rect 28900 5554 28912 6296
rect 28946 5554 28958 6296
rect 28900 5504 28958 5554
rect 27766 5492 28958 5504
rect 27766 5458 27874 5492
rect 28850 5458 28958 5492
rect 27766 5446 28958 5458
rect 27766 5376 28950 5388
rect 27766 5342 27874 5376
rect 28842 5342 28950 5376
rect 27766 5330 28950 5342
rect 27766 5280 27824 5330
rect 27766 4234 27778 5280
rect 27812 4234 27824 5280
rect 28892 5280 28950 5330
rect 27766 4184 27824 4234
rect 28892 4234 28904 5280
rect 28938 4234 28950 5280
rect 28892 4184 28950 4234
rect 27766 4172 28950 4184
rect 27766 4138 27874 4172
rect 28842 4138 28950 4172
rect 27766 4126 28950 4138
rect -174 -8036 1324 -8024
rect -174 -8070 -66 -8036
rect 1216 -8070 1324 -8036
rect -174 -8082 1324 -8070
rect -174 -8132 -116 -8082
rect -174 -8500 -162 -8132
rect -128 -8500 -116 -8132
rect 1266 -8132 1324 -8082
rect -174 -8550 -116 -8500
rect 1266 -8500 1278 -8132
rect 1312 -8500 1324 -8132
rect 1266 -8550 1324 -8500
rect -174 -8562 1324 -8550
rect -174 -8596 -66 -8562
rect 1216 -8596 1324 -8562
rect -174 -8608 1324 -8596
rect -174 -8658 -116 -8608
rect -174 -9626 -162 -8658
rect -128 -9626 -116 -8658
rect 1266 -8658 1324 -8608
rect -174 -9676 -116 -9626
rect 1266 -9626 1278 -8658
rect 1312 -9626 1324 -8658
rect 1266 -9676 1324 -9626
rect -174 -9688 1324 -9676
rect -174 -9722 -66 -9688
rect 1216 -9722 1324 -9688
rect -174 -9734 1324 -9722
rect 1426 -8036 2924 -8024
rect 1426 -8070 1534 -8036
rect 2816 -8070 2924 -8036
rect 1426 -8082 2924 -8070
rect 1426 -8132 1484 -8082
rect 1426 -8500 1438 -8132
rect 1472 -8500 1484 -8132
rect 2866 -8132 2924 -8082
rect 1426 -8550 1484 -8500
rect 2866 -8500 2878 -8132
rect 2912 -8500 2924 -8132
rect 2866 -8550 2924 -8500
rect 1426 -8562 2924 -8550
rect 1426 -8596 1534 -8562
rect 2816 -8596 2924 -8562
rect 1426 -8608 2924 -8596
rect 1426 -8658 1484 -8608
rect 1426 -9626 1438 -8658
rect 1472 -9626 1484 -8658
rect 2866 -8658 2924 -8608
rect 1426 -9676 1484 -9626
rect 2866 -9626 2878 -8658
rect 2912 -9626 2924 -8658
rect 2866 -9676 2924 -9626
rect 1426 -9688 2924 -9676
rect 1426 -9722 1534 -9688
rect 2816 -9722 2924 -9688
rect 1426 -9734 2924 -9722
rect 3026 -8036 4524 -8024
rect 3026 -8070 3134 -8036
rect 4416 -8070 4524 -8036
rect 3026 -8082 4524 -8070
rect 3026 -8132 3084 -8082
rect 3026 -8500 3038 -8132
rect 3072 -8500 3084 -8132
rect 4466 -8132 4524 -8082
rect 3026 -8550 3084 -8500
rect 4466 -8500 4478 -8132
rect 4512 -8500 4524 -8132
rect 4466 -8550 4524 -8500
rect 3026 -8562 4524 -8550
rect 3026 -8596 3134 -8562
rect 4416 -8596 4524 -8562
rect 3026 -8608 4524 -8596
rect 3026 -8658 3084 -8608
rect 3026 -9626 3038 -8658
rect 3072 -9626 3084 -8658
rect 4466 -8658 4524 -8608
rect 3026 -9676 3084 -9626
rect 4466 -9626 4478 -8658
rect 4512 -9626 4524 -8658
rect 4466 -9676 4524 -9626
rect 3026 -9688 4524 -9676
rect 3026 -9722 3134 -9688
rect 4416 -9722 4524 -9688
rect 3026 -9734 4524 -9722
rect 4626 -8036 6124 -8024
rect 4626 -8070 4734 -8036
rect 6016 -8070 6124 -8036
rect 4626 -8082 6124 -8070
rect 4626 -8132 4684 -8082
rect 4626 -8500 4638 -8132
rect 4672 -8500 4684 -8132
rect 6066 -8132 6124 -8082
rect 4626 -8550 4684 -8500
rect 6066 -8500 6078 -8132
rect 6112 -8500 6124 -8132
rect 6066 -8550 6124 -8500
rect 4626 -8562 6124 -8550
rect 4626 -8596 4734 -8562
rect 6016 -8596 6124 -8562
rect 4626 -8608 6124 -8596
rect 4626 -8658 4684 -8608
rect 4626 -9626 4638 -8658
rect 4672 -9626 4684 -8658
rect 6066 -8658 6124 -8608
rect 4626 -9676 4684 -9626
rect 6066 -9626 6078 -8658
rect 6112 -9626 6124 -8658
rect 6066 -9676 6124 -9626
rect 4626 -9688 6124 -9676
rect 4626 -9722 4734 -9688
rect 6016 -9722 6124 -9688
rect 4626 -9734 6124 -9722
rect 6226 -8036 7724 -8024
rect 6226 -8070 6334 -8036
rect 7616 -8070 7724 -8036
rect 6226 -8082 7724 -8070
rect 6226 -8132 6284 -8082
rect 6226 -8500 6238 -8132
rect 6272 -8500 6284 -8132
rect 7666 -8132 7724 -8082
rect 6226 -8550 6284 -8500
rect 7666 -8500 7678 -8132
rect 7712 -8500 7724 -8132
rect 7666 -8550 7724 -8500
rect 6226 -8562 7724 -8550
rect 6226 -8596 6334 -8562
rect 7616 -8596 7724 -8562
rect 6226 -8608 7724 -8596
rect 6226 -8658 6284 -8608
rect 6226 -9626 6238 -8658
rect 6272 -9626 6284 -8658
rect 7666 -8658 7724 -8608
rect 6226 -9676 6284 -9626
rect 7666 -9626 7678 -8658
rect 7712 -9626 7724 -8658
rect 7666 -9676 7724 -9626
rect 6226 -9688 7724 -9676
rect 6226 -9722 6334 -9688
rect 7616 -9722 7724 -9688
rect 6226 -9734 7724 -9722
rect 7826 -8036 9324 -8024
rect 7826 -8070 7934 -8036
rect 9216 -8070 9324 -8036
rect 7826 -8082 9324 -8070
rect 7826 -8132 7884 -8082
rect 7826 -8500 7838 -8132
rect 7872 -8500 7884 -8132
rect 9266 -8132 9324 -8082
rect 7826 -8550 7884 -8500
rect 9266 -8500 9278 -8132
rect 9312 -8500 9324 -8132
rect 9266 -8550 9324 -8500
rect 7826 -8562 9324 -8550
rect 7826 -8596 7934 -8562
rect 9216 -8596 9324 -8562
rect 7826 -8608 9324 -8596
rect 7826 -8658 7884 -8608
rect 7826 -9626 7838 -8658
rect 7872 -9626 7884 -8658
rect 9266 -8658 9324 -8608
rect 7826 -9676 7884 -9626
rect 9266 -9626 9278 -8658
rect 9312 -9626 9324 -8658
rect 9266 -9676 9324 -9626
rect 7826 -9688 9324 -9676
rect 7826 -9722 7934 -9688
rect 9216 -9722 9324 -9688
rect 7826 -9734 9324 -9722
rect 9426 -8036 10924 -8024
rect 9426 -8070 9534 -8036
rect 10816 -8070 10924 -8036
rect 9426 -8082 10924 -8070
rect 9426 -8132 9484 -8082
rect 9426 -8500 9438 -8132
rect 9472 -8500 9484 -8132
rect 10866 -8132 10924 -8082
rect 9426 -8550 9484 -8500
rect 10866 -8500 10878 -8132
rect 10912 -8500 10924 -8132
rect 10866 -8550 10924 -8500
rect 9426 -8562 10924 -8550
rect 9426 -8596 9534 -8562
rect 10816 -8596 10924 -8562
rect 9426 -8608 10924 -8596
rect 9426 -8658 9484 -8608
rect 9426 -9626 9438 -8658
rect 9472 -9626 9484 -8658
rect 10866 -8658 10924 -8608
rect 9426 -9676 9484 -9626
rect 10866 -9626 10878 -8658
rect 10912 -9626 10924 -8658
rect 10866 -9676 10924 -9626
rect 9426 -9688 10924 -9676
rect 9426 -9722 9534 -9688
rect 10816 -9722 10924 -9688
rect 9426 -9734 10924 -9722
rect 11026 -8036 12524 -8024
rect 11026 -8070 11134 -8036
rect 12416 -8070 12524 -8036
rect 11026 -8082 12524 -8070
rect 11026 -8132 11084 -8082
rect 11026 -8500 11038 -8132
rect 11072 -8500 11084 -8132
rect 12466 -8132 12524 -8082
rect 11026 -8550 11084 -8500
rect 12466 -8500 12478 -8132
rect 12512 -8500 12524 -8132
rect 12466 -8550 12524 -8500
rect 11026 -8562 12524 -8550
rect 11026 -8596 11134 -8562
rect 12416 -8596 12524 -8562
rect 11026 -8608 12524 -8596
rect 11026 -8658 11084 -8608
rect 11026 -9626 11038 -8658
rect 11072 -9626 11084 -8658
rect 12466 -8658 12524 -8608
rect 11026 -9676 11084 -9626
rect 12466 -9626 12478 -8658
rect 12512 -9626 12524 -8658
rect 12466 -9676 12524 -9626
rect 11026 -9688 12524 -9676
rect 11026 -9722 11134 -9688
rect 12416 -9722 12524 -9688
rect 11026 -9734 12524 -9722
rect 12626 -8036 14124 -8024
rect 12626 -8070 12734 -8036
rect 14016 -8070 14124 -8036
rect 12626 -8082 14124 -8070
rect 12626 -8132 12684 -8082
rect 12626 -8500 12638 -8132
rect 12672 -8500 12684 -8132
rect 14066 -8132 14124 -8082
rect 12626 -8550 12684 -8500
rect 14066 -8500 14078 -8132
rect 14112 -8500 14124 -8132
rect 14066 -8550 14124 -8500
rect 12626 -8562 14124 -8550
rect 12626 -8596 12734 -8562
rect 14016 -8596 14124 -8562
rect 12626 -8608 14124 -8596
rect 12626 -8658 12684 -8608
rect 12626 -9626 12638 -8658
rect 12672 -9626 12684 -8658
rect 14066 -8658 14124 -8608
rect 12626 -9676 12684 -9626
rect 14066 -9626 14078 -8658
rect 14112 -9626 14124 -8658
rect 14066 -9676 14124 -9626
rect 12626 -9688 14124 -9676
rect 12626 -9722 12734 -9688
rect 14016 -9722 14124 -9688
rect 12626 -9734 14124 -9722
rect 14226 -8036 15724 -8024
rect 14226 -8070 14334 -8036
rect 15616 -8070 15724 -8036
rect 14226 -8082 15724 -8070
rect 14226 -8132 14284 -8082
rect 14226 -8500 14238 -8132
rect 14272 -8500 14284 -8132
rect 15666 -8132 15724 -8082
rect 14226 -8550 14284 -8500
rect 15666 -8500 15678 -8132
rect 15712 -8500 15724 -8132
rect 15666 -8550 15724 -8500
rect 14226 -8562 15724 -8550
rect 14226 -8596 14334 -8562
rect 15616 -8596 15724 -8562
rect 14226 -8608 15724 -8596
rect 14226 -8658 14284 -8608
rect 14226 -9626 14238 -8658
rect 14272 -9626 14284 -8658
rect 15666 -8658 15724 -8608
rect 14226 -9676 14284 -9626
rect 15666 -9626 15678 -8658
rect 15712 -9626 15724 -8658
rect 15666 -9676 15724 -9626
rect 14226 -9688 15724 -9676
rect 14226 -9722 14334 -9688
rect 15616 -9722 15724 -9688
rect 14226 -9734 15724 -9722
rect 15826 -8036 17324 -8024
rect 15826 -8070 15934 -8036
rect 17216 -8070 17324 -8036
rect 15826 -8082 17324 -8070
rect 15826 -8132 15884 -8082
rect 15826 -8500 15838 -8132
rect 15872 -8500 15884 -8132
rect 17266 -8132 17324 -8082
rect 15826 -8550 15884 -8500
rect 17266 -8500 17278 -8132
rect 17312 -8500 17324 -8132
rect 17266 -8550 17324 -8500
rect 15826 -8562 17324 -8550
rect 15826 -8596 15934 -8562
rect 17216 -8596 17324 -8562
rect 15826 -8608 17324 -8596
rect 15826 -8658 15884 -8608
rect 15826 -9626 15838 -8658
rect 15872 -9626 15884 -8658
rect 17266 -8658 17324 -8608
rect 15826 -9676 15884 -9626
rect 17266 -9626 17278 -8658
rect 17312 -9626 17324 -8658
rect 17266 -9676 17324 -9626
rect 15826 -9688 17324 -9676
rect 15826 -9722 15934 -9688
rect 17216 -9722 17324 -9688
rect 15826 -9734 17324 -9722
rect 17426 -8036 18924 -8024
rect 17426 -8070 17534 -8036
rect 18816 -8070 18924 -8036
rect 17426 -8082 18924 -8070
rect 17426 -8132 17484 -8082
rect 17426 -8500 17438 -8132
rect 17472 -8500 17484 -8132
rect 18866 -8132 18924 -8082
rect 17426 -8550 17484 -8500
rect 18866 -8500 18878 -8132
rect 18912 -8500 18924 -8132
rect 18866 -8550 18924 -8500
rect 17426 -8562 18924 -8550
rect 17426 -8596 17534 -8562
rect 18816 -8596 18924 -8562
rect 17426 -8608 18924 -8596
rect 17426 -8658 17484 -8608
rect 17426 -9626 17438 -8658
rect 17472 -9626 17484 -8658
rect 18866 -8658 18924 -8608
rect 17426 -9676 17484 -9626
rect 18866 -9626 18878 -8658
rect 18912 -9626 18924 -8658
rect 18866 -9676 18924 -9626
rect 17426 -9688 18924 -9676
rect 17426 -9722 17534 -9688
rect 18816 -9722 18924 -9688
rect 17426 -9734 18924 -9722
rect 19026 -8036 20524 -8024
rect 19026 -8070 19134 -8036
rect 20416 -8070 20524 -8036
rect 19026 -8082 20524 -8070
rect 19026 -8132 19084 -8082
rect 19026 -8500 19038 -8132
rect 19072 -8500 19084 -8132
rect 20466 -8132 20524 -8082
rect 19026 -8550 19084 -8500
rect 20466 -8500 20478 -8132
rect 20512 -8500 20524 -8132
rect 20466 -8550 20524 -8500
rect 19026 -8562 20524 -8550
rect 19026 -8596 19134 -8562
rect 20416 -8596 20524 -8562
rect 19026 -8608 20524 -8596
rect 19026 -8658 19084 -8608
rect 19026 -9626 19038 -8658
rect 19072 -9626 19084 -8658
rect 20466 -8658 20524 -8608
rect 19026 -9676 19084 -9626
rect 20466 -9626 20478 -8658
rect 20512 -9626 20524 -8658
rect 20466 -9676 20524 -9626
rect 19026 -9688 20524 -9676
rect 19026 -9722 19134 -9688
rect 20416 -9722 20524 -9688
rect 19026 -9734 20524 -9722
rect 20626 -8036 22124 -8024
rect 20626 -8070 20734 -8036
rect 22016 -8070 22124 -8036
rect 20626 -8082 22124 -8070
rect 20626 -8132 20684 -8082
rect 20626 -8500 20638 -8132
rect 20672 -8500 20684 -8132
rect 22066 -8132 22124 -8082
rect 20626 -8550 20684 -8500
rect 22066 -8500 22078 -8132
rect 22112 -8500 22124 -8132
rect 22066 -8550 22124 -8500
rect 20626 -8562 22124 -8550
rect 20626 -8596 20734 -8562
rect 22016 -8596 22124 -8562
rect 20626 -8608 22124 -8596
rect 20626 -8658 20684 -8608
rect 20626 -9626 20638 -8658
rect 20672 -9626 20684 -8658
rect 22066 -8658 22124 -8608
rect 20626 -9676 20684 -9626
rect 22066 -9626 22078 -8658
rect 22112 -9626 22124 -8658
rect 22066 -9676 22124 -9626
rect 20626 -9688 22124 -9676
rect 20626 -9722 20734 -9688
rect 22016 -9722 22124 -9688
rect 20626 -9734 22124 -9722
rect 22226 -8036 23724 -8024
rect 22226 -8070 22334 -8036
rect 23616 -8070 23724 -8036
rect 22226 -8082 23724 -8070
rect 22226 -8132 22284 -8082
rect 22226 -8500 22238 -8132
rect 22272 -8500 22284 -8132
rect 23666 -8132 23724 -8082
rect 22226 -8550 22284 -8500
rect 23666 -8500 23678 -8132
rect 23712 -8500 23724 -8132
rect 23666 -8550 23724 -8500
rect 22226 -8562 23724 -8550
rect 22226 -8596 22334 -8562
rect 23616 -8596 23724 -8562
rect 22226 -8608 23724 -8596
rect 22226 -8658 22284 -8608
rect 22226 -9626 22238 -8658
rect 22272 -9626 22284 -8658
rect 23666 -8658 23724 -8608
rect 22226 -9676 22284 -9626
rect 23666 -9626 23678 -8658
rect 23712 -9626 23724 -8658
rect 23666 -9676 23724 -9626
rect 22226 -9688 23724 -9676
rect 22226 -9722 22334 -9688
rect 23616 -9722 23724 -9688
rect 22226 -9734 23724 -9722
rect 23826 -8036 25324 -8024
rect 23826 -8070 23934 -8036
rect 25216 -8070 25324 -8036
rect 23826 -8082 25324 -8070
rect 23826 -8132 23884 -8082
rect 23826 -8500 23838 -8132
rect 23872 -8500 23884 -8132
rect 25266 -8132 25324 -8082
rect 23826 -8550 23884 -8500
rect 25266 -8500 25278 -8132
rect 25312 -8500 25324 -8132
rect 25266 -8550 25324 -8500
rect 23826 -8562 25324 -8550
rect 23826 -8596 23934 -8562
rect 25216 -8596 25324 -8562
rect 23826 -8608 25324 -8596
rect 23826 -8658 23884 -8608
rect 23826 -9626 23838 -8658
rect 23872 -9626 23884 -8658
rect 25266 -8658 25324 -8608
rect 23826 -9676 23884 -9626
rect 25266 -9626 25278 -8658
rect 25312 -9626 25324 -8658
rect 25266 -9676 25324 -9626
rect 23826 -9688 25324 -9676
rect 23826 -9722 23934 -9688
rect 25216 -9722 25324 -9688
rect 23826 -9734 25324 -9722
rect 25426 -8036 26924 -8024
rect 25426 -8070 25534 -8036
rect 26816 -8070 26924 -8036
rect 25426 -8082 26924 -8070
rect 25426 -8132 25484 -8082
rect 25426 -8500 25438 -8132
rect 25472 -8500 25484 -8132
rect 26866 -8132 26924 -8082
rect 25426 -8550 25484 -8500
rect 26866 -8500 26878 -8132
rect 26912 -8500 26924 -8132
rect 26866 -8550 26924 -8500
rect 25426 -8562 26924 -8550
rect 25426 -8596 25534 -8562
rect 26816 -8596 26924 -8562
rect 25426 -8608 26924 -8596
rect 25426 -8658 25484 -8608
rect 25426 -9626 25438 -8658
rect 25472 -9626 25484 -8658
rect 26866 -8658 26924 -8608
rect 25426 -9676 25484 -9626
rect 26866 -9626 26878 -8658
rect 26912 -9626 26924 -8658
rect 26866 -9676 26924 -9626
rect 25426 -9688 26924 -9676
rect 25426 -9722 25534 -9688
rect 26816 -9722 26924 -9688
rect 25426 -9734 26924 -9722
rect 27026 -8036 28524 -8024
rect 27026 -8070 27134 -8036
rect 28416 -8070 28524 -8036
rect 27026 -8082 28524 -8070
rect 27026 -8132 27084 -8082
rect 27026 -8500 27038 -8132
rect 27072 -8500 27084 -8132
rect 28466 -8132 28524 -8082
rect 27026 -8550 27084 -8500
rect 28466 -8500 28478 -8132
rect 28512 -8500 28524 -8132
rect 28466 -8550 28524 -8500
rect 27026 -8562 28524 -8550
rect 27026 -8596 27134 -8562
rect 28416 -8596 28524 -8562
rect 27026 -8608 28524 -8596
rect 27026 -8658 27084 -8608
rect 27026 -9626 27038 -8658
rect 27072 -9626 27084 -8658
rect 28466 -8658 28524 -8608
rect 27026 -9676 27084 -9626
rect 28466 -9626 28478 -8658
rect 28512 -9626 28524 -8658
rect 28466 -9676 28524 -9626
rect 27026 -9688 28524 -9676
rect 27026 -9722 27134 -9688
rect 28416 -9722 28524 -9688
rect 27026 -9734 28524 -9722
rect 28626 -8036 30124 -8024
rect 28626 -8070 28734 -8036
rect 30016 -8070 30124 -8036
rect 28626 -8082 30124 -8070
rect 28626 -8132 28684 -8082
rect 28626 -8500 28638 -8132
rect 28672 -8500 28684 -8132
rect 30066 -8132 30124 -8082
rect 28626 -8550 28684 -8500
rect 30066 -8500 30078 -8132
rect 30112 -8500 30124 -8132
rect 30066 -8550 30124 -8500
rect 28626 -8562 30124 -8550
rect 28626 -8596 28734 -8562
rect 30016 -8596 30124 -8562
rect 28626 -8608 30124 -8596
rect 28626 -8658 28684 -8608
rect 28626 -9626 28638 -8658
rect 28672 -9626 28684 -8658
rect 30066 -8658 30124 -8608
rect 28626 -9676 28684 -9626
rect 30066 -9626 30078 -8658
rect 30112 -9626 30124 -8658
rect 30066 -9676 30124 -9626
rect 28626 -9688 30124 -9676
rect 28626 -9722 28734 -9688
rect 30016 -9722 30124 -9688
rect 28626 -9734 30124 -9722
rect 30226 -8036 31724 -8024
rect 30226 -8070 30334 -8036
rect 31616 -8070 31724 -8036
rect 30226 -8082 31724 -8070
rect 30226 -8132 30284 -8082
rect 30226 -8500 30238 -8132
rect 30272 -8500 30284 -8132
rect 31666 -8132 31724 -8082
rect 30226 -8550 30284 -8500
rect 31666 -8500 31678 -8132
rect 31712 -8500 31724 -8132
rect 31666 -8550 31724 -8500
rect 30226 -8562 31724 -8550
rect 30226 -8596 30334 -8562
rect 31616 -8596 31724 -8562
rect 30226 -8608 31724 -8596
rect 30226 -8658 30284 -8608
rect 30226 -9626 30238 -8658
rect 30272 -9626 30284 -8658
rect 31666 -8658 31724 -8608
rect 30226 -9676 30284 -9626
rect 31666 -9626 31678 -8658
rect 31712 -9626 31724 -8658
rect 31666 -9676 31724 -9626
rect 30226 -9688 31724 -9676
rect 30226 -9722 30334 -9688
rect 31616 -9722 31724 -9688
rect 30226 -9734 31724 -9722
rect 31826 -8036 33324 -8024
rect 31826 -8070 31934 -8036
rect 33216 -8070 33324 -8036
rect 31826 -8082 33324 -8070
rect 31826 -8132 31884 -8082
rect 31826 -8500 31838 -8132
rect 31872 -8500 31884 -8132
rect 33266 -8132 33324 -8082
rect 31826 -8550 31884 -8500
rect 33266 -8500 33278 -8132
rect 33312 -8500 33324 -8132
rect 33266 -8550 33324 -8500
rect 31826 -8562 33324 -8550
rect 31826 -8596 31934 -8562
rect 33216 -8596 33324 -8562
rect 31826 -8608 33324 -8596
rect 31826 -8658 31884 -8608
rect 31826 -9626 31838 -8658
rect 31872 -9626 31884 -8658
rect 33266 -8658 33324 -8608
rect 31826 -9676 31884 -9626
rect 33266 -9626 33278 -8658
rect 33312 -9626 33324 -8658
rect 33266 -9676 33324 -9626
rect 31826 -9688 33324 -9676
rect 31826 -9722 31934 -9688
rect 33216 -9722 33324 -9688
rect 31826 -9734 33324 -9722
rect 33426 -8036 34924 -8024
rect 33426 -8070 33534 -8036
rect 34816 -8070 34924 -8036
rect 33426 -8082 34924 -8070
rect 33426 -8132 33484 -8082
rect 33426 -8500 33438 -8132
rect 33472 -8500 33484 -8132
rect 34866 -8132 34924 -8082
rect 33426 -8550 33484 -8500
rect 34866 -8500 34878 -8132
rect 34912 -8500 34924 -8132
rect 34866 -8550 34924 -8500
rect 33426 -8562 34924 -8550
rect 33426 -8596 33534 -8562
rect 34816 -8596 34924 -8562
rect 33426 -8608 34924 -8596
rect 33426 -8658 33484 -8608
rect 33426 -9626 33438 -8658
rect 33472 -9626 33484 -8658
rect 34866 -8658 34924 -8608
rect 33426 -9676 33484 -9626
rect 34866 -9626 34878 -8658
rect 34912 -9626 34924 -8658
rect 34866 -9676 34924 -9626
rect 33426 -9688 34924 -9676
rect 33426 -9722 33534 -9688
rect 34816 -9722 34924 -9688
rect 33426 -9734 34924 -9722
rect 35026 -8036 36524 -8024
rect 35026 -8070 35134 -8036
rect 36416 -8070 36524 -8036
rect 35026 -8082 36524 -8070
rect 35026 -8132 35084 -8082
rect 35026 -8500 35038 -8132
rect 35072 -8500 35084 -8132
rect 36466 -8132 36524 -8082
rect 35026 -8550 35084 -8500
rect 36466 -8500 36478 -8132
rect 36512 -8500 36524 -8132
rect 36466 -8550 36524 -8500
rect 35026 -8562 36524 -8550
rect 35026 -8596 35134 -8562
rect 36416 -8596 36524 -8562
rect 35026 -8608 36524 -8596
rect 35026 -8658 35084 -8608
rect 35026 -9626 35038 -8658
rect 35072 -9626 35084 -8658
rect 36466 -8658 36524 -8608
rect 35026 -9676 35084 -9626
rect 36466 -9626 36478 -8658
rect 36512 -9626 36524 -8658
rect 36466 -9676 36524 -9626
rect 35026 -9688 36524 -9676
rect 35026 -9722 35134 -9688
rect 36416 -9722 36524 -9688
rect 35026 -9734 36524 -9722
rect 36626 -8036 38124 -8024
rect 36626 -8070 36734 -8036
rect 38016 -8070 38124 -8036
rect 36626 -8082 38124 -8070
rect 36626 -8132 36684 -8082
rect 36626 -8500 36638 -8132
rect 36672 -8500 36684 -8132
rect 38066 -8132 38124 -8082
rect 36626 -8550 36684 -8500
rect 38066 -8500 38078 -8132
rect 38112 -8500 38124 -8132
rect 38066 -8550 38124 -8500
rect 36626 -8562 38124 -8550
rect 36626 -8596 36734 -8562
rect 38016 -8596 38124 -8562
rect 36626 -8608 38124 -8596
rect 36626 -8658 36684 -8608
rect 36626 -9626 36638 -8658
rect 36672 -9626 36684 -8658
rect 38066 -8658 38124 -8608
rect 36626 -9676 36684 -9626
rect 38066 -9626 38078 -8658
rect 38112 -9626 38124 -8658
rect 38066 -9676 38124 -9626
rect 36626 -9688 38124 -9676
rect 36626 -9722 36734 -9688
rect 38016 -9722 38124 -9688
rect 36626 -9734 38124 -9722
rect -174 -9836 1324 -9824
rect -174 -9870 -66 -9836
rect 1216 -9870 1324 -9836
rect -174 -9882 1324 -9870
rect -174 -9932 -116 -9882
rect -174 -10300 -162 -9932
rect -128 -10300 -116 -9932
rect 1266 -9932 1324 -9882
rect -174 -10350 -116 -10300
rect 1266 -10300 1278 -9932
rect 1312 -10300 1324 -9932
rect 1266 -10350 1324 -10300
rect -174 -10362 1324 -10350
rect -174 -10396 -66 -10362
rect 1216 -10396 1324 -10362
rect -174 -10408 1324 -10396
rect -174 -10458 -116 -10408
rect -174 -11426 -162 -10458
rect -128 -11426 -116 -10458
rect 1266 -10458 1324 -10408
rect -174 -11476 -116 -11426
rect 1266 -11426 1278 -10458
rect 1312 -11426 1324 -10458
rect 1266 -11476 1324 -11426
rect -174 -11488 1324 -11476
rect -174 -11522 -66 -11488
rect 1216 -11522 1324 -11488
rect -174 -11534 1324 -11522
rect 1426 -9836 2924 -9824
rect 1426 -9870 1534 -9836
rect 2816 -9870 2924 -9836
rect 1426 -9882 2924 -9870
rect 1426 -9932 1484 -9882
rect 1426 -10300 1438 -9932
rect 1472 -10300 1484 -9932
rect 2866 -9932 2924 -9882
rect 1426 -10350 1484 -10300
rect 2866 -10300 2878 -9932
rect 2912 -10300 2924 -9932
rect 2866 -10350 2924 -10300
rect 1426 -10362 2924 -10350
rect 1426 -10396 1534 -10362
rect 2816 -10396 2924 -10362
rect 1426 -10408 2924 -10396
rect 1426 -10458 1484 -10408
rect 1426 -11426 1438 -10458
rect 1472 -11426 1484 -10458
rect 2866 -10458 2924 -10408
rect 1426 -11476 1484 -11426
rect 2866 -11426 2878 -10458
rect 2912 -11426 2924 -10458
rect 2866 -11476 2924 -11426
rect 1426 -11488 2924 -11476
rect 1426 -11522 1534 -11488
rect 2816 -11522 2924 -11488
rect 1426 -11534 2924 -11522
rect 3026 -9836 4524 -9824
rect 3026 -9870 3134 -9836
rect 4416 -9870 4524 -9836
rect 3026 -9882 4524 -9870
rect 3026 -9932 3084 -9882
rect 3026 -10300 3038 -9932
rect 3072 -10300 3084 -9932
rect 4466 -9932 4524 -9882
rect 3026 -10350 3084 -10300
rect 4466 -10300 4478 -9932
rect 4512 -10300 4524 -9932
rect 4466 -10350 4524 -10300
rect 3026 -10362 4524 -10350
rect 3026 -10396 3134 -10362
rect 4416 -10396 4524 -10362
rect 3026 -10408 4524 -10396
rect 3026 -10458 3084 -10408
rect 3026 -11426 3038 -10458
rect 3072 -11426 3084 -10458
rect 4466 -10458 4524 -10408
rect 3026 -11476 3084 -11426
rect 4466 -11426 4478 -10458
rect 4512 -11426 4524 -10458
rect 4466 -11476 4524 -11426
rect 3026 -11488 4524 -11476
rect 3026 -11522 3134 -11488
rect 4416 -11522 4524 -11488
rect 3026 -11534 4524 -11522
rect 4626 -9836 6124 -9824
rect 4626 -9870 4734 -9836
rect 6016 -9870 6124 -9836
rect 4626 -9882 6124 -9870
rect 4626 -9932 4684 -9882
rect 4626 -10300 4638 -9932
rect 4672 -10300 4684 -9932
rect 6066 -9932 6124 -9882
rect 4626 -10350 4684 -10300
rect 6066 -10300 6078 -9932
rect 6112 -10300 6124 -9932
rect 6066 -10350 6124 -10300
rect 4626 -10362 6124 -10350
rect 4626 -10396 4734 -10362
rect 6016 -10396 6124 -10362
rect 4626 -10408 6124 -10396
rect 4626 -10458 4684 -10408
rect 4626 -11426 4638 -10458
rect 4672 -11426 4684 -10458
rect 6066 -10458 6124 -10408
rect 4626 -11476 4684 -11426
rect 6066 -11426 6078 -10458
rect 6112 -11426 6124 -10458
rect 6066 -11476 6124 -11426
rect 4626 -11488 6124 -11476
rect 4626 -11522 4734 -11488
rect 6016 -11522 6124 -11488
rect 4626 -11534 6124 -11522
rect 6226 -9836 7724 -9824
rect 6226 -9870 6334 -9836
rect 7616 -9870 7724 -9836
rect 6226 -9882 7724 -9870
rect 6226 -9932 6284 -9882
rect 6226 -10300 6238 -9932
rect 6272 -10300 6284 -9932
rect 7666 -9932 7724 -9882
rect 6226 -10350 6284 -10300
rect 7666 -10300 7678 -9932
rect 7712 -10300 7724 -9932
rect 7666 -10350 7724 -10300
rect 6226 -10362 7724 -10350
rect 6226 -10396 6334 -10362
rect 7616 -10396 7724 -10362
rect 6226 -10408 7724 -10396
rect 6226 -10458 6284 -10408
rect 6226 -11426 6238 -10458
rect 6272 -11426 6284 -10458
rect 7666 -10458 7724 -10408
rect 6226 -11476 6284 -11426
rect 7666 -11426 7678 -10458
rect 7712 -11426 7724 -10458
rect 7666 -11476 7724 -11426
rect 6226 -11488 7724 -11476
rect 6226 -11522 6334 -11488
rect 7616 -11522 7724 -11488
rect 6226 -11534 7724 -11522
rect 7826 -9836 9324 -9824
rect 7826 -9870 7934 -9836
rect 9216 -9870 9324 -9836
rect 7826 -9882 9324 -9870
rect 7826 -9932 7884 -9882
rect 7826 -10300 7838 -9932
rect 7872 -10300 7884 -9932
rect 9266 -9932 9324 -9882
rect 7826 -10350 7884 -10300
rect 9266 -10300 9278 -9932
rect 9312 -10300 9324 -9932
rect 9266 -10350 9324 -10300
rect 7826 -10362 9324 -10350
rect 7826 -10396 7934 -10362
rect 9216 -10396 9324 -10362
rect 7826 -10408 9324 -10396
rect 7826 -10458 7884 -10408
rect 7826 -11426 7838 -10458
rect 7872 -11426 7884 -10458
rect 9266 -10458 9324 -10408
rect 7826 -11476 7884 -11426
rect 9266 -11426 9278 -10458
rect 9312 -11426 9324 -10458
rect 9266 -11476 9324 -11426
rect 7826 -11488 9324 -11476
rect 7826 -11522 7934 -11488
rect 9216 -11522 9324 -11488
rect 7826 -11534 9324 -11522
rect 9426 -9836 10924 -9824
rect 9426 -9870 9534 -9836
rect 10816 -9870 10924 -9836
rect 9426 -9882 10924 -9870
rect 9426 -9932 9484 -9882
rect 9426 -10300 9438 -9932
rect 9472 -10300 9484 -9932
rect 10866 -9932 10924 -9882
rect 9426 -10350 9484 -10300
rect 10866 -10300 10878 -9932
rect 10912 -10300 10924 -9932
rect 10866 -10350 10924 -10300
rect 9426 -10362 10924 -10350
rect 9426 -10396 9534 -10362
rect 10816 -10396 10924 -10362
rect 9426 -10408 10924 -10396
rect 9426 -10458 9484 -10408
rect 9426 -11426 9438 -10458
rect 9472 -11426 9484 -10458
rect 10866 -10458 10924 -10408
rect 9426 -11476 9484 -11426
rect 10866 -11426 10878 -10458
rect 10912 -11426 10924 -10458
rect 10866 -11476 10924 -11426
rect 9426 -11488 10924 -11476
rect 9426 -11522 9534 -11488
rect 10816 -11522 10924 -11488
rect 9426 -11534 10924 -11522
rect 11026 -9836 12524 -9824
rect 11026 -9870 11134 -9836
rect 12416 -9870 12524 -9836
rect 11026 -9882 12524 -9870
rect 11026 -9932 11084 -9882
rect 11026 -10300 11038 -9932
rect 11072 -10300 11084 -9932
rect 12466 -9932 12524 -9882
rect 11026 -10350 11084 -10300
rect 12466 -10300 12478 -9932
rect 12512 -10300 12524 -9932
rect 12466 -10350 12524 -10300
rect 11026 -10362 12524 -10350
rect 11026 -10396 11134 -10362
rect 12416 -10396 12524 -10362
rect 11026 -10408 12524 -10396
rect 11026 -10458 11084 -10408
rect 11026 -11426 11038 -10458
rect 11072 -11426 11084 -10458
rect 12466 -10458 12524 -10408
rect 11026 -11476 11084 -11426
rect 12466 -11426 12478 -10458
rect 12512 -11426 12524 -10458
rect 12466 -11476 12524 -11426
rect 11026 -11488 12524 -11476
rect 11026 -11522 11134 -11488
rect 12416 -11522 12524 -11488
rect 11026 -11534 12524 -11522
rect 12626 -9836 14124 -9824
rect 12626 -9870 12734 -9836
rect 14016 -9870 14124 -9836
rect 12626 -9882 14124 -9870
rect 12626 -9932 12684 -9882
rect 12626 -10300 12638 -9932
rect 12672 -10300 12684 -9932
rect 14066 -9932 14124 -9882
rect 12626 -10350 12684 -10300
rect 14066 -10300 14078 -9932
rect 14112 -10300 14124 -9932
rect 14066 -10350 14124 -10300
rect 12626 -10362 14124 -10350
rect 12626 -10396 12734 -10362
rect 14016 -10396 14124 -10362
rect 12626 -10408 14124 -10396
rect 12626 -10458 12684 -10408
rect 12626 -11426 12638 -10458
rect 12672 -11426 12684 -10458
rect 14066 -10458 14124 -10408
rect 12626 -11476 12684 -11426
rect 14066 -11426 14078 -10458
rect 14112 -11426 14124 -10458
rect 14066 -11476 14124 -11426
rect 12626 -11488 14124 -11476
rect 12626 -11522 12734 -11488
rect 14016 -11522 14124 -11488
rect 12626 -11534 14124 -11522
rect 14226 -9836 15724 -9824
rect 14226 -9870 14334 -9836
rect 15616 -9870 15724 -9836
rect 14226 -9882 15724 -9870
rect 14226 -9932 14284 -9882
rect 14226 -10300 14238 -9932
rect 14272 -10300 14284 -9932
rect 15666 -9932 15724 -9882
rect 14226 -10350 14284 -10300
rect 15666 -10300 15678 -9932
rect 15712 -10300 15724 -9932
rect 15666 -10350 15724 -10300
rect 14226 -10362 15724 -10350
rect 14226 -10396 14334 -10362
rect 15616 -10396 15724 -10362
rect 14226 -10408 15724 -10396
rect 14226 -10458 14284 -10408
rect 14226 -11426 14238 -10458
rect 14272 -11426 14284 -10458
rect 15666 -10458 15724 -10408
rect 14226 -11476 14284 -11426
rect 15666 -11426 15678 -10458
rect 15712 -11426 15724 -10458
rect 15666 -11476 15724 -11426
rect 14226 -11488 15724 -11476
rect 14226 -11522 14334 -11488
rect 15616 -11522 15724 -11488
rect 14226 -11534 15724 -11522
rect 15826 -9836 17324 -9824
rect 15826 -9870 15934 -9836
rect 17216 -9870 17324 -9836
rect 15826 -9882 17324 -9870
rect 15826 -9932 15884 -9882
rect 15826 -10300 15838 -9932
rect 15872 -10300 15884 -9932
rect 17266 -9932 17324 -9882
rect 15826 -10350 15884 -10300
rect 17266 -10300 17278 -9932
rect 17312 -10300 17324 -9932
rect 17266 -10350 17324 -10300
rect 15826 -10362 17324 -10350
rect 15826 -10396 15934 -10362
rect 17216 -10396 17324 -10362
rect 15826 -10408 17324 -10396
rect 15826 -10458 15884 -10408
rect 15826 -11426 15838 -10458
rect 15872 -11426 15884 -10458
rect 17266 -10458 17324 -10408
rect 15826 -11476 15884 -11426
rect 17266 -11426 17278 -10458
rect 17312 -11426 17324 -10458
rect 17266 -11476 17324 -11426
rect 15826 -11488 17324 -11476
rect 15826 -11522 15934 -11488
rect 17216 -11522 17324 -11488
rect 15826 -11534 17324 -11522
rect 17426 -9836 18924 -9824
rect 17426 -9870 17534 -9836
rect 18816 -9870 18924 -9836
rect 17426 -9882 18924 -9870
rect 17426 -9932 17484 -9882
rect 17426 -10300 17438 -9932
rect 17472 -10300 17484 -9932
rect 18866 -9932 18924 -9882
rect 17426 -10350 17484 -10300
rect 18866 -10300 18878 -9932
rect 18912 -10300 18924 -9932
rect 18866 -10350 18924 -10300
rect 17426 -10362 18924 -10350
rect 17426 -10396 17534 -10362
rect 18816 -10396 18924 -10362
rect 17426 -10408 18924 -10396
rect 17426 -10458 17484 -10408
rect 17426 -11426 17438 -10458
rect 17472 -11426 17484 -10458
rect 18866 -10458 18924 -10408
rect 17426 -11476 17484 -11426
rect 18866 -11426 18878 -10458
rect 18912 -11426 18924 -10458
rect 18866 -11476 18924 -11426
rect 17426 -11488 18924 -11476
rect 17426 -11522 17534 -11488
rect 18816 -11522 18924 -11488
rect 17426 -11534 18924 -11522
rect 19026 -9836 20524 -9824
rect 19026 -9870 19134 -9836
rect 20416 -9870 20524 -9836
rect 19026 -9882 20524 -9870
rect 19026 -9932 19084 -9882
rect 19026 -10300 19038 -9932
rect 19072 -10300 19084 -9932
rect 20466 -9932 20524 -9882
rect 19026 -10350 19084 -10300
rect 20466 -10300 20478 -9932
rect 20512 -10300 20524 -9932
rect 20466 -10350 20524 -10300
rect 19026 -10362 20524 -10350
rect 19026 -10396 19134 -10362
rect 20416 -10396 20524 -10362
rect 19026 -10408 20524 -10396
rect 19026 -10458 19084 -10408
rect 19026 -11426 19038 -10458
rect 19072 -11426 19084 -10458
rect 20466 -10458 20524 -10408
rect 19026 -11476 19084 -11426
rect 20466 -11426 20478 -10458
rect 20512 -11426 20524 -10458
rect 20466 -11476 20524 -11426
rect 19026 -11488 20524 -11476
rect 19026 -11522 19134 -11488
rect 20416 -11522 20524 -11488
rect 19026 -11534 20524 -11522
rect 20626 -9836 22124 -9824
rect 20626 -9870 20734 -9836
rect 22016 -9870 22124 -9836
rect 20626 -9882 22124 -9870
rect 20626 -9932 20684 -9882
rect 20626 -10300 20638 -9932
rect 20672 -10300 20684 -9932
rect 22066 -9932 22124 -9882
rect 20626 -10350 20684 -10300
rect 22066 -10300 22078 -9932
rect 22112 -10300 22124 -9932
rect 22066 -10350 22124 -10300
rect 20626 -10362 22124 -10350
rect 20626 -10396 20734 -10362
rect 22016 -10396 22124 -10362
rect 20626 -10408 22124 -10396
rect 20626 -10458 20684 -10408
rect 20626 -11426 20638 -10458
rect 20672 -11426 20684 -10458
rect 22066 -10458 22124 -10408
rect 20626 -11476 20684 -11426
rect 22066 -11426 22078 -10458
rect 22112 -11426 22124 -10458
rect 22066 -11476 22124 -11426
rect 20626 -11488 22124 -11476
rect 20626 -11522 20734 -11488
rect 22016 -11522 22124 -11488
rect 20626 -11534 22124 -11522
rect 22226 -9836 23724 -9824
rect 22226 -9870 22334 -9836
rect 23616 -9870 23724 -9836
rect 22226 -9882 23724 -9870
rect 22226 -9932 22284 -9882
rect 22226 -10300 22238 -9932
rect 22272 -10300 22284 -9932
rect 23666 -9932 23724 -9882
rect 22226 -10350 22284 -10300
rect 23666 -10300 23678 -9932
rect 23712 -10300 23724 -9932
rect 23666 -10350 23724 -10300
rect 22226 -10362 23724 -10350
rect 22226 -10396 22334 -10362
rect 23616 -10396 23724 -10362
rect 22226 -10408 23724 -10396
rect 22226 -10458 22284 -10408
rect 22226 -11426 22238 -10458
rect 22272 -11426 22284 -10458
rect 23666 -10458 23724 -10408
rect 22226 -11476 22284 -11426
rect 23666 -11426 23678 -10458
rect 23712 -11426 23724 -10458
rect 23666 -11476 23724 -11426
rect 22226 -11488 23724 -11476
rect 22226 -11522 22334 -11488
rect 23616 -11522 23724 -11488
rect 22226 -11534 23724 -11522
rect 23826 -9836 25324 -9824
rect 23826 -9870 23934 -9836
rect 25216 -9870 25324 -9836
rect 23826 -9882 25324 -9870
rect 23826 -9932 23884 -9882
rect 23826 -10300 23838 -9932
rect 23872 -10300 23884 -9932
rect 25266 -9932 25324 -9882
rect 23826 -10350 23884 -10300
rect 25266 -10300 25278 -9932
rect 25312 -10300 25324 -9932
rect 25266 -10350 25324 -10300
rect 23826 -10362 25324 -10350
rect 23826 -10396 23934 -10362
rect 25216 -10396 25324 -10362
rect 23826 -10408 25324 -10396
rect 23826 -10458 23884 -10408
rect 23826 -11426 23838 -10458
rect 23872 -11426 23884 -10458
rect 25266 -10458 25324 -10408
rect 23826 -11476 23884 -11426
rect 25266 -11426 25278 -10458
rect 25312 -11426 25324 -10458
rect 25266 -11476 25324 -11426
rect 23826 -11488 25324 -11476
rect 23826 -11522 23934 -11488
rect 25216 -11522 25324 -11488
rect 23826 -11534 25324 -11522
rect 25426 -9836 26924 -9824
rect 25426 -9870 25534 -9836
rect 26816 -9870 26924 -9836
rect 25426 -9882 26924 -9870
rect 25426 -9932 25484 -9882
rect 25426 -10300 25438 -9932
rect 25472 -10300 25484 -9932
rect 26866 -9932 26924 -9882
rect 25426 -10350 25484 -10300
rect 26866 -10300 26878 -9932
rect 26912 -10300 26924 -9932
rect 26866 -10350 26924 -10300
rect 25426 -10362 26924 -10350
rect 25426 -10396 25534 -10362
rect 26816 -10396 26924 -10362
rect 25426 -10408 26924 -10396
rect 25426 -10458 25484 -10408
rect 25426 -11426 25438 -10458
rect 25472 -11426 25484 -10458
rect 26866 -10458 26924 -10408
rect 25426 -11476 25484 -11426
rect 26866 -11426 26878 -10458
rect 26912 -11426 26924 -10458
rect 26866 -11476 26924 -11426
rect 25426 -11488 26924 -11476
rect 25426 -11522 25534 -11488
rect 26816 -11522 26924 -11488
rect 25426 -11534 26924 -11522
rect 27026 -9836 28524 -9824
rect 27026 -9870 27134 -9836
rect 28416 -9870 28524 -9836
rect 27026 -9882 28524 -9870
rect 27026 -9932 27084 -9882
rect 27026 -10300 27038 -9932
rect 27072 -10300 27084 -9932
rect 28466 -9932 28524 -9882
rect 27026 -10350 27084 -10300
rect 28466 -10300 28478 -9932
rect 28512 -10300 28524 -9932
rect 28466 -10350 28524 -10300
rect 27026 -10362 28524 -10350
rect 27026 -10396 27134 -10362
rect 28416 -10396 28524 -10362
rect 27026 -10408 28524 -10396
rect 27026 -10458 27084 -10408
rect 27026 -11426 27038 -10458
rect 27072 -11426 27084 -10458
rect 28466 -10458 28524 -10408
rect 27026 -11476 27084 -11426
rect 28466 -11426 28478 -10458
rect 28512 -11426 28524 -10458
rect 28466 -11476 28524 -11426
rect 27026 -11488 28524 -11476
rect 27026 -11522 27134 -11488
rect 28416 -11522 28524 -11488
rect 27026 -11534 28524 -11522
rect 28626 -9836 30124 -9824
rect 28626 -9870 28734 -9836
rect 30016 -9870 30124 -9836
rect 28626 -9882 30124 -9870
rect 28626 -9932 28684 -9882
rect 28626 -10300 28638 -9932
rect 28672 -10300 28684 -9932
rect 30066 -9932 30124 -9882
rect 28626 -10350 28684 -10300
rect 30066 -10300 30078 -9932
rect 30112 -10300 30124 -9932
rect 30066 -10350 30124 -10300
rect 28626 -10362 30124 -10350
rect 28626 -10396 28734 -10362
rect 30016 -10396 30124 -10362
rect 28626 -10408 30124 -10396
rect 28626 -10458 28684 -10408
rect 28626 -11426 28638 -10458
rect 28672 -11426 28684 -10458
rect 30066 -10458 30124 -10408
rect 28626 -11476 28684 -11426
rect 30066 -11426 30078 -10458
rect 30112 -11426 30124 -10458
rect 30066 -11476 30124 -11426
rect 28626 -11488 30124 -11476
rect 28626 -11522 28734 -11488
rect 30016 -11522 30124 -11488
rect 28626 -11534 30124 -11522
rect 30226 -9836 31724 -9824
rect 30226 -9870 30334 -9836
rect 31616 -9870 31724 -9836
rect 30226 -9882 31724 -9870
rect 30226 -9932 30284 -9882
rect 30226 -10300 30238 -9932
rect 30272 -10300 30284 -9932
rect 31666 -9932 31724 -9882
rect 30226 -10350 30284 -10300
rect 31666 -10300 31678 -9932
rect 31712 -10300 31724 -9932
rect 31666 -10350 31724 -10300
rect 30226 -10362 31724 -10350
rect 30226 -10396 30334 -10362
rect 31616 -10396 31724 -10362
rect 30226 -10408 31724 -10396
rect 30226 -10458 30284 -10408
rect 30226 -11426 30238 -10458
rect 30272 -11426 30284 -10458
rect 31666 -10458 31724 -10408
rect 30226 -11476 30284 -11426
rect 31666 -11426 31678 -10458
rect 31712 -11426 31724 -10458
rect 31666 -11476 31724 -11426
rect 30226 -11488 31724 -11476
rect 30226 -11522 30334 -11488
rect 31616 -11522 31724 -11488
rect 30226 -11534 31724 -11522
rect 31826 -9836 33324 -9824
rect 31826 -9870 31934 -9836
rect 33216 -9870 33324 -9836
rect 31826 -9882 33324 -9870
rect 31826 -9932 31884 -9882
rect 31826 -10300 31838 -9932
rect 31872 -10300 31884 -9932
rect 33266 -9932 33324 -9882
rect 31826 -10350 31884 -10300
rect 33266 -10300 33278 -9932
rect 33312 -10300 33324 -9932
rect 33266 -10350 33324 -10300
rect 31826 -10362 33324 -10350
rect 31826 -10396 31934 -10362
rect 33216 -10396 33324 -10362
rect 31826 -10408 33324 -10396
rect 31826 -10458 31884 -10408
rect 31826 -11426 31838 -10458
rect 31872 -11426 31884 -10458
rect 33266 -10458 33324 -10408
rect 31826 -11476 31884 -11426
rect 33266 -11426 33278 -10458
rect 33312 -11426 33324 -10458
rect 33266 -11476 33324 -11426
rect 31826 -11488 33324 -11476
rect 31826 -11522 31934 -11488
rect 33216 -11522 33324 -11488
rect 31826 -11534 33324 -11522
rect 33426 -9836 34924 -9824
rect 33426 -9870 33534 -9836
rect 34816 -9870 34924 -9836
rect 33426 -9882 34924 -9870
rect 33426 -9932 33484 -9882
rect 33426 -10300 33438 -9932
rect 33472 -10300 33484 -9932
rect 34866 -9932 34924 -9882
rect 33426 -10350 33484 -10300
rect 34866 -10300 34878 -9932
rect 34912 -10300 34924 -9932
rect 34866 -10350 34924 -10300
rect 33426 -10362 34924 -10350
rect 33426 -10396 33534 -10362
rect 34816 -10396 34924 -10362
rect 33426 -10408 34924 -10396
rect 33426 -10458 33484 -10408
rect 33426 -11426 33438 -10458
rect 33472 -11426 33484 -10458
rect 34866 -10458 34924 -10408
rect 33426 -11476 33484 -11426
rect 34866 -11426 34878 -10458
rect 34912 -11426 34924 -10458
rect 34866 -11476 34924 -11426
rect 33426 -11488 34924 -11476
rect 33426 -11522 33534 -11488
rect 34816 -11522 34924 -11488
rect 33426 -11534 34924 -11522
rect 35026 -9836 36524 -9824
rect 35026 -9870 35134 -9836
rect 36416 -9870 36524 -9836
rect 35026 -9882 36524 -9870
rect 35026 -9932 35084 -9882
rect 35026 -10300 35038 -9932
rect 35072 -10300 35084 -9932
rect 36466 -9932 36524 -9882
rect 35026 -10350 35084 -10300
rect 36466 -10300 36478 -9932
rect 36512 -10300 36524 -9932
rect 36466 -10350 36524 -10300
rect 35026 -10362 36524 -10350
rect 35026 -10396 35134 -10362
rect 36416 -10396 36524 -10362
rect 35026 -10408 36524 -10396
rect 35026 -10458 35084 -10408
rect 35026 -11426 35038 -10458
rect 35072 -11426 35084 -10458
rect 36466 -10458 36524 -10408
rect 35026 -11476 35084 -11426
rect 36466 -11426 36478 -10458
rect 36512 -11426 36524 -10458
rect 36466 -11476 36524 -11426
rect 35026 -11488 36524 -11476
rect 35026 -11522 35134 -11488
rect 36416 -11522 36524 -11488
rect 35026 -11534 36524 -11522
rect 36626 -9836 38124 -9824
rect 36626 -9870 36734 -9836
rect 38016 -9870 38124 -9836
rect 36626 -9882 38124 -9870
rect 36626 -9932 36684 -9882
rect 36626 -10300 36638 -9932
rect 36672 -10300 36684 -9932
rect 38066 -9932 38124 -9882
rect 36626 -10350 36684 -10300
rect 38066 -10300 38078 -9932
rect 38112 -10300 38124 -9932
rect 38066 -10350 38124 -10300
rect 36626 -10362 38124 -10350
rect 36626 -10396 36734 -10362
rect 38016 -10396 38124 -10362
rect 36626 -10408 38124 -10396
rect 36626 -10458 36684 -10408
rect 36626 -11426 36638 -10458
rect 36672 -11426 36684 -10458
rect 38066 -10458 38124 -10408
rect 36626 -11476 36684 -11426
rect 38066 -11426 38078 -10458
rect 38112 -11426 38124 -10458
rect 38066 -11476 38124 -11426
rect 36626 -11488 38124 -11476
rect 36626 -11522 36734 -11488
rect 38016 -11522 38124 -11488
rect 36626 -11534 38124 -11522
rect -174 -11636 1324 -11624
rect -174 -11670 -66 -11636
rect 1216 -11670 1324 -11636
rect -174 -11682 1324 -11670
rect -174 -11732 -116 -11682
rect -174 -12100 -162 -11732
rect -128 -12100 -116 -11732
rect 1266 -11732 1324 -11682
rect -174 -12150 -116 -12100
rect 1266 -12100 1278 -11732
rect 1312 -12100 1324 -11732
rect 1266 -12150 1324 -12100
rect -174 -12162 1324 -12150
rect -174 -12196 -66 -12162
rect 1216 -12196 1324 -12162
rect -174 -12208 1324 -12196
rect -174 -12258 -116 -12208
rect -174 -13226 -162 -12258
rect -128 -13226 -116 -12258
rect 1266 -12258 1324 -12208
rect -174 -13276 -116 -13226
rect 1266 -13226 1278 -12258
rect 1312 -13226 1324 -12258
rect 1266 -13276 1324 -13226
rect -174 -13288 1324 -13276
rect -174 -13322 -66 -13288
rect 1216 -13322 1324 -13288
rect -174 -13334 1324 -13322
rect 1426 -11636 2924 -11624
rect 1426 -11670 1534 -11636
rect 2816 -11670 2924 -11636
rect 1426 -11682 2924 -11670
rect 1426 -11732 1484 -11682
rect 1426 -12100 1438 -11732
rect 1472 -12100 1484 -11732
rect 2866 -11732 2924 -11682
rect 1426 -12150 1484 -12100
rect 2866 -12100 2878 -11732
rect 2912 -12100 2924 -11732
rect 2866 -12150 2924 -12100
rect 1426 -12162 2924 -12150
rect 1426 -12196 1534 -12162
rect 2816 -12196 2924 -12162
rect 1426 -12208 2924 -12196
rect 1426 -12258 1484 -12208
rect 1426 -13226 1438 -12258
rect 1472 -13226 1484 -12258
rect 2866 -12258 2924 -12208
rect 1426 -13276 1484 -13226
rect 2866 -13226 2878 -12258
rect 2912 -13226 2924 -12258
rect 2866 -13276 2924 -13226
rect 1426 -13288 2924 -13276
rect 1426 -13322 1534 -13288
rect 2816 -13322 2924 -13288
rect 1426 -13334 2924 -13322
rect 3026 -11636 4524 -11624
rect 3026 -11670 3134 -11636
rect 4416 -11670 4524 -11636
rect 3026 -11682 4524 -11670
rect 3026 -11732 3084 -11682
rect 3026 -12100 3038 -11732
rect 3072 -12100 3084 -11732
rect 4466 -11732 4524 -11682
rect 3026 -12150 3084 -12100
rect 4466 -12100 4478 -11732
rect 4512 -12100 4524 -11732
rect 4466 -12150 4524 -12100
rect 3026 -12162 4524 -12150
rect 3026 -12196 3134 -12162
rect 4416 -12196 4524 -12162
rect 3026 -12208 4524 -12196
rect 3026 -12258 3084 -12208
rect 3026 -13226 3038 -12258
rect 3072 -13226 3084 -12258
rect 4466 -12258 4524 -12208
rect 3026 -13276 3084 -13226
rect 4466 -13226 4478 -12258
rect 4512 -13226 4524 -12258
rect 4466 -13276 4524 -13226
rect 3026 -13288 4524 -13276
rect 3026 -13322 3134 -13288
rect 4416 -13322 4524 -13288
rect 3026 -13334 4524 -13322
rect 4626 -11636 6124 -11624
rect 4626 -11670 4734 -11636
rect 6016 -11670 6124 -11636
rect 4626 -11682 6124 -11670
rect 4626 -11732 4684 -11682
rect 4626 -12100 4638 -11732
rect 4672 -12100 4684 -11732
rect 6066 -11732 6124 -11682
rect 4626 -12150 4684 -12100
rect 6066 -12100 6078 -11732
rect 6112 -12100 6124 -11732
rect 6066 -12150 6124 -12100
rect 4626 -12162 6124 -12150
rect 4626 -12196 4734 -12162
rect 6016 -12196 6124 -12162
rect 4626 -12208 6124 -12196
rect 4626 -12258 4684 -12208
rect 4626 -13226 4638 -12258
rect 4672 -13226 4684 -12258
rect 6066 -12258 6124 -12208
rect 4626 -13276 4684 -13226
rect 6066 -13226 6078 -12258
rect 6112 -13226 6124 -12258
rect 6066 -13276 6124 -13226
rect 4626 -13288 6124 -13276
rect 4626 -13322 4734 -13288
rect 6016 -13322 6124 -13288
rect 4626 -13334 6124 -13322
rect 6226 -11636 7724 -11624
rect 6226 -11670 6334 -11636
rect 7616 -11670 7724 -11636
rect 6226 -11682 7724 -11670
rect 6226 -11732 6284 -11682
rect 6226 -12100 6238 -11732
rect 6272 -12100 6284 -11732
rect 7666 -11732 7724 -11682
rect 6226 -12150 6284 -12100
rect 7666 -12100 7678 -11732
rect 7712 -12100 7724 -11732
rect 7666 -12150 7724 -12100
rect 6226 -12162 7724 -12150
rect 6226 -12196 6334 -12162
rect 7616 -12196 7724 -12162
rect 6226 -12208 7724 -12196
rect 6226 -12258 6284 -12208
rect 6226 -13226 6238 -12258
rect 6272 -13226 6284 -12258
rect 7666 -12258 7724 -12208
rect 6226 -13276 6284 -13226
rect 7666 -13226 7678 -12258
rect 7712 -13226 7724 -12258
rect 7666 -13276 7724 -13226
rect 6226 -13288 7724 -13276
rect 6226 -13322 6334 -13288
rect 7616 -13322 7724 -13288
rect 6226 -13334 7724 -13322
rect 7826 -11636 9324 -11624
rect 7826 -11670 7934 -11636
rect 9216 -11670 9324 -11636
rect 7826 -11682 9324 -11670
rect 7826 -11732 7884 -11682
rect 7826 -12100 7838 -11732
rect 7872 -12100 7884 -11732
rect 9266 -11732 9324 -11682
rect 7826 -12150 7884 -12100
rect 9266 -12100 9278 -11732
rect 9312 -12100 9324 -11732
rect 9266 -12150 9324 -12100
rect 7826 -12162 9324 -12150
rect 7826 -12196 7934 -12162
rect 9216 -12196 9324 -12162
rect 7826 -12208 9324 -12196
rect 7826 -12258 7884 -12208
rect 7826 -13226 7838 -12258
rect 7872 -13226 7884 -12258
rect 9266 -12258 9324 -12208
rect 7826 -13276 7884 -13226
rect 9266 -13226 9278 -12258
rect 9312 -13226 9324 -12258
rect 9266 -13276 9324 -13226
rect 7826 -13288 9324 -13276
rect 7826 -13322 7934 -13288
rect 9216 -13322 9324 -13288
rect 7826 -13334 9324 -13322
rect 9426 -11636 10924 -11624
rect 9426 -11670 9534 -11636
rect 10816 -11670 10924 -11636
rect 9426 -11682 10924 -11670
rect 9426 -11732 9484 -11682
rect 9426 -12100 9438 -11732
rect 9472 -12100 9484 -11732
rect 10866 -11732 10924 -11682
rect 9426 -12150 9484 -12100
rect 10866 -12100 10878 -11732
rect 10912 -12100 10924 -11732
rect 10866 -12150 10924 -12100
rect 9426 -12162 10924 -12150
rect 9426 -12196 9534 -12162
rect 10816 -12196 10924 -12162
rect 9426 -12208 10924 -12196
rect 9426 -12258 9484 -12208
rect 9426 -13226 9438 -12258
rect 9472 -13226 9484 -12258
rect 10866 -12258 10924 -12208
rect 9426 -13276 9484 -13226
rect 10866 -13226 10878 -12258
rect 10912 -13226 10924 -12258
rect 10866 -13276 10924 -13226
rect 9426 -13288 10924 -13276
rect 9426 -13322 9534 -13288
rect 10816 -13322 10924 -13288
rect 9426 -13334 10924 -13322
rect 11026 -11636 12524 -11624
rect 11026 -11670 11134 -11636
rect 12416 -11670 12524 -11636
rect 11026 -11682 12524 -11670
rect 11026 -11732 11084 -11682
rect 11026 -12100 11038 -11732
rect 11072 -12100 11084 -11732
rect 12466 -11732 12524 -11682
rect 11026 -12150 11084 -12100
rect 12466 -12100 12478 -11732
rect 12512 -12100 12524 -11732
rect 12466 -12150 12524 -12100
rect 11026 -12162 12524 -12150
rect 11026 -12196 11134 -12162
rect 12416 -12196 12524 -12162
rect 11026 -12208 12524 -12196
rect 11026 -12258 11084 -12208
rect 11026 -13226 11038 -12258
rect 11072 -13226 11084 -12258
rect 12466 -12258 12524 -12208
rect 11026 -13276 11084 -13226
rect 12466 -13226 12478 -12258
rect 12512 -13226 12524 -12258
rect 12466 -13276 12524 -13226
rect 11026 -13288 12524 -13276
rect 11026 -13322 11134 -13288
rect 12416 -13322 12524 -13288
rect 11026 -13334 12524 -13322
rect 12626 -11636 14124 -11624
rect 12626 -11670 12734 -11636
rect 14016 -11670 14124 -11636
rect 12626 -11682 14124 -11670
rect 12626 -11732 12684 -11682
rect 12626 -12100 12638 -11732
rect 12672 -12100 12684 -11732
rect 14066 -11732 14124 -11682
rect 12626 -12150 12684 -12100
rect 14066 -12100 14078 -11732
rect 14112 -12100 14124 -11732
rect 14066 -12150 14124 -12100
rect 12626 -12162 14124 -12150
rect 12626 -12196 12734 -12162
rect 14016 -12196 14124 -12162
rect 12626 -12208 14124 -12196
rect 12626 -12258 12684 -12208
rect 12626 -13226 12638 -12258
rect 12672 -13226 12684 -12258
rect 14066 -12258 14124 -12208
rect 12626 -13276 12684 -13226
rect 14066 -13226 14078 -12258
rect 14112 -13226 14124 -12258
rect 14066 -13276 14124 -13226
rect 12626 -13288 14124 -13276
rect 12626 -13322 12734 -13288
rect 14016 -13322 14124 -13288
rect 12626 -13334 14124 -13322
rect 14226 -11636 15724 -11624
rect 14226 -11670 14334 -11636
rect 15616 -11670 15724 -11636
rect 14226 -11682 15724 -11670
rect 14226 -11732 14284 -11682
rect 14226 -12100 14238 -11732
rect 14272 -12100 14284 -11732
rect 15666 -11732 15724 -11682
rect 14226 -12150 14284 -12100
rect 15666 -12100 15678 -11732
rect 15712 -12100 15724 -11732
rect 15666 -12150 15724 -12100
rect 14226 -12162 15724 -12150
rect 14226 -12196 14334 -12162
rect 15616 -12196 15724 -12162
rect 14226 -12208 15724 -12196
rect 14226 -12258 14284 -12208
rect 14226 -13226 14238 -12258
rect 14272 -13226 14284 -12258
rect 15666 -12258 15724 -12208
rect 14226 -13276 14284 -13226
rect 15666 -13226 15678 -12258
rect 15712 -13226 15724 -12258
rect 15666 -13276 15724 -13226
rect 14226 -13288 15724 -13276
rect 14226 -13322 14334 -13288
rect 15616 -13322 15724 -13288
rect 14226 -13334 15724 -13322
rect 15826 -11636 17324 -11624
rect 15826 -11670 15934 -11636
rect 17216 -11670 17324 -11636
rect 15826 -11682 17324 -11670
rect 15826 -11732 15884 -11682
rect 15826 -12100 15838 -11732
rect 15872 -12100 15884 -11732
rect 17266 -11732 17324 -11682
rect 15826 -12150 15884 -12100
rect 17266 -12100 17278 -11732
rect 17312 -12100 17324 -11732
rect 17266 -12150 17324 -12100
rect 15826 -12162 17324 -12150
rect 15826 -12196 15934 -12162
rect 17216 -12196 17324 -12162
rect 15826 -12208 17324 -12196
rect 15826 -12258 15884 -12208
rect 15826 -13226 15838 -12258
rect 15872 -13226 15884 -12258
rect 17266 -12258 17324 -12208
rect 15826 -13276 15884 -13226
rect 17266 -13226 17278 -12258
rect 17312 -13226 17324 -12258
rect 17266 -13276 17324 -13226
rect 15826 -13288 17324 -13276
rect 15826 -13322 15934 -13288
rect 17216 -13322 17324 -13288
rect 15826 -13334 17324 -13322
rect 17426 -11636 18924 -11624
rect 17426 -11670 17534 -11636
rect 18816 -11670 18924 -11636
rect 17426 -11682 18924 -11670
rect 17426 -11732 17484 -11682
rect 17426 -12100 17438 -11732
rect 17472 -12100 17484 -11732
rect 18866 -11732 18924 -11682
rect 17426 -12150 17484 -12100
rect 18866 -12100 18878 -11732
rect 18912 -12100 18924 -11732
rect 18866 -12150 18924 -12100
rect 17426 -12162 18924 -12150
rect 17426 -12196 17534 -12162
rect 18816 -12196 18924 -12162
rect 17426 -12208 18924 -12196
rect 17426 -12258 17484 -12208
rect 17426 -13226 17438 -12258
rect 17472 -13226 17484 -12258
rect 18866 -12258 18924 -12208
rect 17426 -13276 17484 -13226
rect 18866 -13226 18878 -12258
rect 18912 -13226 18924 -12258
rect 18866 -13276 18924 -13226
rect 17426 -13288 18924 -13276
rect 17426 -13322 17534 -13288
rect 18816 -13322 18924 -13288
rect 17426 -13334 18924 -13322
rect 19026 -11636 20524 -11624
rect 19026 -11670 19134 -11636
rect 20416 -11670 20524 -11636
rect 19026 -11682 20524 -11670
rect 19026 -11732 19084 -11682
rect 19026 -12100 19038 -11732
rect 19072 -12100 19084 -11732
rect 20466 -11732 20524 -11682
rect 19026 -12150 19084 -12100
rect 20466 -12100 20478 -11732
rect 20512 -12100 20524 -11732
rect 20466 -12150 20524 -12100
rect 19026 -12162 20524 -12150
rect 19026 -12196 19134 -12162
rect 20416 -12196 20524 -12162
rect 19026 -12208 20524 -12196
rect 19026 -12258 19084 -12208
rect 19026 -13226 19038 -12258
rect 19072 -13226 19084 -12258
rect 20466 -12258 20524 -12208
rect 19026 -13276 19084 -13226
rect 20466 -13226 20478 -12258
rect 20512 -13226 20524 -12258
rect 20466 -13276 20524 -13226
rect 19026 -13288 20524 -13276
rect 19026 -13322 19134 -13288
rect 20416 -13322 20524 -13288
rect 19026 -13334 20524 -13322
rect 20626 -11636 22124 -11624
rect 20626 -11670 20734 -11636
rect 22016 -11670 22124 -11636
rect 20626 -11682 22124 -11670
rect 20626 -11732 20684 -11682
rect 20626 -12100 20638 -11732
rect 20672 -12100 20684 -11732
rect 22066 -11732 22124 -11682
rect 20626 -12150 20684 -12100
rect 22066 -12100 22078 -11732
rect 22112 -12100 22124 -11732
rect 22066 -12150 22124 -12100
rect 20626 -12162 22124 -12150
rect 20626 -12196 20734 -12162
rect 22016 -12196 22124 -12162
rect 20626 -12208 22124 -12196
rect 20626 -12258 20684 -12208
rect 20626 -13226 20638 -12258
rect 20672 -13226 20684 -12258
rect 22066 -12258 22124 -12208
rect 20626 -13276 20684 -13226
rect 22066 -13226 22078 -12258
rect 22112 -13226 22124 -12258
rect 22066 -13276 22124 -13226
rect 20626 -13288 22124 -13276
rect 20626 -13322 20734 -13288
rect 22016 -13322 22124 -13288
rect 20626 -13334 22124 -13322
rect 22226 -11636 23724 -11624
rect 22226 -11670 22334 -11636
rect 23616 -11670 23724 -11636
rect 22226 -11682 23724 -11670
rect 22226 -11732 22284 -11682
rect 22226 -12100 22238 -11732
rect 22272 -12100 22284 -11732
rect 23666 -11732 23724 -11682
rect 22226 -12150 22284 -12100
rect 23666 -12100 23678 -11732
rect 23712 -12100 23724 -11732
rect 23666 -12150 23724 -12100
rect 22226 -12162 23724 -12150
rect 22226 -12196 22334 -12162
rect 23616 -12196 23724 -12162
rect 22226 -12208 23724 -12196
rect 22226 -12258 22284 -12208
rect 22226 -13226 22238 -12258
rect 22272 -13226 22284 -12258
rect 23666 -12258 23724 -12208
rect 22226 -13276 22284 -13226
rect 23666 -13226 23678 -12258
rect 23712 -13226 23724 -12258
rect 23666 -13276 23724 -13226
rect 22226 -13288 23724 -13276
rect 22226 -13322 22334 -13288
rect 23616 -13322 23724 -13288
rect 22226 -13334 23724 -13322
rect 23826 -11636 25324 -11624
rect 23826 -11670 23934 -11636
rect 25216 -11670 25324 -11636
rect 23826 -11682 25324 -11670
rect 23826 -11732 23884 -11682
rect 23826 -12100 23838 -11732
rect 23872 -12100 23884 -11732
rect 25266 -11732 25324 -11682
rect 23826 -12150 23884 -12100
rect 25266 -12100 25278 -11732
rect 25312 -12100 25324 -11732
rect 25266 -12150 25324 -12100
rect 23826 -12162 25324 -12150
rect 23826 -12196 23934 -12162
rect 25216 -12196 25324 -12162
rect 23826 -12208 25324 -12196
rect 23826 -12258 23884 -12208
rect 23826 -13226 23838 -12258
rect 23872 -13226 23884 -12258
rect 25266 -12258 25324 -12208
rect 23826 -13276 23884 -13226
rect 25266 -13226 25278 -12258
rect 25312 -13226 25324 -12258
rect 25266 -13276 25324 -13226
rect 23826 -13288 25324 -13276
rect 23826 -13322 23934 -13288
rect 25216 -13322 25324 -13288
rect 23826 -13334 25324 -13322
rect 25426 -11636 26924 -11624
rect 25426 -11670 25534 -11636
rect 26816 -11670 26924 -11636
rect 25426 -11682 26924 -11670
rect 25426 -11732 25484 -11682
rect 25426 -12100 25438 -11732
rect 25472 -12100 25484 -11732
rect 26866 -11732 26924 -11682
rect 25426 -12150 25484 -12100
rect 26866 -12100 26878 -11732
rect 26912 -12100 26924 -11732
rect 26866 -12150 26924 -12100
rect 25426 -12162 26924 -12150
rect 25426 -12196 25534 -12162
rect 26816 -12196 26924 -12162
rect 25426 -12208 26924 -12196
rect 25426 -12258 25484 -12208
rect 25426 -13226 25438 -12258
rect 25472 -13226 25484 -12258
rect 26866 -12258 26924 -12208
rect 25426 -13276 25484 -13226
rect 26866 -13226 26878 -12258
rect 26912 -13226 26924 -12258
rect 26866 -13276 26924 -13226
rect 25426 -13288 26924 -13276
rect 25426 -13322 25534 -13288
rect 26816 -13322 26924 -13288
rect 25426 -13334 26924 -13322
rect 27026 -11636 28524 -11624
rect 27026 -11670 27134 -11636
rect 28416 -11670 28524 -11636
rect 27026 -11682 28524 -11670
rect 27026 -11732 27084 -11682
rect 27026 -12100 27038 -11732
rect 27072 -12100 27084 -11732
rect 28466 -11732 28524 -11682
rect 27026 -12150 27084 -12100
rect 28466 -12100 28478 -11732
rect 28512 -12100 28524 -11732
rect 28466 -12150 28524 -12100
rect 27026 -12162 28524 -12150
rect 27026 -12196 27134 -12162
rect 28416 -12196 28524 -12162
rect 27026 -12208 28524 -12196
rect 27026 -12258 27084 -12208
rect 27026 -13226 27038 -12258
rect 27072 -13226 27084 -12258
rect 28466 -12258 28524 -12208
rect 27026 -13276 27084 -13226
rect 28466 -13226 28478 -12258
rect 28512 -13226 28524 -12258
rect 28466 -13276 28524 -13226
rect 27026 -13288 28524 -13276
rect 27026 -13322 27134 -13288
rect 28416 -13322 28524 -13288
rect 27026 -13334 28524 -13322
rect 28626 -11636 30124 -11624
rect 28626 -11670 28734 -11636
rect 30016 -11670 30124 -11636
rect 28626 -11682 30124 -11670
rect 28626 -11732 28684 -11682
rect 28626 -12100 28638 -11732
rect 28672 -12100 28684 -11732
rect 30066 -11732 30124 -11682
rect 28626 -12150 28684 -12100
rect 30066 -12100 30078 -11732
rect 30112 -12100 30124 -11732
rect 30066 -12150 30124 -12100
rect 28626 -12162 30124 -12150
rect 28626 -12196 28734 -12162
rect 30016 -12196 30124 -12162
rect 28626 -12208 30124 -12196
rect 28626 -12258 28684 -12208
rect 28626 -13226 28638 -12258
rect 28672 -13226 28684 -12258
rect 30066 -12258 30124 -12208
rect 28626 -13276 28684 -13226
rect 30066 -13226 30078 -12258
rect 30112 -13226 30124 -12258
rect 30066 -13276 30124 -13226
rect 28626 -13288 30124 -13276
rect 28626 -13322 28734 -13288
rect 30016 -13322 30124 -13288
rect 28626 -13334 30124 -13322
rect 30226 -11636 31724 -11624
rect 30226 -11670 30334 -11636
rect 31616 -11670 31724 -11636
rect 30226 -11682 31724 -11670
rect 30226 -11732 30284 -11682
rect 30226 -12100 30238 -11732
rect 30272 -12100 30284 -11732
rect 31666 -11732 31724 -11682
rect 30226 -12150 30284 -12100
rect 31666 -12100 31678 -11732
rect 31712 -12100 31724 -11732
rect 31666 -12150 31724 -12100
rect 30226 -12162 31724 -12150
rect 30226 -12196 30334 -12162
rect 31616 -12196 31724 -12162
rect 30226 -12208 31724 -12196
rect 30226 -12258 30284 -12208
rect 30226 -13226 30238 -12258
rect 30272 -13226 30284 -12258
rect 31666 -12258 31724 -12208
rect 30226 -13276 30284 -13226
rect 31666 -13226 31678 -12258
rect 31712 -13226 31724 -12258
rect 31666 -13276 31724 -13226
rect 30226 -13288 31724 -13276
rect 30226 -13322 30334 -13288
rect 31616 -13322 31724 -13288
rect 30226 -13334 31724 -13322
rect 31826 -11636 33324 -11624
rect 31826 -11670 31934 -11636
rect 33216 -11670 33324 -11636
rect 31826 -11682 33324 -11670
rect 31826 -11732 31884 -11682
rect 31826 -12100 31838 -11732
rect 31872 -12100 31884 -11732
rect 33266 -11732 33324 -11682
rect 31826 -12150 31884 -12100
rect 33266 -12100 33278 -11732
rect 33312 -12100 33324 -11732
rect 33266 -12150 33324 -12100
rect 31826 -12162 33324 -12150
rect 31826 -12196 31934 -12162
rect 33216 -12196 33324 -12162
rect 31826 -12208 33324 -12196
rect 31826 -12258 31884 -12208
rect 31826 -13226 31838 -12258
rect 31872 -13226 31884 -12258
rect 33266 -12258 33324 -12208
rect 31826 -13276 31884 -13226
rect 33266 -13226 33278 -12258
rect 33312 -13226 33324 -12258
rect 33266 -13276 33324 -13226
rect 31826 -13288 33324 -13276
rect 31826 -13322 31934 -13288
rect 33216 -13322 33324 -13288
rect 31826 -13334 33324 -13322
rect 33426 -11636 34924 -11624
rect 33426 -11670 33534 -11636
rect 34816 -11670 34924 -11636
rect 33426 -11682 34924 -11670
rect 33426 -11732 33484 -11682
rect 33426 -12100 33438 -11732
rect 33472 -12100 33484 -11732
rect 34866 -11732 34924 -11682
rect 33426 -12150 33484 -12100
rect 34866 -12100 34878 -11732
rect 34912 -12100 34924 -11732
rect 34866 -12150 34924 -12100
rect 33426 -12162 34924 -12150
rect 33426 -12196 33534 -12162
rect 34816 -12196 34924 -12162
rect 33426 -12208 34924 -12196
rect 33426 -12258 33484 -12208
rect 33426 -13226 33438 -12258
rect 33472 -13226 33484 -12258
rect 34866 -12258 34924 -12208
rect 33426 -13276 33484 -13226
rect 34866 -13226 34878 -12258
rect 34912 -13226 34924 -12258
rect 34866 -13276 34924 -13226
rect 33426 -13288 34924 -13276
rect 33426 -13322 33534 -13288
rect 34816 -13322 34924 -13288
rect 33426 -13334 34924 -13322
rect 35026 -11636 36524 -11624
rect 35026 -11670 35134 -11636
rect 36416 -11670 36524 -11636
rect 35026 -11682 36524 -11670
rect 35026 -11732 35084 -11682
rect 35026 -12100 35038 -11732
rect 35072 -12100 35084 -11732
rect 36466 -11732 36524 -11682
rect 35026 -12150 35084 -12100
rect 36466 -12100 36478 -11732
rect 36512 -12100 36524 -11732
rect 36466 -12150 36524 -12100
rect 35026 -12162 36524 -12150
rect 35026 -12196 35134 -12162
rect 36416 -12196 36524 -12162
rect 35026 -12208 36524 -12196
rect 35026 -12258 35084 -12208
rect 35026 -13226 35038 -12258
rect 35072 -13226 35084 -12258
rect 36466 -12258 36524 -12208
rect 35026 -13276 35084 -13226
rect 36466 -13226 36478 -12258
rect 36512 -13226 36524 -12258
rect 36466 -13276 36524 -13226
rect 35026 -13288 36524 -13276
rect 35026 -13322 35134 -13288
rect 36416 -13322 36524 -13288
rect 35026 -13334 36524 -13322
rect 36626 -11636 38124 -11624
rect 36626 -11670 36734 -11636
rect 38016 -11670 38124 -11636
rect 36626 -11682 38124 -11670
rect 36626 -11732 36684 -11682
rect 36626 -12100 36638 -11732
rect 36672 -12100 36684 -11732
rect 38066 -11732 38124 -11682
rect 36626 -12150 36684 -12100
rect 38066 -12100 38078 -11732
rect 38112 -12100 38124 -11732
rect 38066 -12150 38124 -12100
rect 36626 -12162 38124 -12150
rect 36626 -12196 36734 -12162
rect 38016 -12196 38124 -12162
rect 36626 -12208 38124 -12196
rect 36626 -12258 36684 -12208
rect 36626 -13226 36638 -12258
rect 36672 -13226 36684 -12258
rect 38066 -12258 38124 -12208
rect 36626 -13276 36684 -13226
rect 38066 -13226 38078 -12258
rect 38112 -13226 38124 -12258
rect 38066 -13276 38124 -13226
rect 36626 -13288 38124 -13276
rect 36626 -13322 36734 -13288
rect 38016 -13322 38124 -13288
rect 36626 -13334 38124 -13322
rect -174 -13436 1324 -13424
rect -174 -13470 -66 -13436
rect 1216 -13470 1324 -13436
rect -174 -13482 1324 -13470
rect -174 -13532 -116 -13482
rect -174 -13900 -162 -13532
rect -128 -13900 -116 -13532
rect 1266 -13532 1324 -13482
rect -174 -13950 -116 -13900
rect 1266 -13900 1278 -13532
rect 1312 -13900 1324 -13532
rect 1266 -13950 1324 -13900
rect -174 -13962 1324 -13950
rect -174 -13996 -66 -13962
rect 1216 -13996 1324 -13962
rect -174 -14008 1324 -13996
rect -174 -14058 -116 -14008
rect -174 -15026 -162 -14058
rect -128 -15026 -116 -14058
rect 1266 -14058 1324 -14008
rect -174 -15076 -116 -15026
rect 1266 -15026 1278 -14058
rect 1312 -15026 1324 -14058
rect 1266 -15076 1324 -15026
rect -174 -15088 1324 -15076
rect -174 -15122 -66 -15088
rect 1216 -15122 1324 -15088
rect -174 -15134 1324 -15122
rect 1426 -13436 2924 -13424
rect 1426 -13470 1534 -13436
rect 2816 -13470 2924 -13436
rect 1426 -13482 2924 -13470
rect 1426 -13532 1484 -13482
rect 1426 -13900 1438 -13532
rect 1472 -13900 1484 -13532
rect 2866 -13532 2924 -13482
rect 1426 -13950 1484 -13900
rect 2866 -13900 2878 -13532
rect 2912 -13900 2924 -13532
rect 2866 -13950 2924 -13900
rect 1426 -13962 2924 -13950
rect 1426 -13996 1534 -13962
rect 2816 -13996 2924 -13962
rect 1426 -14008 2924 -13996
rect 1426 -14058 1484 -14008
rect 1426 -15026 1438 -14058
rect 1472 -15026 1484 -14058
rect 2866 -14058 2924 -14008
rect 1426 -15076 1484 -15026
rect 2866 -15026 2878 -14058
rect 2912 -15026 2924 -14058
rect 2866 -15076 2924 -15026
rect 1426 -15088 2924 -15076
rect 1426 -15122 1534 -15088
rect 2816 -15122 2924 -15088
rect 1426 -15134 2924 -15122
rect 3026 -13436 4524 -13424
rect 3026 -13470 3134 -13436
rect 4416 -13470 4524 -13436
rect 3026 -13482 4524 -13470
rect 3026 -13532 3084 -13482
rect 3026 -13900 3038 -13532
rect 3072 -13900 3084 -13532
rect 4466 -13532 4524 -13482
rect 3026 -13950 3084 -13900
rect 4466 -13900 4478 -13532
rect 4512 -13900 4524 -13532
rect 4466 -13950 4524 -13900
rect 3026 -13962 4524 -13950
rect 3026 -13996 3134 -13962
rect 4416 -13996 4524 -13962
rect 3026 -14008 4524 -13996
rect 3026 -14058 3084 -14008
rect 3026 -15026 3038 -14058
rect 3072 -15026 3084 -14058
rect 4466 -14058 4524 -14008
rect 3026 -15076 3084 -15026
rect 4466 -15026 4478 -14058
rect 4512 -15026 4524 -14058
rect 4466 -15076 4524 -15026
rect 3026 -15088 4524 -15076
rect 3026 -15122 3134 -15088
rect 4416 -15122 4524 -15088
rect 3026 -15134 4524 -15122
rect 4626 -13436 6124 -13424
rect 4626 -13470 4734 -13436
rect 6016 -13470 6124 -13436
rect 4626 -13482 6124 -13470
rect 4626 -13532 4684 -13482
rect 4626 -13900 4638 -13532
rect 4672 -13900 4684 -13532
rect 6066 -13532 6124 -13482
rect 4626 -13950 4684 -13900
rect 6066 -13900 6078 -13532
rect 6112 -13900 6124 -13532
rect 6066 -13950 6124 -13900
rect 4626 -13962 6124 -13950
rect 4626 -13996 4734 -13962
rect 6016 -13996 6124 -13962
rect 4626 -14008 6124 -13996
rect 4626 -14058 4684 -14008
rect 4626 -15026 4638 -14058
rect 4672 -15026 4684 -14058
rect 6066 -14058 6124 -14008
rect 4626 -15076 4684 -15026
rect 6066 -15026 6078 -14058
rect 6112 -15026 6124 -14058
rect 6066 -15076 6124 -15026
rect 4626 -15088 6124 -15076
rect 4626 -15122 4734 -15088
rect 6016 -15122 6124 -15088
rect 4626 -15134 6124 -15122
rect 6226 -13436 7724 -13424
rect 6226 -13470 6334 -13436
rect 7616 -13470 7724 -13436
rect 6226 -13482 7724 -13470
rect 6226 -13532 6284 -13482
rect 6226 -13900 6238 -13532
rect 6272 -13900 6284 -13532
rect 7666 -13532 7724 -13482
rect 6226 -13950 6284 -13900
rect 7666 -13900 7678 -13532
rect 7712 -13900 7724 -13532
rect 7666 -13950 7724 -13900
rect 6226 -13962 7724 -13950
rect 6226 -13996 6334 -13962
rect 7616 -13996 7724 -13962
rect 6226 -14008 7724 -13996
rect 6226 -14058 6284 -14008
rect 6226 -15026 6238 -14058
rect 6272 -15026 6284 -14058
rect 7666 -14058 7724 -14008
rect 6226 -15076 6284 -15026
rect 7666 -15026 7678 -14058
rect 7712 -15026 7724 -14058
rect 7666 -15076 7724 -15026
rect 6226 -15088 7724 -15076
rect 6226 -15122 6334 -15088
rect 7616 -15122 7724 -15088
rect 6226 -15134 7724 -15122
rect 7826 -13436 9324 -13424
rect 7826 -13470 7934 -13436
rect 9216 -13470 9324 -13436
rect 7826 -13482 9324 -13470
rect 7826 -13532 7884 -13482
rect 7826 -13900 7838 -13532
rect 7872 -13900 7884 -13532
rect 9266 -13532 9324 -13482
rect 7826 -13950 7884 -13900
rect 9266 -13900 9278 -13532
rect 9312 -13900 9324 -13532
rect 9266 -13950 9324 -13900
rect 7826 -13962 9324 -13950
rect 7826 -13996 7934 -13962
rect 9216 -13996 9324 -13962
rect 7826 -14008 9324 -13996
rect 7826 -14058 7884 -14008
rect 7826 -15026 7838 -14058
rect 7872 -15026 7884 -14058
rect 9266 -14058 9324 -14008
rect 7826 -15076 7884 -15026
rect 9266 -15026 9278 -14058
rect 9312 -15026 9324 -14058
rect 9266 -15076 9324 -15026
rect 7826 -15088 9324 -15076
rect 7826 -15122 7934 -15088
rect 9216 -15122 9324 -15088
rect 7826 -15134 9324 -15122
rect 9426 -13436 10924 -13424
rect 9426 -13470 9534 -13436
rect 10816 -13470 10924 -13436
rect 9426 -13482 10924 -13470
rect 9426 -13532 9484 -13482
rect 9426 -13900 9438 -13532
rect 9472 -13900 9484 -13532
rect 10866 -13532 10924 -13482
rect 9426 -13950 9484 -13900
rect 10866 -13900 10878 -13532
rect 10912 -13900 10924 -13532
rect 10866 -13950 10924 -13900
rect 9426 -13962 10924 -13950
rect 9426 -13996 9534 -13962
rect 10816 -13996 10924 -13962
rect 9426 -14008 10924 -13996
rect 9426 -14058 9484 -14008
rect 9426 -15026 9438 -14058
rect 9472 -15026 9484 -14058
rect 10866 -14058 10924 -14008
rect 9426 -15076 9484 -15026
rect 10866 -15026 10878 -14058
rect 10912 -15026 10924 -14058
rect 10866 -15076 10924 -15026
rect 9426 -15088 10924 -15076
rect 9426 -15122 9534 -15088
rect 10816 -15122 10924 -15088
rect 9426 -15134 10924 -15122
rect 11026 -13436 12524 -13424
rect 11026 -13470 11134 -13436
rect 12416 -13470 12524 -13436
rect 11026 -13482 12524 -13470
rect 11026 -13532 11084 -13482
rect 11026 -13900 11038 -13532
rect 11072 -13900 11084 -13532
rect 12466 -13532 12524 -13482
rect 11026 -13950 11084 -13900
rect 12466 -13900 12478 -13532
rect 12512 -13900 12524 -13532
rect 12466 -13950 12524 -13900
rect 11026 -13962 12524 -13950
rect 11026 -13996 11134 -13962
rect 12416 -13996 12524 -13962
rect 11026 -14008 12524 -13996
rect 11026 -14058 11084 -14008
rect 11026 -15026 11038 -14058
rect 11072 -15026 11084 -14058
rect 12466 -14058 12524 -14008
rect 11026 -15076 11084 -15026
rect 12466 -15026 12478 -14058
rect 12512 -15026 12524 -14058
rect 12466 -15076 12524 -15026
rect 11026 -15088 12524 -15076
rect 11026 -15122 11134 -15088
rect 12416 -15122 12524 -15088
rect 11026 -15134 12524 -15122
rect 12626 -13436 14124 -13424
rect 12626 -13470 12734 -13436
rect 14016 -13470 14124 -13436
rect 12626 -13482 14124 -13470
rect 12626 -13532 12684 -13482
rect 12626 -13900 12638 -13532
rect 12672 -13900 12684 -13532
rect 14066 -13532 14124 -13482
rect 12626 -13950 12684 -13900
rect 14066 -13900 14078 -13532
rect 14112 -13900 14124 -13532
rect 14066 -13950 14124 -13900
rect 12626 -13962 14124 -13950
rect 12626 -13996 12734 -13962
rect 14016 -13996 14124 -13962
rect 12626 -14008 14124 -13996
rect 12626 -14058 12684 -14008
rect 12626 -15026 12638 -14058
rect 12672 -15026 12684 -14058
rect 14066 -14058 14124 -14008
rect 12626 -15076 12684 -15026
rect 14066 -15026 14078 -14058
rect 14112 -15026 14124 -14058
rect 14066 -15076 14124 -15026
rect 12626 -15088 14124 -15076
rect 12626 -15122 12734 -15088
rect 14016 -15122 14124 -15088
rect 12626 -15134 14124 -15122
rect 14226 -13436 15724 -13424
rect 14226 -13470 14334 -13436
rect 15616 -13470 15724 -13436
rect 14226 -13482 15724 -13470
rect 14226 -13532 14284 -13482
rect 14226 -13900 14238 -13532
rect 14272 -13900 14284 -13532
rect 15666 -13532 15724 -13482
rect 14226 -13950 14284 -13900
rect 15666 -13900 15678 -13532
rect 15712 -13900 15724 -13532
rect 15666 -13950 15724 -13900
rect 14226 -13962 15724 -13950
rect 14226 -13996 14334 -13962
rect 15616 -13996 15724 -13962
rect 14226 -14008 15724 -13996
rect 14226 -14058 14284 -14008
rect 14226 -15026 14238 -14058
rect 14272 -15026 14284 -14058
rect 15666 -14058 15724 -14008
rect 14226 -15076 14284 -15026
rect 15666 -15026 15678 -14058
rect 15712 -15026 15724 -14058
rect 15666 -15076 15724 -15026
rect 14226 -15088 15724 -15076
rect 14226 -15122 14334 -15088
rect 15616 -15122 15724 -15088
rect 14226 -15134 15724 -15122
rect 15826 -13436 17324 -13424
rect 15826 -13470 15934 -13436
rect 17216 -13470 17324 -13436
rect 15826 -13482 17324 -13470
rect 15826 -13532 15884 -13482
rect 15826 -13900 15838 -13532
rect 15872 -13900 15884 -13532
rect 17266 -13532 17324 -13482
rect 15826 -13950 15884 -13900
rect 17266 -13900 17278 -13532
rect 17312 -13900 17324 -13532
rect 17266 -13950 17324 -13900
rect 15826 -13962 17324 -13950
rect 15826 -13996 15934 -13962
rect 17216 -13996 17324 -13962
rect 15826 -14008 17324 -13996
rect 15826 -14058 15884 -14008
rect 15826 -15026 15838 -14058
rect 15872 -15026 15884 -14058
rect 17266 -14058 17324 -14008
rect 15826 -15076 15884 -15026
rect 17266 -15026 17278 -14058
rect 17312 -15026 17324 -14058
rect 17266 -15076 17324 -15026
rect 15826 -15088 17324 -15076
rect 15826 -15122 15934 -15088
rect 17216 -15122 17324 -15088
rect 15826 -15134 17324 -15122
rect 17426 -13436 18924 -13424
rect 17426 -13470 17534 -13436
rect 18816 -13470 18924 -13436
rect 17426 -13482 18924 -13470
rect 17426 -13532 17484 -13482
rect 17426 -13900 17438 -13532
rect 17472 -13900 17484 -13532
rect 18866 -13532 18924 -13482
rect 17426 -13950 17484 -13900
rect 18866 -13900 18878 -13532
rect 18912 -13900 18924 -13532
rect 18866 -13950 18924 -13900
rect 17426 -13962 18924 -13950
rect 17426 -13996 17534 -13962
rect 18816 -13996 18924 -13962
rect 17426 -14008 18924 -13996
rect 17426 -14058 17484 -14008
rect 17426 -15026 17438 -14058
rect 17472 -15026 17484 -14058
rect 18866 -14058 18924 -14008
rect 17426 -15076 17484 -15026
rect 18866 -15026 18878 -14058
rect 18912 -15026 18924 -14058
rect 18866 -15076 18924 -15026
rect 17426 -15088 18924 -15076
rect 17426 -15122 17534 -15088
rect 18816 -15122 18924 -15088
rect 17426 -15134 18924 -15122
rect 19026 -13436 20524 -13424
rect 19026 -13470 19134 -13436
rect 20416 -13470 20524 -13436
rect 19026 -13482 20524 -13470
rect 19026 -13532 19084 -13482
rect 19026 -13900 19038 -13532
rect 19072 -13900 19084 -13532
rect 20466 -13532 20524 -13482
rect 19026 -13950 19084 -13900
rect 20466 -13900 20478 -13532
rect 20512 -13900 20524 -13532
rect 20466 -13950 20524 -13900
rect 19026 -13962 20524 -13950
rect 19026 -13996 19134 -13962
rect 20416 -13996 20524 -13962
rect 19026 -14008 20524 -13996
rect 19026 -14058 19084 -14008
rect 19026 -15026 19038 -14058
rect 19072 -15026 19084 -14058
rect 20466 -14058 20524 -14008
rect 19026 -15076 19084 -15026
rect 20466 -15026 20478 -14058
rect 20512 -15026 20524 -14058
rect 20466 -15076 20524 -15026
rect 19026 -15088 20524 -15076
rect 19026 -15122 19134 -15088
rect 20416 -15122 20524 -15088
rect 19026 -15134 20524 -15122
rect 20626 -13436 22124 -13424
rect 20626 -13470 20734 -13436
rect 22016 -13470 22124 -13436
rect 20626 -13482 22124 -13470
rect 20626 -13532 20684 -13482
rect 20626 -13900 20638 -13532
rect 20672 -13900 20684 -13532
rect 22066 -13532 22124 -13482
rect 20626 -13950 20684 -13900
rect 22066 -13900 22078 -13532
rect 22112 -13900 22124 -13532
rect 22066 -13950 22124 -13900
rect 20626 -13962 22124 -13950
rect 20626 -13996 20734 -13962
rect 22016 -13996 22124 -13962
rect 20626 -14008 22124 -13996
rect 20626 -14058 20684 -14008
rect 20626 -15026 20638 -14058
rect 20672 -15026 20684 -14058
rect 22066 -14058 22124 -14008
rect 20626 -15076 20684 -15026
rect 22066 -15026 22078 -14058
rect 22112 -15026 22124 -14058
rect 22066 -15076 22124 -15026
rect 20626 -15088 22124 -15076
rect 20626 -15122 20734 -15088
rect 22016 -15122 22124 -15088
rect 20626 -15134 22124 -15122
rect 22226 -13436 23724 -13424
rect 22226 -13470 22334 -13436
rect 23616 -13470 23724 -13436
rect 22226 -13482 23724 -13470
rect 22226 -13532 22284 -13482
rect 22226 -13900 22238 -13532
rect 22272 -13900 22284 -13532
rect 23666 -13532 23724 -13482
rect 22226 -13950 22284 -13900
rect 23666 -13900 23678 -13532
rect 23712 -13900 23724 -13532
rect 23666 -13950 23724 -13900
rect 22226 -13962 23724 -13950
rect 22226 -13996 22334 -13962
rect 23616 -13996 23724 -13962
rect 22226 -14008 23724 -13996
rect 22226 -14058 22284 -14008
rect 22226 -15026 22238 -14058
rect 22272 -15026 22284 -14058
rect 23666 -14058 23724 -14008
rect 22226 -15076 22284 -15026
rect 23666 -15026 23678 -14058
rect 23712 -15026 23724 -14058
rect 23666 -15076 23724 -15026
rect 22226 -15088 23724 -15076
rect 22226 -15122 22334 -15088
rect 23616 -15122 23724 -15088
rect 22226 -15134 23724 -15122
rect 23826 -13436 25324 -13424
rect 23826 -13470 23934 -13436
rect 25216 -13470 25324 -13436
rect 23826 -13482 25324 -13470
rect 23826 -13532 23884 -13482
rect 23826 -13900 23838 -13532
rect 23872 -13900 23884 -13532
rect 25266 -13532 25324 -13482
rect 23826 -13950 23884 -13900
rect 25266 -13900 25278 -13532
rect 25312 -13900 25324 -13532
rect 25266 -13950 25324 -13900
rect 23826 -13962 25324 -13950
rect 23826 -13996 23934 -13962
rect 25216 -13996 25324 -13962
rect 23826 -14008 25324 -13996
rect 23826 -14058 23884 -14008
rect 23826 -15026 23838 -14058
rect 23872 -15026 23884 -14058
rect 25266 -14058 25324 -14008
rect 23826 -15076 23884 -15026
rect 25266 -15026 25278 -14058
rect 25312 -15026 25324 -14058
rect 25266 -15076 25324 -15026
rect 23826 -15088 25324 -15076
rect 23826 -15122 23934 -15088
rect 25216 -15122 25324 -15088
rect 23826 -15134 25324 -15122
rect 25426 -13436 26924 -13424
rect 25426 -13470 25534 -13436
rect 26816 -13470 26924 -13436
rect 25426 -13482 26924 -13470
rect 25426 -13532 25484 -13482
rect 25426 -13900 25438 -13532
rect 25472 -13900 25484 -13532
rect 26866 -13532 26924 -13482
rect 25426 -13950 25484 -13900
rect 26866 -13900 26878 -13532
rect 26912 -13900 26924 -13532
rect 26866 -13950 26924 -13900
rect 25426 -13962 26924 -13950
rect 25426 -13996 25534 -13962
rect 26816 -13996 26924 -13962
rect 25426 -14008 26924 -13996
rect 25426 -14058 25484 -14008
rect 25426 -15026 25438 -14058
rect 25472 -15026 25484 -14058
rect 26866 -14058 26924 -14008
rect 25426 -15076 25484 -15026
rect 26866 -15026 26878 -14058
rect 26912 -15026 26924 -14058
rect 26866 -15076 26924 -15026
rect 25426 -15088 26924 -15076
rect 25426 -15122 25534 -15088
rect 26816 -15122 26924 -15088
rect 25426 -15134 26924 -15122
rect 27026 -13436 28524 -13424
rect 27026 -13470 27134 -13436
rect 28416 -13470 28524 -13436
rect 27026 -13482 28524 -13470
rect 27026 -13532 27084 -13482
rect 27026 -13900 27038 -13532
rect 27072 -13900 27084 -13532
rect 28466 -13532 28524 -13482
rect 27026 -13950 27084 -13900
rect 28466 -13900 28478 -13532
rect 28512 -13900 28524 -13532
rect 28466 -13950 28524 -13900
rect 27026 -13962 28524 -13950
rect 27026 -13996 27134 -13962
rect 28416 -13996 28524 -13962
rect 27026 -14008 28524 -13996
rect 27026 -14058 27084 -14008
rect 27026 -15026 27038 -14058
rect 27072 -15026 27084 -14058
rect 28466 -14058 28524 -14008
rect 27026 -15076 27084 -15026
rect 28466 -15026 28478 -14058
rect 28512 -15026 28524 -14058
rect 28466 -15076 28524 -15026
rect 27026 -15088 28524 -15076
rect 27026 -15122 27134 -15088
rect 28416 -15122 28524 -15088
rect 27026 -15134 28524 -15122
rect 28626 -13436 30124 -13424
rect 28626 -13470 28734 -13436
rect 30016 -13470 30124 -13436
rect 28626 -13482 30124 -13470
rect 28626 -13532 28684 -13482
rect 28626 -13900 28638 -13532
rect 28672 -13900 28684 -13532
rect 30066 -13532 30124 -13482
rect 28626 -13950 28684 -13900
rect 30066 -13900 30078 -13532
rect 30112 -13900 30124 -13532
rect 30066 -13950 30124 -13900
rect 28626 -13962 30124 -13950
rect 28626 -13996 28734 -13962
rect 30016 -13996 30124 -13962
rect 28626 -14008 30124 -13996
rect 28626 -14058 28684 -14008
rect 28626 -15026 28638 -14058
rect 28672 -15026 28684 -14058
rect 30066 -14058 30124 -14008
rect 28626 -15076 28684 -15026
rect 30066 -15026 30078 -14058
rect 30112 -15026 30124 -14058
rect 30066 -15076 30124 -15026
rect 28626 -15088 30124 -15076
rect 28626 -15122 28734 -15088
rect 30016 -15122 30124 -15088
rect 28626 -15134 30124 -15122
rect 30226 -13436 31724 -13424
rect 30226 -13470 30334 -13436
rect 31616 -13470 31724 -13436
rect 30226 -13482 31724 -13470
rect 30226 -13532 30284 -13482
rect 30226 -13900 30238 -13532
rect 30272 -13900 30284 -13532
rect 31666 -13532 31724 -13482
rect 30226 -13950 30284 -13900
rect 31666 -13900 31678 -13532
rect 31712 -13900 31724 -13532
rect 31666 -13950 31724 -13900
rect 30226 -13962 31724 -13950
rect 30226 -13996 30334 -13962
rect 31616 -13996 31724 -13962
rect 30226 -14008 31724 -13996
rect 30226 -14058 30284 -14008
rect 30226 -15026 30238 -14058
rect 30272 -15026 30284 -14058
rect 31666 -14058 31724 -14008
rect 30226 -15076 30284 -15026
rect 31666 -15026 31678 -14058
rect 31712 -15026 31724 -14058
rect 31666 -15076 31724 -15026
rect 30226 -15088 31724 -15076
rect 30226 -15122 30334 -15088
rect 31616 -15122 31724 -15088
rect 30226 -15134 31724 -15122
rect 31826 -13436 33324 -13424
rect 31826 -13470 31934 -13436
rect 33216 -13470 33324 -13436
rect 31826 -13482 33324 -13470
rect 31826 -13532 31884 -13482
rect 31826 -13900 31838 -13532
rect 31872 -13900 31884 -13532
rect 33266 -13532 33324 -13482
rect 31826 -13950 31884 -13900
rect 33266 -13900 33278 -13532
rect 33312 -13900 33324 -13532
rect 33266 -13950 33324 -13900
rect 31826 -13962 33324 -13950
rect 31826 -13996 31934 -13962
rect 33216 -13996 33324 -13962
rect 31826 -14008 33324 -13996
rect 31826 -14058 31884 -14008
rect 31826 -15026 31838 -14058
rect 31872 -15026 31884 -14058
rect 33266 -14058 33324 -14008
rect 31826 -15076 31884 -15026
rect 33266 -15026 33278 -14058
rect 33312 -15026 33324 -14058
rect 33266 -15076 33324 -15026
rect 31826 -15088 33324 -15076
rect 31826 -15122 31934 -15088
rect 33216 -15122 33324 -15088
rect 31826 -15134 33324 -15122
rect 33426 -13436 34924 -13424
rect 33426 -13470 33534 -13436
rect 34816 -13470 34924 -13436
rect 33426 -13482 34924 -13470
rect 33426 -13532 33484 -13482
rect 33426 -13900 33438 -13532
rect 33472 -13900 33484 -13532
rect 34866 -13532 34924 -13482
rect 33426 -13950 33484 -13900
rect 34866 -13900 34878 -13532
rect 34912 -13900 34924 -13532
rect 34866 -13950 34924 -13900
rect 33426 -13962 34924 -13950
rect 33426 -13996 33534 -13962
rect 34816 -13996 34924 -13962
rect 33426 -14008 34924 -13996
rect 33426 -14058 33484 -14008
rect 33426 -15026 33438 -14058
rect 33472 -15026 33484 -14058
rect 34866 -14058 34924 -14008
rect 33426 -15076 33484 -15026
rect 34866 -15026 34878 -14058
rect 34912 -15026 34924 -14058
rect 34866 -15076 34924 -15026
rect 33426 -15088 34924 -15076
rect 33426 -15122 33534 -15088
rect 34816 -15122 34924 -15088
rect 33426 -15134 34924 -15122
rect 35026 -13436 36524 -13424
rect 35026 -13470 35134 -13436
rect 36416 -13470 36524 -13436
rect 35026 -13482 36524 -13470
rect 35026 -13532 35084 -13482
rect 35026 -13900 35038 -13532
rect 35072 -13900 35084 -13532
rect 36466 -13532 36524 -13482
rect 35026 -13950 35084 -13900
rect 36466 -13900 36478 -13532
rect 36512 -13900 36524 -13532
rect 36466 -13950 36524 -13900
rect 35026 -13962 36524 -13950
rect 35026 -13996 35134 -13962
rect 36416 -13996 36524 -13962
rect 35026 -14008 36524 -13996
rect 35026 -14058 35084 -14008
rect 35026 -15026 35038 -14058
rect 35072 -15026 35084 -14058
rect 36466 -14058 36524 -14008
rect 35026 -15076 35084 -15026
rect 36466 -15026 36478 -14058
rect 36512 -15026 36524 -14058
rect 36466 -15076 36524 -15026
rect 35026 -15088 36524 -15076
rect 35026 -15122 35134 -15088
rect 36416 -15122 36524 -15088
rect 35026 -15134 36524 -15122
rect 36626 -13436 38124 -13424
rect 36626 -13470 36734 -13436
rect 38016 -13470 38124 -13436
rect 36626 -13482 38124 -13470
rect 36626 -13532 36684 -13482
rect 36626 -13900 36638 -13532
rect 36672 -13900 36684 -13532
rect 38066 -13532 38124 -13482
rect 36626 -13950 36684 -13900
rect 38066 -13900 38078 -13532
rect 38112 -13900 38124 -13532
rect 38066 -13950 38124 -13900
rect 36626 -13962 38124 -13950
rect 36626 -13996 36734 -13962
rect 38016 -13996 38124 -13962
rect 36626 -14008 38124 -13996
rect 36626 -14058 36684 -14008
rect 36626 -15026 36638 -14058
rect 36672 -15026 36684 -14058
rect 38066 -14058 38124 -14008
rect 36626 -15076 36684 -15026
rect 38066 -15026 38078 -14058
rect 38112 -15026 38124 -14058
rect 38066 -15076 38124 -15026
rect 36626 -15088 38124 -15076
rect 36626 -15122 36734 -15088
rect 38016 -15122 38124 -15088
rect 36626 -15134 38124 -15122
rect -174 -15236 1324 -15224
rect -174 -15270 -66 -15236
rect 1216 -15270 1324 -15236
rect -174 -15282 1324 -15270
rect -174 -15332 -116 -15282
rect -174 -15700 -162 -15332
rect -128 -15700 -116 -15332
rect 1266 -15332 1324 -15282
rect -174 -15750 -116 -15700
rect 1266 -15700 1278 -15332
rect 1312 -15700 1324 -15332
rect 1266 -15750 1324 -15700
rect -174 -15762 1324 -15750
rect -174 -15796 -66 -15762
rect 1216 -15796 1324 -15762
rect -174 -15808 1324 -15796
rect -174 -15858 -116 -15808
rect -174 -16826 -162 -15858
rect -128 -16826 -116 -15858
rect 1266 -15858 1324 -15808
rect -174 -16876 -116 -16826
rect 1266 -16826 1278 -15858
rect 1312 -16826 1324 -15858
rect 1266 -16876 1324 -16826
rect -174 -16888 1324 -16876
rect -174 -16922 -66 -16888
rect 1216 -16922 1324 -16888
rect -174 -16934 1324 -16922
rect 1426 -15236 2924 -15224
rect 1426 -15270 1534 -15236
rect 2816 -15270 2924 -15236
rect 1426 -15282 2924 -15270
rect 1426 -15332 1484 -15282
rect 1426 -15700 1438 -15332
rect 1472 -15700 1484 -15332
rect 2866 -15332 2924 -15282
rect 1426 -15750 1484 -15700
rect 2866 -15700 2878 -15332
rect 2912 -15700 2924 -15332
rect 2866 -15750 2924 -15700
rect 1426 -15762 2924 -15750
rect 1426 -15796 1534 -15762
rect 2816 -15796 2924 -15762
rect 1426 -15808 2924 -15796
rect 1426 -15858 1484 -15808
rect 1426 -16826 1438 -15858
rect 1472 -16826 1484 -15858
rect 2866 -15858 2924 -15808
rect 1426 -16876 1484 -16826
rect 2866 -16826 2878 -15858
rect 2912 -16826 2924 -15858
rect 2866 -16876 2924 -16826
rect 1426 -16888 2924 -16876
rect 1426 -16922 1534 -16888
rect 2816 -16922 2924 -16888
rect 1426 -16934 2924 -16922
rect 3026 -15236 4524 -15224
rect 3026 -15270 3134 -15236
rect 4416 -15270 4524 -15236
rect 3026 -15282 4524 -15270
rect 3026 -15332 3084 -15282
rect 3026 -15700 3038 -15332
rect 3072 -15700 3084 -15332
rect 4466 -15332 4524 -15282
rect 3026 -15750 3084 -15700
rect 4466 -15700 4478 -15332
rect 4512 -15700 4524 -15332
rect 4466 -15750 4524 -15700
rect 3026 -15762 4524 -15750
rect 3026 -15796 3134 -15762
rect 4416 -15796 4524 -15762
rect 3026 -15808 4524 -15796
rect 3026 -15858 3084 -15808
rect 3026 -16826 3038 -15858
rect 3072 -16826 3084 -15858
rect 4466 -15858 4524 -15808
rect 3026 -16876 3084 -16826
rect 4466 -16826 4478 -15858
rect 4512 -16826 4524 -15858
rect 4466 -16876 4524 -16826
rect 3026 -16888 4524 -16876
rect 3026 -16922 3134 -16888
rect 4416 -16922 4524 -16888
rect 3026 -16934 4524 -16922
rect 4626 -15236 6124 -15224
rect 4626 -15270 4734 -15236
rect 6016 -15270 6124 -15236
rect 4626 -15282 6124 -15270
rect 4626 -15332 4684 -15282
rect 4626 -15700 4638 -15332
rect 4672 -15700 4684 -15332
rect 6066 -15332 6124 -15282
rect 4626 -15750 4684 -15700
rect 6066 -15700 6078 -15332
rect 6112 -15700 6124 -15332
rect 6066 -15750 6124 -15700
rect 4626 -15762 6124 -15750
rect 4626 -15796 4734 -15762
rect 6016 -15796 6124 -15762
rect 4626 -15808 6124 -15796
rect 4626 -15858 4684 -15808
rect 4626 -16826 4638 -15858
rect 4672 -16826 4684 -15858
rect 6066 -15858 6124 -15808
rect 4626 -16876 4684 -16826
rect 6066 -16826 6078 -15858
rect 6112 -16826 6124 -15858
rect 6066 -16876 6124 -16826
rect 4626 -16888 6124 -16876
rect 4626 -16922 4734 -16888
rect 6016 -16922 6124 -16888
rect 4626 -16934 6124 -16922
rect 6226 -15236 7724 -15224
rect 6226 -15270 6334 -15236
rect 7616 -15270 7724 -15236
rect 6226 -15282 7724 -15270
rect 6226 -15332 6284 -15282
rect 6226 -15700 6238 -15332
rect 6272 -15700 6284 -15332
rect 7666 -15332 7724 -15282
rect 6226 -15750 6284 -15700
rect 7666 -15700 7678 -15332
rect 7712 -15700 7724 -15332
rect 7666 -15750 7724 -15700
rect 6226 -15762 7724 -15750
rect 6226 -15796 6334 -15762
rect 7616 -15796 7724 -15762
rect 6226 -15808 7724 -15796
rect 6226 -15858 6284 -15808
rect 6226 -16826 6238 -15858
rect 6272 -16826 6284 -15858
rect 7666 -15858 7724 -15808
rect 6226 -16876 6284 -16826
rect 7666 -16826 7678 -15858
rect 7712 -16826 7724 -15858
rect 7666 -16876 7724 -16826
rect 6226 -16888 7724 -16876
rect 6226 -16922 6334 -16888
rect 7616 -16922 7724 -16888
rect 6226 -16934 7724 -16922
rect 7826 -15236 9324 -15224
rect 7826 -15270 7934 -15236
rect 9216 -15270 9324 -15236
rect 7826 -15282 9324 -15270
rect 7826 -15332 7884 -15282
rect 7826 -15700 7838 -15332
rect 7872 -15700 7884 -15332
rect 9266 -15332 9324 -15282
rect 7826 -15750 7884 -15700
rect 9266 -15700 9278 -15332
rect 9312 -15700 9324 -15332
rect 9266 -15750 9324 -15700
rect 7826 -15762 9324 -15750
rect 7826 -15796 7934 -15762
rect 9216 -15796 9324 -15762
rect 7826 -15808 9324 -15796
rect 7826 -15858 7884 -15808
rect 7826 -16826 7838 -15858
rect 7872 -16826 7884 -15858
rect 9266 -15858 9324 -15808
rect 7826 -16876 7884 -16826
rect 9266 -16826 9278 -15858
rect 9312 -16826 9324 -15858
rect 9266 -16876 9324 -16826
rect 7826 -16888 9324 -16876
rect 7826 -16922 7934 -16888
rect 9216 -16922 9324 -16888
rect 7826 -16934 9324 -16922
rect 9426 -15236 10924 -15224
rect 9426 -15270 9534 -15236
rect 10816 -15270 10924 -15236
rect 9426 -15282 10924 -15270
rect 9426 -15332 9484 -15282
rect 9426 -15700 9438 -15332
rect 9472 -15700 9484 -15332
rect 10866 -15332 10924 -15282
rect 9426 -15750 9484 -15700
rect 10866 -15700 10878 -15332
rect 10912 -15700 10924 -15332
rect 10866 -15750 10924 -15700
rect 9426 -15762 10924 -15750
rect 9426 -15796 9534 -15762
rect 10816 -15796 10924 -15762
rect 9426 -15808 10924 -15796
rect 9426 -15858 9484 -15808
rect 9426 -16826 9438 -15858
rect 9472 -16826 9484 -15858
rect 10866 -15858 10924 -15808
rect 9426 -16876 9484 -16826
rect 10866 -16826 10878 -15858
rect 10912 -16826 10924 -15858
rect 10866 -16876 10924 -16826
rect 9426 -16888 10924 -16876
rect 9426 -16922 9534 -16888
rect 10816 -16922 10924 -16888
rect 9426 -16934 10924 -16922
rect 11026 -15236 12524 -15224
rect 11026 -15270 11134 -15236
rect 12416 -15270 12524 -15236
rect 11026 -15282 12524 -15270
rect 11026 -15332 11084 -15282
rect 11026 -15700 11038 -15332
rect 11072 -15700 11084 -15332
rect 12466 -15332 12524 -15282
rect 11026 -15750 11084 -15700
rect 12466 -15700 12478 -15332
rect 12512 -15700 12524 -15332
rect 12466 -15750 12524 -15700
rect 11026 -15762 12524 -15750
rect 11026 -15796 11134 -15762
rect 12416 -15796 12524 -15762
rect 11026 -15808 12524 -15796
rect 11026 -15858 11084 -15808
rect 11026 -16826 11038 -15858
rect 11072 -16826 11084 -15858
rect 12466 -15858 12524 -15808
rect 11026 -16876 11084 -16826
rect 12466 -16826 12478 -15858
rect 12512 -16826 12524 -15858
rect 12466 -16876 12524 -16826
rect 11026 -16888 12524 -16876
rect 11026 -16922 11134 -16888
rect 12416 -16922 12524 -16888
rect 11026 -16934 12524 -16922
rect 12626 -15236 14124 -15224
rect 12626 -15270 12734 -15236
rect 14016 -15270 14124 -15236
rect 12626 -15282 14124 -15270
rect 12626 -15332 12684 -15282
rect 12626 -15700 12638 -15332
rect 12672 -15700 12684 -15332
rect 14066 -15332 14124 -15282
rect 12626 -15750 12684 -15700
rect 14066 -15700 14078 -15332
rect 14112 -15700 14124 -15332
rect 14066 -15750 14124 -15700
rect 12626 -15762 14124 -15750
rect 12626 -15796 12734 -15762
rect 14016 -15796 14124 -15762
rect 12626 -15808 14124 -15796
rect 12626 -15858 12684 -15808
rect 12626 -16826 12638 -15858
rect 12672 -16826 12684 -15858
rect 14066 -15858 14124 -15808
rect 12626 -16876 12684 -16826
rect 14066 -16826 14078 -15858
rect 14112 -16826 14124 -15858
rect 14066 -16876 14124 -16826
rect 12626 -16888 14124 -16876
rect 12626 -16922 12734 -16888
rect 14016 -16922 14124 -16888
rect 12626 -16934 14124 -16922
rect 14226 -15236 15724 -15224
rect 14226 -15270 14334 -15236
rect 15616 -15270 15724 -15236
rect 14226 -15282 15724 -15270
rect 14226 -15332 14284 -15282
rect 14226 -15700 14238 -15332
rect 14272 -15700 14284 -15332
rect 15666 -15332 15724 -15282
rect 14226 -15750 14284 -15700
rect 15666 -15700 15678 -15332
rect 15712 -15700 15724 -15332
rect 15666 -15750 15724 -15700
rect 14226 -15762 15724 -15750
rect 14226 -15796 14334 -15762
rect 15616 -15796 15724 -15762
rect 14226 -15808 15724 -15796
rect 14226 -15858 14284 -15808
rect 14226 -16826 14238 -15858
rect 14272 -16826 14284 -15858
rect 15666 -15858 15724 -15808
rect 14226 -16876 14284 -16826
rect 15666 -16826 15678 -15858
rect 15712 -16826 15724 -15858
rect 15666 -16876 15724 -16826
rect 14226 -16888 15724 -16876
rect 14226 -16922 14334 -16888
rect 15616 -16922 15724 -16888
rect 14226 -16934 15724 -16922
rect 15826 -15236 17324 -15224
rect 15826 -15270 15934 -15236
rect 17216 -15270 17324 -15236
rect 15826 -15282 17324 -15270
rect 15826 -15332 15884 -15282
rect 15826 -15700 15838 -15332
rect 15872 -15700 15884 -15332
rect 17266 -15332 17324 -15282
rect 15826 -15750 15884 -15700
rect 17266 -15700 17278 -15332
rect 17312 -15700 17324 -15332
rect 17266 -15750 17324 -15700
rect 15826 -15762 17324 -15750
rect 15826 -15796 15934 -15762
rect 17216 -15796 17324 -15762
rect 15826 -15808 17324 -15796
rect 15826 -15858 15884 -15808
rect 15826 -16826 15838 -15858
rect 15872 -16826 15884 -15858
rect 17266 -15858 17324 -15808
rect 15826 -16876 15884 -16826
rect 17266 -16826 17278 -15858
rect 17312 -16826 17324 -15858
rect 17266 -16876 17324 -16826
rect 15826 -16888 17324 -16876
rect 15826 -16922 15934 -16888
rect 17216 -16922 17324 -16888
rect 15826 -16934 17324 -16922
rect 17426 -15236 18924 -15224
rect 17426 -15270 17534 -15236
rect 18816 -15270 18924 -15236
rect 17426 -15282 18924 -15270
rect 17426 -15332 17484 -15282
rect 17426 -15700 17438 -15332
rect 17472 -15700 17484 -15332
rect 18866 -15332 18924 -15282
rect 17426 -15750 17484 -15700
rect 18866 -15700 18878 -15332
rect 18912 -15700 18924 -15332
rect 18866 -15750 18924 -15700
rect 17426 -15762 18924 -15750
rect 17426 -15796 17534 -15762
rect 18816 -15796 18924 -15762
rect 17426 -15808 18924 -15796
rect 17426 -15858 17484 -15808
rect 17426 -16826 17438 -15858
rect 17472 -16826 17484 -15858
rect 18866 -15858 18924 -15808
rect 17426 -16876 17484 -16826
rect 18866 -16826 18878 -15858
rect 18912 -16826 18924 -15858
rect 18866 -16876 18924 -16826
rect 17426 -16888 18924 -16876
rect 17426 -16922 17534 -16888
rect 18816 -16922 18924 -16888
rect 17426 -16934 18924 -16922
rect 19026 -15236 20524 -15224
rect 19026 -15270 19134 -15236
rect 20416 -15270 20524 -15236
rect 19026 -15282 20524 -15270
rect 19026 -15332 19084 -15282
rect 19026 -15700 19038 -15332
rect 19072 -15700 19084 -15332
rect 20466 -15332 20524 -15282
rect 19026 -15750 19084 -15700
rect 20466 -15700 20478 -15332
rect 20512 -15700 20524 -15332
rect 20466 -15750 20524 -15700
rect 19026 -15762 20524 -15750
rect 19026 -15796 19134 -15762
rect 20416 -15796 20524 -15762
rect 19026 -15808 20524 -15796
rect 19026 -15858 19084 -15808
rect 19026 -16826 19038 -15858
rect 19072 -16826 19084 -15858
rect 20466 -15858 20524 -15808
rect 19026 -16876 19084 -16826
rect 20466 -16826 20478 -15858
rect 20512 -16826 20524 -15858
rect 20466 -16876 20524 -16826
rect 19026 -16888 20524 -16876
rect 19026 -16922 19134 -16888
rect 20416 -16922 20524 -16888
rect 19026 -16934 20524 -16922
rect 20626 -15236 22124 -15224
rect 20626 -15270 20734 -15236
rect 22016 -15270 22124 -15236
rect 20626 -15282 22124 -15270
rect 20626 -15332 20684 -15282
rect 20626 -15700 20638 -15332
rect 20672 -15700 20684 -15332
rect 22066 -15332 22124 -15282
rect 20626 -15750 20684 -15700
rect 22066 -15700 22078 -15332
rect 22112 -15700 22124 -15332
rect 22066 -15750 22124 -15700
rect 20626 -15762 22124 -15750
rect 20626 -15796 20734 -15762
rect 22016 -15796 22124 -15762
rect 20626 -15808 22124 -15796
rect 20626 -15858 20684 -15808
rect 20626 -16826 20638 -15858
rect 20672 -16826 20684 -15858
rect 22066 -15858 22124 -15808
rect 20626 -16876 20684 -16826
rect 22066 -16826 22078 -15858
rect 22112 -16826 22124 -15858
rect 22066 -16876 22124 -16826
rect 20626 -16888 22124 -16876
rect 20626 -16922 20734 -16888
rect 22016 -16922 22124 -16888
rect 20626 -16934 22124 -16922
rect 22226 -15236 23724 -15224
rect 22226 -15270 22334 -15236
rect 23616 -15270 23724 -15236
rect 22226 -15282 23724 -15270
rect 22226 -15332 22284 -15282
rect 22226 -15700 22238 -15332
rect 22272 -15700 22284 -15332
rect 23666 -15332 23724 -15282
rect 22226 -15750 22284 -15700
rect 23666 -15700 23678 -15332
rect 23712 -15700 23724 -15332
rect 23666 -15750 23724 -15700
rect 22226 -15762 23724 -15750
rect 22226 -15796 22334 -15762
rect 23616 -15796 23724 -15762
rect 22226 -15808 23724 -15796
rect 22226 -15858 22284 -15808
rect 22226 -16826 22238 -15858
rect 22272 -16826 22284 -15858
rect 23666 -15858 23724 -15808
rect 22226 -16876 22284 -16826
rect 23666 -16826 23678 -15858
rect 23712 -16826 23724 -15858
rect 23666 -16876 23724 -16826
rect 22226 -16888 23724 -16876
rect 22226 -16922 22334 -16888
rect 23616 -16922 23724 -16888
rect 22226 -16934 23724 -16922
rect 23826 -15236 25324 -15224
rect 23826 -15270 23934 -15236
rect 25216 -15270 25324 -15236
rect 23826 -15282 25324 -15270
rect 23826 -15332 23884 -15282
rect 23826 -15700 23838 -15332
rect 23872 -15700 23884 -15332
rect 25266 -15332 25324 -15282
rect 23826 -15750 23884 -15700
rect 25266 -15700 25278 -15332
rect 25312 -15700 25324 -15332
rect 25266 -15750 25324 -15700
rect 23826 -15762 25324 -15750
rect 23826 -15796 23934 -15762
rect 25216 -15796 25324 -15762
rect 23826 -15808 25324 -15796
rect 23826 -15858 23884 -15808
rect 23826 -16826 23838 -15858
rect 23872 -16826 23884 -15858
rect 25266 -15858 25324 -15808
rect 23826 -16876 23884 -16826
rect 25266 -16826 25278 -15858
rect 25312 -16826 25324 -15858
rect 25266 -16876 25324 -16826
rect 23826 -16888 25324 -16876
rect 23826 -16922 23934 -16888
rect 25216 -16922 25324 -16888
rect 23826 -16934 25324 -16922
rect 25426 -15236 26924 -15224
rect 25426 -15270 25534 -15236
rect 26816 -15270 26924 -15236
rect 25426 -15282 26924 -15270
rect 25426 -15332 25484 -15282
rect 25426 -15700 25438 -15332
rect 25472 -15700 25484 -15332
rect 26866 -15332 26924 -15282
rect 25426 -15750 25484 -15700
rect 26866 -15700 26878 -15332
rect 26912 -15700 26924 -15332
rect 26866 -15750 26924 -15700
rect 25426 -15762 26924 -15750
rect 25426 -15796 25534 -15762
rect 26816 -15796 26924 -15762
rect 25426 -15808 26924 -15796
rect 25426 -15858 25484 -15808
rect 25426 -16826 25438 -15858
rect 25472 -16826 25484 -15858
rect 26866 -15858 26924 -15808
rect 25426 -16876 25484 -16826
rect 26866 -16826 26878 -15858
rect 26912 -16826 26924 -15858
rect 26866 -16876 26924 -16826
rect 25426 -16888 26924 -16876
rect 25426 -16922 25534 -16888
rect 26816 -16922 26924 -16888
rect 25426 -16934 26924 -16922
rect 27026 -15236 28524 -15224
rect 27026 -15270 27134 -15236
rect 28416 -15270 28524 -15236
rect 27026 -15282 28524 -15270
rect 27026 -15332 27084 -15282
rect 27026 -15700 27038 -15332
rect 27072 -15700 27084 -15332
rect 28466 -15332 28524 -15282
rect 27026 -15750 27084 -15700
rect 28466 -15700 28478 -15332
rect 28512 -15700 28524 -15332
rect 28466 -15750 28524 -15700
rect 27026 -15762 28524 -15750
rect 27026 -15796 27134 -15762
rect 28416 -15796 28524 -15762
rect 27026 -15808 28524 -15796
rect 27026 -15858 27084 -15808
rect 27026 -16826 27038 -15858
rect 27072 -16826 27084 -15858
rect 28466 -15858 28524 -15808
rect 27026 -16876 27084 -16826
rect 28466 -16826 28478 -15858
rect 28512 -16826 28524 -15858
rect 28466 -16876 28524 -16826
rect 27026 -16888 28524 -16876
rect 27026 -16922 27134 -16888
rect 28416 -16922 28524 -16888
rect 27026 -16934 28524 -16922
rect 28626 -15236 30124 -15224
rect 28626 -15270 28734 -15236
rect 30016 -15270 30124 -15236
rect 28626 -15282 30124 -15270
rect 28626 -15332 28684 -15282
rect 28626 -15700 28638 -15332
rect 28672 -15700 28684 -15332
rect 30066 -15332 30124 -15282
rect 28626 -15750 28684 -15700
rect 30066 -15700 30078 -15332
rect 30112 -15700 30124 -15332
rect 30066 -15750 30124 -15700
rect 28626 -15762 30124 -15750
rect 28626 -15796 28734 -15762
rect 30016 -15796 30124 -15762
rect 28626 -15808 30124 -15796
rect 28626 -15858 28684 -15808
rect 28626 -16826 28638 -15858
rect 28672 -16826 28684 -15858
rect 30066 -15858 30124 -15808
rect 28626 -16876 28684 -16826
rect 30066 -16826 30078 -15858
rect 30112 -16826 30124 -15858
rect 30066 -16876 30124 -16826
rect 28626 -16888 30124 -16876
rect 28626 -16922 28734 -16888
rect 30016 -16922 30124 -16888
rect 28626 -16934 30124 -16922
rect 30226 -15236 31724 -15224
rect 30226 -15270 30334 -15236
rect 31616 -15270 31724 -15236
rect 30226 -15282 31724 -15270
rect 30226 -15332 30284 -15282
rect 30226 -15700 30238 -15332
rect 30272 -15700 30284 -15332
rect 31666 -15332 31724 -15282
rect 30226 -15750 30284 -15700
rect 31666 -15700 31678 -15332
rect 31712 -15700 31724 -15332
rect 31666 -15750 31724 -15700
rect 30226 -15762 31724 -15750
rect 30226 -15796 30334 -15762
rect 31616 -15796 31724 -15762
rect 30226 -15808 31724 -15796
rect 30226 -15858 30284 -15808
rect 30226 -16826 30238 -15858
rect 30272 -16826 30284 -15858
rect 31666 -15858 31724 -15808
rect 30226 -16876 30284 -16826
rect 31666 -16826 31678 -15858
rect 31712 -16826 31724 -15858
rect 31666 -16876 31724 -16826
rect 30226 -16888 31724 -16876
rect 30226 -16922 30334 -16888
rect 31616 -16922 31724 -16888
rect 30226 -16934 31724 -16922
rect 31826 -15236 33324 -15224
rect 31826 -15270 31934 -15236
rect 33216 -15270 33324 -15236
rect 31826 -15282 33324 -15270
rect 31826 -15332 31884 -15282
rect 31826 -15700 31838 -15332
rect 31872 -15700 31884 -15332
rect 33266 -15332 33324 -15282
rect 31826 -15750 31884 -15700
rect 33266 -15700 33278 -15332
rect 33312 -15700 33324 -15332
rect 33266 -15750 33324 -15700
rect 31826 -15762 33324 -15750
rect 31826 -15796 31934 -15762
rect 33216 -15796 33324 -15762
rect 31826 -15808 33324 -15796
rect 31826 -15858 31884 -15808
rect 31826 -16826 31838 -15858
rect 31872 -16826 31884 -15858
rect 33266 -15858 33324 -15808
rect 31826 -16876 31884 -16826
rect 33266 -16826 33278 -15858
rect 33312 -16826 33324 -15858
rect 33266 -16876 33324 -16826
rect 31826 -16888 33324 -16876
rect 31826 -16922 31934 -16888
rect 33216 -16922 33324 -16888
rect 31826 -16934 33324 -16922
rect 33426 -15236 34924 -15224
rect 33426 -15270 33534 -15236
rect 34816 -15270 34924 -15236
rect 33426 -15282 34924 -15270
rect 33426 -15332 33484 -15282
rect 33426 -15700 33438 -15332
rect 33472 -15700 33484 -15332
rect 34866 -15332 34924 -15282
rect 33426 -15750 33484 -15700
rect 34866 -15700 34878 -15332
rect 34912 -15700 34924 -15332
rect 34866 -15750 34924 -15700
rect 33426 -15762 34924 -15750
rect 33426 -15796 33534 -15762
rect 34816 -15796 34924 -15762
rect 33426 -15808 34924 -15796
rect 33426 -15858 33484 -15808
rect 33426 -16826 33438 -15858
rect 33472 -16826 33484 -15858
rect 34866 -15858 34924 -15808
rect 33426 -16876 33484 -16826
rect 34866 -16826 34878 -15858
rect 34912 -16826 34924 -15858
rect 34866 -16876 34924 -16826
rect 33426 -16888 34924 -16876
rect 33426 -16922 33534 -16888
rect 34816 -16922 34924 -16888
rect 33426 -16934 34924 -16922
rect 35026 -15236 36524 -15224
rect 35026 -15270 35134 -15236
rect 36416 -15270 36524 -15236
rect 35026 -15282 36524 -15270
rect 35026 -15332 35084 -15282
rect 35026 -15700 35038 -15332
rect 35072 -15700 35084 -15332
rect 36466 -15332 36524 -15282
rect 35026 -15750 35084 -15700
rect 36466 -15700 36478 -15332
rect 36512 -15700 36524 -15332
rect 36466 -15750 36524 -15700
rect 35026 -15762 36524 -15750
rect 35026 -15796 35134 -15762
rect 36416 -15796 36524 -15762
rect 35026 -15808 36524 -15796
rect 35026 -15858 35084 -15808
rect 35026 -16826 35038 -15858
rect 35072 -16826 35084 -15858
rect 36466 -15858 36524 -15808
rect 35026 -16876 35084 -16826
rect 36466 -16826 36478 -15858
rect 36512 -16826 36524 -15858
rect 36466 -16876 36524 -16826
rect 35026 -16888 36524 -16876
rect 35026 -16922 35134 -16888
rect 36416 -16922 36524 -16888
rect 35026 -16934 36524 -16922
rect 36626 -15236 38124 -15224
rect 36626 -15270 36734 -15236
rect 38016 -15270 38124 -15236
rect 36626 -15282 38124 -15270
rect 36626 -15332 36684 -15282
rect 36626 -15700 36638 -15332
rect 36672 -15700 36684 -15332
rect 38066 -15332 38124 -15282
rect 36626 -15750 36684 -15700
rect 38066 -15700 38078 -15332
rect 38112 -15700 38124 -15332
rect 38066 -15750 38124 -15700
rect 36626 -15762 38124 -15750
rect 36626 -15796 36734 -15762
rect 38016 -15796 38124 -15762
rect 36626 -15808 38124 -15796
rect 36626 -15858 36684 -15808
rect 36626 -16826 36638 -15858
rect 36672 -16826 36684 -15858
rect 38066 -15858 38124 -15808
rect 36626 -16876 36684 -16826
rect 38066 -16826 38078 -15858
rect 38112 -16826 38124 -15858
rect 38066 -16876 38124 -16826
rect 36626 -16888 38124 -16876
rect 36626 -16922 36734 -16888
rect 38016 -16922 38124 -16888
rect 36626 -16934 38124 -16922
rect -174 -17036 1324 -17024
rect -174 -17070 -66 -17036
rect 1216 -17070 1324 -17036
rect -174 -17082 1324 -17070
rect -174 -17132 -116 -17082
rect -174 -17500 -162 -17132
rect -128 -17500 -116 -17132
rect 1266 -17132 1324 -17082
rect -174 -17550 -116 -17500
rect 1266 -17500 1278 -17132
rect 1312 -17500 1324 -17132
rect 1266 -17550 1324 -17500
rect -174 -17562 1324 -17550
rect -174 -17596 -66 -17562
rect 1216 -17596 1324 -17562
rect -174 -17608 1324 -17596
rect -174 -17658 -116 -17608
rect -174 -18626 -162 -17658
rect -128 -18626 -116 -17658
rect 1266 -17658 1324 -17608
rect -174 -18676 -116 -18626
rect 1266 -18626 1278 -17658
rect 1312 -18626 1324 -17658
rect 1266 -18676 1324 -18626
rect -174 -18688 1324 -18676
rect -174 -18722 -66 -18688
rect 1216 -18722 1324 -18688
rect -174 -18734 1324 -18722
rect 1426 -17036 2924 -17024
rect 1426 -17070 1534 -17036
rect 2816 -17070 2924 -17036
rect 1426 -17082 2924 -17070
rect 1426 -17132 1484 -17082
rect 1426 -17500 1438 -17132
rect 1472 -17500 1484 -17132
rect 2866 -17132 2924 -17082
rect 1426 -17550 1484 -17500
rect 2866 -17500 2878 -17132
rect 2912 -17500 2924 -17132
rect 2866 -17550 2924 -17500
rect 1426 -17562 2924 -17550
rect 1426 -17596 1534 -17562
rect 2816 -17596 2924 -17562
rect 1426 -17608 2924 -17596
rect 1426 -17658 1484 -17608
rect 1426 -18626 1438 -17658
rect 1472 -18626 1484 -17658
rect 2866 -17658 2924 -17608
rect 1426 -18676 1484 -18626
rect 2866 -18626 2878 -17658
rect 2912 -18626 2924 -17658
rect 2866 -18676 2924 -18626
rect 1426 -18688 2924 -18676
rect 1426 -18722 1534 -18688
rect 2816 -18722 2924 -18688
rect 1426 -18734 2924 -18722
rect 3026 -17036 4524 -17024
rect 3026 -17070 3134 -17036
rect 4416 -17070 4524 -17036
rect 3026 -17082 4524 -17070
rect 3026 -17132 3084 -17082
rect 3026 -17500 3038 -17132
rect 3072 -17500 3084 -17132
rect 4466 -17132 4524 -17082
rect 3026 -17550 3084 -17500
rect 4466 -17500 4478 -17132
rect 4512 -17500 4524 -17132
rect 4466 -17550 4524 -17500
rect 3026 -17562 4524 -17550
rect 3026 -17596 3134 -17562
rect 4416 -17596 4524 -17562
rect 3026 -17608 4524 -17596
rect 3026 -17658 3084 -17608
rect 3026 -18626 3038 -17658
rect 3072 -18626 3084 -17658
rect 4466 -17658 4524 -17608
rect 3026 -18676 3084 -18626
rect 4466 -18626 4478 -17658
rect 4512 -18626 4524 -17658
rect 4466 -18676 4524 -18626
rect 3026 -18688 4524 -18676
rect 3026 -18722 3134 -18688
rect 4416 -18722 4524 -18688
rect 3026 -18734 4524 -18722
rect 4626 -17036 6124 -17024
rect 4626 -17070 4734 -17036
rect 6016 -17070 6124 -17036
rect 4626 -17082 6124 -17070
rect 4626 -17132 4684 -17082
rect 4626 -17500 4638 -17132
rect 4672 -17500 4684 -17132
rect 6066 -17132 6124 -17082
rect 4626 -17550 4684 -17500
rect 6066 -17500 6078 -17132
rect 6112 -17500 6124 -17132
rect 6066 -17550 6124 -17500
rect 4626 -17562 6124 -17550
rect 4626 -17596 4734 -17562
rect 6016 -17596 6124 -17562
rect 4626 -17608 6124 -17596
rect 4626 -17658 4684 -17608
rect 4626 -18626 4638 -17658
rect 4672 -18626 4684 -17658
rect 6066 -17658 6124 -17608
rect 4626 -18676 4684 -18626
rect 6066 -18626 6078 -17658
rect 6112 -18626 6124 -17658
rect 6066 -18676 6124 -18626
rect 4626 -18688 6124 -18676
rect 4626 -18722 4734 -18688
rect 6016 -18722 6124 -18688
rect 4626 -18734 6124 -18722
rect 6226 -17036 7724 -17024
rect 6226 -17070 6334 -17036
rect 7616 -17070 7724 -17036
rect 6226 -17082 7724 -17070
rect 6226 -17132 6284 -17082
rect 6226 -17500 6238 -17132
rect 6272 -17500 6284 -17132
rect 7666 -17132 7724 -17082
rect 6226 -17550 6284 -17500
rect 7666 -17500 7678 -17132
rect 7712 -17500 7724 -17132
rect 7666 -17550 7724 -17500
rect 6226 -17562 7724 -17550
rect 6226 -17596 6334 -17562
rect 7616 -17596 7724 -17562
rect 6226 -17608 7724 -17596
rect 6226 -17658 6284 -17608
rect 6226 -18626 6238 -17658
rect 6272 -18626 6284 -17658
rect 7666 -17658 7724 -17608
rect 6226 -18676 6284 -18626
rect 7666 -18626 7678 -17658
rect 7712 -18626 7724 -17658
rect 7666 -18676 7724 -18626
rect 6226 -18688 7724 -18676
rect 6226 -18722 6334 -18688
rect 7616 -18722 7724 -18688
rect 6226 -18734 7724 -18722
rect 7826 -17036 9324 -17024
rect 7826 -17070 7934 -17036
rect 9216 -17070 9324 -17036
rect 7826 -17082 9324 -17070
rect 7826 -17132 7884 -17082
rect 7826 -17500 7838 -17132
rect 7872 -17500 7884 -17132
rect 9266 -17132 9324 -17082
rect 7826 -17550 7884 -17500
rect 9266 -17500 9278 -17132
rect 9312 -17500 9324 -17132
rect 9266 -17550 9324 -17500
rect 7826 -17562 9324 -17550
rect 7826 -17596 7934 -17562
rect 9216 -17596 9324 -17562
rect 7826 -17608 9324 -17596
rect 7826 -17658 7884 -17608
rect 7826 -18626 7838 -17658
rect 7872 -18626 7884 -17658
rect 9266 -17658 9324 -17608
rect 7826 -18676 7884 -18626
rect 9266 -18626 9278 -17658
rect 9312 -18626 9324 -17658
rect 9266 -18676 9324 -18626
rect 7826 -18688 9324 -18676
rect 7826 -18722 7934 -18688
rect 9216 -18722 9324 -18688
rect 7826 -18734 9324 -18722
rect 9426 -17036 10924 -17024
rect 9426 -17070 9534 -17036
rect 10816 -17070 10924 -17036
rect 9426 -17082 10924 -17070
rect 9426 -17132 9484 -17082
rect 9426 -17500 9438 -17132
rect 9472 -17500 9484 -17132
rect 10866 -17132 10924 -17082
rect 9426 -17550 9484 -17500
rect 10866 -17500 10878 -17132
rect 10912 -17500 10924 -17132
rect 10866 -17550 10924 -17500
rect 9426 -17562 10924 -17550
rect 9426 -17596 9534 -17562
rect 10816 -17596 10924 -17562
rect 9426 -17608 10924 -17596
rect 9426 -17658 9484 -17608
rect 9426 -18626 9438 -17658
rect 9472 -18626 9484 -17658
rect 10866 -17658 10924 -17608
rect 9426 -18676 9484 -18626
rect 10866 -18626 10878 -17658
rect 10912 -18626 10924 -17658
rect 10866 -18676 10924 -18626
rect 9426 -18688 10924 -18676
rect 9426 -18722 9534 -18688
rect 10816 -18722 10924 -18688
rect 9426 -18734 10924 -18722
rect 11026 -17036 12524 -17024
rect 11026 -17070 11134 -17036
rect 12416 -17070 12524 -17036
rect 11026 -17082 12524 -17070
rect 11026 -17132 11084 -17082
rect 11026 -17500 11038 -17132
rect 11072 -17500 11084 -17132
rect 12466 -17132 12524 -17082
rect 11026 -17550 11084 -17500
rect 12466 -17500 12478 -17132
rect 12512 -17500 12524 -17132
rect 12466 -17550 12524 -17500
rect 11026 -17562 12524 -17550
rect 11026 -17596 11134 -17562
rect 12416 -17596 12524 -17562
rect 11026 -17608 12524 -17596
rect 11026 -17658 11084 -17608
rect 11026 -18626 11038 -17658
rect 11072 -18626 11084 -17658
rect 12466 -17658 12524 -17608
rect 11026 -18676 11084 -18626
rect 12466 -18626 12478 -17658
rect 12512 -18626 12524 -17658
rect 12466 -18676 12524 -18626
rect 11026 -18688 12524 -18676
rect 11026 -18722 11134 -18688
rect 12416 -18722 12524 -18688
rect 11026 -18734 12524 -18722
rect 12626 -17036 14124 -17024
rect 12626 -17070 12734 -17036
rect 14016 -17070 14124 -17036
rect 12626 -17082 14124 -17070
rect 12626 -17132 12684 -17082
rect 12626 -17500 12638 -17132
rect 12672 -17500 12684 -17132
rect 14066 -17132 14124 -17082
rect 12626 -17550 12684 -17500
rect 14066 -17500 14078 -17132
rect 14112 -17500 14124 -17132
rect 14066 -17550 14124 -17500
rect 12626 -17562 14124 -17550
rect 12626 -17596 12734 -17562
rect 14016 -17596 14124 -17562
rect 12626 -17608 14124 -17596
rect 12626 -17658 12684 -17608
rect 12626 -18626 12638 -17658
rect 12672 -18626 12684 -17658
rect 14066 -17658 14124 -17608
rect 12626 -18676 12684 -18626
rect 14066 -18626 14078 -17658
rect 14112 -18626 14124 -17658
rect 14066 -18676 14124 -18626
rect 12626 -18688 14124 -18676
rect 12626 -18722 12734 -18688
rect 14016 -18722 14124 -18688
rect 12626 -18734 14124 -18722
rect 14226 -17036 15724 -17024
rect 14226 -17070 14334 -17036
rect 15616 -17070 15724 -17036
rect 14226 -17082 15724 -17070
rect 14226 -17132 14284 -17082
rect 14226 -17500 14238 -17132
rect 14272 -17500 14284 -17132
rect 15666 -17132 15724 -17082
rect 14226 -17550 14284 -17500
rect 15666 -17500 15678 -17132
rect 15712 -17500 15724 -17132
rect 15666 -17550 15724 -17500
rect 14226 -17562 15724 -17550
rect 14226 -17596 14334 -17562
rect 15616 -17596 15724 -17562
rect 14226 -17608 15724 -17596
rect 14226 -17658 14284 -17608
rect 14226 -18626 14238 -17658
rect 14272 -18626 14284 -17658
rect 15666 -17658 15724 -17608
rect 14226 -18676 14284 -18626
rect 15666 -18626 15678 -17658
rect 15712 -18626 15724 -17658
rect 15666 -18676 15724 -18626
rect 14226 -18688 15724 -18676
rect 14226 -18722 14334 -18688
rect 15616 -18722 15724 -18688
rect 14226 -18734 15724 -18722
rect 15826 -17036 17324 -17024
rect 15826 -17070 15934 -17036
rect 17216 -17070 17324 -17036
rect 15826 -17082 17324 -17070
rect 15826 -17132 15884 -17082
rect 15826 -17500 15838 -17132
rect 15872 -17500 15884 -17132
rect 17266 -17132 17324 -17082
rect 15826 -17550 15884 -17500
rect 17266 -17500 17278 -17132
rect 17312 -17500 17324 -17132
rect 17266 -17550 17324 -17500
rect 15826 -17562 17324 -17550
rect 15826 -17596 15934 -17562
rect 17216 -17596 17324 -17562
rect 15826 -17608 17324 -17596
rect 15826 -17658 15884 -17608
rect 15826 -18626 15838 -17658
rect 15872 -18626 15884 -17658
rect 17266 -17658 17324 -17608
rect 15826 -18676 15884 -18626
rect 17266 -18626 17278 -17658
rect 17312 -18626 17324 -17658
rect 17266 -18676 17324 -18626
rect 15826 -18688 17324 -18676
rect 15826 -18722 15934 -18688
rect 17216 -18722 17324 -18688
rect 15826 -18734 17324 -18722
rect 17426 -17036 18924 -17024
rect 17426 -17070 17534 -17036
rect 18816 -17070 18924 -17036
rect 17426 -17082 18924 -17070
rect 17426 -17132 17484 -17082
rect 17426 -17500 17438 -17132
rect 17472 -17500 17484 -17132
rect 18866 -17132 18924 -17082
rect 17426 -17550 17484 -17500
rect 18866 -17500 18878 -17132
rect 18912 -17500 18924 -17132
rect 18866 -17550 18924 -17500
rect 17426 -17562 18924 -17550
rect 17426 -17596 17534 -17562
rect 18816 -17596 18924 -17562
rect 17426 -17608 18924 -17596
rect 17426 -17658 17484 -17608
rect 17426 -18626 17438 -17658
rect 17472 -18626 17484 -17658
rect 18866 -17658 18924 -17608
rect 17426 -18676 17484 -18626
rect 18866 -18626 18878 -17658
rect 18912 -18626 18924 -17658
rect 18866 -18676 18924 -18626
rect 17426 -18688 18924 -18676
rect 17426 -18722 17534 -18688
rect 18816 -18722 18924 -18688
rect 17426 -18734 18924 -18722
rect 19026 -17036 20524 -17024
rect 19026 -17070 19134 -17036
rect 20416 -17070 20524 -17036
rect 19026 -17082 20524 -17070
rect 19026 -17132 19084 -17082
rect 19026 -17500 19038 -17132
rect 19072 -17500 19084 -17132
rect 20466 -17132 20524 -17082
rect 19026 -17550 19084 -17500
rect 20466 -17500 20478 -17132
rect 20512 -17500 20524 -17132
rect 20466 -17550 20524 -17500
rect 19026 -17562 20524 -17550
rect 19026 -17596 19134 -17562
rect 20416 -17596 20524 -17562
rect 19026 -17608 20524 -17596
rect 19026 -17658 19084 -17608
rect 19026 -18626 19038 -17658
rect 19072 -18626 19084 -17658
rect 20466 -17658 20524 -17608
rect 19026 -18676 19084 -18626
rect 20466 -18626 20478 -17658
rect 20512 -18626 20524 -17658
rect 20466 -18676 20524 -18626
rect 19026 -18688 20524 -18676
rect 19026 -18722 19134 -18688
rect 20416 -18722 20524 -18688
rect 19026 -18734 20524 -18722
rect 20626 -17036 22124 -17024
rect 20626 -17070 20734 -17036
rect 22016 -17070 22124 -17036
rect 20626 -17082 22124 -17070
rect 20626 -17132 20684 -17082
rect 20626 -17500 20638 -17132
rect 20672 -17500 20684 -17132
rect 22066 -17132 22124 -17082
rect 20626 -17550 20684 -17500
rect 22066 -17500 22078 -17132
rect 22112 -17500 22124 -17132
rect 22066 -17550 22124 -17500
rect 20626 -17562 22124 -17550
rect 20626 -17596 20734 -17562
rect 22016 -17596 22124 -17562
rect 20626 -17608 22124 -17596
rect 20626 -17658 20684 -17608
rect 20626 -18626 20638 -17658
rect 20672 -18626 20684 -17658
rect 22066 -17658 22124 -17608
rect 20626 -18676 20684 -18626
rect 22066 -18626 22078 -17658
rect 22112 -18626 22124 -17658
rect 22066 -18676 22124 -18626
rect 20626 -18688 22124 -18676
rect 20626 -18722 20734 -18688
rect 22016 -18722 22124 -18688
rect 20626 -18734 22124 -18722
rect 22226 -17036 23724 -17024
rect 22226 -17070 22334 -17036
rect 23616 -17070 23724 -17036
rect 22226 -17082 23724 -17070
rect 22226 -17132 22284 -17082
rect 22226 -17500 22238 -17132
rect 22272 -17500 22284 -17132
rect 23666 -17132 23724 -17082
rect 22226 -17550 22284 -17500
rect 23666 -17500 23678 -17132
rect 23712 -17500 23724 -17132
rect 23666 -17550 23724 -17500
rect 22226 -17562 23724 -17550
rect 22226 -17596 22334 -17562
rect 23616 -17596 23724 -17562
rect 22226 -17608 23724 -17596
rect 22226 -17658 22284 -17608
rect 22226 -18626 22238 -17658
rect 22272 -18626 22284 -17658
rect 23666 -17658 23724 -17608
rect 22226 -18676 22284 -18626
rect 23666 -18626 23678 -17658
rect 23712 -18626 23724 -17658
rect 23666 -18676 23724 -18626
rect 22226 -18688 23724 -18676
rect 22226 -18722 22334 -18688
rect 23616 -18722 23724 -18688
rect 22226 -18734 23724 -18722
rect 23826 -17036 25324 -17024
rect 23826 -17070 23934 -17036
rect 25216 -17070 25324 -17036
rect 23826 -17082 25324 -17070
rect 23826 -17132 23884 -17082
rect 23826 -17500 23838 -17132
rect 23872 -17500 23884 -17132
rect 25266 -17132 25324 -17082
rect 23826 -17550 23884 -17500
rect 25266 -17500 25278 -17132
rect 25312 -17500 25324 -17132
rect 25266 -17550 25324 -17500
rect 23826 -17562 25324 -17550
rect 23826 -17596 23934 -17562
rect 25216 -17596 25324 -17562
rect 23826 -17608 25324 -17596
rect 23826 -17658 23884 -17608
rect 23826 -18626 23838 -17658
rect 23872 -18626 23884 -17658
rect 25266 -17658 25324 -17608
rect 23826 -18676 23884 -18626
rect 25266 -18626 25278 -17658
rect 25312 -18626 25324 -17658
rect 25266 -18676 25324 -18626
rect 23826 -18688 25324 -18676
rect 23826 -18722 23934 -18688
rect 25216 -18722 25324 -18688
rect 23826 -18734 25324 -18722
rect 25426 -17036 26924 -17024
rect 25426 -17070 25534 -17036
rect 26816 -17070 26924 -17036
rect 25426 -17082 26924 -17070
rect 25426 -17132 25484 -17082
rect 25426 -17500 25438 -17132
rect 25472 -17500 25484 -17132
rect 26866 -17132 26924 -17082
rect 25426 -17550 25484 -17500
rect 26866 -17500 26878 -17132
rect 26912 -17500 26924 -17132
rect 26866 -17550 26924 -17500
rect 25426 -17562 26924 -17550
rect 25426 -17596 25534 -17562
rect 26816 -17596 26924 -17562
rect 25426 -17608 26924 -17596
rect 25426 -17658 25484 -17608
rect 25426 -18626 25438 -17658
rect 25472 -18626 25484 -17658
rect 26866 -17658 26924 -17608
rect 25426 -18676 25484 -18626
rect 26866 -18626 26878 -17658
rect 26912 -18626 26924 -17658
rect 26866 -18676 26924 -18626
rect 25426 -18688 26924 -18676
rect 25426 -18722 25534 -18688
rect 26816 -18722 26924 -18688
rect 25426 -18734 26924 -18722
rect 27026 -17036 28524 -17024
rect 27026 -17070 27134 -17036
rect 28416 -17070 28524 -17036
rect 27026 -17082 28524 -17070
rect 27026 -17132 27084 -17082
rect 27026 -17500 27038 -17132
rect 27072 -17500 27084 -17132
rect 28466 -17132 28524 -17082
rect 27026 -17550 27084 -17500
rect 28466 -17500 28478 -17132
rect 28512 -17500 28524 -17132
rect 28466 -17550 28524 -17500
rect 27026 -17562 28524 -17550
rect 27026 -17596 27134 -17562
rect 28416 -17596 28524 -17562
rect 27026 -17608 28524 -17596
rect 27026 -17658 27084 -17608
rect 27026 -18626 27038 -17658
rect 27072 -18626 27084 -17658
rect 28466 -17658 28524 -17608
rect 27026 -18676 27084 -18626
rect 28466 -18626 28478 -17658
rect 28512 -18626 28524 -17658
rect 28466 -18676 28524 -18626
rect 27026 -18688 28524 -18676
rect 27026 -18722 27134 -18688
rect 28416 -18722 28524 -18688
rect 27026 -18734 28524 -18722
rect 28626 -17036 30124 -17024
rect 28626 -17070 28734 -17036
rect 30016 -17070 30124 -17036
rect 28626 -17082 30124 -17070
rect 28626 -17132 28684 -17082
rect 28626 -17500 28638 -17132
rect 28672 -17500 28684 -17132
rect 30066 -17132 30124 -17082
rect 28626 -17550 28684 -17500
rect 30066 -17500 30078 -17132
rect 30112 -17500 30124 -17132
rect 30066 -17550 30124 -17500
rect 28626 -17562 30124 -17550
rect 28626 -17596 28734 -17562
rect 30016 -17596 30124 -17562
rect 28626 -17608 30124 -17596
rect 28626 -17658 28684 -17608
rect 28626 -18626 28638 -17658
rect 28672 -18626 28684 -17658
rect 30066 -17658 30124 -17608
rect 28626 -18676 28684 -18626
rect 30066 -18626 30078 -17658
rect 30112 -18626 30124 -17658
rect 30066 -18676 30124 -18626
rect 28626 -18688 30124 -18676
rect 28626 -18722 28734 -18688
rect 30016 -18722 30124 -18688
rect 28626 -18734 30124 -18722
rect 30226 -17036 31724 -17024
rect 30226 -17070 30334 -17036
rect 31616 -17070 31724 -17036
rect 30226 -17082 31724 -17070
rect 30226 -17132 30284 -17082
rect 30226 -17500 30238 -17132
rect 30272 -17500 30284 -17132
rect 31666 -17132 31724 -17082
rect 30226 -17550 30284 -17500
rect 31666 -17500 31678 -17132
rect 31712 -17500 31724 -17132
rect 31666 -17550 31724 -17500
rect 30226 -17562 31724 -17550
rect 30226 -17596 30334 -17562
rect 31616 -17596 31724 -17562
rect 30226 -17608 31724 -17596
rect 30226 -17658 30284 -17608
rect 30226 -18626 30238 -17658
rect 30272 -18626 30284 -17658
rect 31666 -17658 31724 -17608
rect 30226 -18676 30284 -18626
rect 31666 -18626 31678 -17658
rect 31712 -18626 31724 -17658
rect 31666 -18676 31724 -18626
rect 30226 -18688 31724 -18676
rect 30226 -18722 30334 -18688
rect 31616 -18722 31724 -18688
rect 30226 -18734 31724 -18722
rect 31826 -17036 33324 -17024
rect 31826 -17070 31934 -17036
rect 33216 -17070 33324 -17036
rect 31826 -17082 33324 -17070
rect 31826 -17132 31884 -17082
rect 31826 -17500 31838 -17132
rect 31872 -17500 31884 -17132
rect 33266 -17132 33324 -17082
rect 31826 -17550 31884 -17500
rect 33266 -17500 33278 -17132
rect 33312 -17500 33324 -17132
rect 33266 -17550 33324 -17500
rect 31826 -17562 33324 -17550
rect 31826 -17596 31934 -17562
rect 33216 -17596 33324 -17562
rect 31826 -17608 33324 -17596
rect 31826 -17658 31884 -17608
rect 31826 -18626 31838 -17658
rect 31872 -18626 31884 -17658
rect 33266 -17658 33324 -17608
rect 31826 -18676 31884 -18626
rect 33266 -18626 33278 -17658
rect 33312 -18626 33324 -17658
rect 33266 -18676 33324 -18626
rect 31826 -18688 33324 -18676
rect 31826 -18722 31934 -18688
rect 33216 -18722 33324 -18688
rect 31826 -18734 33324 -18722
rect 33426 -17036 34924 -17024
rect 33426 -17070 33534 -17036
rect 34816 -17070 34924 -17036
rect 33426 -17082 34924 -17070
rect 33426 -17132 33484 -17082
rect 33426 -17500 33438 -17132
rect 33472 -17500 33484 -17132
rect 34866 -17132 34924 -17082
rect 33426 -17550 33484 -17500
rect 34866 -17500 34878 -17132
rect 34912 -17500 34924 -17132
rect 34866 -17550 34924 -17500
rect 33426 -17562 34924 -17550
rect 33426 -17596 33534 -17562
rect 34816 -17596 34924 -17562
rect 33426 -17608 34924 -17596
rect 33426 -17658 33484 -17608
rect 33426 -18626 33438 -17658
rect 33472 -18626 33484 -17658
rect 34866 -17658 34924 -17608
rect 33426 -18676 33484 -18626
rect 34866 -18626 34878 -17658
rect 34912 -18626 34924 -17658
rect 34866 -18676 34924 -18626
rect 33426 -18688 34924 -18676
rect 33426 -18722 33534 -18688
rect 34816 -18722 34924 -18688
rect 33426 -18734 34924 -18722
rect 35026 -17036 36524 -17024
rect 35026 -17070 35134 -17036
rect 36416 -17070 36524 -17036
rect 35026 -17082 36524 -17070
rect 35026 -17132 35084 -17082
rect 35026 -17500 35038 -17132
rect 35072 -17500 35084 -17132
rect 36466 -17132 36524 -17082
rect 35026 -17550 35084 -17500
rect 36466 -17500 36478 -17132
rect 36512 -17500 36524 -17132
rect 36466 -17550 36524 -17500
rect 35026 -17562 36524 -17550
rect 35026 -17596 35134 -17562
rect 36416 -17596 36524 -17562
rect 35026 -17608 36524 -17596
rect 35026 -17658 35084 -17608
rect 35026 -18626 35038 -17658
rect 35072 -18626 35084 -17658
rect 36466 -17658 36524 -17608
rect 35026 -18676 35084 -18626
rect 36466 -18626 36478 -17658
rect 36512 -18626 36524 -17658
rect 36466 -18676 36524 -18626
rect 35026 -18688 36524 -18676
rect 35026 -18722 35134 -18688
rect 36416 -18722 36524 -18688
rect 35026 -18734 36524 -18722
rect 36626 -17036 38124 -17024
rect 36626 -17070 36734 -17036
rect 38016 -17070 38124 -17036
rect 36626 -17082 38124 -17070
rect 36626 -17132 36684 -17082
rect 36626 -17500 36638 -17132
rect 36672 -17500 36684 -17132
rect 38066 -17132 38124 -17082
rect 36626 -17550 36684 -17500
rect 38066 -17500 38078 -17132
rect 38112 -17500 38124 -17132
rect 38066 -17550 38124 -17500
rect 36626 -17562 38124 -17550
rect 36626 -17596 36734 -17562
rect 38016 -17596 38124 -17562
rect 36626 -17608 38124 -17596
rect 36626 -17658 36684 -17608
rect 36626 -18626 36638 -17658
rect 36672 -18626 36684 -17658
rect 38066 -17658 38124 -17608
rect 36626 -18676 36684 -18626
rect 38066 -18626 38078 -17658
rect 38112 -18626 38124 -17658
rect 38066 -18676 38124 -18626
rect 36626 -18688 38124 -18676
rect 36626 -18722 36734 -18688
rect 38016 -18722 38124 -18688
rect 36626 -18734 38124 -18722
rect -174 -18836 1324 -18824
rect -174 -18870 -66 -18836
rect 1216 -18870 1324 -18836
rect -174 -18882 1324 -18870
rect -174 -18932 -116 -18882
rect -174 -19300 -162 -18932
rect -128 -19300 -116 -18932
rect 1266 -18932 1324 -18882
rect -174 -19350 -116 -19300
rect 1266 -19300 1278 -18932
rect 1312 -19300 1324 -18932
rect 1266 -19350 1324 -19300
rect -174 -19362 1324 -19350
rect -174 -19396 -66 -19362
rect 1216 -19396 1324 -19362
rect -174 -19408 1324 -19396
rect -174 -19458 -116 -19408
rect -174 -20426 -162 -19458
rect -128 -20426 -116 -19458
rect 1266 -19458 1324 -19408
rect -174 -20476 -116 -20426
rect 1266 -20426 1278 -19458
rect 1312 -20426 1324 -19458
rect 1266 -20476 1324 -20426
rect -174 -20488 1324 -20476
rect -174 -20522 -66 -20488
rect 1216 -20522 1324 -20488
rect -174 -20534 1324 -20522
rect 1426 -18836 2924 -18824
rect 1426 -18870 1534 -18836
rect 2816 -18870 2924 -18836
rect 1426 -18882 2924 -18870
rect 1426 -18932 1484 -18882
rect 1426 -19300 1438 -18932
rect 1472 -19300 1484 -18932
rect 2866 -18932 2924 -18882
rect 1426 -19350 1484 -19300
rect 2866 -19300 2878 -18932
rect 2912 -19300 2924 -18932
rect 2866 -19350 2924 -19300
rect 1426 -19362 2924 -19350
rect 1426 -19396 1534 -19362
rect 2816 -19396 2924 -19362
rect 1426 -19408 2924 -19396
rect 1426 -19458 1484 -19408
rect 1426 -20426 1438 -19458
rect 1472 -20426 1484 -19458
rect 2866 -19458 2924 -19408
rect 1426 -20476 1484 -20426
rect 2866 -20426 2878 -19458
rect 2912 -20426 2924 -19458
rect 2866 -20476 2924 -20426
rect 1426 -20488 2924 -20476
rect 1426 -20522 1534 -20488
rect 2816 -20522 2924 -20488
rect 1426 -20534 2924 -20522
rect 3026 -18836 4524 -18824
rect 3026 -18870 3134 -18836
rect 4416 -18870 4524 -18836
rect 3026 -18882 4524 -18870
rect 3026 -18932 3084 -18882
rect 3026 -19300 3038 -18932
rect 3072 -19300 3084 -18932
rect 4466 -18932 4524 -18882
rect 3026 -19350 3084 -19300
rect 4466 -19300 4478 -18932
rect 4512 -19300 4524 -18932
rect 4466 -19350 4524 -19300
rect 3026 -19362 4524 -19350
rect 3026 -19396 3134 -19362
rect 4416 -19396 4524 -19362
rect 3026 -19408 4524 -19396
rect 3026 -19458 3084 -19408
rect 3026 -20426 3038 -19458
rect 3072 -20426 3084 -19458
rect 4466 -19458 4524 -19408
rect 3026 -20476 3084 -20426
rect 4466 -20426 4478 -19458
rect 4512 -20426 4524 -19458
rect 4466 -20476 4524 -20426
rect 3026 -20488 4524 -20476
rect 3026 -20522 3134 -20488
rect 4416 -20522 4524 -20488
rect 3026 -20534 4524 -20522
rect 4626 -18836 6124 -18824
rect 4626 -18870 4734 -18836
rect 6016 -18870 6124 -18836
rect 4626 -18882 6124 -18870
rect 4626 -18932 4684 -18882
rect 4626 -19300 4638 -18932
rect 4672 -19300 4684 -18932
rect 6066 -18932 6124 -18882
rect 4626 -19350 4684 -19300
rect 6066 -19300 6078 -18932
rect 6112 -19300 6124 -18932
rect 6066 -19350 6124 -19300
rect 4626 -19362 6124 -19350
rect 4626 -19396 4734 -19362
rect 6016 -19396 6124 -19362
rect 4626 -19408 6124 -19396
rect 4626 -19458 4684 -19408
rect 4626 -20426 4638 -19458
rect 4672 -20426 4684 -19458
rect 6066 -19458 6124 -19408
rect 4626 -20476 4684 -20426
rect 6066 -20426 6078 -19458
rect 6112 -20426 6124 -19458
rect 6066 -20476 6124 -20426
rect 4626 -20488 6124 -20476
rect 4626 -20522 4734 -20488
rect 6016 -20522 6124 -20488
rect 4626 -20534 6124 -20522
rect 6226 -18836 7724 -18824
rect 6226 -18870 6334 -18836
rect 7616 -18870 7724 -18836
rect 6226 -18882 7724 -18870
rect 6226 -18932 6284 -18882
rect 6226 -19300 6238 -18932
rect 6272 -19300 6284 -18932
rect 7666 -18932 7724 -18882
rect 6226 -19350 6284 -19300
rect 7666 -19300 7678 -18932
rect 7712 -19300 7724 -18932
rect 7666 -19350 7724 -19300
rect 6226 -19362 7724 -19350
rect 6226 -19396 6334 -19362
rect 7616 -19396 7724 -19362
rect 6226 -19408 7724 -19396
rect 6226 -19458 6284 -19408
rect 6226 -20426 6238 -19458
rect 6272 -20426 6284 -19458
rect 7666 -19458 7724 -19408
rect 6226 -20476 6284 -20426
rect 7666 -20426 7678 -19458
rect 7712 -20426 7724 -19458
rect 7666 -20476 7724 -20426
rect 6226 -20488 7724 -20476
rect 6226 -20522 6334 -20488
rect 7616 -20522 7724 -20488
rect 6226 -20534 7724 -20522
rect 7826 -18836 9324 -18824
rect 7826 -18870 7934 -18836
rect 9216 -18870 9324 -18836
rect 7826 -18882 9324 -18870
rect 7826 -18932 7884 -18882
rect 7826 -19300 7838 -18932
rect 7872 -19300 7884 -18932
rect 9266 -18932 9324 -18882
rect 7826 -19350 7884 -19300
rect 9266 -19300 9278 -18932
rect 9312 -19300 9324 -18932
rect 9266 -19350 9324 -19300
rect 7826 -19362 9324 -19350
rect 7826 -19396 7934 -19362
rect 9216 -19396 9324 -19362
rect 7826 -19408 9324 -19396
rect 7826 -19458 7884 -19408
rect 7826 -20426 7838 -19458
rect 7872 -20426 7884 -19458
rect 9266 -19458 9324 -19408
rect 7826 -20476 7884 -20426
rect 9266 -20426 9278 -19458
rect 9312 -20426 9324 -19458
rect 9266 -20476 9324 -20426
rect 7826 -20488 9324 -20476
rect 7826 -20522 7934 -20488
rect 9216 -20522 9324 -20488
rect 7826 -20534 9324 -20522
rect 9426 -18836 10924 -18824
rect 9426 -18870 9534 -18836
rect 10816 -18870 10924 -18836
rect 9426 -18882 10924 -18870
rect 9426 -18932 9484 -18882
rect 9426 -19300 9438 -18932
rect 9472 -19300 9484 -18932
rect 10866 -18932 10924 -18882
rect 9426 -19350 9484 -19300
rect 10866 -19300 10878 -18932
rect 10912 -19300 10924 -18932
rect 10866 -19350 10924 -19300
rect 9426 -19362 10924 -19350
rect 9426 -19396 9534 -19362
rect 10816 -19396 10924 -19362
rect 9426 -19408 10924 -19396
rect 9426 -19458 9484 -19408
rect 9426 -20426 9438 -19458
rect 9472 -20426 9484 -19458
rect 10866 -19458 10924 -19408
rect 9426 -20476 9484 -20426
rect 10866 -20426 10878 -19458
rect 10912 -20426 10924 -19458
rect 10866 -20476 10924 -20426
rect 9426 -20488 10924 -20476
rect 9426 -20522 9534 -20488
rect 10816 -20522 10924 -20488
rect 9426 -20534 10924 -20522
rect 11026 -18836 12524 -18824
rect 11026 -18870 11134 -18836
rect 12416 -18870 12524 -18836
rect 11026 -18882 12524 -18870
rect 11026 -18932 11084 -18882
rect 11026 -19300 11038 -18932
rect 11072 -19300 11084 -18932
rect 12466 -18932 12524 -18882
rect 11026 -19350 11084 -19300
rect 12466 -19300 12478 -18932
rect 12512 -19300 12524 -18932
rect 12466 -19350 12524 -19300
rect 11026 -19362 12524 -19350
rect 11026 -19396 11134 -19362
rect 12416 -19396 12524 -19362
rect 11026 -19408 12524 -19396
rect 11026 -19458 11084 -19408
rect 11026 -20426 11038 -19458
rect 11072 -20426 11084 -19458
rect 12466 -19458 12524 -19408
rect 11026 -20476 11084 -20426
rect 12466 -20426 12478 -19458
rect 12512 -20426 12524 -19458
rect 12466 -20476 12524 -20426
rect 11026 -20488 12524 -20476
rect 11026 -20522 11134 -20488
rect 12416 -20522 12524 -20488
rect 11026 -20534 12524 -20522
rect 12626 -18836 14124 -18824
rect 12626 -18870 12734 -18836
rect 14016 -18870 14124 -18836
rect 12626 -18882 14124 -18870
rect 12626 -18932 12684 -18882
rect 12626 -19300 12638 -18932
rect 12672 -19300 12684 -18932
rect 14066 -18932 14124 -18882
rect 12626 -19350 12684 -19300
rect 14066 -19300 14078 -18932
rect 14112 -19300 14124 -18932
rect 14066 -19350 14124 -19300
rect 12626 -19362 14124 -19350
rect 12626 -19396 12734 -19362
rect 14016 -19396 14124 -19362
rect 12626 -19408 14124 -19396
rect 12626 -19458 12684 -19408
rect 12626 -20426 12638 -19458
rect 12672 -20426 12684 -19458
rect 14066 -19458 14124 -19408
rect 12626 -20476 12684 -20426
rect 14066 -20426 14078 -19458
rect 14112 -20426 14124 -19458
rect 14066 -20476 14124 -20426
rect 12626 -20488 14124 -20476
rect 12626 -20522 12734 -20488
rect 14016 -20522 14124 -20488
rect 12626 -20534 14124 -20522
rect 14226 -18836 15724 -18824
rect 14226 -18870 14334 -18836
rect 15616 -18870 15724 -18836
rect 14226 -18882 15724 -18870
rect 14226 -18932 14284 -18882
rect 14226 -19300 14238 -18932
rect 14272 -19300 14284 -18932
rect 15666 -18932 15724 -18882
rect 14226 -19350 14284 -19300
rect 15666 -19300 15678 -18932
rect 15712 -19300 15724 -18932
rect 15666 -19350 15724 -19300
rect 14226 -19362 15724 -19350
rect 14226 -19396 14334 -19362
rect 15616 -19396 15724 -19362
rect 14226 -19408 15724 -19396
rect 14226 -19458 14284 -19408
rect 14226 -20426 14238 -19458
rect 14272 -20426 14284 -19458
rect 15666 -19458 15724 -19408
rect 14226 -20476 14284 -20426
rect 15666 -20426 15678 -19458
rect 15712 -20426 15724 -19458
rect 15666 -20476 15724 -20426
rect 14226 -20488 15724 -20476
rect 14226 -20522 14334 -20488
rect 15616 -20522 15724 -20488
rect 14226 -20534 15724 -20522
rect 15826 -18836 17324 -18824
rect 15826 -18870 15934 -18836
rect 17216 -18870 17324 -18836
rect 15826 -18882 17324 -18870
rect 15826 -18932 15884 -18882
rect 15826 -19300 15838 -18932
rect 15872 -19300 15884 -18932
rect 17266 -18932 17324 -18882
rect 15826 -19350 15884 -19300
rect 17266 -19300 17278 -18932
rect 17312 -19300 17324 -18932
rect 17266 -19350 17324 -19300
rect 15826 -19362 17324 -19350
rect 15826 -19396 15934 -19362
rect 17216 -19396 17324 -19362
rect 15826 -19408 17324 -19396
rect 15826 -19458 15884 -19408
rect 15826 -20426 15838 -19458
rect 15872 -20426 15884 -19458
rect 17266 -19458 17324 -19408
rect 15826 -20476 15884 -20426
rect 17266 -20426 17278 -19458
rect 17312 -20426 17324 -19458
rect 17266 -20476 17324 -20426
rect 15826 -20488 17324 -20476
rect 15826 -20522 15934 -20488
rect 17216 -20522 17324 -20488
rect 15826 -20534 17324 -20522
rect 17426 -18836 18924 -18824
rect 17426 -18870 17534 -18836
rect 18816 -18870 18924 -18836
rect 17426 -18882 18924 -18870
rect 17426 -18932 17484 -18882
rect 17426 -19300 17438 -18932
rect 17472 -19300 17484 -18932
rect 18866 -18932 18924 -18882
rect 17426 -19350 17484 -19300
rect 18866 -19300 18878 -18932
rect 18912 -19300 18924 -18932
rect 18866 -19350 18924 -19300
rect 17426 -19362 18924 -19350
rect 17426 -19396 17534 -19362
rect 18816 -19396 18924 -19362
rect 17426 -19408 18924 -19396
rect 17426 -19458 17484 -19408
rect 17426 -20426 17438 -19458
rect 17472 -20426 17484 -19458
rect 18866 -19458 18924 -19408
rect 17426 -20476 17484 -20426
rect 18866 -20426 18878 -19458
rect 18912 -20426 18924 -19458
rect 18866 -20476 18924 -20426
rect 17426 -20488 18924 -20476
rect 17426 -20522 17534 -20488
rect 18816 -20522 18924 -20488
rect 17426 -20534 18924 -20522
rect 19026 -18836 20524 -18824
rect 19026 -18870 19134 -18836
rect 20416 -18870 20524 -18836
rect 19026 -18882 20524 -18870
rect 19026 -18932 19084 -18882
rect 19026 -19300 19038 -18932
rect 19072 -19300 19084 -18932
rect 20466 -18932 20524 -18882
rect 19026 -19350 19084 -19300
rect 20466 -19300 20478 -18932
rect 20512 -19300 20524 -18932
rect 20466 -19350 20524 -19300
rect 19026 -19362 20524 -19350
rect 19026 -19396 19134 -19362
rect 20416 -19396 20524 -19362
rect 19026 -19408 20524 -19396
rect 19026 -19458 19084 -19408
rect 19026 -20426 19038 -19458
rect 19072 -20426 19084 -19458
rect 20466 -19458 20524 -19408
rect 19026 -20476 19084 -20426
rect 20466 -20426 20478 -19458
rect 20512 -20426 20524 -19458
rect 20466 -20476 20524 -20426
rect 19026 -20488 20524 -20476
rect 19026 -20522 19134 -20488
rect 20416 -20522 20524 -20488
rect 19026 -20534 20524 -20522
rect 20626 -18836 22124 -18824
rect 20626 -18870 20734 -18836
rect 22016 -18870 22124 -18836
rect 20626 -18882 22124 -18870
rect 20626 -18932 20684 -18882
rect 20626 -19300 20638 -18932
rect 20672 -19300 20684 -18932
rect 22066 -18932 22124 -18882
rect 20626 -19350 20684 -19300
rect 22066 -19300 22078 -18932
rect 22112 -19300 22124 -18932
rect 22066 -19350 22124 -19300
rect 20626 -19362 22124 -19350
rect 20626 -19396 20734 -19362
rect 22016 -19396 22124 -19362
rect 20626 -19408 22124 -19396
rect 20626 -19458 20684 -19408
rect 20626 -20426 20638 -19458
rect 20672 -20426 20684 -19458
rect 22066 -19458 22124 -19408
rect 20626 -20476 20684 -20426
rect 22066 -20426 22078 -19458
rect 22112 -20426 22124 -19458
rect 22066 -20476 22124 -20426
rect 20626 -20488 22124 -20476
rect 20626 -20522 20734 -20488
rect 22016 -20522 22124 -20488
rect 20626 -20534 22124 -20522
rect 22226 -18836 23724 -18824
rect 22226 -18870 22334 -18836
rect 23616 -18870 23724 -18836
rect 22226 -18882 23724 -18870
rect 22226 -18932 22284 -18882
rect 22226 -19300 22238 -18932
rect 22272 -19300 22284 -18932
rect 23666 -18932 23724 -18882
rect 22226 -19350 22284 -19300
rect 23666 -19300 23678 -18932
rect 23712 -19300 23724 -18932
rect 23666 -19350 23724 -19300
rect 22226 -19362 23724 -19350
rect 22226 -19396 22334 -19362
rect 23616 -19396 23724 -19362
rect 22226 -19408 23724 -19396
rect 22226 -19458 22284 -19408
rect 22226 -20426 22238 -19458
rect 22272 -20426 22284 -19458
rect 23666 -19458 23724 -19408
rect 22226 -20476 22284 -20426
rect 23666 -20426 23678 -19458
rect 23712 -20426 23724 -19458
rect 23666 -20476 23724 -20426
rect 22226 -20488 23724 -20476
rect 22226 -20522 22334 -20488
rect 23616 -20522 23724 -20488
rect 22226 -20534 23724 -20522
rect 23826 -18836 25324 -18824
rect 23826 -18870 23934 -18836
rect 25216 -18870 25324 -18836
rect 23826 -18882 25324 -18870
rect 23826 -18932 23884 -18882
rect 23826 -19300 23838 -18932
rect 23872 -19300 23884 -18932
rect 25266 -18932 25324 -18882
rect 23826 -19350 23884 -19300
rect 25266 -19300 25278 -18932
rect 25312 -19300 25324 -18932
rect 25266 -19350 25324 -19300
rect 23826 -19362 25324 -19350
rect 23826 -19396 23934 -19362
rect 25216 -19396 25324 -19362
rect 23826 -19408 25324 -19396
rect 23826 -19458 23884 -19408
rect 23826 -20426 23838 -19458
rect 23872 -20426 23884 -19458
rect 25266 -19458 25324 -19408
rect 23826 -20476 23884 -20426
rect 25266 -20426 25278 -19458
rect 25312 -20426 25324 -19458
rect 25266 -20476 25324 -20426
rect 23826 -20488 25324 -20476
rect 23826 -20522 23934 -20488
rect 25216 -20522 25324 -20488
rect 23826 -20534 25324 -20522
rect 25426 -18836 26924 -18824
rect 25426 -18870 25534 -18836
rect 26816 -18870 26924 -18836
rect 25426 -18882 26924 -18870
rect 25426 -18932 25484 -18882
rect 25426 -19300 25438 -18932
rect 25472 -19300 25484 -18932
rect 26866 -18932 26924 -18882
rect 25426 -19350 25484 -19300
rect 26866 -19300 26878 -18932
rect 26912 -19300 26924 -18932
rect 26866 -19350 26924 -19300
rect 25426 -19362 26924 -19350
rect 25426 -19396 25534 -19362
rect 26816 -19396 26924 -19362
rect 25426 -19408 26924 -19396
rect 25426 -19458 25484 -19408
rect 25426 -20426 25438 -19458
rect 25472 -20426 25484 -19458
rect 26866 -19458 26924 -19408
rect 25426 -20476 25484 -20426
rect 26866 -20426 26878 -19458
rect 26912 -20426 26924 -19458
rect 26866 -20476 26924 -20426
rect 25426 -20488 26924 -20476
rect 25426 -20522 25534 -20488
rect 26816 -20522 26924 -20488
rect 25426 -20534 26924 -20522
rect 27026 -18836 28524 -18824
rect 27026 -18870 27134 -18836
rect 28416 -18870 28524 -18836
rect 27026 -18882 28524 -18870
rect 27026 -18932 27084 -18882
rect 27026 -19300 27038 -18932
rect 27072 -19300 27084 -18932
rect 28466 -18932 28524 -18882
rect 27026 -19350 27084 -19300
rect 28466 -19300 28478 -18932
rect 28512 -19300 28524 -18932
rect 28466 -19350 28524 -19300
rect 27026 -19362 28524 -19350
rect 27026 -19396 27134 -19362
rect 28416 -19396 28524 -19362
rect 27026 -19408 28524 -19396
rect 27026 -19458 27084 -19408
rect 27026 -20426 27038 -19458
rect 27072 -20426 27084 -19458
rect 28466 -19458 28524 -19408
rect 27026 -20476 27084 -20426
rect 28466 -20426 28478 -19458
rect 28512 -20426 28524 -19458
rect 28466 -20476 28524 -20426
rect 27026 -20488 28524 -20476
rect 27026 -20522 27134 -20488
rect 28416 -20522 28524 -20488
rect 27026 -20534 28524 -20522
rect 28626 -18836 30124 -18824
rect 28626 -18870 28734 -18836
rect 30016 -18870 30124 -18836
rect 28626 -18882 30124 -18870
rect 28626 -18932 28684 -18882
rect 28626 -19300 28638 -18932
rect 28672 -19300 28684 -18932
rect 30066 -18932 30124 -18882
rect 28626 -19350 28684 -19300
rect 30066 -19300 30078 -18932
rect 30112 -19300 30124 -18932
rect 30066 -19350 30124 -19300
rect 28626 -19362 30124 -19350
rect 28626 -19396 28734 -19362
rect 30016 -19396 30124 -19362
rect 28626 -19408 30124 -19396
rect 28626 -19458 28684 -19408
rect 28626 -20426 28638 -19458
rect 28672 -20426 28684 -19458
rect 30066 -19458 30124 -19408
rect 28626 -20476 28684 -20426
rect 30066 -20426 30078 -19458
rect 30112 -20426 30124 -19458
rect 30066 -20476 30124 -20426
rect 28626 -20488 30124 -20476
rect 28626 -20522 28734 -20488
rect 30016 -20522 30124 -20488
rect 28626 -20534 30124 -20522
rect 30226 -18836 31724 -18824
rect 30226 -18870 30334 -18836
rect 31616 -18870 31724 -18836
rect 30226 -18882 31724 -18870
rect 30226 -18932 30284 -18882
rect 30226 -19300 30238 -18932
rect 30272 -19300 30284 -18932
rect 31666 -18932 31724 -18882
rect 30226 -19350 30284 -19300
rect 31666 -19300 31678 -18932
rect 31712 -19300 31724 -18932
rect 31666 -19350 31724 -19300
rect 30226 -19362 31724 -19350
rect 30226 -19396 30334 -19362
rect 31616 -19396 31724 -19362
rect 30226 -19408 31724 -19396
rect 30226 -19458 30284 -19408
rect 30226 -20426 30238 -19458
rect 30272 -20426 30284 -19458
rect 31666 -19458 31724 -19408
rect 30226 -20476 30284 -20426
rect 31666 -20426 31678 -19458
rect 31712 -20426 31724 -19458
rect 31666 -20476 31724 -20426
rect 30226 -20488 31724 -20476
rect 30226 -20522 30334 -20488
rect 31616 -20522 31724 -20488
rect 30226 -20534 31724 -20522
rect 31826 -18836 33324 -18824
rect 31826 -18870 31934 -18836
rect 33216 -18870 33324 -18836
rect 31826 -18882 33324 -18870
rect 31826 -18932 31884 -18882
rect 31826 -19300 31838 -18932
rect 31872 -19300 31884 -18932
rect 33266 -18932 33324 -18882
rect 31826 -19350 31884 -19300
rect 33266 -19300 33278 -18932
rect 33312 -19300 33324 -18932
rect 33266 -19350 33324 -19300
rect 31826 -19362 33324 -19350
rect 31826 -19396 31934 -19362
rect 33216 -19396 33324 -19362
rect 31826 -19408 33324 -19396
rect 31826 -19458 31884 -19408
rect 31826 -20426 31838 -19458
rect 31872 -20426 31884 -19458
rect 33266 -19458 33324 -19408
rect 31826 -20476 31884 -20426
rect 33266 -20426 33278 -19458
rect 33312 -20426 33324 -19458
rect 33266 -20476 33324 -20426
rect 31826 -20488 33324 -20476
rect 31826 -20522 31934 -20488
rect 33216 -20522 33324 -20488
rect 31826 -20534 33324 -20522
rect 33426 -18836 34924 -18824
rect 33426 -18870 33534 -18836
rect 34816 -18870 34924 -18836
rect 33426 -18882 34924 -18870
rect 33426 -18932 33484 -18882
rect 33426 -19300 33438 -18932
rect 33472 -19300 33484 -18932
rect 34866 -18932 34924 -18882
rect 33426 -19350 33484 -19300
rect 34866 -19300 34878 -18932
rect 34912 -19300 34924 -18932
rect 34866 -19350 34924 -19300
rect 33426 -19362 34924 -19350
rect 33426 -19396 33534 -19362
rect 34816 -19396 34924 -19362
rect 33426 -19408 34924 -19396
rect 33426 -19458 33484 -19408
rect 33426 -20426 33438 -19458
rect 33472 -20426 33484 -19458
rect 34866 -19458 34924 -19408
rect 33426 -20476 33484 -20426
rect 34866 -20426 34878 -19458
rect 34912 -20426 34924 -19458
rect 34866 -20476 34924 -20426
rect 33426 -20488 34924 -20476
rect 33426 -20522 33534 -20488
rect 34816 -20522 34924 -20488
rect 33426 -20534 34924 -20522
rect 35026 -18836 36524 -18824
rect 35026 -18870 35134 -18836
rect 36416 -18870 36524 -18836
rect 35026 -18882 36524 -18870
rect 35026 -18932 35084 -18882
rect 35026 -19300 35038 -18932
rect 35072 -19300 35084 -18932
rect 36466 -18932 36524 -18882
rect 35026 -19350 35084 -19300
rect 36466 -19300 36478 -18932
rect 36512 -19300 36524 -18932
rect 36466 -19350 36524 -19300
rect 35026 -19362 36524 -19350
rect 35026 -19396 35134 -19362
rect 36416 -19396 36524 -19362
rect 35026 -19408 36524 -19396
rect 35026 -19458 35084 -19408
rect 35026 -20426 35038 -19458
rect 35072 -20426 35084 -19458
rect 36466 -19458 36524 -19408
rect 35026 -20476 35084 -20426
rect 36466 -20426 36478 -19458
rect 36512 -20426 36524 -19458
rect 36466 -20476 36524 -20426
rect 35026 -20488 36524 -20476
rect 35026 -20522 35134 -20488
rect 36416 -20522 36524 -20488
rect 35026 -20534 36524 -20522
rect 36626 -18836 38124 -18824
rect 36626 -18870 36734 -18836
rect 38016 -18870 38124 -18836
rect 36626 -18882 38124 -18870
rect 36626 -18932 36684 -18882
rect 36626 -19300 36638 -18932
rect 36672 -19300 36684 -18932
rect 38066 -18932 38124 -18882
rect 36626 -19350 36684 -19300
rect 38066 -19300 38078 -18932
rect 38112 -19300 38124 -18932
rect 38066 -19350 38124 -19300
rect 36626 -19362 38124 -19350
rect 36626 -19396 36734 -19362
rect 38016 -19396 38124 -19362
rect 36626 -19408 38124 -19396
rect 36626 -19458 36684 -19408
rect 36626 -20426 36638 -19458
rect 36672 -20426 36684 -19458
rect 38066 -19458 38124 -19408
rect 36626 -20476 36684 -20426
rect 38066 -20426 38078 -19458
rect 38112 -20426 38124 -19458
rect 38066 -20476 38124 -20426
rect 36626 -20488 38124 -20476
rect 36626 -20522 36734 -20488
rect 38016 -20522 38124 -20488
rect 36626 -20534 38124 -20522
rect -174 -20636 1324 -20624
rect -174 -20670 -66 -20636
rect 1216 -20670 1324 -20636
rect -174 -20682 1324 -20670
rect -174 -20732 -116 -20682
rect -174 -21100 -162 -20732
rect -128 -21100 -116 -20732
rect 1266 -20732 1324 -20682
rect -174 -21150 -116 -21100
rect 1266 -21100 1278 -20732
rect 1312 -21100 1324 -20732
rect 1266 -21150 1324 -21100
rect -174 -21162 1324 -21150
rect -174 -21196 -66 -21162
rect 1216 -21196 1324 -21162
rect -174 -21208 1324 -21196
rect -174 -21258 -116 -21208
rect -174 -22226 -162 -21258
rect -128 -22226 -116 -21258
rect 1266 -21258 1324 -21208
rect -174 -22276 -116 -22226
rect 1266 -22226 1278 -21258
rect 1312 -22226 1324 -21258
rect 1266 -22276 1324 -22226
rect -174 -22288 1324 -22276
rect -174 -22322 -66 -22288
rect 1216 -22322 1324 -22288
rect -174 -22334 1324 -22322
rect 1426 -20636 2924 -20624
rect 1426 -20670 1534 -20636
rect 2816 -20670 2924 -20636
rect 1426 -20682 2924 -20670
rect 1426 -20732 1484 -20682
rect 1426 -21100 1438 -20732
rect 1472 -21100 1484 -20732
rect 2866 -20732 2924 -20682
rect 1426 -21150 1484 -21100
rect 2866 -21100 2878 -20732
rect 2912 -21100 2924 -20732
rect 2866 -21150 2924 -21100
rect 1426 -21162 2924 -21150
rect 1426 -21196 1534 -21162
rect 2816 -21196 2924 -21162
rect 1426 -21208 2924 -21196
rect 1426 -21258 1484 -21208
rect 1426 -22226 1438 -21258
rect 1472 -22226 1484 -21258
rect 2866 -21258 2924 -21208
rect 1426 -22276 1484 -22226
rect 2866 -22226 2878 -21258
rect 2912 -22226 2924 -21258
rect 2866 -22276 2924 -22226
rect 1426 -22288 2924 -22276
rect 1426 -22322 1534 -22288
rect 2816 -22322 2924 -22288
rect 1426 -22334 2924 -22322
rect 3026 -20636 4524 -20624
rect 3026 -20670 3134 -20636
rect 4416 -20670 4524 -20636
rect 3026 -20682 4524 -20670
rect 3026 -20732 3084 -20682
rect 3026 -21100 3038 -20732
rect 3072 -21100 3084 -20732
rect 4466 -20732 4524 -20682
rect 3026 -21150 3084 -21100
rect 4466 -21100 4478 -20732
rect 4512 -21100 4524 -20732
rect 4466 -21150 4524 -21100
rect 3026 -21162 4524 -21150
rect 3026 -21196 3134 -21162
rect 4416 -21196 4524 -21162
rect 3026 -21208 4524 -21196
rect 3026 -21258 3084 -21208
rect 3026 -22226 3038 -21258
rect 3072 -22226 3084 -21258
rect 4466 -21258 4524 -21208
rect 3026 -22276 3084 -22226
rect 4466 -22226 4478 -21258
rect 4512 -22226 4524 -21258
rect 4466 -22276 4524 -22226
rect 3026 -22288 4524 -22276
rect 3026 -22322 3134 -22288
rect 4416 -22322 4524 -22288
rect 3026 -22334 4524 -22322
rect 4626 -20636 6124 -20624
rect 4626 -20670 4734 -20636
rect 6016 -20670 6124 -20636
rect 4626 -20682 6124 -20670
rect 4626 -20732 4684 -20682
rect 4626 -21100 4638 -20732
rect 4672 -21100 4684 -20732
rect 6066 -20732 6124 -20682
rect 4626 -21150 4684 -21100
rect 6066 -21100 6078 -20732
rect 6112 -21100 6124 -20732
rect 6066 -21150 6124 -21100
rect 4626 -21162 6124 -21150
rect 4626 -21196 4734 -21162
rect 6016 -21196 6124 -21162
rect 4626 -21208 6124 -21196
rect 4626 -21258 4684 -21208
rect 4626 -22226 4638 -21258
rect 4672 -22226 4684 -21258
rect 6066 -21258 6124 -21208
rect 4626 -22276 4684 -22226
rect 6066 -22226 6078 -21258
rect 6112 -22226 6124 -21258
rect 6066 -22276 6124 -22226
rect 4626 -22288 6124 -22276
rect 4626 -22322 4734 -22288
rect 6016 -22322 6124 -22288
rect 4626 -22334 6124 -22322
rect 6226 -20636 7724 -20624
rect 6226 -20670 6334 -20636
rect 7616 -20670 7724 -20636
rect 6226 -20682 7724 -20670
rect 6226 -20732 6284 -20682
rect 6226 -21100 6238 -20732
rect 6272 -21100 6284 -20732
rect 7666 -20732 7724 -20682
rect 6226 -21150 6284 -21100
rect 7666 -21100 7678 -20732
rect 7712 -21100 7724 -20732
rect 7666 -21150 7724 -21100
rect 6226 -21162 7724 -21150
rect 6226 -21196 6334 -21162
rect 7616 -21196 7724 -21162
rect 6226 -21208 7724 -21196
rect 6226 -21258 6284 -21208
rect 6226 -22226 6238 -21258
rect 6272 -22226 6284 -21258
rect 7666 -21258 7724 -21208
rect 6226 -22276 6284 -22226
rect 7666 -22226 7678 -21258
rect 7712 -22226 7724 -21258
rect 7666 -22276 7724 -22226
rect 6226 -22288 7724 -22276
rect 6226 -22322 6334 -22288
rect 7616 -22322 7724 -22288
rect 6226 -22334 7724 -22322
rect 7826 -20636 9324 -20624
rect 7826 -20670 7934 -20636
rect 9216 -20670 9324 -20636
rect 7826 -20682 9324 -20670
rect 7826 -20732 7884 -20682
rect 7826 -21100 7838 -20732
rect 7872 -21100 7884 -20732
rect 9266 -20732 9324 -20682
rect 7826 -21150 7884 -21100
rect 9266 -21100 9278 -20732
rect 9312 -21100 9324 -20732
rect 9266 -21150 9324 -21100
rect 7826 -21162 9324 -21150
rect 7826 -21196 7934 -21162
rect 9216 -21196 9324 -21162
rect 7826 -21208 9324 -21196
rect 7826 -21258 7884 -21208
rect 7826 -22226 7838 -21258
rect 7872 -22226 7884 -21258
rect 9266 -21258 9324 -21208
rect 7826 -22276 7884 -22226
rect 9266 -22226 9278 -21258
rect 9312 -22226 9324 -21258
rect 9266 -22276 9324 -22226
rect 7826 -22288 9324 -22276
rect 7826 -22322 7934 -22288
rect 9216 -22322 9324 -22288
rect 7826 -22334 9324 -22322
rect 9426 -20636 10924 -20624
rect 9426 -20670 9534 -20636
rect 10816 -20670 10924 -20636
rect 9426 -20682 10924 -20670
rect 9426 -20732 9484 -20682
rect 9426 -21100 9438 -20732
rect 9472 -21100 9484 -20732
rect 10866 -20732 10924 -20682
rect 9426 -21150 9484 -21100
rect 10866 -21100 10878 -20732
rect 10912 -21100 10924 -20732
rect 10866 -21150 10924 -21100
rect 9426 -21162 10924 -21150
rect 9426 -21196 9534 -21162
rect 10816 -21196 10924 -21162
rect 9426 -21208 10924 -21196
rect 9426 -21258 9484 -21208
rect 9426 -22226 9438 -21258
rect 9472 -22226 9484 -21258
rect 10866 -21258 10924 -21208
rect 9426 -22276 9484 -22226
rect 10866 -22226 10878 -21258
rect 10912 -22226 10924 -21258
rect 10866 -22276 10924 -22226
rect 9426 -22288 10924 -22276
rect 9426 -22322 9534 -22288
rect 10816 -22322 10924 -22288
rect 9426 -22334 10924 -22322
rect 11026 -20636 12524 -20624
rect 11026 -20670 11134 -20636
rect 12416 -20670 12524 -20636
rect 11026 -20682 12524 -20670
rect 11026 -20732 11084 -20682
rect 11026 -21100 11038 -20732
rect 11072 -21100 11084 -20732
rect 12466 -20732 12524 -20682
rect 11026 -21150 11084 -21100
rect 12466 -21100 12478 -20732
rect 12512 -21100 12524 -20732
rect 12466 -21150 12524 -21100
rect 11026 -21162 12524 -21150
rect 11026 -21196 11134 -21162
rect 12416 -21196 12524 -21162
rect 11026 -21208 12524 -21196
rect 11026 -21258 11084 -21208
rect 11026 -22226 11038 -21258
rect 11072 -22226 11084 -21258
rect 12466 -21258 12524 -21208
rect 11026 -22276 11084 -22226
rect 12466 -22226 12478 -21258
rect 12512 -22226 12524 -21258
rect 12466 -22276 12524 -22226
rect 11026 -22288 12524 -22276
rect 11026 -22322 11134 -22288
rect 12416 -22322 12524 -22288
rect 11026 -22334 12524 -22322
rect 12626 -20636 14124 -20624
rect 12626 -20670 12734 -20636
rect 14016 -20670 14124 -20636
rect 12626 -20682 14124 -20670
rect 12626 -20732 12684 -20682
rect 12626 -21100 12638 -20732
rect 12672 -21100 12684 -20732
rect 14066 -20732 14124 -20682
rect 12626 -21150 12684 -21100
rect 14066 -21100 14078 -20732
rect 14112 -21100 14124 -20732
rect 14066 -21150 14124 -21100
rect 12626 -21162 14124 -21150
rect 12626 -21196 12734 -21162
rect 14016 -21196 14124 -21162
rect 12626 -21208 14124 -21196
rect 12626 -21258 12684 -21208
rect 12626 -22226 12638 -21258
rect 12672 -22226 12684 -21258
rect 14066 -21258 14124 -21208
rect 12626 -22276 12684 -22226
rect 14066 -22226 14078 -21258
rect 14112 -22226 14124 -21258
rect 14066 -22276 14124 -22226
rect 12626 -22288 14124 -22276
rect 12626 -22322 12734 -22288
rect 14016 -22322 14124 -22288
rect 12626 -22334 14124 -22322
rect 14226 -20636 15724 -20624
rect 14226 -20670 14334 -20636
rect 15616 -20670 15724 -20636
rect 14226 -20682 15724 -20670
rect 14226 -20732 14284 -20682
rect 14226 -21100 14238 -20732
rect 14272 -21100 14284 -20732
rect 15666 -20732 15724 -20682
rect 14226 -21150 14284 -21100
rect 15666 -21100 15678 -20732
rect 15712 -21100 15724 -20732
rect 15666 -21150 15724 -21100
rect 14226 -21162 15724 -21150
rect 14226 -21196 14334 -21162
rect 15616 -21196 15724 -21162
rect 14226 -21208 15724 -21196
rect 14226 -21258 14284 -21208
rect 14226 -22226 14238 -21258
rect 14272 -22226 14284 -21258
rect 15666 -21258 15724 -21208
rect 14226 -22276 14284 -22226
rect 15666 -22226 15678 -21258
rect 15712 -22226 15724 -21258
rect 15666 -22276 15724 -22226
rect 14226 -22288 15724 -22276
rect 14226 -22322 14334 -22288
rect 15616 -22322 15724 -22288
rect 14226 -22334 15724 -22322
rect 15826 -20636 17324 -20624
rect 15826 -20670 15934 -20636
rect 17216 -20670 17324 -20636
rect 15826 -20682 17324 -20670
rect 15826 -20732 15884 -20682
rect 15826 -21100 15838 -20732
rect 15872 -21100 15884 -20732
rect 17266 -20732 17324 -20682
rect 15826 -21150 15884 -21100
rect 17266 -21100 17278 -20732
rect 17312 -21100 17324 -20732
rect 17266 -21150 17324 -21100
rect 15826 -21162 17324 -21150
rect 15826 -21196 15934 -21162
rect 17216 -21196 17324 -21162
rect 15826 -21208 17324 -21196
rect 15826 -21258 15884 -21208
rect 15826 -22226 15838 -21258
rect 15872 -22226 15884 -21258
rect 17266 -21258 17324 -21208
rect 15826 -22276 15884 -22226
rect 17266 -22226 17278 -21258
rect 17312 -22226 17324 -21258
rect 17266 -22276 17324 -22226
rect 15826 -22288 17324 -22276
rect 15826 -22322 15934 -22288
rect 17216 -22322 17324 -22288
rect 15826 -22334 17324 -22322
rect 17426 -20636 18924 -20624
rect 17426 -20670 17534 -20636
rect 18816 -20670 18924 -20636
rect 17426 -20682 18924 -20670
rect 17426 -20732 17484 -20682
rect 17426 -21100 17438 -20732
rect 17472 -21100 17484 -20732
rect 18866 -20732 18924 -20682
rect 17426 -21150 17484 -21100
rect 18866 -21100 18878 -20732
rect 18912 -21100 18924 -20732
rect 18866 -21150 18924 -21100
rect 17426 -21162 18924 -21150
rect 17426 -21196 17534 -21162
rect 18816 -21196 18924 -21162
rect 17426 -21208 18924 -21196
rect 17426 -21258 17484 -21208
rect 17426 -22226 17438 -21258
rect 17472 -22226 17484 -21258
rect 18866 -21258 18924 -21208
rect 17426 -22276 17484 -22226
rect 18866 -22226 18878 -21258
rect 18912 -22226 18924 -21258
rect 18866 -22276 18924 -22226
rect 17426 -22288 18924 -22276
rect 17426 -22322 17534 -22288
rect 18816 -22322 18924 -22288
rect 17426 -22334 18924 -22322
rect 19026 -20636 20524 -20624
rect 19026 -20670 19134 -20636
rect 20416 -20670 20524 -20636
rect 19026 -20682 20524 -20670
rect 19026 -20732 19084 -20682
rect 19026 -21100 19038 -20732
rect 19072 -21100 19084 -20732
rect 20466 -20732 20524 -20682
rect 19026 -21150 19084 -21100
rect 20466 -21100 20478 -20732
rect 20512 -21100 20524 -20732
rect 20466 -21150 20524 -21100
rect 19026 -21162 20524 -21150
rect 19026 -21196 19134 -21162
rect 20416 -21196 20524 -21162
rect 19026 -21208 20524 -21196
rect 19026 -21258 19084 -21208
rect 19026 -22226 19038 -21258
rect 19072 -22226 19084 -21258
rect 20466 -21258 20524 -21208
rect 19026 -22276 19084 -22226
rect 20466 -22226 20478 -21258
rect 20512 -22226 20524 -21258
rect 20466 -22276 20524 -22226
rect 19026 -22288 20524 -22276
rect 19026 -22322 19134 -22288
rect 20416 -22322 20524 -22288
rect 19026 -22334 20524 -22322
rect 20626 -20636 22124 -20624
rect 20626 -20670 20734 -20636
rect 22016 -20670 22124 -20636
rect 20626 -20682 22124 -20670
rect 20626 -20732 20684 -20682
rect 20626 -21100 20638 -20732
rect 20672 -21100 20684 -20732
rect 22066 -20732 22124 -20682
rect 20626 -21150 20684 -21100
rect 22066 -21100 22078 -20732
rect 22112 -21100 22124 -20732
rect 22066 -21150 22124 -21100
rect 20626 -21162 22124 -21150
rect 20626 -21196 20734 -21162
rect 22016 -21196 22124 -21162
rect 20626 -21208 22124 -21196
rect 20626 -21258 20684 -21208
rect 20626 -22226 20638 -21258
rect 20672 -22226 20684 -21258
rect 22066 -21258 22124 -21208
rect 20626 -22276 20684 -22226
rect 22066 -22226 22078 -21258
rect 22112 -22226 22124 -21258
rect 22066 -22276 22124 -22226
rect 20626 -22288 22124 -22276
rect 20626 -22322 20734 -22288
rect 22016 -22322 22124 -22288
rect 20626 -22334 22124 -22322
rect 22226 -20636 23724 -20624
rect 22226 -20670 22334 -20636
rect 23616 -20670 23724 -20636
rect 22226 -20682 23724 -20670
rect 22226 -20732 22284 -20682
rect 22226 -21100 22238 -20732
rect 22272 -21100 22284 -20732
rect 23666 -20732 23724 -20682
rect 22226 -21150 22284 -21100
rect 23666 -21100 23678 -20732
rect 23712 -21100 23724 -20732
rect 23666 -21150 23724 -21100
rect 22226 -21162 23724 -21150
rect 22226 -21196 22334 -21162
rect 23616 -21196 23724 -21162
rect 22226 -21208 23724 -21196
rect 22226 -21258 22284 -21208
rect 22226 -22226 22238 -21258
rect 22272 -22226 22284 -21258
rect 23666 -21258 23724 -21208
rect 22226 -22276 22284 -22226
rect 23666 -22226 23678 -21258
rect 23712 -22226 23724 -21258
rect 23666 -22276 23724 -22226
rect 22226 -22288 23724 -22276
rect 22226 -22322 22334 -22288
rect 23616 -22322 23724 -22288
rect 22226 -22334 23724 -22322
rect 23826 -20636 25324 -20624
rect 23826 -20670 23934 -20636
rect 25216 -20670 25324 -20636
rect 23826 -20682 25324 -20670
rect 23826 -20732 23884 -20682
rect 23826 -21100 23838 -20732
rect 23872 -21100 23884 -20732
rect 25266 -20732 25324 -20682
rect 23826 -21150 23884 -21100
rect 25266 -21100 25278 -20732
rect 25312 -21100 25324 -20732
rect 25266 -21150 25324 -21100
rect 23826 -21162 25324 -21150
rect 23826 -21196 23934 -21162
rect 25216 -21196 25324 -21162
rect 23826 -21208 25324 -21196
rect 23826 -21258 23884 -21208
rect 23826 -22226 23838 -21258
rect 23872 -22226 23884 -21258
rect 25266 -21258 25324 -21208
rect 23826 -22276 23884 -22226
rect 25266 -22226 25278 -21258
rect 25312 -22226 25324 -21258
rect 25266 -22276 25324 -22226
rect 23826 -22288 25324 -22276
rect 23826 -22322 23934 -22288
rect 25216 -22322 25324 -22288
rect 23826 -22334 25324 -22322
rect 25426 -20636 26924 -20624
rect 25426 -20670 25534 -20636
rect 26816 -20670 26924 -20636
rect 25426 -20682 26924 -20670
rect 25426 -20732 25484 -20682
rect 25426 -21100 25438 -20732
rect 25472 -21100 25484 -20732
rect 26866 -20732 26924 -20682
rect 25426 -21150 25484 -21100
rect 26866 -21100 26878 -20732
rect 26912 -21100 26924 -20732
rect 26866 -21150 26924 -21100
rect 25426 -21162 26924 -21150
rect 25426 -21196 25534 -21162
rect 26816 -21196 26924 -21162
rect 25426 -21208 26924 -21196
rect 25426 -21258 25484 -21208
rect 25426 -22226 25438 -21258
rect 25472 -22226 25484 -21258
rect 26866 -21258 26924 -21208
rect 25426 -22276 25484 -22226
rect 26866 -22226 26878 -21258
rect 26912 -22226 26924 -21258
rect 26866 -22276 26924 -22226
rect 25426 -22288 26924 -22276
rect 25426 -22322 25534 -22288
rect 26816 -22322 26924 -22288
rect 25426 -22334 26924 -22322
rect 27026 -20636 28524 -20624
rect 27026 -20670 27134 -20636
rect 28416 -20670 28524 -20636
rect 27026 -20682 28524 -20670
rect 27026 -20732 27084 -20682
rect 27026 -21100 27038 -20732
rect 27072 -21100 27084 -20732
rect 28466 -20732 28524 -20682
rect 27026 -21150 27084 -21100
rect 28466 -21100 28478 -20732
rect 28512 -21100 28524 -20732
rect 28466 -21150 28524 -21100
rect 27026 -21162 28524 -21150
rect 27026 -21196 27134 -21162
rect 28416 -21196 28524 -21162
rect 27026 -21208 28524 -21196
rect 27026 -21258 27084 -21208
rect 27026 -22226 27038 -21258
rect 27072 -22226 27084 -21258
rect 28466 -21258 28524 -21208
rect 27026 -22276 27084 -22226
rect 28466 -22226 28478 -21258
rect 28512 -22226 28524 -21258
rect 28466 -22276 28524 -22226
rect 27026 -22288 28524 -22276
rect 27026 -22322 27134 -22288
rect 28416 -22322 28524 -22288
rect 27026 -22334 28524 -22322
rect 28626 -20636 30124 -20624
rect 28626 -20670 28734 -20636
rect 30016 -20670 30124 -20636
rect 28626 -20682 30124 -20670
rect 28626 -20732 28684 -20682
rect 28626 -21100 28638 -20732
rect 28672 -21100 28684 -20732
rect 30066 -20732 30124 -20682
rect 28626 -21150 28684 -21100
rect 30066 -21100 30078 -20732
rect 30112 -21100 30124 -20732
rect 30066 -21150 30124 -21100
rect 28626 -21162 30124 -21150
rect 28626 -21196 28734 -21162
rect 30016 -21196 30124 -21162
rect 28626 -21208 30124 -21196
rect 28626 -21258 28684 -21208
rect 28626 -22226 28638 -21258
rect 28672 -22226 28684 -21258
rect 30066 -21258 30124 -21208
rect 28626 -22276 28684 -22226
rect 30066 -22226 30078 -21258
rect 30112 -22226 30124 -21258
rect 30066 -22276 30124 -22226
rect 28626 -22288 30124 -22276
rect 28626 -22322 28734 -22288
rect 30016 -22322 30124 -22288
rect 28626 -22334 30124 -22322
rect 30226 -20636 31724 -20624
rect 30226 -20670 30334 -20636
rect 31616 -20670 31724 -20636
rect 30226 -20682 31724 -20670
rect 30226 -20732 30284 -20682
rect 30226 -21100 30238 -20732
rect 30272 -21100 30284 -20732
rect 31666 -20732 31724 -20682
rect 30226 -21150 30284 -21100
rect 31666 -21100 31678 -20732
rect 31712 -21100 31724 -20732
rect 31666 -21150 31724 -21100
rect 30226 -21162 31724 -21150
rect 30226 -21196 30334 -21162
rect 31616 -21196 31724 -21162
rect 30226 -21208 31724 -21196
rect 30226 -21258 30284 -21208
rect 30226 -22226 30238 -21258
rect 30272 -22226 30284 -21258
rect 31666 -21258 31724 -21208
rect 30226 -22276 30284 -22226
rect 31666 -22226 31678 -21258
rect 31712 -22226 31724 -21258
rect 31666 -22276 31724 -22226
rect 30226 -22288 31724 -22276
rect 30226 -22322 30334 -22288
rect 31616 -22322 31724 -22288
rect 30226 -22334 31724 -22322
rect 31826 -20636 33324 -20624
rect 31826 -20670 31934 -20636
rect 33216 -20670 33324 -20636
rect 31826 -20682 33324 -20670
rect 31826 -20732 31884 -20682
rect 31826 -21100 31838 -20732
rect 31872 -21100 31884 -20732
rect 33266 -20732 33324 -20682
rect 31826 -21150 31884 -21100
rect 33266 -21100 33278 -20732
rect 33312 -21100 33324 -20732
rect 33266 -21150 33324 -21100
rect 31826 -21162 33324 -21150
rect 31826 -21196 31934 -21162
rect 33216 -21196 33324 -21162
rect 31826 -21208 33324 -21196
rect 31826 -21258 31884 -21208
rect 31826 -22226 31838 -21258
rect 31872 -22226 31884 -21258
rect 33266 -21258 33324 -21208
rect 31826 -22276 31884 -22226
rect 33266 -22226 33278 -21258
rect 33312 -22226 33324 -21258
rect 33266 -22276 33324 -22226
rect 31826 -22288 33324 -22276
rect 31826 -22322 31934 -22288
rect 33216 -22322 33324 -22288
rect 31826 -22334 33324 -22322
rect 33426 -20636 34924 -20624
rect 33426 -20670 33534 -20636
rect 34816 -20670 34924 -20636
rect 33426 -20682 34924 -20670
rect 33426 -20732 33484 -20682
rect 33426 -21100 33438 -20732
rect 33472 -21100 33484 -20732
rect 34866 -20732 34924 -20682
rect 33426 -21150 33484 -21100
rect 34866 -21100 34878 -20732
rect 34912 -21100 34924 -20732
rect 34866 -21150 34924 -21100
rect 33426 -21162 34924 -21150
rect 33426 -21196 33534 -21162
rect 34816 -21196 34924 -21162
rect 33426 -21208 34924 -21196
rect 33426 -21258 33484 -21208
rect 33426 -22226 33438 -21258
rect 33472 -22226 33484 -21258
rect 34866 -21258 34924 -21208
rect 33426 -22276 33484 -22226
rect 34866 -22226 34878 -21258
rect 34912 -22226 34924 -21258
rect 34866 -22276 34924 -22226
rect 33426 -22288 34924 -22276
rect 33426 -22322 33534 -22288
rect 34816 -22322 34924 -22288
rect 33426 -22334 34924 -22322
rect 35026 -20636 36524 -20624
rect 35026 -20670 35134 -20636
rect 36416 -20670 36524 -20636
rect 35026 -20682 36524 -20670
rect 35026 -20732 35084 -20682
rect 35026 -21100 35038 -20732
rect 35072 -21100 35084 -20732
rect 36466 -20732 36524 -20682
rect 35026 -21150 35084 -21100
rect 36466 -21100 36478 -20732
rect 36512 -21100 36524 -20732
rect 36466 -21150 36524 -21100
rect 35026 -21162 36524 -21150
rect 35026 -21196 35134 -21162
rect 36416 -21196 36524 -21162
rect 35026 -21208 36524 -21196
rect 35026 -21258 35084 -21208
rect 35026 -22226 35038 -21258
rect 35072 -22226 35084 -21258
rect 36466 -21258 36524 -21208
rect 35026 -22276 35084 -22226
rect 36466 -22226 36478 -21258
rect 36512 -22226 36524 -21258
rect 36466 -22276 36524 -22226
rect 35026 -22288 36524 -22276
rect 35026 -22322 35134 -22288
rect 36416 -22322 36524 -22288
rect 35026 -22334 36524 -22322
rect 36626 -20636 38124 -20624
rect 36626 -20670 36734 -20636
rect 38016 -20670 38124 -20636
rect 36626 -20682 38124 -20670
rect 36626 -20732 36684 -20682
rect 36626 -21100 36638 -20732
rect 36672 -21100 36684 -20732
rect 38066 -20732 38124 -20682
rect 36626 -21150 36684 -21100
rect 38066 -21100 38078 -20732
rect 38112 -21100 38124 -20732
rect 38066 -21150 38124 -21100
rect 36626 -21162 38124 -21150
rect 36626 -21196 36734 -21162
rect 38016 -21196 38124 -21162
rect 36626 -21208 38124 -21196
rect 36626 -21258 36684 -21208
rect 36626 -22226 36638 -21258
rect 36672 -22226 36684 -21258
rect 38066 -21258 38124 -21208
rect 36626 -22276 36684 -22226
rect 38066 -22226 38078 -21258
rect 38112 -22226 38124 -21258
rect 38066 -22276 38124 -22226
rect 36626 -22288 38124 -22276
rect 36626 -22322 36734 -22288
rect 38016 -22322 38124 -22288
rect 36626 -22334 38124 -22322
rect 32486 -22404 33444 -22392
rect 32486 -22438 32594 -22404
rect 33336 -22438 33444 -22404
rect 32486 -22450 33444 -22438
rect 32486 -22500 32544 -22450
rect 28206 -22524 29164 -22512
rect 28206 -22558 28314 -22524
rect 29056 -22558 29164 -22524
rect 28206 -22570 29164 -22558
rect 28206 -22620 28264 -22570
rect 28206 -23596 28218 -22620
rect 28252 -23596 28264 -22620
rect 29106 -22620 29164 -22570
rect 28206 -23646 28264 -23596
rect 29106 -23596 29118 -22620
rect 29152 -23596 29164 -22620
rect 32486 -23146 32498 -22500
rect 32532 -23146 32544 -22500
rect 33386 -22500 33444 -22450
rect 32486 -23196 32544 -23146
rect 33386 -23146 33398 -22500
rect 33432 -23146 33444 -22500
rect 33386 -23196 33444 -23146
rect 32486 -23208 33444 -23196
rect 32486 -23242 32594 -23208
rect 33336 -23242 33444 -23208
rect 32486 -23254 33444 -23242
rect 33856 -22424 34498 -22412
rect 33856 -22458 33964 -22424
rect 34390 -22458 34498 -22424
rect 33856 -22470 34498 -22458
rect 33856 -22520 33914 -22470
rect 33856 -23166 33868 -22520
rect 33902 -23166 33914 -22520
rect 34440 -22520 34498 -22470
rect 33856 -23216 33914 -23166
rect 34440 -23166 34452 -22520
rect 34486 -23166 34498 -22520
rect 34440 -23216 34498 -23166
rect 33856 -23228 34498 -23216
rect 33856 -23262 33964 -23228
rect 34390 -23262 34498 -23228
rect 33856 -23274 34498 -23262
rect 29106 -23646 29164 -23596
rect 28206 -23658 29164 -23646
rect 28206 -23692 28314 -23658
rect 29056 -23692 29164 -23658
rect 28206 -23704 29164 -23692
rect 33024 -23546 34298 -23534
rect 33024 -23580 33132 -23546
rect 34190 -23580 34298 -23546
rect 33024 -23592 34298 -23580
rect 33024 -23642 33082 -23592
rect 36 -24172 2098 -24160
rect 36 -24206 144 -24172
rect 1990 -24206 2098 -24172
rect 36 -24218 2098 -24206
rect 36 -24268 94 -24218
rect 36 -24736 48 -24268
rect 82 -24736 94 -24268
rect 2040 -24268 2098 -24218
rect 36 -24786 94 -24736
rect 2040 -24736 2052 -24268
rect 2086 -24736 2098 -24268
rect 2040 -24786 2098 -24736
rect 36 -24798 2098 -24786
rect 36 -24832 144 -24798
rect 1990 -24832 2098 -24798
rect 36 -24844 2098 -24832
rect 2236 -24172 4298 -24160
rect 2236 -24206 2344 -24172
rect 4190 -24206 4298 -24172
rect 2236 -24218 4298 -24206
rect 2236 -24268 2294 -24218
rect 2236 -24736 2248 -24268
rect 2282 -24736 2294 -24268
rect 4240 -24268 4298 -24218
rect 2236 -24786 2294 -24736
rect 4240 -24736 4252 -24268
rect 4286 -24736 4298 -24268
rect 4240 -24786 4298 -24736
rect 2236 -24798 4298 -24786
rect 2236 -24832 2344 -24798
rect 4190 -24832 4298 -24798
rect 2236 -24844 4298 -24832
rect 4436 -24172 6498 -24160
rect 4436 -24206 4544 -24172
rect 6390 -24206 6498 -24172
rect 4436 -24218 6498 -24206
rect 4436 -24268 4494 -24218
rect 4436 -24736 4448 -24268
rect 4482 -24736 4494 -24268
rect 6440 -24268 6498 -24218
rect 4436 -24786 4494 -24736
rect 6440 -24736 6452 -24268
rect 6486 -24736 6498 -24268
rect 6440 -24786 6498 -24736
rect 4436 -24798 6498 -24786
rect 4436 -24832 4544 -24798
rect 6390 -24832 6498 -24798
rect 4436 -24844 6498 -24832
rect 6636 -24172 8698 -24160
rect 6636 -24206 6744 -24172
rect 8590 -24206 8698 -24172
rect 6636 -24218 8698 -24206
rect 6636 -24268 6694 -24218
rect 6636 -24736 6648 -24268
rect 6682 -24736 6694 -24268
rect 8640 -24268 8698 -24218
rect 6636 -24786 6694 -24736
rect 8640 -24736 8652 -24268
rect 8686 -24736 8698 -24268
rect 8640 -24786 8698 -24736
rect 6636 -24798 8698 -24786
rect 6636 -24832 6744 -24798
rect 8590 -24832 8698 -24798
rect 6636 -24844 8698 -24832
rect 8836 -24172 10898 -24160
rect 8836 -24206 8944 -24172
rect 10790 -24206 10898 -24172
rect 8836 -24218 10898 -24206
rect 8836 -24268 8894 -24218
rect 8836 -24736 8848 -24268
rect 8882 -24736 8894 -24268
rect 10840 -24268 10898 -24218
rect 8836 -24786 8894 -24736
rect 10840 -24736 10852 -24268
rect 10886 -24736 10898 -24268
rect 10840 -24786 10898 -24736
rect 8836 -24798 10898 -24786
rect 8836 -24832 8944 -24798
rect 10790 -24832 10898 -24798
rect 8836 -24844 10898 -24832
rect 11036 -24172 13098 -24160
rect 11036 -24206 11144 -24172
rect 12990 -24206 13098 -24172
rect 11036 -24218 13098 -24206
rect 11036 -24268 11094 -24218
rect 11036 -24736 11048 -24268
rect 11082 -24736 11094 -24268
rect 13040 -24268 13098 -24218
rect 11036 -24786 11094 -24736
rect 13040 -24736 13052 -24268
rect 13086 -24736 13098 -24268
rect 13040 -24786 13098 -24736
rect 11036 -24798 13098 -24786
rect 11036 -24832 11144 -24798
rect 12990 -24832 13098 -24798
rect 11036 -24844 13098 -24832
rect 13236 -24172 15298 -24160
rect 13236 -24206 13344 -24172
rect 15190 -24206 15298 -24172
rect 13236 -24218 15298 -24206
rect 13236 -24268 13294 -24218
rect 13236 -24736 13248 -24268
rect 13282 -24736 13294 -24268
rect 15240 -24268 15298 -24218
rect 13236 -24786 13294 -24736
rect 15240 -24736 15252 -24268
rect 15286 -24736 15298 -24268
rect 15240 -24786 15298 -24736
rect 13236 -24798 15298 -24786
rect 13236 -24832 13344 -24798
rect 15190 -24832 15298 -24798
rect 13236 -24844 15298 -24832
rect 15436 -24172 17498 -24160
rect 15436 -24206 15544 -24172
rect 17390 -24206 17498 -24172
rect 15436 -24218 17498 -24206
rect 15436 -24268 15494 -24218
rect 15436 -24736 15448 -24268
rect 15482 -24736 15494 -24268
rect 17440 -24268 17498 -24218
rect 15436 -24786 15494 -24736
rect 17440 -24736 17452 -24268
rect 17486 -24736 17498 -24268
rect 17440 -24786 17498 -24736
rect 15436 -24798 17498 -24786
rect 15436 -24832 15544 -24798
rect 17390 -24832 17498 -24798
rect 15436 -24844 17498 -24832
rect 17636 -24172 19698 -24160
rect 17636 -24206 17744 -24172
rect 19590 -24206 19698 -24172
rect 17636 -24218 19698 -24206
rect 17636 -24268 17694 -24218
rect 17636 -24736 17648 -24268
rect 17682 -24736 17694 -24268
rect 19640 -24268 19698 -24218
rect 17636 -24786 17694 -24736
rect 19640 -24736 19652 -24268
rect 19686 -24736 19698 -24268
rect 19640 -24786 19698 -24736
rect 17636 -24798 19698 -24786
rect 17636 -24832 17744 -24798
rect 19590 -24832 19698 -24798
rect 17636 -24844 19698 -24832
rect 19836 -24172 21898 -24160
rect 19836 -24206 19944 -24172
rect 21790 -24206 21898 -24172
rect 19836 -24218 21898 -24206
rect 19836 -24268 19894 -24218
rect 19836 -24736 19848 -24268
rect 19882 -24736 19894 -24268
rect 21840 -24268 21898 -24218
rect 19836 -24786 19894 -24736
rect 21840 -24736 21852 -24268
rect 21886 -24736 21898 -24268
rect 33024 -24288 33036 -23642
rect 33070 -24288 33082 -23642
rect 34240 -23642 34298 -23592
rect 33024 -24338 33082 -24288
rect 34240 -24288 34252 -23642
rect 34286 -24288 34298 -23642
rect 34240 -24338 34298 -24288
rect 33024 -24350 34298 -24338
rect 33024 -24384 33132 -24350
rect 34190 -24384 34298 -24350
rect 33024 -24396 34298 -24384
rect 34396 -23544 37250 -23532
rect 34396 -23578 34504 -23544
rect 37142 -23578 37250 -23544
rect 34396 -23590 37250 -23578
rect 34396 -23640 34454 -23590
rect 34396 -24286 34408 -23640
rect 34442 -24286 34454 -23640
rect 37192 -23640 37250 -23590
rect 34396 -24336 34454 -24286
rect 37192 -24286 37204 -23640
rect 37238 -24286 37250 -23640
rect 37192 -24336 37250 -24286
rect 34396 -24348 37250 -24336
rect 34396 -24382 34504 -24348
rect 37142 -24382 37250 -24348
rect 34396 -24394 37250 -24382
rect 21840 -24786 21898 -24736
rect 19836 -24798 21898 -24786
rect 19836 -24832 19944 -24798
rect 21790 -24832 21898 -24798
rect 19836 -24844 21898 -24832
rect 22184 -24514 27076 -24502
rect 22184 -24548 22292 -24514
rect 26968 -24548 27076 -24514
rect 22184 -24560 27076 -24548
rect 22184 -24610 22242 -24560
rect 36 -24972 2098 -24960
rect 36 -25006 144 -24972
rect 1990 -25006 2098 -24972
rect 36 -25018 2098 -25006
rect 36 -25068 94 -25018
rect 36 -25536 48 -25068
rect 82 -25536 94 -25068
rect 2040 -25068 2098 -25018
rect 36 -25586 94 -25536
rect 2040 -25536 2052 -25068
rect 2086 -25536 2098 -25068
rect 2040 -25586 2098 -25536
rect 36 -25598 2098 -25586
rect 36 -25632 144 -25598
rect 1990 -25632 2098 -25598
rect 36 -25644 2098 -25632
rect 2236 -24972 4298 -24960
rect 2236 -25006 2344 -24972
rect 4190 -25006 4298 -24972
rect 2236 -25018 4298 -25006
rect 2236 -25068 2294 -25018
rect 2236 -25536 2248 -25068
rect 2282 -25536 2294 -25068
rect 4240 -25068 4298 -25018
rect 2236 -25586 2294 -25536
rect 4240 -25536 4252 -25068
rect 4286 -25536 4298 -25068
rect 4240 -25586 4298 -25536
rect 2236 -25598 4298 -25586
rect 2236 -25632 2344 -25598
rect 4190 -25632 4298 -25598
rect 2236 -25644 4298 -25632
rect 4436 -24972 6498 -24960
rect 4436 -25006 4544 -24972
rect 6390 -25006 6498 -24972
rect 4436 -25018 6498 -25006
rect 4436 -25068 4494 -25018
rect 4436 -25536 4448 -25068
rect 4482 -25536 4494 -25068
rect 6440 -25068 6498 -25018
rect 4436 -25586 4494 -25536
rect 6440 -25536 6452 -25068
rect 6486 -25536 6498 -25068
rect 6440 -25586 6498 -25536
rect 4436 -25598 6498 -25586
rect 4436 -25632 4544 -25598
rect 6390 -25632 6498 -25598
rect 4436 -25644 6498 -25632
rect 6636 -24972 8698 -24960
rect 6636 -25006 6744 -24972
rect 8590 -25006 8698 -24972
rect 6636 -25018 8698 -25006
rect 6636 -25068 6694 -25018
rect 6636 -25536 6648 -25068
rect 6682 -25536 6694 -25068
rect 8640 -25068 8698 -25018
rect 6636 -25586 6694 -25536
rect 8640 -25536 8652 -25068
rect 8686 -25536 8698 -25068
rect 8640 -25586 8698 -25536
rect 6636 -25598 8698 -25586
rect 6636 -25632 6744 -25598
rect 8590 -25632 8698 -25598
rect 6636 -25644 8698 -25632
rect 8836 -24972 10898 -24960
rect 8836 -25006 8944 -24972
rect 10790 -25006 10898 -24972
rect 8836 -25018 10898 -25006
rect 8836 -25068 8894 -25018
rect 8836 -25536 8848 -25068
rect 8882 -25536 8894 -25068
rect 10840 -25068 10898 -25018
rect 8836 -25586 8894 -25536
rect 10840 -25536 10852 -25068
rect 10886 -25536 10898 -25068
rect 10840 -25586 10898 -25536
rect 8836 -25598 10898 -25586
rect 8836 -25632 8944 -25598
rect 10790 -25632 10898 -25598
rect 8836 -25644 10898 -25632
rect 11036 -24972 13098 -24960
rect 11036 -25006 11144 -24972
rect 12990 -25006 13098 -24972
rect 11036 -25018 13098 -25006
rect 11036 -25068 11094 -25018
rect 11036 -25536 11048 -25068
rect 11082 -25536 11094 -25068
rect 13040 -25068 13098 -25018
rect 11036 -25586 11094 -25536
rect 13040 -25536 13052 -25068
rect 13086 -25536 13098 -25068
rect 13040 -25586 13098 -25536
rect 11036 -25598 13098 -25586
rect 11036 -25632 11144 -25598
rect 12990 -25632 13098 -25598
rect 11036 -25644 13098 -25632
rect 13236 -24972 15298 -24960
rect 13236 -25006 13344 -24972
rect 15190 -25006 15298 -24972
rect 13236 -25018 15298 -25006
rect 13236 -25068 13294 -25018
rect 13236 -25536 13248 -25068
rect 13282 -25536 13294 -25068
rect 15240 -25068 15298 -25018
rect 13236 -25586 13294 -25536
rect 15240 -25536 15252 -25068
rect 15286 -25536 15298 -25068
rect 15240 -25586 15298 -25536
rect 13236 -25598 15298 -25586
rect 13236 -25632 13344 -25598
rect 15190 -25632 15298 -25598
rect 13236 -25644 15298 -25632
rect 15436 -24972 17498 -24960
rect 15436 -25006 15544 -24972
rect 17390 -25006 17498 -24972
rect 15436 -25018 17498 -25006
rect 15436 -25068 15494 -25018
rect 15436 -25536 15448 -25068
rect 15482 -25536 15494 -25068
rect 17440 -25068 17498 -25018
rect 15436 -25586 15494 -25536
rect 17440 -25536 17452 -25068
rect 17486 -25536 17498 -25068
rect 17440 -25586 17498 -25536
rect 15436 -25598 17498 -25586
rect 15436 -25632 15544 -25598
rect 17390 -25632 17498 -25598
rect 15436 -25644 17498 -25632
rect 17636 -24972 19698 -24960
rect 17636 -25006 17744 -24972
rect 19590 -25006 19698 -24972
rect 17636 -25018 19698 -25006
rect 17636 -25068 17694 -25018
rect 17636 -25536 17648 -25068
rect 17682 -25536 17694 -25068
rect 19640 -25068 19698 -25018
rect 17636 -25586 17694 -25536
rect 19640 -25536 19652 -25068
rect 19686 -25536 19698 -25068
rect 19640 -25586 19698 -25536
rect 17636 -25598 19698 -25586
rect 17636 -25632 17744 -25598
rect 19590 -25632 19698 -25598
rect 17636 -25644 19698 -25632
rect 19836 -24972 21898 -24960
rect 19836 -25006 19944 -24972
rect 21790 -25006 21898 -24972
rect 19836 -25018 21898 -25006
rect 19836 -25068 19894 -25018
rect 19836 -25536 19848 -25068
rect 19882 -25536 19894 -25068
rect 21840 -25068 21898 -25018
rect 19836 -25586 19894 -25536
rect 21840 -25536 21852 -25068
rect 21886 -25536 21898 -25068
rect 21840 -25586 21898 -25536
rect 19836 -25598 21898 -25586
rect 19836 -25632 19944 -25598
rect 21790 -25632 21898 -25598
rect 19836 -25644 21898 -25632
rect 36 -25772 2098 -25760
rect 36 -25806 144 -25772
rect 1990 -25806 2098 -25772
rect 36 -25818 2098 -25806
rect 36 -25868 94 -25818
rect 36 -26336 48 -25868
rect 82 -26336 94 -25868
rect 2040 -25868 2098 -25818
rect 36 -26386 94 -26336
rect 2040 -26336 2052 -25868
rect 2086 -26336 2098 -25868
rect 2040 -26386 2098 -26336
rect 36 -26398 2098 -26386
rect 36 -26432 144 -26398
rect 1990 -26432 2098 -26398
rect 36 -26444 2098 -26432
rect 2236 -25772 4298 -25760
rect 2236 -25806 2344 -25772
rect 4190 -25806 4298 -25772
rect 2236 -25818 4298 -25806
rect 2236 -25868 2294 -25818
rect 2236 -26336 2248 -25868
rect 2282 -26336 2294 -25868
rect 4240 -25868 4298 -25818
rect 2236 -26386 2294 -26336
rect 4240 -26336 4252 -25868
rect 4286 -26336 4298 -25868
rect 4240 -26386 4298 -26336
rect 2236 -26398 4298 -26386
rect 2236 -26432 2344 -26398
rect 4190 -26432 4298 -26398
rect 2236 -26444 4298 -26432
rect 4436 -25772 6498 -25760
rect 4436 -25806 4544 -25772
rect 6390 -25806 6498 -25772
rect 4436 -25818 6498 -25806
rect 4436 -25868 4494 -25818
rect 4436 -26336 4448 -25868
rect 4482 -26336 4494 -25868
rect 6440 -25868 6498 -25818
rect 4436 -26386 4494 -26336
rect 6440 -26336 6452 -25868
rect 6486 -26336 6498 -25868
rect 6440 -26386 6498 -26336
rect 4436 -26398 6498 -26386
rect 4436 -26432 4544 -26398
rect 6390 -26432 6498 -26398
rect 4436 -26444 6498 -26432
rect 6636 -25772 8698 -25760
rect 6636 -25806 6744 -25772
rect 8590 -25806 8698 -25772
rect 6636 -25818 8698 -25806
rect 6636 -25868 6694 -25818
rect 6636 -26336 6648 -25868
rect 6682 -26336 6694 -25868
rect 8640 -25868 8698 -25818
rect 6636 -26386 6694 -26336
rect 8640 -26336 8652 -25868
rect 8686 -26336 8698 -25868
rect 8640 -26386 8698 -26336
rect 6636 -26398 8698 -26386
rect 6636 -26432 6744 -26398
rect 8590 -26432 8698 -26398
rect 6636 -26444 8698 -26432
rect 8836 -25772 10898 -25760
rect 8836 -25806 8944 -25772
rect 10790 -25806 10898 -25772
rect 8836 -25818 10898 -25806
rect 8836 -25868 8894 -25818
rect 8836 -26336 8848 -25868
rect 8882 -26336 8894 -25868
rect 10840 -25868 10898 -25818
rect 8836 -26386 8894 -26336
rect 10840 -26336 10852 -25868
rect 10886 -26336 10898 -25868
rect 10840 -26386 10898 -26336
rect 8836 -26398 10898 -26386
rect 8836 -26432 8944 -26398
rect 10790 -26432 10898 -26398
rect 8836 -26444 10898 -26432
rect 11036 -25772 13098 -25760
rect 11036 -25806 11144 -25772
rect 12990 -25806 13098 -25772
rect 11036 -25818 13098 -25806
rect 11036 -25868 11094 -25818
rect 11036 -26336 11048 -25868
rect 11082 -26336 11094 -25868
rect 13040 -25868 13098 -25818
rect 11036 -26386 11094 -26336
rect 13040 -26336 13052 -25868
rect 13086 -26336 13098 -25868
rect 13040 -26386 13098 -26336
rect 11036 -26398 13098 -26386
rect 11036 -26432 11144 -26398
rect 12990 -26432 13098 -26398
rect 11036 -26444 13098 -26432
rect 13236 -25772 15298 -25760
rect 13236 -25806 13344 -25772
rect 15190 -25806 15298 -25772
rect 13236 -25818 15298 -25806
rect 13236 -25868 13294 -25818
rect 13236 -26336 13248 -25868
rect 13282 -26336 13294 -25868
rect 15240 -25868 15298 -25818
rect 13236 -26386 13294 -26336
rect 15240 -26336 15252 -25868
rect 15286 -26336 15298 -25868
rect 15240 -26386 15298 -26336
rect 13236 -26398 15298 -26386
rect 13236 -26432 13344 -26398
rect 15190 -26432 15298 -26398
rect 13236 -26444 15298 -26432
rect 15436 -25772 17498 -25760
rect 15436 -25806 15544 -25772
rect 17390 -25806 17498 -25772
rect 15436 -25818 17498 -25806
rect 15436 -25868 15494 -25818
rect 15436 -26336 15448 -25868
rect 15482 -26336 15494 -25868
rect 17440 -25868 17498 -25818
rect 15436 -26386 15494 -26336
rect 17440 -26336 17452 -25868
rect 17486 -26336 17498 -25868
rect 17440 -26386 17498 -26336
rect 15436 -26398 17498 -26386
rect 15436 -26432 15544 -26398
rect 17390 -26432 17498 -26398
rect 15436 -26444 17498 -26432
rect 17636 -25772 19698 -25760
rect 17636 -25806 17744 -25772
rect 19590 -25806 19698 -25772
rect 17636 -25818 19698 -25806
rect 17636 -25868 17694 -25818
rect 17636 -26336 17648 -25868
rect 17682 -26336 17694 -25868
rect 19640 -25868 19698 -25818
rect 17636 -26386 17694 -26336
rect 19640 -26336 19652 -25868
rect 19686 -26336 19698 -25868
rect 19640 -26386 19698 -26336
rect 17636 -26398 19698 -26386
rect 17636 -26432 17744 -26398
rect 19590 -26432 19698 -26398
rect 17636 -26444 19698 -26432
rect 19836 -25772 21898 -25760
rect 19836 -25806 19944 -25772
rect 21790 -25806 21898 -25772
rect 19836 -25818 21898 -25806
rect 19836 -25868 19894 -25818
rect 19836 -26336 19848 -25868
rect 19882 -26336 19894 -25868
rect 21840 -25868 21898 -25818
rect 19836 -26386 19894 -26336
rect 21840 -26336 21852 -25868
rect 21886 -26336 21898 -25868
rect 21840 -26386 21898 -26336
rect 19836 -26398 21898 -26386
rect 19836 -26432 19944 -26398
rect 21790 -26432 21898 -26398
rect 19836 -26444 21898 -26432
rect 36 -26572 2098 -26560
rect 36 -26606 144 -26572
rect 1990 -26606 2098 -26572
rect 36 -26618 2098 -26606
rect 36 -26668 94 -26618
rect 36 -27136 48 -26668
rect 82 -27136 94 -26668
rect 2040 -26668 2098 -26618
rect 36 -27186 94 -27136
rect 2040 -27136 2052 -26668
rect 2086 -27136 2098 -26668
rect 2040 -27186 2098 -27136
rect 36 -27198 2098 -27186
rect 36 -27232 144 -27198
rect 1990 -27232 2098 -27198
rect 36 -27244 2098 -27232
rect 2236 -26572 4298 -26560
rect 2236 -26606 2344 -26572
rect 4190 -26606 4298 -26572
rect 2236 -26618 4298 -26606
rect 2236 -26668 2294 -26618
rect 2236 -27136 2248 -26668
rect 2282 -27136 2294 -26668
rect 4240 -26668 4298 -26618
rect 2236 -27186 2294 -27136
rect 4240 -27136 4252 -26668
rect 4286 -27136 4298 -26668
rect 4240 -27186 4298 -27136
rect 2236 -27198 4298 -27186
rect 2236 -27232 2344 -27198
rect 4190 -27232 4298 -27198
rect 2236 -27244 4298 -27232
rect 4436 -26572 6498 -26560
rect 4436 -26606 4544 -26572
rect 6390 -26606 6498 -26572
rect 4436 -26618 6498 -26606
rect 4436 -26668 4494 -26618
rect 4436 -27136 4448 -26668
rect 4482 -27136 4494 -26668
rect 6440 -26668 6498 -26618
rect 4436 -27186 4494 -27136
rect 6440 -27136 6452 -26668
rect 6486 -27136 6498 -26668
rect 6440 -27186 6498 -27136
rect 4436 -27198 6498 -27186
rect 4436 -27232 4544 -27198
rect 6390 -27232 6498 -27198
rect 4436 -27244 6498 -27232
rect 6636 -26572 8698 -26560
rect 6636 -26606 6744 -26572
rect 8590 -26606 8698 -26572
rect 6636 -26618 8698 -26606
rect 6636 -26668 6694 -26618
rect 6636 -27136 6648 -26668
rect 6682 -27136 6694 -26668
rect 8640 -26668 8698 -26618
rect 6636 -27186 6694 -27136
rect 8640 -27136 8652 -26668
rect 8686 -27136 8698 -26668
rect 8640 -27186 8698 -27136
rect 6636 -27198 8698 -27186
rect 6636 -27232 6744 -27198
rect 8590 -27232 8698 -27198
rect 6636 -27244 8698 -27232
rect 8836 -26572 10898 -26560
rect 8836 -26606 8944 -26572
rect 10790 -26606 10898 -26572
rect 8836 -26618 10898 -26606
rect 8836 -26668 8894 -26618
rect 8836 -27136 8848 -26668
rect 8882 -27136 8894 -26668
rect 10840 -26668 10898 -26618
rect 8836 -27186 8894 -27136
rect 10840 -27136 10852 -26668
rect 10886 -27136 10898 -26668
rect 10840 -27186 10898 -27136
rect 8836 -27198 10898 -27186
rect 8836 -27232 8944 -27198
rect 10790 -27232 10898 -27198
rect 8836 -27244 10898 -27232
rect 11036 -26572 13098 -26560
rect 11036 -26606 11144 -26572
rect 12990 -26606 13098 -26572
rect 11036 -26618 13098 -26606
rect 11036 -26668 11094 -26618
rect 11036 -27136 11048 -26668
rect 11082 -27136 11094 -26668
rect 13040 -26668 13098 -26618
rect 11036 -27186 11094 -27136
rect 13040 -27136 13052 -26668
rect 13086 -27136 13098 -26668
rect 13040 -27186 13098 -27136
rect 11036 -27198 13098 -27186
rect 11036 -27232 11144 -27198
rect 12990 -27232 13098 -27198
rect 11036 -27244 13098 -27232
rect 13236 -26572 15298 -26560
rect 13236 -26606 13344 -26572
rect 15190 -26606 15298 -26572
rect 13236 -26618 15298 -26606
rect 13236 -26668 13294 -26618
rect 13236 -27136 13248 -26668
rect 13282 -27136 13294 -26668
rect 15240 -26668 15298 -26618
rect 13236 -27186 13294 -27136
rect 15240 -27136 15252 -26668
rect 15286 -27136 15298 -26668
rect 15240 -27186 15298 -27136
rect 13236 -27198 15298 -27186
rect 13236 -27232 13344 -27198
rect 15190 -27232 15298 -27198
rect 13236 -27244 15298 -27232
rect 15436 -26572 17498 -26560
rect 15436 -26606 15544 -26572
rect 17390 -26606 17498 -26572
rect 15436 -26618 17498 -26606
rect 15436 -26668 15494 -26618
rect 15436 -27136 15448 -26668
rect 15482 -27136 15494 -26668
rect 17440 -26668 17498 -26618
rect 15436 -27186 15494 -27136
rect 17440 -27136 17452 -26668
rect 17486 -27136 17498 -26668
rect 17440 -27186 17498 -27136
rect 15436 -27198 17498 -27186
rect 15436 -27232 15544 -27198
rect 17390 -27232 17498 -27198
rect 15436 -27244 17498 -27232
rect 17636 -26572 19698 -26560
rect 17636 -26606 17744 -26572
rect 19590 -26606 19698 -26572
rect 17636 -26618 19698 -26606
rect 17636 -26668 17694 -26618
rect 17636 -27136 17648 -26668
rect 17682 -27136 17694 -26668
rect 19640 -26668 19698 -26618
rect 17636 -27186 17694 -27136
rect 19640 -27136 19652 -26668
rect 19686 -27136 19698 -26668
rect 19640 -27186 19698 -27136
rect 17636 -27198 19698 -27186
rect 17636 -27232 17744 -27198
rect 19590 -27232 19698 -27198
rect 17636 -27244 19698 -27232
rect 19836 -26572 21898 -26560
rect 19836 -26606 19944 -26572
rect 21790 -26606 21898 -26572
rect 19836 -26618 21898 -26606
rect 19836 -26668 19894 -26618
rect 19836 -27136 19848 -26668
rect 19882 -27136 19894 -26668
rect 21840 -26668 21898 -26618
rect 19836 -27186 19894 -27136
rect 21840 -27136 21852 -26668
rect 21886 -27136 21898 -26668
rect 21840 -27186 21898 -27136
rect 19836 -27198 21898 -27186
rect 19836 -27232 19944 -27198
rect 21790 -27232 21898 -27198
rect 19836 -27244 21898 -27232
rect 36 -27372 2098 -27360
rect 36 -27406 144 -27372
rect 1990 -27406 2098 -27372
rect 36 -27418 2098 -27406
rect 36 -27468 94 -27418
rect 36 -27936 48 -27468
rect 82 -27936 94 -27468
rect 2040 -27468 2098 -27418
rect 36 -27986 94 -27936
rect 2040 -27936 2052 -27468
rect 2086 -27936 2098 -27468
rect 2040 -27986 2098 -27936
rect 36 -27998 2098 -27986
rect 36 -28032 144 -27998
rect 1990 -28032 2098 -27998
rect 36 -28044 2098 -28032
rect 2236 -27372 4298 -27360
rect 2236 -27406 2344 -27372
rect 4190 -27406 4298 -27372
rect 2236 -27418 4298 -27406
rect 2236 -27468 2294 -27418
rect 2236 -27936 2248 -27468
rect 2282 -27936 2294 -27468
rect 4240 -27468 4298 -27418
rect 2236 -27986 2294 -27936
rect 4240 -27936 4252 -27468
rect 4286 -27936 4298 -27468
rect 4240 -27986 4298 -27936
rect 2236 -27998 4298 -27986
rect 2236 -28032 2344 -27998
rect 4190 -28032 4298 -27998
rect 2236 -28044 4298 -28032
rect 4436 -27372 6498 -27360
rect 4436 -27406 4544 -27372
rect 6390 -27406 6498 -27372
rect 4436 -27418 6498 -27406
rect 4436 -27468 4494 -27418
rect 4436 -27936 4448 -27468
rect 4482 -27936 4494 -27468
rect 6440 -27468 6498 -27418
rect 4436 -27986 4494 -27936
rect 6440 -27936 6452 -27468
rect 6486 -27936 6498 -27468
rect 6440 -27986 6498 -27936
rect 4436 -27998 6498 -27986
rect 4436 -28032 4544 -27998
rect 6390 -28032 6498 -27998
rect 4436 -28044 6498 -28032
rect 6636 -27372 8698 -27360
rect 6636 -27406 6744 -27372
rect 8590 -27406 8698 -27372
rect 6636 -27418 8698 -27406
rect 6636 -27468 6694 -27418
rect 6636 -27936 6648 -27468
rect 6682 -27936 6694 -27468
rect 8640 -27468 8698 -27418
rect 6636 -27986 6694 -27936
rect 8640 -27936 8652 -27468
rect 8686 -27936 8698 -27468
rect 8640 -27986 8698 -27936
rect 6636 -27998 8698 -27986
rect 6636 -28032 6744 -27998
rect 8590 -28032 8698 -27998
rect 6636 -28044 8698 -28032
rect 8836 -27372 10898 -27360
rect 8836 -27406 8944 -27372
rect 10790 -27406 10898 -27372
rect 8836 -27418 10898 -27406
rect 8836 -27468 8894 -27418
rect 8836 -27936 8848 -27468
rect 8882 -27936 8894 -27468
rect 10840 -27468 10898 -27418
rect 8836 -27986 8894 -27936
rect 10840 -27936 10852 -27468
rect 10886 -27936 10898 -27468
rect 10840 -27986 10898 -27936
rect 8836 -27998 10898 -27986
rect 8836 -28032 8944 -27998
rect 10790 -28032 10898 -27998
rect 8836 -28044 10898 -28032
rect 11036 -27372 13098 -27360
rect 11036 -27406 11144 -27372
rect 12990 -27406 13098 -27372
rect 11036 -27418 13098 -27406
rect 11036 -27468 11094 -27418
rect 11036 -27936 11048 -27468
rect 11082 -27936 11094 -27468
rect 13040 -27468 13098 -27418
rect 11036 -27986 11094 -27936
rect 13040 -27936 13052 -27468
rect 13086 -27936 13098 -27468
rect 13040 -27986 13098 -27936
rect 11036 -27998 13098 -27986
rect 11036 -28032 11144 -27998
rect 12990 -28032 13098 -27998
rect 11036 -28044 13098 -28032
rect 13236 -27372 15298 -27360
rect 13236 -27406 13344 -27372
rect 15190 -27406 15298 -27372
rect 13236 -27418 15298 -27406
rect 13236 -27468 13294 -27418
rect 13236 -27936 13248 -27468
rect 13282 -27936 13294 -27468
rect 15240 -27468 15298 -27418
rect 13236 -27986 13294 -27936
rect 15240 -27936 15252 -27468
rect 15286 -27936 15298 -27468
rect 15240 -27986 15298 -27936
rect 13236 -27998 15298 -27986
rect 13236 -28032 13344 -27998
rect 15190 -28032 15298 -27998
rect 13236 -28044 15298 -28032
rect 15436 -27372 17498 -27360
rect 15436 -27406 15544 -27372
rect 17390 -27406 17498 -27372
rect 15436 -27418 17498 -27406
rect 15436 -27468 15494 -27418
rect 15436 -27936 15448 -27468
rect 15482 -27936 15494 -27468
rect 17440 -27468 17498 -27418
rect 15436 -27986 15494 -27936
rect 17440 -27936 17452 -27468
rect 17486 -27936 17498 -27468
rect 17440 -27986 17498 -27936
rect 15436 -27998 17498 -27986
rect 15436 -28032 15544 -27998
rect 17390 -28032 17498 -27998
rect 15436 -28044 17498 -28032
rect 17636 -27372 19698 -27360
rect 17636 -27406 17744 -27372
rect 19590 -27406 19698 -27372
rect 17636 -27418 19698 -27406
rect 17636 -27468 17694 -27418
rect 17636 -27936 17648 -27468
rect 17682 -27936 17694 -27468
rect 19640 -27468 19698 -27418
rect 17636 -27986 17694 -27936
rect 19640 -27936 19652 -27468
rect 19686 -27936 19698 -27468
rect 19640 -27986 19698 -27936
rect 17636 -27998 19698 -27986
rect 17636 -28032 17744 -27998
rect 19590 -28032 19698 -27998
rect 17636 -28044 19698 -28032
rect 19836 -27372 21898 -27360
rect 19836 -27406 19944 -27372
rect 21790 -27406 21898 -27372
rect 19836 -27418 21898 -27406
rect 19836 -27468 19894 -27418
rect 19836 -27936 19848 -27468
rect 19882 -27936 19894 -27468
rect 21840 -27468 21898 -27418
rect 19836 -27986 19894 -27936
rect 21840 -27936 21852 -27468
rect 21886 -27936 21898 -27468
rect 21840 -27986 21898 -27936
rect 19836 -27998 21898 -27986
rect 19836 -28032 19944 -27998
rect 21790 -28032 21898 -27998
rect 19836 -28044 21898 -28032
rect 36 -28172 2098 -28160
rect 36 -28206 144 -28172
rect 1990 -28206 2098 -28172
rect 36 -28218 2098 -28206
rect 36 -28268 94 -28218
rect 36 -28736 48 -28268
rect 82 -28736 94 -28268
rect 2040 -28268 2098 -28218
rect 36 -28786 94 -28736
rect 2040 -28736 2052 -28268
rect 2086 -28736 2098 -28268
rect 2040 -28786 2098 -28736
rect 36 -28798 2098 -28786
rect 36 -28832 144 -28798
rect 1990 -28832 2098 -28798
rect 36 -28844 2098 -28832
rect 2236 -28172 4298 -28160
rect 2236 -28206 2344 -28172
rect 4190 -28206 4298 -28172
rect 2236 -28218 4298 -28206
rect 2236 -28268 2294 -28218
rect 2236 -28736 2248 -28268
rect 2282 -28736 2294 -28268
rect 4240 -28268 4298 -28218
rect 2236 -28786 2294 -28736
rect 4240 -28736 4252 -28268
rect 4286 -28736 4298 -28268
rect 4240 -28786 4298 -28736
rect 2236 -28798 4298 -28786
rect 2236 -28832 2344 -28798
rect 4190 -28832 4298 -28798
rect 2236 -28844 4298 -28832
rect 4436 -28172 6498 -28160
rect 4436 -28206 4544 -28172
rect 6390 -28206 6498 -28172
rect 4436 -28218 6498 -28206
rect 4436 -28268 4494 -28218
rect 4436 -28736 4448 -28268
rect 4482 -28736 4494 -28268
rect 6440 -28268 6498 -28218
rect 4436 -28786 4494 -28736
rect 6440 -28736 6452 -28268
rect 6486 -28736 6498 -28268
rect 6440 -28786 6498 -28736
rect 4436 -28798 6498 -28786
rect 4436 -28832 4544 -28798
rect 6390 -28832 6498 -28798
rect 4436 -28844 6498 -28832
rect 6636 -28172 8698 -28160
rect 6636 -28206 6744 -28172
rect 8590 -28206 8698 -28172
rect 6636 -28218 8698 -28206
rect 6636 -28268 6694 -28218
rect 6636 -28736 6648 -28268
rect 6682 -28736 6694 -28268
rect 8640 -28268 8698 -28218
rect 6636 -28786 6694 -28736
rect 8640 -28736 8652 -28268
rect 8686 -28736 8698 -28268
rect 8640 -28786 8698 -28736
rect 6636 -28798 8698 -28786
rect 6636 -28832 6744 -28798
rect 8590 -28832 8698 -28798
rect 6636 -28844 8698 -28832
rect 8836 -28172 10898 -28160
rect 8836 -28206 8944 -28172
rect 10790 -28206 10898 -28172
rect 8836 -28218 10898 -28206
rect 8836 -28268 8894 -28218
rect 8836 -28736 8848 -28268
rect 8882 -28736 8894 -28268
rect 10840 -28268 10898 -28218
rect 8836 -28786 8894 -28736
rect 10840 -28736 10852 -28268
rect 10886 -28736 10898 -28268
rect 10840 -28786 10898 -28736
rect 8836 -28798 10898 -28786
rect 8836 -28832 8944 -28798
rect 10790 -28832 10898 -28798
rect 8836 -28844 10898 -28832
rect 11036 -28172 13098 -28160
rect 11036 -28206 11144 -28172
rect 12990 -28206 13098 -28172
rect 11036 -28218 13098 -28206
rect 11036 -28268 11094 -28218
rect 11036 -28736 11048 -28268
rect 11082 -28736 11094 -28268
rect 13040 -28268 13098 -28218
rect 11036 -28786 11094 -28736
rect 13040 -28736 13052 -28268
rect 13086 -28736 13098 -28268
rect 13040 -28786 13098 -28736
rect 11036 -28798 13098 -28786
rect 11036 -28832 11144 -28798
rect 12990 -28832 13098 -28798
rect 11036 -28844 13098 -28832
rect 13236 -28172 15298 -28160
rect 13236 -28206 13344 -28172
rect 15190 -28206 15298 -28172
rect 13236 -28218 15298 -28206
rect 13236 -28268 13294 -28218
rect 13236 -28736 13248 -28268
rect 13282 -28736 13294 -28268
rect 15240 -28268 15298 -28218
rect 13236 -28786 13294 -28736
rect 15240 -28736 15252 -28268
rect 15286 -28736 15298 -28268
rect 15240 -28786 15298 -28736
rect 13236 -28798 15298 -28786
rect 13236 -28832 13344 -28798
rect 15190 -28832 15298 -28798
rect 13236 -28844 15298 -28832
rect 15436 -28172 17498 -28160
rect 15436 -28206 15544 -28172
rect 17390 -28206 17498 -28172
rect 15436 -28218 17498 -28206
rect 15436 -28268 15494 -28218
rect 15436 -28736 15448 -28268
rect 15482 -28736 15494 -28268
rect 17440 -28268 17498 -28218
rect 15436 -28786 15494 -28736
rect 17440 -28736 17452 -28268
rect 17486 -28736 17498 -28268
rect 17440 -28786 17498 -28736
rect 15436 -28798 17498 -28786
rect 15436 -28832 15544 -28798
rect 17390 -28832 17498 -28798
rect 15436 -28844 17498 -28832
rect 17636 -28172 19698 -28160
rect 17636 -28206 17744 -28172
rect 19590 -28206 19698 -28172
rect 17636 -28218 19698 -28206
rect 17636 -28268 17694 -28218
rect 17636 -28736 17648 -28268
rect 17682 -28736 17694 -28268
rect 19640 -28268 19698 -28218
rect 17636 -28786 17694 -28736
rect 19640 -28736 19652 -28268
rect 19686 -28736 19698 -28268
rect 19640 -28786 19698 -28736
rect 17636 -28798 19698 -28786
rect 17636 -28832 17744 -28798
rect 19590 -28832 19698 -28798
rect 17636 -28844 19698 -28832
rect 19836 -28172 21898 -28160
rect 19836 -28206 19944 -28172
rect 21790 -28206 21898 -28172
rect 19836 -28218 21898 -28206
rect 19836 -28268 19894 -28218
rect 19836 -28736 19848 -28268
rect 19882 -28736 19894 -28268
rect 21840 -28268 21898 -28218
rect 19836 -28786 19894 -28736
rect 21840 -28736 21852 -28268
rect 21886 -28736 21898 -28268
rect 21840 -28786 21898 -28736
rect 19836 -28798 21898 -28786
rect 19836 -28832 19944 -28798
rect 21790 -28832 21898 -28798
rect 19836 -28844 21898 -28832
rect 36 -28972 2098 -28960
rect 36 -29006 144 -28972
rect 1990 -29006 2098 -28972
rect 36 -29018 2098 -29006
rect 36 -29068 94 -29018
rect 36 -29536 48 -29068
rect 82 -29536 94 -29068
rect 2040 -29068 2098 -29018
rect 36 -29586 94 -29536
rect 2040 -29536 2052 -29068
rect 2086 -29536 2098 -29068
rect 2040 -29586 2098 -29536
rect 36 -29598 2098 -29586
rect 36 -29632 144 -29598
rect 1990 -29632 2098 -29598
rect 36 -29644 2098 -29632
rect 2236 -28972 4298 -28960
rect 2236 -29006 2344 -28972
rect 4190 -29006 4298 -28972
rect 2236 -29018 4298 -29006
rect 2236 -29068 2294 -29018
rect 2236 -29536 2248 -29068
rect 2282 -29536 2294 -29068
rect 4240 -29068 4298 -29018
rect 2236 -29586 2294 -29536
rect 4240 -29536 4252 -29068
rect 4286 -29536 4298 -29068
rect 4240 -29586 4298 -29536
rect 2236 -29598 4298 -29586
rect 2236 -29632 2344 -29598
rect 4190 -29632 4298 -29598
rect 2236 -29644 4298 -29632
rect 4436 -28972 6498 -28960
rect 4436 -29006 4544 -28972
rect 6390 -29006 6498 -28972
rect 4436 -29018 6498 -29006
rect 4436 -29068 4494 -29018
rect 4436 -29536 4448 -29068
rect 4482 -29536 4494 -29068
rect 6440 -29068 6498 -29018
rect 4436 -29586 4494 -29536
rect 6440 -29536 6452 -29068
rect 6486 -29536 6498 -29068
rect 6440 -29586 6498 -29536
rect 4436 -29598 6498 -29586
rect 4436 -29632 4544 -29598
rect 6390 -29632 6498 -29598
rect 4436 -29644 6498 -29632
rect 6636 -28972 8698 -28960
rect 6636 -29006 6744 -28972
rect 8590 -29006 8698 -28972
rect 6636 -29018 8698 -29006
rect 6636 -29068 6694 -29018
rect 6636 -29536 6648 -29068
rect 6682 -29536 6694 -29068
rect 8640 -29068 8698 -29018
rect 6636 -29586 6694 -29536
rect 8640 -29536 8652 -29068
rect 8686 -29536 8698 -29068
rect 8640 -29586 8698 -29536
rect 6636 -29598 8698 -29586
rect 6636 -29632 6744 -29598
rect 8590 -29632 8698 -29598
rect 6636 -29644 8698 -29632
rect 8836 -28972 10898 -28960
rect 8836 -29006 8944 -28972
rect 10790 -29006 10898 -28972
rect 8836 -29018 10898 -29006
rect 8836 -29068 8894 -29018
rect 8836 -29536 8848 -29068
rect 8882 -29536 8894 -29068
rect 10840 -29068 10898 -29018
rect 8836 -29586 8894 -29536
rect 10840 -29536 10852 -29068
rect 10886 -29536 10898 -29068
rect 10840 -29586 10898 -29536
rect 8836 -29598 10898 -29586
rect 8836 -29632 8944 -29598
rect 10790 -29632 10898 -29598
rect 8836 -29644 10898 -29632
rect 11036 -28972 13098 -28960
rect 11036 -29006 11144 -28972
rect 12990 -29006 13098 -28972
rect 11036 -29018 13098 -29006
rect 11036 -29068 11094 -29018
rect 11036 -29536 11048 -29068
rect 11082 -29536 11094 -29068
rect 13040 -29068 13098 -29018
rect 11036 -29586 11094 -29536
rect 13040 -29536 13052 -29068
rect 13086 -29536 13098 -29068
rect 13040 -29586 13098 -29536
rect 11036 -29598 13098 -29586
rect 11036 -29632 11144 -29598
rect 12990 -29632 13098 -29598
rect 11036 -29644 13098 -29632
rect 13236 -28972 15298 -28960
rect 13236 -29006 13344 -28972
rect 15190 -29006 15298 -28972
rect 13236 -29018 15298 -29006
rect 13236 -29068 13294 -29018
rect 13236 -29536 13248 -29068
rect 13282 -29536 13294 -29068
rect 15240 -29068 15298 -29018
rect 13236 -29586 13294 -29536
rect 15240 -29536 15252 -29068
rect 15286 -29536 15298 -29068
rect 15240 -29586 15298 -29536
rect 13236 -29598 15298 -29586
rect 13236 -29632 13344 -29598
rect 15190 -29632 15298 -29598
rect 13236 -29644 15298 -29632
rect 15436 -28972 17498 -28960
rect 15436 -29006 15544 -28972
rect 17390 -29006 17498 -28972
rect 15436 -29018 17498 -29006
rect 15436 -29068 15494 -29018
rect 15436 -29536 15448 -29068
rect 15482 -29536 15494 -29068
rect 17440 -29068 17498 -29018
rect 15436 -29586 15494 -29536
rect 17440 -29536 17452 -29068
rect 17486 -29536 17498 -29068
rect 17440 -29586 17498 -29536
rect 15436 -29598 17498 -29586
rect 15436 -29632 15544 -29598
rect 17390 -29632 17498 -29598
rect 15436 -29644 17498 -29632
rect 17636 -28972 19698 -28960
rect 17636 -29006 17744 -28972
rect 19590 -29006 19698 -28972
rect 17636 -29018 19698 -29006
rect 17636 -29068 17694 -29018
rect 17636 -29536 17648 -29068
rect 17682 -29536 17694 -29068
rect 19640 -29068 19698 -29018
rect 17636 -29586 17694 -29536
rect 19640 -29536 19652 -29068
rect 19686 -29536 19698 -29068
rect 19640 -29586 19698 -29536
rect 17636 -29598 19698 -29586
rect 17636 -29632 17744 -29598
rect 19590 -29632 19698 -29598
rect 17636 -29644 19698 -29632
rect 19836 -28972 21898 -28960
rect 19836 -29006 19944 -28972
rect 21790 -29006 21898 -28972
rect 19836 -29018 21898 -29006
rect 19836 -29068 19894 -29018
rect 19836 -29536 19848 -29068
rect 19882 -29536 19894 -29068
rect 21840 -29068 21898 -29018
rect 19836 -29586 19894 -29536
rect 21840 -29536 21852 -29068
rect 21886 -29536 21898 -29068
rect 21840 -29586 21898 -29536
rect 19836 -29598 21898 -29586
rect 19836 -29632 19944 -29598
rect 21790 -29632 21898 -29598
rect 19836 -29644 21898 -29632
rect 36 -29772 2098 -29760
rect 36 -29806 144 -29772
rect 1990 -29806 2098 -29772
rect 36 -29818 2098 -29806
rect 36 -29868 94 -29818
rect 36 -30336 48 -29868
rect 82 -30336 94 -29868
rect 2040 -29868 2098 -29818
rect 36 -30386 94 -30336
rect 2040 -30336 2052 -29868
rect 2086 -30336 2098 -29868
rect 2040 -30386 2098 -30336
rect 36 -30398 2098 -30386
rect 36 -30432 144 -30398
rect 1990 -30432 2098 -30398
rect 36 -30444 2098 -30432
rect 2236 -29772 4298 -29760
rect 2236 -29806 2344 -29772
rect 4190 -29806 4298 -29772
rect 2236 -29818 4298 -29806
rect 2236 -29868 2294 -29818
rect 2236 -30336 2248 -29868
rect 2282 -30336 2294 -29868
rect 4240 -29868 4298 -29818
rect 2236 -30386 2294 -30336
rect 4240 -30336 4252 -29868
rect 4286 -30336 4298 -29868
rect 4240 -30386 4298 -30336
rect 2236 -30398 4298 -30386
rect 2236 -30432 2344 -30398
rect 4190 -30432 4298 -30398
rect 2236 -30444 4298 -30432
rect 4436 -29772 6498 -29760
rect 4436 -29806 4544 -29772
rect 6390 -29806 6498 -29772
rect 4436 -29818 6498 -29806
rect 4436 -29868 4494 -29818
rect 4436 -30336 4448 -29868
rect 4482 -30336 4494 -29868
rect 6440 -29868 6498 -29818
rect 4436 -30386 4494 -30336
rect 6440 -30336 6452 -29868
rect 6486 -30336 6498 -29868
rect 6440 -30386 6498 -30336
rect 4436 -30398 6498 -30386
rect 4436 -30432 4544 -30398
rect 6390 -30432 6498 -30398
rect 4436 -30444 6498 -30432
rect 6636 -29772 8698 -29760
rect 6636 -29806 6744 -29772
rect 8590 -29806 8698 -29772
rect 6636 -29818 8698 -29806
rect 6636 -29868 6694 -29818
rect 6636 -30336 6648 -29868
rect 6682 -30336 6694 -29868
rect 8640 -29868 8698 -29818
rect 6636 -30386 6694 -30336
rect 8640 -30336 8652 -29868
rect 8686 -30336 8698 -29868
rect 8640 -30386 8698 -30336
rect 6636 -30398 8698 -30386
rect 6636 -30432 6744 -30398
rect 8590 -30432 8698 -30398
rect 6636 -30444 8698 -30432
rect 8836 -29772 10898 -29760
rect 8836 -29806 8944 -29772
rect 10790 -29806 10898 -29772
rect 8836 -29818 10898 -29806
rect 8836 -29868 8894 -29818
rect 8836 -30336 8848 -29868
rect 8882 -30336 8894 -29868
rect 10840 -29868 10898 -29818
rect 8836 -30386 8894 -30336
rect 10840 -30336 10852 -29868
rect 10886 -30336 10898 -29868
rect 10840 -30386 10898 -30336
rect 8836 -30398 10898 -30386
rect 8836 -30432 8944 -30398
rect 10790 -30432 10898 -30398
rect 8836 -30444 10898 -30432
rect 11036 -29772 13098 -29760
rect 11036 -29806 11144 -29772
rect 12990 -29806 13098 -29772
rect 11036 -29818 13098 -29806
rect 11036 -29868 11094 -29818
rect 11036 -30336 11048 -29868
rect 11082 -30336 11094 -29868
rect 13040 -29868 13098 -29818
rect 11036 -30386 11094 -30336
rect 13040 -30336 13052 -29868
rect 13086 -30336 13098 -29868
rect 13040 -30386 13098 -30336
rect 11036 -30398 13098 -30386
rect 11036 -30432 11144 -30398
rect 12990 -30432 13098 -30398
rect 11036 -30444 13098 -30432
rect 13236 -29772 15298 -29760
rect 13236 -29806 13344 -29772
rect 15190 -29806 15298 -29772
rect 13236 -29818 15298 -29806
rect 13236 -29868 13294 -29818
rect 13236 -30336 13248 -29868
rect 13282 -30336 13294 -29868
rect 15240 -29868 15298 -29818
rect 13236 -30386 13294 -30336
rect 15240 -30336 15252 -29868
rect 15286 -30336 15298 -29868
rect 15240 -30386 15298 -30336
rect 13236 -30398 15298 -30386
rect 13236 -30432 13344 -30398
rect 15190 -30432 15298 -30398
rect 13236 -30444 15298 -30432
rect 15436 -29772 17498 -29760
rect 15436 -29806 15544 -29772
rect 17390 -29806 17498 -29772
rect 15436 -29818 17498 -29806
rect 15436 -29868 15494 -29818
rect 15436 -30336 15448 -29868
rect 15482 -30336 15494 -29868
rect 17440 -29868 17498 -29818
rect 15436 -30386 15494 -30336
rect 17440 -30336 17452 -29868
rect 17486 -30336 17498 -29868
rect 17440 -30386 17498 -30336
rect 15436 -30398 17498 -30386
rect 15436 -30432 15544 -30398
rect 17390 -30432 17498 -30398
rect 15436 -30444 17498 -30432
rect 17636 -29772 19698 -29760
rect 17636 -29806 17744 -29772
rect 19590 -29806 19698 -29772
rect 17636 -29818 19698 -29806
rect 17636 -29868 17694 -29818
rect 17636 -30336 17648 -29868
rect 17682 -30336 17694 -29868
rect 19640 -29868 19698 -29818
rect 17636 -30386 17694 -30336
rect 19640 -30336 19652 -29868
rect 19686 -30336 19698 -29868
rect 19640 -30386 19698 -30336
rect 17636 -30398 19698 -30386
rect 17636 -30432 17744 -30398
rect 19590 -30432 19698 -30398
rect 17636 -30444 19698 -30432
rect 19836 -29772 21898 -29760
rect 19836 -29806 19944 -29772
rect 21790 -29806 21898 -29772
rect 19836 -29818 21898 -29806
rect 19836 -29868 19894 -29818
rect 19836 -30336 19848 -29868
rect 19882 -30336 19894 -29868
rect 21840 -29868 21898 -29818
rect 19836 -30386 19894 -30336
rect 21840 -30336 21852 -29868
rect 21886 -30336 21898 -29868
rect 21840 -30386 21898 -30336
rect 19836 -30398 21898 -30386
rect 19836 -30432 19944 -30398
rect 21790 -30432 21898 -30398
rect 19836 -30444 21898 -30432
rect 36 -30572 2098 -30560
rect 36 -30606 144 -30572
rect 1990 -30606 2098 -30572
rect 36 -30618 2098 -30606
rect 36 -30668 94 -30618
rect 36 -31136 48 -30668
rect 82 -31136 94 -30668
rect 2040 -30668 2098 -30618
rect 36 -31186 94 -31136
rect 2040 -31136 2052 -30668
rect 2086 -31136 2098 -30668
rect 2040 -31186 2098 -31136
rect 36 -31198 2098 -31186
rect 36 -31232 144 -31198
rect 1990 -31232 2098 -31198
rect 36 -31244 2098 -31232
rect 2236 -30572 4298 -30560
rect 2236 -30606 2344 -30572
rect 4190 -30606 4298 -30572
rect 2236 -30618 4298 -30606
rect 2236 -30668 2294 -30618
rect 2236 -31136 2248 -30668
rect 2282 -31136 2294 -30668
rect 4240 -30668 4298 -30618
rect 2236 -31186 2294 -31136
rect 4240 -31136 4252 -30668
rect 4286 -31136 4298 -30668
rect 4240 -31186 4298 -31136
rect 2236 -31198 4298 -31186
rect 2236 -31232 2344 -31198
rect 4190 -31232 4298 -31198
rect 2236 -31244 4298 -31232
rect 4436 -30572 6498 -30560
rect 4436 -30606 4544 -30572
rect 6390 -30606 6498 -30572
rect 4436 -30618 6498 -30606
rect 4436 -30668 4494 -30618
rect 4436 -31136 4448 -30668
rect 4482 -31136 4494 -30668
rect 6440 -30668 6498 -30618
rect 4436 -31186 4494 -31136
rect 6440 -31136 6452 -30668
rect 6486 -31136 6498 -30668
rect 6440 -31186 6498 -31136
rect 4436 -31198 6498 -31186
rect 4436 -31232 4544 -31198
rect 6390 -31232 6498 -31198
rect 4436 -31244 6498 -31232
rect 6636 -30572 8698 -30560
rect 6636 -30606 6744 -30572
rect 8590 -30606 8698 -30572
rect 6636 -30618 8698 -30606
rect 6636 -30668 6694 -30618
rect 6636 -31136 6648 -30668
rect 6682 -31136 6694 -30668
rect 8640 -30668 8698 -30618
rect 6636 -31186 6694 -31136
rect 8640 -31136 8652 -30668
rect 8686 -31136 8698 -30668
rect 8640 -31186 8698 -31136
rect 6636 -31198 8698 -31186
rect 6636 -31232 6744 -31198
rect 8590 -31232 8698 -31198
rect 6636 -31244 8698 -31232
rect 8836 -30572 10898 -30560
rect 8836 -30606 8944 -30572
rect 10790 -30606 10898 -30572
rect 8836 -30618 10898 -30606
rect 8836 -30668 8894 -30618
rect 8836 -31136 8848 -30668
rect 8882 -31136 8894 -30668
rect 10840 -30668 10898 -30618
rect 8836 -31186 8894 -31136
rect 10840 -31136 10852 -30668
rect 10886 -31136 10898 -30668
rect 10840 -31186 10898 -31136
rect 8836 -31198 10898 -31186
rect 8836 -31232 8944 -31198
rect 10790 -31232 10898 -31198
rect 8836 -31244 10898 -31232
rect 11036 -30572 13098 -30560
rect 11036 -30606 11144 -30572
rect 12990 -30606 13098 -30572
rect 11036 -30618 13098 -30606
rect 11036 -30668 11094 -30618
rect 11036 -31136 11048 -30668
rect 11082 -31136 11094 -30668
rect 13040 -30668 13098 -30618
rect 11036 -31186 11094 -31136
rect 13040 -31136 13052 -30668
rect 13086 -31136 13098 -30668
rect 13040 -31186 13098 -31136
rect 11036 -31198 13098 -31186
rect 11036 -31232 11144 -31198
rect 12990 -31232 13098 -31198
rect 11036 -31244 13098 -31232
rect 13236 -30572 15298 -30560
rect 13236 -30606 13344 -30572
rect 15190 -30606 15298 -30572
rect 13236 -30618 15298 -30606
rect 13236 -30668 13294 -30618
rect 13236 -31136 13248 -30668
rect 13282 -31136 13294 -30668
rect 15240 -30668 15298 -30618
rect 13236 -31186 13294 -31136
rect 15240 -31136 15252 -30668
rect 15286 -31136 15298 -30668
rect 15240 -31186 15298 -31136
rect 13236 -31198 15298 -31186
rect 13236 -31232 13344 -31198
rect 15190 -31232 15298 -31198
rect 13236 -31244 15298 -31232
rect 15436 -30572 17498 -30560
rect 15436 -30606 15544 -30572
rect 17390 -30606 17498 -30572
rect 15436 -30618 17498 -30606
rect 15436 -30668 15494 -30618
rect 15436 -31136 15448 -30668
rect 15482 -31136 15494 -30668
rect 17440 -30668 17498 -30618
rect 15436 -31186 15494 -31136
rect 17440 -31136 17452 -30668
rect 17486 -31136 17498 -30668
rect 17440 -31186 17498 -31136
rect 15436 -31198 17498 -31186
rect 15436 -31232 15544 -31198
rect 17390 -31232 17498 -31198
rect 15436 -31244 17498 -31232
rect 17636 -30572 19698 -30560
rect 17636 -30606 17744 -30572
rect 19590 -30606 19698 -30572
rect 17636 -30618 19698 -30606
rect 17636 -30668 17694 -30618
rect 17636 -31136 17648 -30668
rect 17682 -31136 17694 -30668
rect 19640 -30668 19698 -30618
rect 17636 -31186 17694 -31136
rect 19640 -31136 19652 -30668
rect 19686 -31136 19698 -30668
rect 19640 -31186 19698 -31136
rect 17636 -31198 19698 -31186
rect 17636 -31232 17744 -31198
rect 19590 -31232 19698 -31198
rect 17636 -31244 19698 -31232
rect 19836 -30572 21898 -30560
rect 19836 -30606 19944 -30572
rect 21790 -30606 21898 -30572
rect 19836 -30618 21898 -30606
rect 19836 -30668 19894 -30618
rect 19836 -31136 19848 -30668
rect 19882 -31136 19894 -30668
rect 21840 -30668 21898 -30618
rect 19836 -31186 19894 -31136
rect 21840 -31136 21852 -30668
rect 21886 -31136 21898 -30668
rect 21840 -31186 21898 -31136
rect 19836 -31198 21898 -31186
rect 19836 -31232 19944 -31198
rect 21790 -31232 21898 -31198
rect 19836 -31244 21898 -31232
rect 36 -31372 2098 -31360
rect 36 -31406 144 -31372
rect 1990 -31406 2098 -31372
rect 36 -31418 2098 -31406
rect 36 -31468 94 -31418
rect 36 -31936 48 -31468
rect 82 -31936 94 -31468
rect 2040 -31468 2098 -31418
rect 36 -31986 94 -31936
rect 2040 -31936 2052 -31468
rect 2086 -31936 2098 -31468
rect 2040 -31986 2098 -31936
rect 36 -31998 2098 -31986
rect 36 -32032 144 -31998
rect 1990 -32032 2098 -31998
rect 36 -32044 2098 -32032
rect 2236 -31372 4298 -31360
rect 2236 -31406 2344 -31372
rect 4190 -31406 4298 -31372
rect 2236 -31418 4298 -31406
rect 2236 -31468 2294 -31418
rect 2236 -31936 2248 -31468
rect 2282 -31936 2294 -31468
rect 4240 -31468 4298 -31418
rect 2236 -31986 2294 -31936
rect 4240 -31936 4252 -31468
rect 4286 -31936 4298 -31468
rect 4240 -31986 4298 -31936
rect 2236 -31998 4298 -31986
rect 2236 -32032 2344 -31998
rect 4190 -32032 4298 -31998
rect 2236 -32044 4298 -32032
rect 4436 -31372 6498 -31360
rect 4436 -31406 4544 -31372
rect 6390 -31406 6498 -31372
rect 4436 -31418 6498 -31406
rect 4436 -31468 4494 -31418
rect 4436 -31936 4448 -31468
rect 4482 -31936 4494 -31468
rect 6440 -31468 6498 -31418
rect 4436 -31986 4494 -31936
rect 6440 -31936 6452 -31468
rect 6486 -31936 6498 -31468
rect 6440 -31986 6498 -31936
rect 4436 -31998 6498 -31986
rect 4436 -32032 4544 -31998
rect 6390 -32032 6498 -31998
rect 4436 -32044 6498 -32032
rect 6636 -31372 8698 -31360
rect 6636 -31406 6744 -31372
rect 8590 -31406 8698 -31372
rect 6636 -31418 8698 -31406
rect 6636 -31468 6694 -31418
rect 6636 -31936 6648 -31468
rect 6682 -31936 6694 -31468
rect 8640 -31468 8698 -31418
rect 6636 -31986 6694 -31936
rect 8640 -31936 8652 -31468
rect 8686 -31936 8698 -31468
rect 8640 -31986 8698 -31936
rect 6636 -31998 8698 -31986
rect 6636 -32032 6744 -31998
rect 8590 -32032 8698 -31998
rect 6636 -32044 8698 -32032
rect 8836 -31372 10898 -31360
rect 8836 -31406 8944 -31372
rect 10790 -31406 10898 -31372
rect 8836 -31418 10898 -31406
rect 8836 -31468 8894 -31418
rect 8836 -31936 8848 -31468
rect 8882 -31936 8894 -31468
rect 10840 -31468 10898 -31418
rect 8836 -31986 8894 -31936
rect 10840 -31936 10852 -31468
rect 10886 -31936 10898 -31468
rect 10840 -31986 10898 -31936
rect 8836 -31998 10898 -31986
rect 8836 -32032 8944 -31998
rect 10790 -32032 10898 -31998
rect 8836 -32044 10898 -32032
rect 11036 -31372 13098 -31360
rect 11036 -31406 11144 -31372
rect 12990 -31406 13098 -31372
rect 11036 -31418 13098 -31406
rect 11036 -31468 11094 -31418
rect 11036 -31936 11048 -31468
rect 11082 -31936 11094 -31468
rect 13040 -31468 13098 -31418
rect 11036 -31986 11094 -31936
rect 13040 -31936 13052 -31468
rect 13086 -31936 13098 -31468
rect 13040 -31986 13098 -31936
rect 11036 -31998 13098 -31986
rect 11036 -32032 11144 -31998
rect 12990 -32032 13098 -31998
rect 11036 -32044 13098 -32032
rect 13236 -31372 15298 -31360
rect 13236 -31406 13344 -31372
rect 15190 -31406 15298 -31372
rect 13236 -31418 15298 -31406
rect 13236 -31468 13294 -31418
rect 13236 -31936 13248 -31468
rect 13282 -31936 13294 -31468
rect 15240 -31468 15298 -31418
rect 13236 -31986 13294 -31936
rect 15240 -31936 15252 -31468
rect 15286 -31936 15298 -31468
rect 15240 -31986 15298 -31936
rect 13236 -31998 15298 -31986
rect 13236 -32032 13344 -31998
rect 15190 -32032 15298 -31998
rect 13236 -32044 15298 -32032
rect 15436 -31372 17498 -31360
rect 15436 -31406 15544 -31372
rect 17390 -31406 17498 -31372
rect 15436 -31418 17498 -31406
rect 15436 -31468 15494 -31418
rect 15436 -31936 15448 -31468
rect 15482 -31936 15494 -31468
rect 17440 -31468 17498 -31418
rect 15436 -31986 15494 -31936
rect 17440 -31936 17452 -31468
rect 17486 -31936 17498 -31468
rect 17440 -31986 17498 -31936
rect 15436 -31998 17498 -31986
rect 15436 -32032 15544 -31998
rect 17390 -32032 17498 -31998
rect 15436 -32044 17498 -32032
rect 17636 -31372 19698 -31360
rect 17636 -31406 17744 -31372
rect 19590 -31406 19698 -31372
rect 17636 -31418 19698 -31406
rect 17636 -31468 17694 -31418
rect 17636 -31936 17648 -31468
rect 17682 -31936 17694 -31468
rect 19640 -31468 19698 -31418
rect 17636 -31986 17694 -31936
rect 19640 -31936 19652 -31468
rect 19686 -31936 19698 -31468
rect 19640 -31986 19698 -31936
rect 17636 -31998 19698 -31986
rect 17636 -32032 17744 -31998
rect 19590 -32032 19698 -31998
rect 17636 -32044 19698 -32032
rect 19836 -31372 21898 -31360
rect 19836 -31406 19944 -31372
rect 21790 -31406 21898 -31372
rect 19836 -31418 21898 -31406
rect 19836 -31468 19894 -31418
rect 19836 -31936 19848 -31468
rect 19882 -31936 19894 -31468
rect 21840 -31468 21898 -31418
rect 19836 -31986 19894 -31936
rect 21840 -31936 21852 -31468
rect 21886 -31936 21898 -31468
rect 21840 -31986 21898 -31936
rect 19836 -31998 21898 -31986
rect 19836 -32032 19944 -31998
rect 21790 -32032 21898 -31998
rect 19836 -32044 21898 -32032
rect 22184 -31968 22196 -24610
rect 22230 -31968 22242 -24610
rect 27018 -24610 27076 -24560
rect 22184 -32018 22242 -31968
rect 27018 -31968 27030 -24610
rect 27064 -31968 27076 -24610
rect 34746 -24696 36008 -24684
rect 34746 -24730 34854 -24696
rect 35900 -24730 36008 -24696
rect 34746 -24742 36008 -24730
rect 34746 -24792 34804 -24742
rect 34746 -26966 34758 -24792
rect 34792 -26966 34804 -24792
rect 35950 -24792 36008 -24742
rect 34746 -27016 34804 -26966
rect 35950 -26966 35962 -24792
rect 35996 -26966 36008 -24792
rect 35950 -27016 36008 -26966
rect 34746 -27028 36008 -27016
rect 34746 -27062 34854 -27028
rect 35900 -27062 36008 -27028
rect 34746 -27074 36008 -27062
rect 36086 -24696 37348 -24684
rect 36086 -24730 36194 -24696
rect 37240 -24730 37348 -24696
rect 36086 -24742 37348 -24730
rect 36086 -24792 36144 -24742
rect 36086 -26966 36098 -24792
rect 36132 -26966 36144 -24792
rect 37290 -24792 37348 -24742
rect 36086 -27016 36144 -26966
rect 37290 -26966 37302 -24792
rect 37336 -26966 37348 -24792
rect 37290 -27016 37348 -26966
rect 36086 -27028 37348 -27016
rect 36086 -27062 36194 -27028
rect 37240 -27062 37348 -27028
rect 36086 -27074 37348 -27062
rect 31666 -28302 33030 -28290
rect 31666 -28336 31774 -28302
rect 32042 -28336 32214 -28302
rect 32482 -28336 32654 -28302
rect 32922 -28336 33030 -28302
rect 31666 -28348 33030 -28336
rect 31666 -28398 31724 -28348
rect 31666 -29044 31678 -28398
rect 31712 -29044 31724 -28398
rect 32092 -28398 32164 -28348
rect 31666 -29094 31724 -29044
rect 32092 -29044 32104 -28398
rect 32138 -29044 32164 -28398
rect 32092 -29094 32164 -29044
rect 32532 -29094 32604 -28348
rect 32972 -28590 33030 -28348
rect 33866 -28302 35230 -28290
rect 33866 -28336 33974 -28302
rect 34242 -28336 34414 -28302
rect 34682 -28336 34854 -28302
rect 35122 -28336 35230 -28302
rect 33866 -28348 35230 -28336
rect 33866 -28398 33924 -28348
rect 32960 -28602 33744 -28590
rect 32960 -28636 33068 -28602
rect 33636 -28636 33744 -28602
rect 32960 -28648 33744 -28636
rect 32960 -28698 33030 -28648
rect 32960 -29044 32972 -28698
rect 33006 -29044 33030 -28698
rect 33686 -28698 33744 -28648
rect 32960 -29094 33030 -29044
rect 33686 -29044 33698 -28698
rect 33732 -29044 33744 -28698
rect 33686 -29094 33744 -29044
rect 31666 -29106 33744 -29094
rect 31666 -29140 31774 -29106
rect 32042 -29140 32214 -29106
rect 32482 -29140 32654 -29106
rect 32922 -29140 33068 -29106
rect 33636 -29140 33744 -29106
rect 31666 -29152 33744 -29140
rect 33866 -29044 33878 -28398
rect 33912 -29044 33924 -28398
rect 34292 -28398 34364 -28348
rect 33866 -29094 33924 -29044
rect 34292 -29044 34304 -28398
rect 34338 -29044 34364 -28398
rect 34292 -29094 34364 -29044
rect 34732 -29094 34804 -28348
rect 35172 -28590 35230 -28348
rect 36066 -28302 37430 -28290
rect 36066 -28336 36174 -28302
rect 36442 -28336 36614 -28302
rect 36882 -28336 37054 -28302
rect 37322 -28336 37430 -28302
rect 36066 -28348 37430 -28336
rect 36066 -28398 36124 -28348
rect 35160 -28602 35944 -28590
rect 35160 -28636 35268 -28602
rect 35836 -28636 35944 -28602
rect 35160 -28648 35944 -28636
rect 35160 -28698 35230 -28648
rect 35160 -29044 35172 -28698
rect 35206 -29044 35230 -28698
rect 35886 -28698 35944 -28648
rect 35160 -29094 35230 -29044
rect 35886 -29044 35898 -28698
rect 35932 -29044 35944 -28698
rect 35886 -29094 35944 -29044
rect 33866 -29106 35944 -29094
rect 33866 -29140 33974 -29106
rect 34242 -29140 34414 -29106
rect 34682 -29140 34854 -29106
rect 35122 -29140 35268 -29106
rect 35836 -29140 35944 -29106
rect 33866 -29152 35944 -29140
rect 36066 -29044 36078 -28398
rect 36112 -29044 36124 -28398
rect 36492 -28398 36564 -28348
rect 36066 -29094 36124 -29044
rect 36492 -29044 36504 -28398
rect 36538 -29044 36564 -28398
rect 36492 -29094 36564 -29044
rect 36932 -29094 37004 -28348
rect 37372 -28590 37430 -28348
rect 37360 -28602 38144 -28590
rect 37360 -28636 37468 -28602
rect 38036 -28636 38144 -28602
rect 37360 -28648 38144 -28636
rect 37360 -28698 37430 -28648
rect 37360 -29044 37372 -28698
rect 37406 -29044 37430 -28698
rect 38086 -28698 38144 -28648
rect 37360 -29094 37430 -29044
rect 38086 -29044 38098 -28698
rect 38132 -29044 38144 -28698
rect 38086 -29094 38144 -29044
rect 36066 -29106 38144 -29094
rect 36066 -29140 36174 -29106
rect 36442 -29140 36614 -29106
rect 36882 -29140 37054 -29106
rect 37322 -29140 37468 -29106
rect 38036 -29140 38144 -29106
rect 36066 -29152 38144 -29140
rect 31678 -30884 33756 -30872
rect 31678 -30918 31786 -30884
rect 32354 -30918 32500 -30884
rect 32768 -30918 32940 -30884
rect 33208 -30918 33380 -30884
rect 33648 -30918 33756 -30884
rect 31678 -30930 33756 -30918
rect 31678 -30980 31736 -30930
rect 31678 -31326 31690 -30980
rect 31724 -31326 31736 -30980
rect 32392 -30980 32462 -30930
rect 31678 -31376 31736 -31326
rect 32392 -31326 32416 -30980
rect 32450 -31326 32462 -30980
rect 32392 -31376 32462 -31326
rect 31678 -31388 32462 -31376
rect 31678 -31422 31786 -31388
rect 32354 -31422 32462 -31388
rect 31678 -31434 32462 -31422
rect 32392 -31676 32450 -31434
rect 32818 -31676 32890 -30930
rect 33258 -30980 33330 -30930
rect 33258 -31626 33284 -30980
rect 33318 -31626 33330 -30980
rect 33698 -30980 33756 -30930
rect 33258 -31676 33330 -31626
rect 33698 -31626 33710 -30980
rect 33744 -31626 33756 -30980
rect 33878 -30884 35956 -30872
rect 33878 -30918 33986 -30884
rect 34554 -30918 34700 -30884
rect 34968 -30918 35140 -30884
rect 35408 -30918 35580 -30884
rect 35848 -30918 35956 -30884
rect 33878 -30930 35956 -30918
rect 33878 -30980 33936 -30930
rect 33878 -31326 33890 -30980
rect 33924 -31326 33936 -30980
rect 34592 -30980 34662 -30930
rect 33878 -31376 33936 -31326
rect 34592 -31326 34616 -30980
rect 34650 -31326 34662 -30980
rect 34592 -31376 34662 -31326
rect 33878 -31388 34662 -31376
rect 33878 -31422 33986 -31388
rect 34554 -31422 34662 -31388
rect 33878 -31434 34662 -31422
rect 33698 -31676 33756 -31626
rect 32392 -31688 33756 -31676
rect 32392 -31722 32500 -31688
rect 32768 -31722 32940 -31688
rect 33208 -31722 33380 -31688
rect 33648 -31722 33756 -31688
rect 32392 -31734 33756 -31722
rect 34592 -31676 34650 -31434
rect 35018 -31676 35090 -30930
rect 35458 -30980 35530 -30930
rect 35458 -31626 35484 -30980
rect 35518 -31626 35530 -30980
rect 35898 -30980 35956 -30930
rect 35458 -31676 35530 -31626
rect 35898 -31626 35910 -30980
rect 35944 -31626 35956 -30980
rect 36078 -30884 38156 -30872
rect 36078 -30918 36186 -30884
rect 36754 -30918 36900 -30884
rect 37168 -30918 37340 -30884
rect 37608 -30918 37780 -30884
rect 38048 -30918 38156 -30884
rect 36078 -30930 38156 -30918
rect 36078 -30980 36136 -30930
rect 36078 -31326 36090 -30980
rect 36124 -31326 36136 -30980
rect 36792 -30980 36862 -30930
rect 36078 -31376 36136 -31326
rect 36792 -31326 36816 -30980
rect 36850 -31326 36862 -30980
rect 36792 -31376 36862 -31326
rect 36078 -31388 36862 -31376
rect 36078 -31422 36186 -31388
rect 36754 -31422 36862 -31388
rect 36078 -31434 36862 -31422
rect 35898 -31676 35956 -31626
rect 34592 -31688 35956 -31676
rect 34592 -31722 34700 -31688
rect 34968 -31722 35140 -31688
rect 35408 -31722 35580 -31688
rect 35848 -31722 35956 -31688
rect 34592 -31734 35956 -31722
rect 36792 -31676 36850 -31434
rect 37218 -31676 37290 -30930
rect 37658 -30980 37730 -30930
rect 37658 -31626 37684 -30980
rect 37718 -31626 37730 -30980
rect 38098 -30980 38156 -30930
rect 37658 -31676 37730 -31626
rect 38098 -31626 38110 -30980
rect 38144 -31626 38156 -30980
rect 38098 -31676 38156 -31626
rect 36792 -31688 38156 -31676
rect 36792 -31722 36900 -31688
rect 37168 -31722 37340 -31688
rect 37608 -31722 37780 -31688
rect 38048 -31722 38156 -31688
rect 36792 -31734 38156 -31722
rect 27018 -32018 27076 -31968
rect 22184 -32030 27076 -32018
rect 22184 -32064 22292 -32030
rect 26968 -32064 27076 -32030
rect 22184 -32076 27076 -32064
<< psubdiffcont >>
rect 22332 11910 26966 11944
rect 22236 4532 22270 11848
rect 27028 4532 27062 11848
rect 34572 7470 34730 7504
rect 34476 7052 34510 7408
rect 34792 7052 34826 7408
rect 34572 6956 34730 6990
rect 34992 7470 35150 7504
rect 34896 7052 34930 7408
rect 35212 7052 35246 7408
rect 34992 6956 35150 6990
rect 35412 7470 35570 7504
rect 35316 7052 35350 7408
rect 35632 7052 35666 7408
rect 35412 6956 35570 6990
rect 22332 4436 26966 4470
<< nsubdiffcont >>
rect 32892 9008 33478 9042
rect 32796 7972 32830 8946
rect 33540 7972 33574 8946
rect 32892 7876 33478 7910
rect 33732 9008 34318 9042
rect 33636 7972 33670 8946
rect 34380 7972 34414 8946
rect 34572 8788 34730 8822
rect 34476 8152 34510 8726
rect 34792 8152 34826 8726
rect 34572 8056 34730 8090
rect 34992 8788 35150 8822
rect 34896 8152 34930 8726
rect 35212 8152 35246 8726
rect 34992 8056 35150 8090
rect 35412 8788 35570 8822
rect 35316 8152 35350 8726
rect 35632 8152 35666 8726
rect 35412 8056 35570 8090
rect 33732 7876 34318 7910
<< mvpsubdiffcont >>
rect 145 11875 1973 11909
rect 49 11345 83 11813
rect 2035 11345 2069 11813
rect 145 11249 1973 11283
rect 2345 11875 4173 11909
rect 2249 11345 2283 11813
rect 4235 11345 4269 11813
rect 2345 11249 4173 11283
rect 4545 11875 6373 11909
rect 4449 11345 4483 11813
rect 6435 11345 6469 11813
rect 4545 11249 6373 11283
rect 6745 11875 8573 11909
rect 6649 11345 6683 11813
rect 8635 11345 8669 11813
rect 6745 11249 8573 11283
rect 8945 11875 10773 11909
rect 8849 11345 8883 11813
rect 10835 11345 10869 11813
rect 8945 11249 10773 11283
rect 11145 11875 12973 11909
rect 11049 11345 11083 11813
rect 13035 11345 13069 11813
rect 11145 11249 12973 11283
rect 13345 11875 15173 11909
rect 13249 11345 13283 11813
rect 15235 11345 15269 11813
rect 13345 11249 15173 11283
rect 15545 11875 17373 11909
rect 15449 11345 15483 11813
rect 17435 11345 17469 11813
rect 15545 11249 17373 11283
rect 17745 11875 19573 11909
rect 17649 11345 17683 11813
rect 19635 11345 19669 11813
rect 17745 11249 19573 11283
rect 19945 11875 21773 11909
rect 19849 11345 19883 11813
rect 21835 11345 21869 11813
rect 19945 11249 21773 11283
rect 145 11075 1973 11109
rect 49 10545 83 11013
rect 2035 10545 2069 11013
rect 145 10449 1973 10483
rect 2344 11074 4172 11108
rect 2248 10544 2282 11012
rect 4234 10544 4268 11012
rect 2344 10448 4172 10482
rect 4544 11074 6372 11108
rect 4448 10544 4482 11012
rect 6434 10544 6468 11012
rect 4544 10448 6372 10482
rect 6744 11074 8572 11108
rect 6648 10544 6682 11012
rect 8634 10544 8668 11012
rect 6744 10448 8572 10482
rect 8944 11074 10772 11108
rect 8848 10544 8882 11012
rect 10834 10544 10868 11012
rect 8944 10448 10772 10482
rect 11144 11074 12972 11108
rect 11048 10544 11082 11012
rect 13034 10544 13068 11012
rect 11144 10448 12972 10482
rect 13344 11074 15172 11108
rect 13248 10544 13282 11012
rect 15234 10544 15268 11012
rect 13344 10448 15172 10482
rect 15544 11074 17372 11108
rect 15448 10544 15482 11012
rect 17434 10544 17468 11012
rect 15544 10448 17372 10482
rect 17744 11074 19572 11108
rect 17648 10544 17682 11012
rect 19634 10544 19668 11012
rect 17744 10448 19572 10482
rect 19945 11075 21773 11109
rect 19849 10545 19883 11013
rect 21835 10545 21869 11013
rect 19945 10449 21773 10483
rect 145 10275 1973 10309
rect 49 9745 83 10213
rect 2035 9745 2069 10213
rect 145 9649 1973 9683
rect 2344 10274 4172 10308
rect 2248 9744 2282 10212
rect 4234 9744 4268 10212
rect 2344 9648 4172 9682
rect 4544 10274 6372 10308
rect 4448 9744 4482 10212
rect 6434 9744 6468 10212
rect 4544 9648 6372 9682
rect 6744 10274 8572 10308
rect 6648 9744 6682 10212
rect 8634 9744 8668 10212
rect 6744 9648 8572 9682
rect 8944 10274 10772 10308
rect 8848 9744 8882 10212
rect 10834 9744 10868 10212
rect 8944 9648 10772 9682
rect 11144 10274 12972 10308
rect 11048 9744 11082 10212
rect 13034 9744 13068 10212
rect 11144 9648 12972 9682
rect 13344 10274 15172 10308
rect 13248 9744 13282 10212
rect 15234 9744 15268 10212
rect 13344 9648 15172 9682
rect 15544 10274 17372 10308
rect 15448 9744 15482 10212
rect 17434 9744 17468 10212
rect 15544 9648 17372 9682
rect 17744 10274 19572 10308
rect 17648 9744 17682 10212
rect 19634 9744 19668 10212
rect 17744 9648 19572 9682
rect 19945 10275 21773 10309
rect 19849 9745 19883 10213
rect 21835 9745 21869 10213
rect 19945 9649 21773 9683
rect 145 9475 1973 9509
rect 49 8945 83 9413
rect 2035 8945 2069 9413
rect 145 8849 1973 8883
rect 2344 9474 4172 9508
rect 2248 8944 2282 9412
rect 4234 8944 4268 9412
rect 2344 8848 4172 8882
rect 4544 9474 6372 9508
rect 4448 8944 4482 9412
rect 6434 8944 6468 9412
rect 4544 8848 6372 8882
rect 6744 9474 8572 9508
rect 6648 8944 6682 9412
rect 8634 8944 8668 9412
rect 6744 8848 8572 8882
rect 8944 9474 10772 9508
rect 8848 8944 8882 9412
rect 10834 8944 10868 9412
rect 8944 8848 10772 8882
rect 11144 9474 12972 9508
rect 11048 8944 11082 9412
rect 13034 8944 13068 9412
rect 11144 8848 12972 8882
rect 13344 9474 15172 9508
rect 13248 8944 13282 9412
rect 15234 8944 15268 9412
rect 13344 8848 15172 8882
rect 15544 9474 17372 9508
rect 15448 8944 15482 9412
rect 17434 8944 17468 9412
rect 15544 8848 17372 8882
rect 17744 9474 19572 9508
rect 17648 8944 17682 9412
rect 19634 8944 19668 9412
rect 17744 8848 19572 8882
rect 19945 9475 21773 9509
rect 19849 8945 19883 9413
rect 21835 8945 21869 9413
rect 19945 8849 21773 8883
rect 145 8675 1973 8709
rect 49 8145 83 8613
rect 2035 8145 2069 8613
rect 145 8049 1973 8083
rect 2344 8674 4172 8708
rect 2248 8144 2282 8612
rect 4234 8144 4268 8612
rect 2344 8048 4172 8082
rect 4544 8674 6372 8708
rect 4448 8144 4482 8612
rect 6434 8144 6468 8612
rect 4544 8048 6372 8082
rect 6744 8674 8572 8708
rect 6648 8144 6682 8612
rect 8634 8144 8668 8612
rect 6744 8048 8572 8082
rect 8944 8674 10772 8708
rect 8848 8144 8882 8612
rect 10834 8144 10868 8612
rect 8944 8048 10772 8082
rect 11144 8674 12972 8708
rect 11048 8144 11082 8612
rect 13034 8144 13068 8612
rect 11144 8048 12972 8082
rect 13344 8674 15172 8708
rect 13248 8144 13282 8612
rect 15234 8144 15268 8612
rect 13344 8048 15172 8082
rect 15544 8674 17372 8708
rect 15448 8144 15482 8612
rect 17434 8144 17468 8612
rect 15544 8048 17372 8082
rect 17744 8674 19572 8708
rect 17648 8144 17682 8612
rect 19634 8144 19668 8612
rect 17744 8048 19572 8082
rect 19945 8675 21773 8709
rect 19849 8145 19883 8613
rect 21835 8145 21869 8613
rect 19945 8049 21773 8083
rect 145 7875 1973 7909
rect 49 7345 83 7813
rect 2035 7345 2069 7813
rect 145 7249 1973 7283
rect 2344 7874 4172 7908
rect 2248 7344 2282 7812
rect 4234 7344 4268 7812
rect 2344 7248 4172 7282
rect 4544 7874 6372 7908
rect 4448 7344 4482 7812
rect 6434 7344 6468 7812
rect 4544 7248 6372 7282
rect 6744 7874 8572 7908
rect 6648 7344 6682 7812
rect 8634 7344 8668 7812
rect 6744 7248 8572 7282
rect 8944 7874 10772 7908
rect 8848 7344 8882 7812
rect 10834 7344 10868 7812
rect 8944 7248 10772 7282
rect 11144 7874 12972 7908
rect 11048 7344 11082 7812
rect 13034 7344 13068 7812
rect 11144 7248 12972 7282
rect 13344 7874 15172 7908
rect 13248 7344 13282 7812
rect 15234 7344 15268 7812
rect 13344 7248 15172 7282
rect 15544 7874 17372 7908
rect 15448 7344 15482 7812
rect 17434 7344 17468 7812
rect 15544 7248 17372 7282
rect 17744 7874 19572 7908
rect 17648 7344 17682 7812
rect 19634 7344 19668 7812
rect 17744 7248 19572 7282
rect 19945 7875 21773 7909
rect 19849 7345 19883 7813
rect 21835 7345 21869 7813
rect 19945 7249 21773 7283
rect 145 7075 1973 7109
rect 49 6545 83 7013
rect 2035 6545 2069 7013
rect 145 6449 1973 6483
rect 2344 7074 4172 7108
rect 2248 6544 2282 7012
rect 4234 6544 4268 7012
rect 2344 6448 4172 6482
rect 4544 7074 6372 7108
rect 4448 6544 4482 7012
rect 6434 6544 6468 7012
rect 4544 6448 6372 6482
rect 6744 7074 8572 7108
rect 6648 6544 6682 7012
rect 8634 6544 8668 7012
rect 6744 6448 8572 6482
rect 8944 7074 10772 7108
rect 8848 6544 8882 7012
rect 10834 6544 10868 7012
rect 8944 6448 10772 6482
rect 11144 7074 12972 7108
rect 11048 6544 11082 7012
rect 13034 6544 13068 7012
rect 11144 6448 12972 6482
rect 13344 7074 15172 7108
rect 13248 6544 13282 7012
rect 15234 6544 15268 7012
rect 13344 6448 15172 6482
rect 15544 7074 17372 7108
rect 15448 6544 15482 7012
rect 17434 6544 17468 7012
rect 15544 6448 17372 6482
rect 17744 7074 19572 7108
rect 17648 6544 17682 7012
rect 19634 6544 19668 7012
rect 17744 6448 19572 6482
rect 19945 7075 21773 7109
rect 19849 6545 19883 7013
rect 21835 6545 21869 7013
rect 19945 6449 21773 6483
rect 145 6275 1973 6309
rect 49 5745 83 6213
rect 2035 5745 2069 6213
rect 145 5649 1973 5683
rect 2344 6274 4172 6308
rect 2248 5744 2282 6212
rect 4234 5744 4268 6212
rect 2344 5648 4172 5682
rect 4544 6274 6372 6308
rect 4448 5744 4482 6212
rect 6434 5744 6468 6212
rect 4544 5648 6372 5682
rect 6744 6274 8572 6308
rect 6648 5744 6682 6212
rect 8634 5744 8668 6212
rect 6744 5648 8572 5682
rect 8944 6274 10772 6308
rect 8848 5744 8882 6212
rect 10834 5744 10868 6212
rect 8944 5648 10772 5682
rect 11144 6274 12972 6308
rect 11048 5744 11082 6212
rect 13034 5744 13068 6212
rect 11144 5648 12972 5682
rect 13344 6274 15172 6308
rect 13248 5744 13282 6212
rect 15234 5744 15268 6212
rect 13344 5648 15172 5682
rect 15544 6274 17372 6308
rect 15448 5744 15482 6212
rect 17434 5744 17468 6212
rect 15544 5648 17372 5682
rect 17744 6274 19572 6308
rect 17648 5744 17682 6212
rect 19634 5744 19668 6212
rect 17744 5648 19572 5682
rect 19945 6275 21773 6309
rect 19849 5745 19883 6213
rect 21835 5745 21869 6213
rect 19945 5649 21773 5683
rect 145 5475 1973 5509
rect 49 4945 83 5413
rect 2035 4945 2069 5413
rect 145 4849 1973 4883
rect 2344 5474 4172 5508
rect 2248 4944 2282 5412
rect 4234 4944 4268 5412
rect 2344 4848 4172 4882
rect 4544 5474 6372 5508
rect 4448 4944 4482 5412
rect 6434 4944 6468 5412
rect 4544 4848 6372 4882
rect 6744 5474 8572 5508
rect 6648 4944 6682 5412
rect 8634 4944 8668 5412
rect 6744 4848 8572 4882
rect 8944 5474 10772 5508
rect 8848 4944 8882 5412
rect 10834 4944 10868 5412
rect 8944 4848 10772 4882
rect 11144 5474 12972 5508
rect 11048 4944 11082 5412
rect 13034 4944 13068 5412
rect 11144 4848 12972 4882
rect 13344 5474 15172 5508
rect 13248 4944 13282 5412
rect 15234 4944 15268 5412
rect 13344 4848 15172 4882
rect 15544 5474 17372 5508
rect 15448 4944 15482 5412
rect 17434 4944 17468 5412
rect 15544 4848 17372 4882
rect 17744 5474 19572 5508
rect 17648 4944 17682 5412
rect 19634 4944 19668 5412
rect 17744 4848 19572 4882
rect 19945 5475 21773 5509
rect 19849 4945 19883 5413
rect 21835 4945 21869 5413
rect 19945 4849 21773 4883
rect 145 4675 1973 4709
rect 49 4145 83 4613
rect 2035 4145 2069 4613
rect 145 4049 1973 4083
rect 2345 4675 4173 4709
rect 2249 4145 2283 4613
rect 4235 4145 4269 4613
rect 2345 4049 4173 4083
rect 4545 4675 6373 4709
rect 4449 4145 4483 4613
rect 6435 4145 6469 4613
rect 4545 4049 6373 4083
rect 6745 4675 8573 4709
rect 6649 4145 6683 4613
rect 8635 4145 8669 4613
rect 6745 4049 8573 4083
rect 8946 4676 10774 4710
rect 8850 4146 8884 4614
rect 10836 4146 10870 4614
rect 8946 4050 10774 4084
rect 11146 4676 12974 4710
rect 11050 4146 11084 4614
rect 13036 4146 13070 4614
rect 11146 4050 12974 4084
rect 13345 4675 15173 4709
rect 13249 4145 13283 4613
rect 15235 4145 15269 4613
rect 13345 4049 15173 4083
rect 15545 4675 17373 4709
rect 15449 4145 15483 4613
rect 17435 4145 17469 4613
rect 15545 4049 17373 4083
rect 17745 4675 19573 4709
rect 17649 4145 17683 4613
rect 19635 4145 19669 4613
rect 17745 4049 19573 4083
rect 19945 4675 21773 4709
rect 19849 4145 19883 4613
rect 21835 4145 21869 4613
rect 30064 11903 30648 11937
rect 30819 11903 31087 11937
rect 31259 11903 31527 11937
rect 31699 11903 31967 11937
rect 29968 11413 30002 11841
rect 30710 11413 30744 11841
rect 31603 11413 31637 11841
rect 32029 11413 32063 11841
rect 30064 11317 30648 11351
rect 30819 11317 31087 11351
rect 31259 11317 31527 11351
rect 31699 11317 31967 11351
rect 32264 11903 32848 11937
rect 33019 11903 33287 11937
rect 33459 11903 33727 11937
rect 33899 11903 34167 11937
rect 32168 11413 32202 11841
rect 32910 11413 32944 11841
rect 33803 11413 33837 11841
rect 34229 11413 34263 11841
rect 32264 11317 32848 11351
rect 33019 11317 33287 11351
rect 33459 11317 33727 11351
rect 33899 11317 34167 11351
rect 34464 11903 35048 11937
rect 35219 11903 35487 11937
rect 35659 11903 35927 11937
rect 36099 11903 36367 11937
rect 34368 11413 34402 11841
rect 35110 11413 35144 11841
rect 36003 11413 36037 11841
rect 36429 11413 36463 11841
rect 34464 11317 35048 11351
rect 35219 11317 35487 11351
rect 35659 11317 35927 11351
rect 36099 11317 36367 11351
rect 33434 7614 34176 7648
rect 33338 6924 33372 7552
rect 34238 6924 34272 7552
rect 33434 6828 34176 6862
rect 29644 6334 30672 6368
rect 29548 5904 29582 6272
rect 30734 5904 30768 6272
rect 29644 5808 30672 5842
rect 30984 6334 32012 6368
rect 30888 5904 30922 6272
rect 32074 5904 32108 6272
rect 30984 5808 32012 5842
rect 36334 6100 36962 6134
rect 37120 6100 37748 6134
rect 29884 5684 30452 5718
rect 29788 5294 29822 5622
rect 30514 5294 30548 5622
rect 29884 5198 30452 5232
rect 31194 5684 31762 5718
rect 31098 5294 31132 5622
rect 31824 5294 31858 5622
rect 31194 5198 31762 5232
rect 29644 5074 30672 5108
rect 29548 4644 29582 5012
rect 30734 4644 30768 5012
rect 29644 4548 30672 4582
rect 30984 5074 32012 5108
rect 30888 4644 30922 5012
rect 32074 4644 32108 5012
rect 30984 4548 32012 4582
rect 32684 4134 34058 4168
rect 19945 4049 21773 4083
rect 17064 3492 17806 3526
rect 16968 2464 17002 3430
rect 17868 2464 17902 3430
rect 32588 3444 32622 4072
rect 34120 3444 34154 4072
rect 32684 3348 34058 3382
rect 34874 4134 35458 4168
rect 34778 3444 34812 4072
rect 35520 3444 35554 4072
rect 36238 3864 36272 6038
rect 37024 3864 37058 6038
rect 37810 3864 37844 6038
rect 36334 3768 36962 3802
rect 37120 3768 37748 3802
rect 34874 3348 35458 3382
rect 32354 3204 32780 3238
rect 32258 2514 32292 3142
rect 32842 2514 32876 3142
rect 32354 2418 32780 2452
rect 33954 3204 34380 3238
rect 33858 2514 33892 3142
rect 34442 2514 34476 3142
rect 33954 2418 34380 2452
rect 35554 3204 35980 3238
rect 35458 2514 35492 3142
rect 36042 2514 36076 3142
rect 35554 2418 35980 2452
rect 17064 2368 17806 2402
rect -55 2195 1191 2229
rect -151 1165 -117 2133
rect 1253 1165 1287 2133
rect -55 1069 1191 1103
rect -151 619 -117 987
rect 1253 619 1287 987
rect 1545 2195 2791 2229
rect 1449 1165 1483 2133
rect 2853 1165 2887 2133
rect 1545 1069 2791 1103
rect 1449 619 1483 987
rect 2853 619 2887 987
rect 3145 2195 4391 2229
rect 3049 1165 3083 2133
rect 4453 1165 4487 2133
rect 3145 1069 4391 1103
rect 3049 619 3083 987
rect 4453 619 4487 987
rect 4745 2195 5991 2229
rect 4649 1165 4683 2133
rect 6053 1165 6087 2133
rect 4745 1069 5991 1103
rect 4649 619 4683 987
rect 6053 619 6087 987
rect 6345 2195 7591 2229
rect 6249 1165 6283 2133
rect 7653 1165 7687 2133
rect 6345 1069 7591 1103
rect 6249 619 6283 987
rect 7653 619 7687 987
rect 7945 2195 9191 2229
rect 7849 1165 7883 2133
rect 9253 1165 9287 2133
rect 7945 1069 9191 1103
rect 7849 619 7883 987
rect 9253 619 9287 987
rect 9545 2195 10791 2229
rect 9449 1165 9483 2133
rect 10853 1165 10887 2133
rect 9545 1069 10791 1103
rect 9449 619 9483 987
rect 10853 619 10887 987
rect 11145 2195 12391 2229
rect 11049 1165 11083 2133
rect 12453 1165 12487 2133
rect 11145 1069 12391 1103
rect 11049 619 11083 987
rect 12453 619 12487 987
rect 12745 2195 13991 2229
rect 12649 1165 12683 2133
rect 14053 1165 14087 2133
rect 12745 1069 13991 1103
rect 12649 619 12683 987
rect 14053 619 14087 987
rect 14345 2195 15591 2229
rect 14249 1165 14283 2133
rect 15653 1165 15687 2133
rect 14345 1069 15591 1103
rect 14249 619 14283 987
rect 15653 619 15687 987
rect 15945 2195 17191 2229
rect 15849 1165 15883 2133
rect 17253 1165 17287 2133
rect 15945 1069 17191 1103
rect 15849 619 15883 987
rect 17253 619 17287 987
rect 17545 2195 18791 2229
rect 17449 1165 17483 2133
rect 18853 1165 18887 2133
rect 17545 1069 18791 1103
rect 17449 619 17483 987
rect 18853 619 18887 987
rect 19145 2195 20391 2229
rect 19049 1165 19083 2133
rect 20453 1165 20487 2133
rect 19145 1069 20391 1103
rect 19049 619 19083 987
rect 20453 619 20487 987
rect 20745 2195 21991 2229
rect 20649 1165 20683 2133
rect 22053 1165 22087 2133
rect 20745 1069 21991 1103
rect 20649 619 20683 987
rect 22053 619 22087 987
rect 22345 2195 23591 2229
rect 22249 1165 22283 2133
rect 23653 1165 23687 2133
rect 22345 1069 23591 1103
rect 22249 619 22283 987
rect 23653 619 23687 987
rect 23945 2195 25191 2229
rect 23849 1165 23883 2133
rect 25253 1165 25287 2133
rect 23945 1069 25191 1103
rect 23849 619 23883 987
rect 25253 619 25287 987
rect 25545 2195 26791 2229
rect 25449 1165 25483 2133
rect 26853 1165 26887 2133
rect 25545 1069 26791 1103
rect 25449 619 25483 987
rect 26853 619 26887 987
rect 27145 2195 28391 2229
rect 27049 1165 27083 2133
rect 28453 1165 28487 2133
rect 27145 1069 28391 1103
rect 27049 619 27083 987
rect 28453 619 28487 987
rect 28745 2195 29991 2229
rect 28649 1165 28683 2133
rect 30053 1165 30087 2133
rect 28745 1069 29991 1103
rect 28649 619 28683 987
rect 30053 619 30087 987
rect 30345 2195 31591 2229
rect 30249 1165 30283 2133
rect 31653 1165 31687 2133
rect 30345 1069 31591 1103
rect 30249 619 30283 987
rect 31653 619 31687 987
rect 31945 2195 33191 2229
rect 31849 1165 31883 2133
rect 33253 1165 33287 2133
rect 31945 1069 33191 1103
rect 31849 619 31883 987
rect 33253 619 33287 987
rect 33545 2195 34791 2229
rect 33449 1165 33483 2133
rect 34853 1165 34887 2133
rect 33545 1069 34791 1103
rect 33449 619 33483 987
rect 34853 619 34887 987
rect 35145 2195 36391 2229
rect 35049 1165 35083 2133
rect 36453 1165 36487 2133
rect 35145 1069 36391 1103
rect 35049 619 35083 987
rect 36453 619 36487 987
rect 36745 2195 37991 2229
rect 36649 1165 36683 2133
rect 38053 1165 38087 2133
rect 36745 1069 37991 1103
rect 36649 619 36683 987
rect 38053 619 38087 987
rect -55 395 1191 429
rect -151 -635 -117 333
rect 1253 -635 1287 333
rect -55 -731 1191 -697
rect -151 -1181 -117 -813
rect 1253 -1181 1287 -813
rect 1545 395 2791 429
rect 1449 -635 1483 333
rect 2853 -635 2887 333
rect 1545 -731 2791 -697
rect 1449 -1181 1483 -813
rect 2853 -1181 2887 -813
rect 3145 395 4391 429
rect 3049 -635 3083 333
rect 4453 -635 4487 333
rect 3145 -731 4391 -697
rect 3049 -1181 3083 -813
rect 4453 -1181 4487 -813
rect 4745 395 5991 429
rect 4649 -635 4683 333
rect 6053 -635 6087 333
rect 4745 -731 5991 -697
rect 4649 -1181 4683 -813
rect 6053 -1181 6087 -813
rect 6345 395 7591 429
rect 6249 -635 6283 333
rect 7653 -635 7687 333
rect 6345 -731 7591 -697
rect 6249 -1181 6283 -813
rect 7653 -1181 7687 -813
rect 7945 395 9191 429
rect 7849 -635 7883 333
rect 9253 -635 9287 333
rect 7945 -731 9191 -697
rect 7849 -1181 7883 -813
rect 9253 -1181 9287 -813
rect 9545 395 10791 429
rect 9449 -635 9483 333
rect 10853 -635 10887 333
rect 9545 -731 10791 -697
rect 9449 -1181 9483 -813
rect 10853 -1181 10887 -813
rect 11145 395 12391 429
rect 11049 -635 11083 333
rect 12453 -635 12487 333
rect 11145 -731 12391 -697
rect 11049 -1181 11083 -813
rect 12453 -1181 12487 -813
rect 12745 395 13991 429
rect 12649 -635 12683 333
rect 14053 -635 14087 333
rect 12745 -731 13991 -697
rect 12649 -1181 12683 -813
rect 14053 -1181 14087 -813
rect 14345 395 15591 429
rect 14249 -635 14283 333
rect 15653 -635 15687 333
rect 14345 -731 15591 -697
rect 14249 -1181 14283 -813
rect 15653 -1181 15687 -813
rect 15945 395 17191 429
rect 15849 -635 15883 333
rect 17253 -635 17287 333
rect 15945 -731 17191 -697
rect 15849 -1181 15883 -813
rect 17253 -1181 17287 -813
rect 17545 395 18791 429
rect 17449 -635 17483 333
rect 18853 -635 18887 333
rect 17545 -731 18791 -697
rect 17449 -1181 17483 -813
rect 18853 -1181 18887 -813
rect 19145 395 20391 429
rect 19049 -635 19083 333
rect 20453 -635 20487 333
rect 19145 -731 20391 -697
rect 19049 -1181 19083 -813
rect 20453 -1181 20487 -813
rect 20745 395 21991 429
rect 20649 -635 20683 333
rect 22053 -635 22087 333
rect 20745 -731 21991 -697
rect 20649 -1181 20683 -813
rect 22053 -1181 22087 -813
rect 22345 395 23591 429
rect 22249 -635 22283 333
rect 23653 -635 23687 333
rect 22345 -731 23591 -697
rect 22249 -1181 22283 -813
rect 23653 -1181 23687 -813
rect 23945 395 25191 429
rect 23849 -635 23883 333
rect 25253 -635 25287 333
rect 23945 -731 25191 -697
rect 23849 -1181 23883 -813
rect 25253 -1181 25287 -813
rect 25545 395 26791 429
rect 25449 -635 25483 333
rect 26853 -635 26887 333
rect 25545 -731 26791 -697
rect 25449 -1181 25483 -813
rect 26853 -1181 26887 -813
rect 27145 395 28391 429
rect 27049 -635 27083 333
rect 28453 -635 28487 333
rect 27145 -731 28391 -697
rect 27049 -1181 27083 -813
rect 28453 -1181 28487 -813
rect 28745 395 29991 429
rect 28649 -635 28683 333
rect 30053 -635 30087 333
rect 28745 -731 29991 -697
rect 28649 -1181 28683 -813
rect 30053 -1181 30087 -813
rect 30345 395 31591 429
rect 30249 -635 30283 333
rect 31653 -635 31687 333
rect 30345 -731 31591 -697
rect 30249 -1181 30283 -813
rect 31653 -1181 31687 -813
rect 31945 395 33191 429
rect 31849 -635 31883 333
rect 33253 -635 33287 333
rect 31945 -731 33191 -697
rect 31849 -1181 31883 -813
rect 33253 -1181 33287 -813
rect 33545 395 34791 429
rect 33449 -635 33483 333
rect 34853 -635 34887 333
rect 33545 -731 34791 -697
rect 33449 -1181 33483 -813
rect 34853 -1181 34887 -813
rect 35145 395 36391 429
rect 35049 -635 35083 333
rect 36453 -635 36487 333
rect 35145 -731 36391 -697
rect 35049 -1181 35083 -813
rect 36453 -1181 36487 -813
rect 36745 395 37991 429
rect 36649 -635 36683 333
rect 38053 -635 38087 333
rect 36745 -731 37991 -697
rect 36649 -1181 36683 -813
rect 38053 -1181 38087 -813
rect -55 -1405 1191 -1371
rect -151 -2435 -117 -1467
rect 1253 -2435 1287 -1467
rect -55 -2531 1191 -2497
rect -151 -2981 -117 -2613
rect 1253 -2981 1287 -2613
rect 1545 -1405 2791 -1371
rect 1449 -2435 1483 -1467
rect 2853 -2435 2887 -1467
rect 1545 -2531 2791 -2497
rect 1449 -2981 1483 -2613
rect 2853 -2981 2887 -2613
rect 3145 -1405 4391 -1371
rect 3049 -2435 3083 -1467
rect 4453 -2435 4487 -1467
rect 3145 -2531 4391 -2497
rect 3049 -2981 3083 -2613
rect 4453 -2981 4487 -2613
rect 4745 -1405 5991 -1371
rect 4649 -2435 4683 -1467
rect 6053 -2435 6087 -1467
rect 4745 -2531 5991 -2497
rect 4649 -2981 4683 -2613
rect 6053 -2981 6087 -2613
rect 6345 -1405 7591 -1371
rect 6249 -2435 6283 -1467
rect 7653 -2435 7687 -1467
rect 6345 -2531 7591 -2497
rect 6249 -2981 6283 -2613
rect 7653 -2981 7687 -2613
rect 7945 -1405 9191 -1371
rect 7849 -2435 7883 -1467
rect 9253 -2435 9287 -1467
rect 7945 -2531 9191 -2497
rect 7849 -2981 7883 -2613
rect 9253 -2981 9287 -2613
rect 9545 -1405 10791 -1371
rect 9449 -2435 9483 -1467
rect 10853 -2435 10887 -1467
rect 9545 -2531 10791 -2497
rect 9449 -2981 9483 -2613
rect 10853 -2981 10887 -2613
rect 11145 -1405 12391 -1371
rect 11049 -2435 11083 -1467
rect 12453 -2435 12487 -1467
rect 11145 -2531 12391 -2497
rect 11049 -2981 11083 -2613
rect 12453 -2981 12487 -2613
rect 12745 -1405 13991 -1371
rect 12649 -2435 12683 -1467
rect 14053 -2435 14087 -1467
rect 12745 -2531 13991 -2497
rect 12649 -2981 12683 -2613
rect 14053 -2981 14087 -2613
rect 14345 -1405 15591 -1371
rect 14249 -2435 14283 -1467
rect 15653 -2435 15687 -1467
rect 14345 -2531 15591 -2497
rect 14249 -2981 14283 -2613
rect 15653 -2981 15687 -2613
rect 15945 -1405 17191 -1371
rect 15849 -2435 15883 -1467
rect 17253 -2435 17287 -1467
rect 15945 -2531 17191 -2497
rect 15849 -2981 15883 -2613
rect 17253 -2981 17287 -2613
rect 17545 -1405 18791 -1371
rect 17449 -2435 17483 -1467
rect 18853 -2435 18887 -1467
rect 17545 -2531 18791 -2497
rect 17449 -2981 17483 -2613
rect 18853 -2981 18887 -2613
rect 19145 -1405 20391 -1371
rect 19049 -2435 19083 -1467
rect 20453 -2435 20487 -1467
rect 19145 -2531 20391 -2497
rect 19049 -2981 19083 -2613
rect 20453 -2981 20487 -2613
rect 20745 -1405 21991 -1371
rect 20649 -2435 20683 -1467
rect 22053 -2435 22087 -1467
rect 20745 -2531 21991 -2497
rect 20649 -2981 20683 -2613
rect 22053 -2981 22087 -2613
rect 22345 -1405 23591 -1371
rect 22249 -2435 22283 -1467
rect 23653 -2435 23687 -1467
rect 22345 -2531 23591 -2497
rect 22249 -2981 22283 -2613
rect 23653 -2981 23687 -2613
rect 23945 -1405 25191 -1371
rect 23849 -2435 23883 -1467
rect 25253 -2435 25287 -1467
rect 23945 -2531 25191 -2497
rect 23849 -2981 23883 -2613
rect 25253 -2981 25287 -2613
rect 25545 -1405 26791 -1371
rect 25449 -2435 25483 -1467
rect 26853 -2435 26887 -1467
rect 25545 -2531 26791 -2497
rect 25449 -2981 25483 -2613
rect 26853 -2981 26887 -2613
rect 27145 -1405 28391 -1371
rect 27049 -2435 27083 -1467
rect 28453 -2435 28487 -1467
rect 27145 -2531 28391 -2497
rect 27049 -2981 27083 -2613
rect 28453 -2981 28487 -2613
rect 28745 -1405 29991 -1371
rect 28649 -2435 28683 -1467
rect 30053 -2435 30087 -1467
rect 28745 -2531 29991 -2497
rect 28649 -2981 28683 -2613
rect 30053 -2981 30087 -2613
rect 30345 -1405 31591 -1371
rect 30249 -2435 30283 -1467
rect 31653 -2435 31687 -1467
rect 30345 -2531 31591 -2497
rect 30249 -2981 30283 -2613
rect 31653 -2981 31687 -2613
rect 31945 -1405 33191 -1371
rect 31849 -2435 31883 -1467
rect 33253 -2435 33287 -1467
rect 31945 -2531 33191 -2497
rect 31849 -2981 31883 -2613
rect 33253 -2981 33287 -2613
rect 33545 -1405 34791 -1371
rect 33449 -2435 33483 -1467
rect 34853 -2435 34887 -1467
rect 33545 -2531 34791 -2497
rect 33449 -2981 33483 -2613
rect 34853 -2981 34887 -2613
rect 35145 -1405 36391 -1371
rect 35049 -2435 35083 -1467
rect 36453 -2435 36487 -1467
rect 35145 -2531 36391 -2497
rect 35049 -2981 35083 -2613
rect 36453 -2981 36487 -2613
rect 36745 -1405 37991 -1371
rect 36649 -2435 36683 -1467
rect 38053 -2435 38087 -1467
rect 36745 -2531 37991 -2497
rect 36649 -2981 36683 -2613
rect 38053 -2981 38087 -2613
rect -55 -3205 1191 -3171
rect -151 -4235 -117 -3267
rect 1253 -4235 1287 -3267
rect -55 -4331 1191 -4297
rect -151 -4781 -117 -4413
rect 1253 -4781 1287 -4413
rect 1545 -3205 2791 -3171
rect 1449 -4235 1483 -3267
rect 2853 -4235 2887 -3267
rect 1545 -4331 2791 -4297
rect 1449 -4781 1483 -4413
rect 2853 -4781 2887 -4413
rect 3145 -3205 4391 -3171
rect 3049 -4235 3083 -3267
rect 4453 -4235 4487 -3267
rect 3145 -4331 4391 -4297
rect 3049 -4781 3083 -4413
rect 4453 -4781 4487 -4413
rect 4745 -3205 5991 -3171
rect 4649 -4235 4683 -3267
rect 6053 -4235 6087 -3267
rect 4745 -4331 5991 -4297
rect 4649 -4781 4683 -4413
rect 6053 -4781 6087 -4413
rect 6345 -3205 7591 -3171
rect 6249 -4235 6283 -3267
rect 7653 -4235 7687 -3267
rect 6345 -4331 7591 -4297
rect 6249 -4781 6283 -4413
rect 7653 -4781 7687 -4413
rect 7945 -3205 9191 -3171
rect 7849 -4235 7883 -3267
rect 9253 -4235 9287 -3267
rect 7945 -4331 9191 -4297
rect 7849 -4781 7883 -4413
rect 9253 -4781 9287 -4413
rect 9545 -3205 10791 -3171
rect 9449 -4235 9483 -3267
rect 10853 -4235 10887 -3267
rect 9545 -4331 10791 -4297
rect 9449 -4781 9483 -4413
rect 10853 -4781 10887 -4413
rect 11145 -3205 12391 -3171
rect 11049 -4235 11083 -3267
rect 12453 -4235 12487 -3267
rect 11145 -4331 12391 -4297
rect 11049 -4781 11083 -4413
rect 12453 -4781 12487 -4413
rect 12745 -3205 13991 -3171
rect 12649 -4235 12683 -3267
rect 14053 -4235 14087 -3267
rect 12745 -4331 13991 -4297
rect 12649 -4781 12683 -4413
rect 14053 -4781 14087 -4413
rect 14345 -3205 15591 -3171
rect 14249 -4235 14283 -3267
rect 15653 -4235 15687 -3267
rect 14345 -4331 15591 -4297
rect 14249 -4781 14283 -4413
rect 15653 -4781 15687 -4413
rect 15945 -3205 17191 -3171
rect 15849 -4235 15883 -3267
rect 17253 -4235 17287 -3267
rect 15945 -4331 17191 -4297
rect 15849 -4781 15883 -4413
rect 17253 -4781 17287 -4413
rect 17545 -3205 18791 -3171
rect 17449 -4235 17483 -3267
rect 18853 -4235 18887 -3267
rect 17545 -4331 18791 -4297
rect 17449 -4781 17483 -4413
rect 18853 -4781 18887 -4413
rect 19145 -3205 20391 -3171
rect 19049 -4235 19083 -3267
rect 20453 -4235 20487 -3267
rect 19145 -4331 20391 -4297
rect 19049 -4781 19083 -4413
rect 20453 -4781 20487 -4413
rect 20745 -3205 21991 -3171
rect 20649 -4235 20683 -3267
rect 22053 -4235 22087 -3267
rect 20745 -4331 21991 -4297
rect 20649 -4781 20683 -4413
rect 22053 -4781 22087 -4413
rect 22345 -3205 23591 -3171
rect 22249 -4235 22283 -3267
rect 23653 -4235 23687 -3267
rect 22345 -4331 23591 -4297
rect 22249 -4781 22283 -4413
rect 23653 -4781 23687 -4413
rect 23945 -3205 25191 -3171
rect 23849 -4235 23883 -3267
rect 25253 -4235 25287 -3267
rect 23945 -4331 25191 -4297
rect 23849 -4781 23883 -4413
rect 25253 -4781 25287 -4413
rect 25545 -3205 26791 -3171
rect 25449 -4235 25483 -3267
rect 26853 -4235 26887 -3267
rect 25545 -4331 26791 -4297
rect 25449 -4781 25483 -4413
rect 26853 -4781 26887 -4413
rect 27145 -3205 28391 -3171
rect 27049 -4235 27083 -3267
rect 28453 -4235 28487 -3267
rect 27145 -4331 28391 -4297
rect 27049 -4781 27083 -4413
rect 28453 -4781 28487 -4413
rect 28745 -3205 29991 -3171
rect 28649 -4235 28683 -3267
rect 30053 -4235 30087 -3267
rect 28745 -4331 29991 -4297
rect 28649 -4781 28683 -4413
rect 30053 -4781 30087 -4413
rect 30345 -3205 31591 -3171
rect 30249 -4235 30283 -3267
rect 31653 -4235 31687 -3267
rect 30345 -4331 31591 -4297
rect 30249 -4781 30283 -4413
rect 31653 -4781 31687 -4413
rect 31945 -3205 33191 -3171
rect 31849 -4235 31883 -3267
rect 33253 -4235 33287 -3267
rect 31945 -4331 33191 -4297
rect 31849 -4781 31883 -4413
rect 33253 -4781 33287 -4413
rect 33545 -3205 34791 -3171
rect 33449 -4235 33483 -3267
rect 34853 -4235 34887 -3267
rect 33545 -4331 34791 -4297
rect 33449 -4781 33483 -4413
rect 34853 -4781 34887 -4413
rect 35145 -3205 36391 -3171
rect 35049 -4235 35083 -3267
rect 36453 -4235 36487 -3267
rect 35145 -4331 36391 -4297
rect 35049 -4781 35083 -4413
rect 36453 -4781 36487 -4413
rect 36745 -3205 37991 -3171
rect 36649 -4235 36683 -3267
rect 38053 -4235 38087 -3267
rect 36745 -4331 37991 -4297
rect 36649 -4781 36683 -4413
rect 38053 -4781 38087 -4413
rect 27884 -24536 28852 -24502
rect 27788 -25226 27822 -24598
rect 28914 -25226 28948 -24598
rect 27884 -25322 28852 -25288
rect 27884 -25442 28850 -25408
rect 27788 -26246 27822 -25504
rect 28912 -26246 28946 -25504
rect 27884 -26342 28850 -26308
rect 27884 -26482 28850 -26448
rect 27788 -27286 27822 -26544
rect 28912 -27286 28946 -26544
rect 27884 -27382 28850 -27348
rect 27884 -27522 28850 -27488
rect 27788 -28326 27822 -27584
rect 28912 -28326 28946 -27584
rect 27884 -28422 28850 -28388
rect 27884 -28562 28850 -28528
rect 27788 -29366 27822 -28624
rect 28912 -29366 28946 -28624
rect 27884 -29462 28850 -29428
rect 31775 -29365 32043 -29331
rect 32215 -29365 32483 -29331
rect 32655 -29365 32923 -29331
rect 33094 -29365 33678 -29331
rect 27884 -29602 28850 -29568
rect 27788 -30406 27822 -29664
rect 28912 -30406 28946 -29664
rect 31679 -29855 31713 -29427
rect 32105 -29855 32139 -29427
rect 32998 -29855 33032 -29427
rect 33740 -29855 33774 -29427
rect 31775 -29951 32043 -29917
rect 32215 -29951 32483 -29917
rect 32655 -29951 32923 -29917
rect 33094 -29951 33678 -29917
rect 33975 -29365 34243 -29331
rect 34415 -29365 34683 -29331
rect 34855 -29365 35123 -29331
rect 35294 -29365 35878 -29331
rect 33879 -29855 33913 -29427
rect 34305 -29855 34339 -29427
rect 35198 -29855 35232 -29427
rect 35940 -29855 35974 -29427
rect 33975 -29951 34243 -29917
rect 34415 -29951 34683 -29917
rect 34855 -29951 35123 -29917
rect 35294 -29951 35878 -29917
rect 36175 -29365 36443 -29331
rect 36615 -29365 36883 -29331
rect 37055 -29365 37323 -29331
rect 37494 -29365 38078 -29331
rect 36079 -29855 36113 -29427
rect 36505 -29855 36539 -29427
rect 37398 -29855 37432 -29427
rect 38140 -29855 38174 -29427
rect 36175 -29951 36443 -29917
rect 36615 -29951 36883 -29917
rect 37055 -29951 37323 -29917
rect 37494 -29951 38078 -29917
rect 27884 -30502 28850 -30468
rect 31744 -30107 32328 -30073
rect 32499 -30107 32767 -30073
rect 32939 -30107 33207 -30073
rect 33379 -30107 33647 -30073
rect 27884 -30642 28850 -30608
rect 27788 -31446 27822 -30704
rect 28912 -31446 28946 -30704
rect 31648 -30597 31682 -30169
rect 32390 -30597 32424 -30169
rect 33283 -30597 33317 -30169
rect 33709 -30597 33743 -30169
rect 31744 -30693 32328 -30659
rect 32499 -30693 32767 -30659
rect 32939 -30693 33207 -30659
rect 33379 -30693 33647 -30659
rect 33944 -30107 34528 -30073
rect 34699 -30107 34967 -30073
rect 35139 -30107 35407 -30073
rect 35579 -30107 35847 -30073
rect 33848 -30597 33882 -30169
rect 34590 -30597 34624 -30169
rect 35483 -30597 35517 -30169
rect 35909 -30597 35943 -30169
rect 33944 -30693 34528 -30659
rect 34699 -30693 34967 -30659
rect 35139 -30693 35407 -30659
rect 35579 -30693 35847 -30659
rect 36144 -30107 36728 -30073
rect 36899 -30107 37167 -30073
rect 37339 -30107 37607 -30073
rect 37779 -30107 38047 -30073
rect 36048 -30597 36082 -30169
rect 36790 -30597 36824 -30169
rect 37683 -30597 37717 -30169
rect 38109 -30597 38143 -30169
rect 36144 -30693 36728 -30659
rect 36899 -30693 37167 -30659
rect 37339 -30693 37607 -30659
rect 37779 -30693 38047 -30659
rect 27884 -31542 28850 -31508
<< mvnsubdiffcont >>
rect 27874 11558 28850 11592
rect 27778 10754 27812 11496
rect 28912 10754 28946 11496
rect 27874 10658 28850 10692
rect 30106 11092 30674 11126
rect 30820 11092 31088 11126
rect 31260 11092 31528 11126
rect 31700 11092 31968 11126
rect 30010 10684 30044 11030
rect 30736 10684 30770 11030
rect 30106 10588 30674 10622
rect 27874 10518 28850 10552
rect 27778 9714 27812 10456
rect 28912 9714 28946 10456
rect 31604 10384 31638 11030
rect 32030 10384 32064 11030
rect 32306 11092 32874 11126
rect 33020 11092 33288 11126
rect 33460 11092 33728 11126
rect 33900 11092 34168 11126
rect 32210 10684 32244 11030
rect 32936 10684 32970 11030
rect 32306 10588 32874 10622
rect 30820 10288 31088 10322
rect 31260 10288 31528 10322
rect 31700 10288 31968 10322
rect 33804 10384 33838 11030
rect 34230 10384 34264 11030
rect 34506 11092 35074 11126
rect 35220 11092 35488 11126
rect 35660 11092 35928 11126
rect 36100 11092 36368 11126
rect 34410 10684 34444 11030
rect 35136 10684 35170 11030
rect 34506 10588 35074 10622
rect 33020 10288 33288 10322
rect 33460 10288 33728 10322
rect 33900 10288 34168 10322
rect 36004 10384 36038 11030
rect 36430 10384 36464 11030
rect 35220 10288 35488 10322
rect 35660 10288 35928 10322
rect 36100 10288 36368 10322
rect 27874 9618 28850 9652
rect 29694 9782 31520 9816
rect 27874 9478 28850 9512
rect 27778 8674 27812 9416
rect 28912 8674 28946 9416
rect 29598 9074 29632 9720
rect 31582 9074 31616 9720
rect 29694 8978 31520 9012
rect 27874 8578 28850 8612
rect 29694 8778 31520 8812
rect 27874 8438 28850 8472
rect 27778 7634 27812 8376
rect 28912 7634 28946 8376
rect 27874 7538 28850 7572
rect 27874 7398 28850 7432
rect 27778 6594 27812 7336
rect 28912 6594 28946 7336
rect 29598 7434 29632 8716
rect 31582 7434 31616 8716
rect 29694 7338 31520 7372
rect 29538 6734 29572 7102
rect 30742 6734 30776 7102
rect 30878 6734 30912 7102
rect 32082 6734 32116 7102
rect 27874 6498 28850 6532
rect 27874 6358 28850 6392
rect 27778 5554 27812 6296
rect 28912 5554 28946 6296
rect 27874 5458 28850 5492
rect 27874 5342 28842 5376
rect 27778 4234 27812 5280
rect 28904 4234 28938 5280
rect 27874 4138 28842 4172
rect -66 -8070 1216 -8036
rect -162 -8500 -128 -8132
rect 1278 -8500 1312 -8132
rect -66 -8596 1216 -8562
rect -162 -9626 -128 -8658
rect 1278 -9626 1312 -8658
rect -66 -9722 1216 -9688
rect 1534 -8070 2816 -8036
rect 1438 -8500 1472 -8132
rect 2878 -8500 2912 -8132
rect 1534 -8596 2816 -8562
rect 1438 -9626 1472 -8658
rect 2878 -9626 2912 -8658
rect 1534 -9722 2816 -9688
rect 3134 -8070 4416 -8036
rect 3038 -8500 3072 -8132
rect 4478 -8500 4512 -8132
rect 3134 -8596 4416 -8562
rect 3038 -9626 3072 -8658
rect 4478 -9626 4512 -8658
rect 3134 -9722 4416 -9688
rect 4734 -8070 6016 -8036
rect 4638 -8500 4672 -8132
rect 6078 -8500 6112 -8132
rect 4734 -8596 6016 -8562
rect 4638 -9626 4672 -8658
rect 6078 -9626 6112 -8658
rect 4734 -9722 6016 -9688
rect 6334 -8070 7616 -8036
rect 6238 -8500 6272 -8132
rect 7678 -8500 7712 -8132
rect 6334 -8596 7616 -8562
rect 6238 -9626 6272 -8658
rect 7678 -9626 7712 -8658
rect 6334 -9722 7616 -9688
rect 7934 -8070 9216 -8036
rect 7838 -8500 7872 -8132
rect 9278 -8500 9312 -8132
rect 7934 -8596 9216 -8562
rect 7838 -9626 7872 -8658
rect 9278 -9626 9312 -8658
rect 7934 -9722 9216 -9688
rect 9534 -8070 10816 -8036
rect 9438 -8500 9472 -8132
rect 10878 -8500 10912 -8132
rect 9534 -8596 10816 -8562
rect 9438 -9626 9472 -8658
rect 10878 -9626 10912 -8658
rect 9534 -9722 10816 -9688
rect 11134 -8070 12416 -8036
rect 11038 -8500 11072 -8132
rect 12478 -8500 12512 -8132
rect 11134 -8596 12416 -8562
rect 11038 -9626 11072 -8658
rect 12478 -9626 12512 -8658
rect 11134 -9722 12416 -9688
rect 12734 -8070 14016 -8036
rect 12638 -8500 12672 -8132
rect 14078 -8500 14112 -8132
rect 12734 -8596 14016 -8562
rect 12638 -9626 12672 -8658
rect 14078 -9626 14112 -8658
rect 12734 -9722 14016 -9688
rect 14334 -8070 15616 -8036
rect 14238 -8500 14272 -8132
rect 15678 -8500 15712 -8132
rect 14334 -8596 15616 -8562
rect 14238 -9626 14272 -8658
rect 15678 -9626 15712 -8658
rect 14334 -9722 15616 -9688
rect 15934 -8070 17216 -8036
rect 15838 -8500 15872 -8132
rect 17278 -8500 17312 -8132
rect 15934 -8596 17216 -8562
rect 15838 -9626 15872 -8658
rect 17278 -9626 17312 -8658
rect 15934 -9722 17216 -9688
rect 17534 -8070 18816 -8036
rect 17438 -8500 17472 -8132
rect 18878 -8500 18912 -8132
rect 17534 -8596 18816 -8562
rect 17438 -9626 17472 -8658
rect 18878 -9626 18912 -8658
rect 17534 -9722 18816 -9688
rect 19134 -8070 20416 -8036
rect 19038 -8500 19072 -8132
rect 20478 -8500 20512 -8132
rect 19134 -8596 20416 -8562
rect 19038 -9626 19072 -8658
rect 20478 -9626 20512 -8658
rect 19134 -9722 20416 -9688
rect 20734 -8070 22016 -8036
rect 20638 -8500 20672 -8132
rect 22078 -8500 22112 -8132
rect 20734 -8596 22016 -8562
rect 20638 -9626 20672 -8658
rect 22078 -9626 22112 -8658
rect 20734 -9722 22016 -9688
rect 22334 -8070 23616 -8036
rect 22238 -8500 22272 -8132
rect 23678 -8500 23712 -8132
rect 22334 -8596 23616 -8562
rect 22238 -9626 22272 -8658
rect 23678 -9626 23712 -8658
rect 22334 -9722 23616 -9688
rect 23934 -8070 25216 -8036
rect 23838 -8500 23872 -8132
rect 25278 -8500 25312 -8132
rect 23934 -8596 25216 -8562
rect 23838 -9626 23872 -8658
rect 25278 -9626 25312 -8658
rect 23934 -9722 25216 -9688
rect 25534 -8070 26816 -8036
rect 25438 -8500 25472 -8132
rect 26878 -8500 26912 -8132
rect 25534 -8596 26816 -8562
rect 25438 -9626 25472 -8658
rect 26878 -9626 26912 -8658
rect 25534 -9722 26816 -9688
rect 27134 -8070 28416 -8036
rect 27038 -8500 27072 -8132
rect 28478 -8500 28512 -8132
rect 27134 -8596 28416 -8562
rect 27038 -9626 27072 -8658
rect 28478 -9626 28512 -8658
rect 27134 -9722 28416 -9688
rect 28734 -8070 30016 -8036
rect 28638 -8500 28672 -8132
rect 30078 -8500 30112 -8132
rect 28734 -8596 30016 -8562
rect 28638 -9626 28672 -8658
rect 30078 -9626 30112 -8658
rect 28734 -9722 30016 -9688
rect 30334 -8070 31616 -8036
rect 30238 -8500 30272 -8132
rect 31678 -8500 31712 -8132
rect 30334 -8596 31616 -8562
rect 30238 -9626 30272 -8658
rect 31678 -9626 31712 -8658
rect 30334 -9722 31616 -9688
rect 31934 -8070 33216 -8036
rect 31838 -8500 31872 -8132
rect 33278 -8500 33312 -8132
rect 31934 -8596 33216 -8562
rect 31838 -9626 31872 -8658
rect 33278 -9626 33312 -8658
rect 31934 -9722 33216 -9688
rect 33534 -8070 34816 -8036
rect 33438 -8500 33472 -8132
rect 34878 -8500 34912 -8132
rect 33534 -8596 34816 -8562
rect 33438 -9626 33472 -8658
rect 34878 -9626 34912 -8658
rect 33534 -9722 34816 -9688
rect 35134 -8070 36416 -8036
rect 35038 -8500 35072 -8132
rect 36478 -8500 36512 -8132
rect 35134 -8596 36416 -8562
rect 35038 -9626 35072 -8658
rect 36478 -9626 36512 -8658
rect 35134 -9722 36416 -9688
rect 36734 -8070 38016 -8036
rect 36638 -8500 36672 -8132
rect 38078 -8500 38112 -8132
rect 36734 -8596 38016 -8562
rect 36638 -9626 36672 -8658
rect 38078 -9626 38112 -8658
rect 36734 -9722 38016 -9688
rect -66 -9870 1216 -9836
rect -162 -10300 -128 -9932
rect 1278 -10300 1312 -9932
rect -66 -10396 1216 -10362
rect -162 -11426 -128 -10458
rect 1278 -11426 1312 -10458
rect -66 -11522 1216 -11488
rect 1534 -9870 2816 -9836
rect 1438 -10300 1472 -9932
rect 2878 -10300 2912 -9932
rect 1534 -10396 2816 -10362
rect 1438 -11426 1472 -10458
rect 2878 -11426 2912 -10458
rect 1534 -11522 2816 -11488
rect 3134 -9870 4416 -9836
rect 3038 -10300 3072 -9932
rect 4478 -10300 4512 -9932
rect 3134 -10396 4416 -10362
rect 3038 -11426 3072 -10458
rect 4478 -11426 4512 -10458
rect 3134 -11522 4416 -11488
rect 4734 -9870 6016 -9836
rect 4638 -10300 4672 -9932
rect 6078 -10300 6112 -9932
rect 4734 -10396 6016 -10362
rect 4638 -11426 4672 -10458
rect 6078 -11426 6112 -10458
rect 4734 -11522 6016 -11488
rect 6334 -9870 7616 -9836
rect 6238 -10300 6272 -9932
rect 7678 -10300 7712 -9932
rect 6334 -10396 7616 -10362
rect 6238 -11426 6272 -10458
rect 7678 -11426 7712 -10458
rect 6334 -11522 7616 -11488
rect 7934 -9870 9216 -9836
rect 7838 -10300 7872 -9932
rect 9278 -10300 9312 -9932
rect 7934 -10396 9216 -10362
rect 7838 -11426 7872 -10458
rect 9278 -11426 9312 -10458
rect 7934 -11522 9216 -11488
rect 9534 -9870 10816 -9836
rect 9438 -10300 9472 -9932
rect 10878 -10300 10912 -9932
rect 9534 -10396 10816 -10362
rect 9438 -11426 9472 -10458
rect 10878 -11426 10912 -10458
rect 9534 -11522 10816 -11488
rect 11134 -9870 12416 -9836
rect 11038 -10300 11072 -9932
rect 12478 -10300 12512 -9932
rect 11134 -10396 12416 -10362
rect 11038 -11426 11072 -10458
rect 12478 -11426 12512 -10458
rect 11134 -11522 12416 -11488
rect 12734 -9870 14016 -9836
rect 12638 -10300 12672 -9932
rect 14078 -10300 14112 -9932
rect 12734 -10396 14016 -10362
rect 12638 -11426 12672 -10458
rect 14078 -11426 14112 -10458
rect 12734 -11522 14016 -11488
rect 14334 -9870 15616 -9836
rect 14238 -10300 14272 -9932
rect 15678 -10300 15712 -9932
rect 14334 -10396 15616 -10362
rect 14238 -11426 14272 -10458
rect 15678 -11426 15712 -10458
rect 14334 -11522 15616 -11488
rect 15934 -9870 17216 -9836
rect 15838 -10300 15872 -9932
rect 17278 -10300 17312 -9932
rect 15934 -10396 17216 -10362
rect 15838 -11426 15872 -10458
rect 17278 -11426 17312 -10458
rect 15934 -11522 17216 -11488
rect 17534 -9870 18816 -9836
rect 17438 -10300 17472 -9932
rect 18878 -10300 18912 -9932
rect 17534 -10396 18816 -10362
rect 17438 -11426 17472 -10458
rect 18878 -11426 18912 -10458
rect 17534 -11522 18816 -11488
rect 19134 -9870 20416 -9836
rect 19038 -10300 19072 -9932
rect 20478 -10300 20512 -9932
rect 19134 -10396 20416 -10362
rect 19038 -11426 19072 -10458
rect 20478 -11426 20512 -10458
rect 19134 -11522 20416 -11488
rect 20734 -9870 22016 -9836
rect 20638 -10300 20672 -9932
rect 22078 -10300 22112 -9932
rect 20734 -10396 22016 -10362
rect 20638 -11426 20672 -10458
rect 22078 -11426 22112 -10458
rect 20734 -11522 22016 -11488
rect 22334 -9870 23616 -9836
rect 22238 -10300 22272 -9932
rect 23678 -10300 23712 -9932
rect 22334 -10396 23616 -10362
rect 22238 -11426 22272 -10458
rect 23678 -11426 23712 -10458
rect 22334 -11522 23616 -11488
rect 23934 -9870 25216 -9836
rect 23838 -10300 23872 -9932
rect 25278 -10300 25312 -9932
rect 23934 -10396 25216 -10362
rect 23838 -11426 23872 -10458
rect 25278 -11426 25312 -10458
rect 23934 -11522 25216 -11488
rect 25534 -9870 26816 -9836
rect 25438 -10300 25472 -9932
rect 26878 -10300 26912 -9932
rect 25534 -10396 26816 -10362
rect 25438 -11426 25472 -10458
rect 26878 -11426 26912 -10458
rect 25534 -11522 26816 -11488
rect 27134 -9870 28416 -9836
rect 27038 -10300 27072 -9932
rect 28478 -10300 28512 -9932
rect 27134 -10396 28416 -10362
rect 27038 -11426 27072 -10458
rect 28478 -11426 28512 -10458
rect 27134 -11522 28416 -11488
rect 28734 -9870 30016 -9836
rect 28638 -10300 28672 -9932
rect 30078 -10300 30112 -9932
rect 28734 -10396 30016 -10362
rect 28638 -11426 28672 -10458
rect 30078 -11426 30112 -10458
rect 28734 -11522 30016 -11488
rect 30334 -9870 31616 -9836
rect 30238 -10300 30272 -9932
rect 31678 -10300 31712 -9932
rect 30334 -10396 31616 -10362
rect 30238 -11426 30272 -10458
rect 31678 -11426 31712 -10458
rect 30334 -11522 31616 -11488
rect 31934 -9870 33216 -9836
rect 31838 -10300 31872 -9932
rect 33278 -10300 33312 -9932
rect 31934 -10396 33216 -10362
rect 31838 -11426 31872 -10458
rect 33278 -11426 33312 -10458
rect 31934 -11522 33216 -11488
rect 33534 -9870 34816 -9836
rect 33438 -10300 33472 -9932
rect 34878 -10300 34912 -9932
rect 33534 -10396 34816 -10362
rect 33438 -11426 33472 -10458
rect 34878 -11426 34912 -10458
rect 33534 -11522 34816 -11488
rect 35134 -9870 36416 -9836
rect 35038 -10300 35072 -9932
rect 36478 -10300 36512 -9932
rect 35134 -10396 36416 -10362
rect 35038 -11426 35072 -10458
rect 36478 -11426 36512 -10458
rect 35134 -11522 36416 -11488
rect 36734 -9870 38016 -9836
rect 36638 -10300 36672 -9932
rect 38078 -10300 38112 -9932
rect 36734 -10396 38016 -10362
rect 36638 -11426 36672 -10458
rect 38078 -11426 38112 -10458
rect 36734 -11522 38016 -11488
rect -66 -11670 1216 -11636
rect -162 -12100 -128 -11732
rect 1278 -12100 1312 -11732
rect -66 -12196 1216 -12162
rect -162 -13226 -128 -12258
rect 1278 -13226 1312 -12258
rect -66 -13322 1216 -13288
rect 1534 -11670 2816 -11636
rect 1438 -12100 1472 -11732
rect 2878 -12100 2912 -11732
rect 1534 -12196 2816 -12162
rect 1438 -13226 1472 -12258
rect 2878 -13226 2912 -12258
rect 1534 -13322 2816 -13288
rect 3134 -11670 4416 -11636
rect 3038 -12100 3072 -11732
rect 4478 -12100 4512 -11732
rect 3134 -12196 4416 -12162
rect 3038 -13226 3072 -12258
rect 4478 -13226 4512 -12258
rect 3134 -13322 4416 -13288
rect 4734 -11670 6016 -11636
rect 4638 -12100 4672 -11732
rect 6078 -12100 6112 -11732
rect 4734 -12196 6016 -12162
rect 4638 -13226 4672 -12258
rect 6078 -13226 6112 -12258
rect 4734 -13322 6016 -13288
rect 6334 -11670 7616 -11636
rect 6238 -12100 6272 -11732
rect 7678 -12100 7712 -11732
rect 6334 -12196 7616 -12162
rect 6238 -13226 6272 -12258
rect 7678 -13226 7712 -12258
rect 6334 -13322 7616 -13288
rect 7934 -11670 9216 -11636
rect 7838 -12100 7872 -11732
rect 9278 -12100 9312 -11732
rect 7934 -12196 9216 -12162
rect 7838 -13226 7872 -12258
rect 9278 -13226 9312 -12258
rect 7934 -13322 9216 -13288
rect 9534 -11670 10816 -11636
rect 9438 -12100 9472 -11732
rect 10878 -12100 10912 -11732
rect 9534 -12196 10816 -12162
rect 9438 -13226 9472 -12258
rect 10878 -13226 10912 -12258
rect 9534 -13322 10816 -13288
rect 11134 -11670 12416 -11636
rect 11038 -12100 11072 -11732
rect 12478 -12100 12512 -11732
rect 11134 -12196 12416 -12162
rect 11038 -13226 11072 -12258
rect 12478 -13226 12512 -12258
rect 11134 -13322 12416 -13288
rect 12734 -11670 14016 -11636
rect 12638 -12100 12672 -11732
rect 14078 -12100 14112 -11732
rect 12734 -12196 14016 -12162
rect 12638 -13226 12672 -12258
rect 14078 -13226 14112 -12258
rect 12734 -13322 14016 -13288
rect 14334 -11670 15616 -11636
rect 14238 -12100 14272 -11732
rect 15678 -12100 15712 -11732
rect 14334 -12196 15616 -12162
rect 14238 -13226 14272 -12258
rect 15678 -13226 15712 -12258
rect 14334 -13322 15616 -13288
rect 15934 -11670 17216 -11636
rect 15838 -12100 15872 -11732
rect 17278 -12100 17312 -11732
rect 15934 -12196 17216 -12162
rect 15838 -13226 15872 -12258
rect 17278 -13226 17312 -12258
rect 15934 -13322 17216 -13288
rect 17534 -11670 18816 -11636
rect 17438 -12100 17472 -11732
rect 18878 -12100 18912 -11732
rect 17534 -12196 18816 -12162
rect 17438 -13226 17472 -12258
rect 18878 -13226 18912 -12258
rect 17534 -13322 18816 -13288
rect 19134 -11670 20416 -11636
rect 19038 -12100 19072 -11732
rect 20478 -12100 20512 -11732
rect 19134 -12196 20416 -12162
rect 19038 -13226 19072 -12258
rect 20478 -13226 20512 -12258
rect 19134 -13322 20416 -13288
rect 20734 -11670 22016 -11636
rect 20638 -12100 20672 -11732
rect 22078 -12100 22112 -11732
rect 20734 -12196 22016 -12162
rect 20638 -13226 20672 -12258
rect 22078 -13226 22112 -12258
rect 20734 -13322 22016 -13288
rect 22334 -11670 23616 -11636
rect 22238 -12100 22272 -11732
rect 23678 -12100 23712 -11732
rect 22334 -12196 23616 -12162
rect 22238 -13226 22272 -12258
rect 23678 -13226 23712 -12258
rect 22334 -13322 23616 -13288
rect 23934 -11670 25216 -11636
rect 23838 -12100 23872 -11732
rect 25278 -12100 25312 -11732
rect 23934 -12196 25216 -12162
rect 23838 -13226 23872 -12258
rect 25278 -13226 25312 -12258
rect 23934 -13322 25216 -13288
rect 25534 -11670 26816 -11636
rect 25438 -12100 25472 -11732
rect 26878 -12100 26912 -11732
rect 25534 -12196 26816 -12162
rect 25438 -13226 25472 -12258
rect 26878 -13226 26912 -12258
rect 25534 -13322 26816 -13288
rect 27134 -11670 28416 -11636
rect 27038 -12100 27072 -11732
rect 28478 -12100 28512 -11732
rect 27134 -12196 28416 -12162
rect 27038 -13226 27072 -12258
rect 28478 -13226 28512 -12258
rect 27134 -13322 28416 -13288
rect 28734 -11670 30016 -11636
rect 28638 -12100 28672 -11732
rect 30078 -12100 30112 -11732
rect 28734 -12196 30016 -12162
rect 28638 -13226 28672 -12258
rect 30078 -13226 30112 -12258
rect 28734 -13322 30016 -13288
rect 30334 -11670 31616 -11636
rect 30238 -12100 30272 -11732
rect 31678 -12100 31712 -11732
rect 30334 -12196 31616 -12162
rect 30238 -13226 30272 -12258
rect 31678 -13226 31712 -12258
rect 30334 -13322 31616 -13288
rect 31934 -11670 33216 -11636
rect 31838 -12100 31872 -11732
rect 33278 -12100 33312 -11732
rect 31934 -12196 33216 -12162
rect 31838 -13226 31872 -12258
rect 33278 -13226 33312 -12258
rect 31934 -13322 33216 -13288
rect 33534 -11670 34816 -11636
rect 33438 -12100 33472 -11732
rect 34878 -12100 34912 -11732
rect 33534 -12196 34816 -12162
rect 33438 -13226 33472 -12258
rect 34878 -13226 34912 -12258
rect 33534 -13322 34816 -13288
rect 35134 -11670 36416 -11636
rect 35038 -12100 35072 -11732
rect 36478 -12100 36512 -11732
rect 35134 -12196 36416 -12162
rect 35038 -13226 35072 -12258
rect 36478 -13226 36512 -12258
rect 35134 -13322 36416 -13288
rect 36734 -11670 38016 -11636
rect 36638 -12100 36672 -11732
rect 38078 -12100 38112 -11732
rect 36734 -12196 38016 -12162
rect 36638 -13226 36672 -12258
rect 38078 -13226 38112 -12258
rect 36734 -13322 38016 -13288
rect -66 -13470 1216 -13436
rect -162 -13900 -128 -13532
rect 1278 -13900 1312 -13532
rect -66 -13996 1216 -13962
rect -162 -15026 -128 -14058
rect 1278 -15026 1312 -14058
rect -66 -15122 1216 -15088
rect 1534 -13470 2816 -13436
rect 1438 -13900 1472 -13532
rect 2878 -13900 2912 -13532
rect 1534 -13996 2816 -13962
rect 1438 -15026 1472 -14058
rect 2878 -15026 2912 -14058
rect 1534 -15122 2816 -15088
rect 3134 -13470 4416 -13436
rect 3038 -13900 3072 -13532
rect 4478 -13900 4512 -13532
rect 3134 -13996 4416 -13962
rect 3038 -15026 3072 -14058
rect 4478 -15026 4512 -14058
rect 3134 -15122 4416 -15088
rect 4734 -13470 6016 -13436
rect 4638 -13900 4672 -13532
rect 6078 -13900 6112 -13532
rect 4734 -13996 6016 -13962
rect 4638 -15026 4672 -14058
rect 6078 -15026 6112 -14058
rect 4734 -15122 6016 -15088
rect 6334 -13470 7616 -13436
rect 6238 -13900 6272 -13532
rect 7678 -13900 7712 -13532
rect 6334 -13996 7616 -13962
rect 6238 -15026 6272 -14058
rect 7678 -15026 7712 -14058
rect 6334 -15122 7616 -15088
rect 7934 -13470 9216 -13436
rect 7838 -13900 7872 -13532
rect 9278 -13900 9312 -13532
rect 7934 -13996 9216 -13962
rect 7838 -15026 7872 -14058
rect 9278 -15026 9312 -14058
rect 7934 -15122 9216 -15088
rect 9534 -13470 10816 -13436
rect 9438 -13900 9472 -13532
rect 10878 -13900 10912 -13532
rect 9534 -13996 10816 -13962
rect 9438 -15026 9472 -14058
rect 10878 -15026 10912 -14058
rect 9534 -15122 10816 -15088
rect 11134 -13470 12416 -13436
rect 11038 -13900 11072 -13532
rect 12478 -13900 12512 -13532
rect 11134 -13996 12416 -13962
rect 11038 -15026 11072 -14058
rect 12478 -15026 12512 -14058
rect 11134 -15122 12416 -15088
rect 12734 -13470 14016 -13436
rect 12638 -13900 12672 -13532
rect 14078 -13900 14112 -13532
rect 12734 -13996 14016 -13962
rect 12638 -15026 12672 -14058
rect 14078 -15026 14112 -14058
rect 12734 -15122 14016 -15088
rect 14334 -13470 15616 -13436
rect 14238 -13900 14272 -13532
rect 15678 -13900 15712 -13532
rect 14334 -13996 15616 -13962
rect 14238 -15026 14272 -14058
rect 15678 -15026 15712 -14058
rect 14334 -15122 15616 -15088
rect 15934 -13470 17216 -13436
rect 15838 -13900 15872 -13532
rect 17278 -13900 17312 -13532
rect 15934 -13996 17216 -13962
rect 15838 -15026 15872 -14058
rect 17278 -15026 17312 -14058
rect 15934 -15122 17216 -15088
rect 17534 -13470 18816 -13436
rect 17438 -13900 17472 -13532
rect 18878 -13900 18912 -13532
rect 17534 -13996 18816 -13962
rect 17438 -15026 17472 -14058
rect 18878 -15026 18912 -14058
rect 17534 -15122 18816 -15088
rect 19134 -13470 20416 -13436
rect 19038 -13900 19072 -13532
rect 20478 -13900 20512 -13532
rect 19134 -13996 20416 -13962
rect 19038 -15026 19072 -14058
rect 20478 -15026 20512 -14058
rect 19134 -15122 20416 -15088
rect 20734 -13470 22016 -13436
rect 20638 -13900 20672 -13532
rect 22078 -13900 22112 -13532
rect 20734 -13996 22016 -13962
rect 20638 -15026 20672 -14058
rect 22078 -15026 22112 -14058
rect 20734 -15122 22016 -15088
rect 22334 -13470 23616 -13436
rect 22238 -13900 22272 -13532
rect 23678 -13900 23712 -13532
rect 22334 -13996 23616 -13962
rect 22238 -15026 22272 -14058
rect 23678 -15026 23712 -14058
rect 22334 -15122 23616 -15088
rect 23934 -13470 25216 -13436
rect 23838 -13900 23872 -13532
rect 25278 -13900 25312 -13532
rect 23934 -13996 25216 -13962
rect 23838 -15026 23872 -14058
rect 25278 -15026 25312 -14058
rect 23934 -15122 25216 -15088
rect 25534 -13470 26816 -13436
rect 25438 -13900 25472 -13532
rect 26878 -13900 26912 -13532
rect 25534 -13996 26816 -13962
rect 25438 -15026 25472 -14058
rect 26878 -15026 26912 -14058
rect 25534 -15122 26816 -15088
rect 27134 -13470 28416 -13436
rect 27038 -13900 27072 -13532
rect 28478 -13900 28512 -13532
rect 27134 -13996 28416 -13962
rect 27038 -15026 27072 -14058
rect 28478 -15026 28512 -14058
rect 27134 -15122 28416 -15088
rect 28734 -13470 30016 -13436
rect 28638 -13900 28672 -13532
rect 30078 -13900 30112 -13532
rect 28734 -13996 30016 -13962
rect 28638 -15026 28672 -14058
rect 30078 -15026 30112 -14058
rect 28734 -15122 30016 -15088
rect 30334 -13470 31616 -13436
rect 30238 -13900 30272 -13532
rect 31678 -13900 31712 -13532
rect 30334 -13996 31616 -13962
rect 30238 -15026 30272 -14058
rect 31678 -15026 31712 -14058
rect 30334 -15122 31616 -15088
rect 31934 -13470 33216 -13436
rect 31838 -13900 31872 -13532
rect 33278 -13900 33312 -13532
rect 31934 -13996 33216 -13962
rect 31838 -15026 31872 -14058
rect 33278 -15026 33312 -14058
rect 31934 -15122 33216 -15088
rect 33534 -13470 34816 -13436
rect 33438 -13900 33472 -13532
rect 34878 -13900 34912 -13532
rect 33534 -13996 34816 -13962
rect 33438 -15026 33472 -14058
rect 34878 -15026 34912 -14058
rect 33534 -15122 34816 -15088
rect 35134 -13470 36416 -13436
rect 35038 -13900 35072 -13532
rect 36478 -13900 36512 -13532
rect 35134 -13996 36416 -13962
rect 35038 -15026 35072 -14058
rect 36478 -15026 36512 -14058
rect 35134 -15122 36416 -15088
rect 36734 -13470 38016 -13436
rect 36638 -13900 36672 -13532
rect 38078 -13900 38112 -13532
rect 36734 -13996 38016 -13962
rect 36638 -15026 36672 -14058
rect 38078 -15026 38112 -14058
rect 36734 -15122 38016 -15088
rect -66 -15270 1216 -15236
rect -162 -15700 -128 -15332
rect 1278 -15700 1312 -15332
rect -66 -15796 1216 -15762
rect -162 -16826 -128 -15858
rect 1278 -16826 1312 -15858
rect -66 -16922 1216 -16888
rect 1534 -15270 2816 -15236
rect 1438 -15700 1472 -15332
rect 2878 -15700 2912 -15332
rect 1534 -15796 2816 -15762
rect 1438 -16826 1472 -15858
rect 2878 -16826 2912 -15858
rect 1534 -16922 2816 -16888
rect 3134 -15270 4416 -15236
rect 3038 -15700 3072 -15332
rect 4478 -15700 4512 -15332
rect 3134 -15796 4416 -15762
rect 3038 -16826 3072 -15858
rect 4478 -16826 4512 -15858
rect 3134 -16922 4416 -16888
rect 4734 -15270 6016 -15236
rect 4638 -15700 4672 -15332
rect 6078 -15700 6112 -15332
rect 4734 -15796 6016 -15762
rect 4638 -16826 4672 -15858
rect 6078 -16826 6112 -15858
rect 4734 -16922 6016 -16888
rect 6334 -15270 7616 -15236
rect 6238 -15700 6272 -15332
rect 7678 -15700 7712 -15332
rect 6334 -15796 7616 -15762
rect 6238 -16826 6272 -15858
rect 7678 -16826 7712 -15858
rect 6334 -16922 7616 -16888
rect 7934 -15270 9216 -15236
rect 7838 -15700 7872 -15332
rect 9278 -15700 9312 -15332
rect 7934 -15796 9216 -15762
rect 7838 -16826 7872 -15858
rect 9278 -16826 9312 -15858
rect 7934 -16922 9216 -16888
rect 9534 -15270 10816 -15236
rect 9438 -15700 9472 -15332
rect 10878 -15700 10912 -15332
rect 9534 -15796 10816 -15762
rect 9438 -16826 9472 -15858
rect 10878 -16826 10912 -15858
rect 9534 -16922 10816 -16888
rect 11134 -15270 12416 -15236
rect 11038 -15700 11072 -15332
rect 12478 -15700 12512 -15332
rect 11134 -15796 12416 -15762
rect 11038 -16826 11072 -15858
rect 12478 -16826 12512 -15858
rect 11134 -16922 12416 -16888
rect 12734 -15270 14016 -15236
rect 12638 -15700 12672 -15332
rect 14078 -15700 14112 -15332
rect 12734 -15796 14016 -15762
rect 12638 -16826 12672 -15858
rect 14078 -16826 14112 -15858
rect 12734 -16922 14016 -16888
rect 14334 -15270 15616 -15236
rect 14238 -15700 14272 -15332
rect 15678 -15700 15712 -15332
rect 14334 -15796 15616 -15762
rect 14238 -16826 14272 -15858
rect 15678 -16826 15712 -15858
rect 14334 -16922 15616 -16888
rect 15934 -15270 17216 -15236
rect 15838 -15700 15872 -15332
rect 17278 -15700 17312 -15332
rect 15934 -15796 17216 -15762
rect 15838 -16826 15872 -15858
rect 17278 -16826 17312 -15858
rect 15934 -16922 17216 -16888
rect 17534 -15270 18816 -15236
rect 17438 -15700 17472 -15332
rect 18878 -15700 18912 -15332
rect 17534 -15796 18816 -15762
rect 17438 -16826 17472 -15858
rect 18878 -16826 18912 -15858
rect 17534 -16922 18816 -16888
rect 19134 -15270 20416 -15236
rect 19038 -15700 19072 -15332
rect 20478 -15700 20512 -15332
rect 19134 -15796 20416 -15762
rect 19038 -16826 19072 -15858
rect 20478 -16826 20512 -15858
rect 19134 -16922 20416 -16888
rect 20734 -15270 22016 -15236
rect 20638 -15700 20672 -15332
rect 22078 -15700 22112 -15332
rect 20734 -15796 22016 -15762
rect 20638 -16826 20672 -15858
rect 22078 -16826 22112 -15858
rect 20734 -16922 22016 -16888
rect 22334 -15270 23616 -15236
rect 22238 -15700 22272 -15332
rect 23678 -15700 23712 -15332
rect 22334 -15796 23616 -15762
rect 22238 -16826 22272 -15858
rect 23678 -16826 23712 -15858
rect 22334 -16922 23616 -16888
rect 23934 -15270 25216 -15236
rect 23838 -15700 23872 -15332
rect 25278 -15700 25312 -15332
rect 23934 -15796 25216 -15762
rect 23838 -16826 23872 -15858
rect 25278 -16826 25312 -15858
rect 23934 -16922 25216 -16888
rect 25534 -15270 26816 -15236
rect 25438 -15700 25472 -15332
rect 26878 -15700 26912 -15332
rect 25534 -15796 26816 -15762
rect 25438 -16826 25472 -15858
rect 26878 -16826 26912 -15858
rect 25534 -16922 26816 -16888
rect 27134 -15270 28416 -15236
rect 27038 -15700 27072 -15332
rect 28478 -15700 28512 -15332
rect 27134 -15796 28416 -15762
rect 27038 -16826 27072 -15858
rect 28478 -16826 28512 -15858
rect 27134 -16922 28416 -16888
rect 28734 -15270 30016 -15236
rect 28638 -15700 28672 -15332
rect 30078 -15700 30112 -15332
rect 28734 -15796 30016 -15762
rect 28638 -16826 28672 -15858
rect 30078 -16826 30112 -15858
rect 28734 -16922 30016 -16888
rect 30334 -15270 31616 -15236
rect 30238 -15700 30272 -15332
rect 31678 -15700 31712 -15332
rect 30334 -15796 31616 -15762
rect 30238 -16826 30272 -15858
rect 31678 -16826 31712 -15858
rect 30334 -16922 31616 -16888
rect 31934 -15270 33216 -15236
rect 31838 -15700 31872 -15332
rect 33278 -15700 33312 -15332
rect 31934 -15796 33216 -15762
rect 31838 -16826 31872 -15858
rect 33278 -16826 33312 -15858
rect 31934 -16922 33216 -16888
rect 33534 -15270 34816 -15236
rect 33438 -15700 33472 -15332
rect 34878 -15700 34912 -15332
rect 33534 -15796 34816 -15762
rect 33438 -16826 33472 -15858
rect 34878 -16826 34912 -15858
rect 33534 -16922 34816 -16888
rect 35134 -15270 36416 -15236
rect 35038 -15700 35072 -15332
rect 36478 -15700 36512 -15332
rect 35134 -15796 36416 -15762
rect 35038 -16826 35072 -15858
rect 36478 -16826 36512 -15858
rect 35134 -16922 36416 -16888
rect 36734 -15270 38016 -15236
rect 36638 -15700 36672 -15332
rect 38078 -15700 38112 -15332
rect 36734 -15796 38016 -15762
rect 36638 -16826 36672 -15858
rect 38078 -16826 38112 -15858
rect 36734 -16922 38016 -16888
rect -66 -17070 1216 -17036
rect -162 -17500 -128 -17132
rect 1278 -17500 1312 -17132
rect -66 -17596 1216 -17562
rect -162 -18626 -128 -17658
rect 1278 -18626 1312 -17658
rect -66 -18722 1216 -18688
rect 1534 -17070 2816 -17036
rect 1438 -17500 1472 -17132
rect 2878 -17500 2912 -17132
rect 1534 -17596 2816 -17562
rect 1438 -18626 1472 -17658
rect 2878 -18626 2912 -17658
rect 1534 -18722 2816 -18688
rect 3134 -17070 4416 -17036
rect 3038 -17500 3072 -17132
rect 4478 -17500 4512 -17132
rect 3134 -17596 4416 -17562
rect 3038 -18626 3072 -17658
rect 4478 -18626 4512 -17658
rect 3134 -18722 4416 -18688
rect 4734 -17070 6016 -17036
rect 4638 -17500 4672 -17132
rect 6078 -17500 6112 -17132
rect 4734 -17596 6016 -17562
rect 4638 -18626 4672 -17658
rect 6078 -18626 6112 -17658
rect 4734 -18722 6016 -18688
rect 6334 -17070 7616 -17036
rect 6238 -17500 6272 -17132
rect 7678 -17500 7712 -17132
rect 6334 -17596 7616 -17562
rect 6238 -18626 6272 -17658
rect 7678 -18626 7712 -17658
rect 6334 -18722 7616 -18688
rect 7934 -17070 9216 -17036
rect 7838 -17500 7872 -17132
rect 9278 -17500 9312 -17132
rect 7934 -17596 9216 -17562
rect 7838 -18626 7872 -17658
rect 9278 -18626 9312 -17658
rect 7934 -18722 9216 -18688
rect 9534 -17070 10816 -17036
rect 9438 -17500 9472 -17132
rect 10878 -17500 10912 -17132
rect 9534 -17596 10816 -17562
rect 9438 -18626 9472 -17658
rect 10878 -18626 10912 -17658
rect 9534 -18722 10816 -18688
rect 11134 -17070 12416 -17036
rect 11038 -17500 11072 -17132
rect 12478 -17500 12512 -17132
rect 11134 -17596 12416 -17562
rect 11038 -18626 11072 -17658
rect 12478 -18626 12512 -17658
rect 11134 -18722 12416 -18688
rect 12734 -17070 14016 -17036
rect 12638 -17500 12672 -17132
rect 14078 -17500 14112 -17132
rect 12734 -17596 14016 -17562
rect 12638 -18626 12672 -17658
rect 14078 -18626 14112 -17658
rect 12734 -18722 14016 -18688
rect 14334 -17070 15616 -17036
rect 14238 -17500 14272 -17132
rect 15678 -17500 15712 -17132
rect 14334 -17596 15616 -17562
rect 14238 -18626 14272 -17658
rect 15678 -18626 15712 -17658
rect 14334 -18722 15616 -18688
rect 15934 -17070 17216 -17036
rect 15838 -17500 15872 -17132
rect 17278 -17500 17312 -17132
rect 15934 -17596 17216 -17562
rect 15838 -18626 15872 -17658
rect 17278 -18626 17312 -17658
rect 15934 -18722 17216 -18688
rect 17534 -17070 18816 -17036
rect 17438 -17500 17472 -17132
rect 18878 -17500 18912 -17132
rect 17534 -17596 18816 -17562
rect 17438 -18626 17472 -17658
rect 18878 -18626 18912 -17658
rect 17534 -18722 18816 -18688
rect 19134 -17070 20416 -17036
rect 19038 -17500 19072 -17132
rect 20478 -17500 20512 -17132
rect 19134 -17596 20416 -17562
rect 19038 -18626 19072 -17658
rect 20478 -18626 20512 -17658
rect 19134 -18722 20416 -18688
rect 20734 -17070 22016 -17036
rect 20638 -17500 20672 -17132
rect 22078 -17500 22112 -17132
rect 20734 -17596 22016 -17562
rect 20638 -18626 20672 -17658
rect 22078 -18626 22112 -17658
rect 20734 -18722 22016 -18688
rect 22334 -17070 23616 -17036
rect 22238 -17500 22272 -17132
rect 23678 -17500 23712 -17132
rect 22334 -17596 23616 -17562
rect 22238 -18626 22272 -17658
rect 23678 -18626 23712 -17658
rect 22334 -18722 23616 -18688
rect 23934 -17070 25216 -17036
rect 23838 -17500 23872 -17132
rect 25278 -17500 25312 -17132
rect 23934 -17596 25216 -17562
rect 23838 -18626 23872 -17658
rect 25278 -18626 25312 -17658
rect 23934 -18722 25216 -18688
rect 25534 -17070 26816 -17036
rect 25438 -17500 25472 -17132
rect 26878 -17500 26912 -17132
rect 25534 -17596 26816 -17562
rect 25438 -18626 25472 -17658
rect 26878 -18626 26912 -17658
rect 25534 -18722 26816 -18688
rect 27134 -17070 28416 -17036
rect 27038 -17500 27072 -17132
rect 28478 -17500 28512 -17132
rect 27134 -17596 28416 -17562
rect 27038 -18626 27072 -17658
rect 28478 -18626 28512 -17658
rect 27134 -18722 28416 -18688
rect 28734 -17070 30016 -17036
rect 28638 -17500 28672 -17132
rect 30078 -17500 30112 -17132
rect 28734 -17596 30016 -17562
rect 28638 -18626 28672 -17658
rect 30078 -18626 30112 -17658
rect 28734 -18722 30016 -18688
rect 30334 -17070 31616 -17036
rect 30238 -17500 30272 -17132
rect 31678 -17500 31712 -17132
rect 30334 -17596 31616 -17562
rect 30238 -18626 30272 -17658
rect 31678 -18626 31712 -17658
rect 30334 -18722 31616 -18688
rect 31934 -17070 33216 -17036
rect 31838 -17500 31872 -17132
rect 33278 -17500 33312 -17132
rect 31934 -17596 33216 -17562
rect 31838 -18626 31872 -17658
rect 33278 -18626 33312 -17658
rect 31934 -18722 33216 -18688
rect 33534 -17070 34816 -17036
rect 33438 -17500 33472 -17132
rect 34878 -17500 34912 -17132
rect 33534 -17596 34816 -17562
rect 33438 -18626 33472 -17658
rect 34878 -18626 34912 -17658
rect 33534 -18722 34816 -18688
rect 35134 -17070 36416 -17036
rect 35038 -17500 35072 -17132
rect 36478 -17500 36512 -17132
rect 35134 -17596 36416 -17562
rect 35038 -18626 35072 -17658
rect 36478 -18626 36512 -17658
rect 35134 -18722 36416 -18688
rect 36734 -17070 38016 -17036
rect 36638 -17500 36672 -17132
rect 38078 -17500 38112 -17132
rect 36734 -17596 38016 -17562
rect 36638 -18626 36672 -17658
rect 38078 -18626 38112 -17658
rect 36734 -18722 38016 -18688
rect -66 -18870 1216 -18836
rect -162 -19300 -128 -18932
rect 1278 -19300 1312 -18932
rect -66 -19396 1216 -19362
rect -162 -20426 -128 -19458
rect 1278 -20426 1312 -19458
rect -66 -20522 1216 -20488
rect 1534 -18870 2816 -18836
rect 1438 -19300 1472 -18932
rect 2878 -19300 2912 -18932
rect 1534 -19396 2816 -19362
rect 1438 -20426 1472 -19458
rect 2878 -20426 2912 -19458
rect 1534 -20522 2816 -20488
rect 3134 -18870 4416 -18836
rect 3038 -19300 3072 -18932
rect 4478 -19300 4512 -18932
rect 3134 -19396 4416 -19362
rect 3038 -20426 3072 -19458
rect 4478 -20426 4512 -19458
rect 3134 -20522 4416 -20488
rect 4734 -18870 6016 -18836
rect 4638 -19300 4672 -18932
rect 6078 -19300 6112 -18932
rect 4734 -19396 6016 -19362
rect 4638 -20426 4672 -19458
rect 6078 -20426 6112 -19458
rect 4734 -20522 6016 -20488
rect 6334 -18870 7616 -18836
rect 6238 -19300 6272 -18932
rect 7678 -19300 7712 -18932
rect 6334 -19396 7616 -19362
rect 6238 -20426 6272 -19458
rect 7678 -20426 7712 -19458
rect 6334 -20522 7616 -20488
rect 7934 -18870 9216 -18836
rect 7838 -19300 7872 -18932
rect 9278 -19300 9312 -18932
rect 7934 -19396 9216 -19362
rect 7838 -20426 7872 -19458
rect 9278 -20426 9312 -19458
rect 7934 -20522 9216 -20488
rect 9534 -18870 10816 -18836
rect 9438 -19300 9472 -18932
rect 10878 -19300 10912 -18932
rect 9534 -19396 10816 -19362
rect 9438 -20426 9472 -19458
rect 10878 -20426 10912 -19458
rect 9534 -20522 10816 -20488
rect 11134 -18870 12416 -18836
rect 11038 -19300 11072 -18932
rect 12478 -19300 12512 -18932
rect 11134 -19396 12416 -19362
rect 11038 -20426 11072 -19458
rect 12478 -20426 12512 -19458
rect 11134 -20522 12416 -20488
rect 12734 -18870 14016 -18836
rect 12638 -19300 12672 -18932
rect 14078 -19300 14112 -18932
rect 12734 -19396 14016 -19362
rect 12638 -20426 12672 -19458
rect 14078 -20426 14112 -19458
rect 12734 -20522 14016 -20488
rect 14334 -18870 15616 -18836
rect 14238 -19300 14272 -18932
rect 15678 -19300 15712 -18932
rect 14334 -19396 15616 -19362
rect 14238 -20426 14272 -19458
rect 15678 -20426 15712 -19458
rect 14334 -20522 15616 -20488
rect 15934 -18870 17216 -18836
rect 15838 -19300 15872 -18932
rect 17278 -19300 17312 -18932
rect 15934 -19396 17216 -19362
rect 15838 -20426 15872 -19458
rect 17278 -20426 17312 -19458
rect 15934 -20522 17216 -20488
rect 17534 -18870 18816 -18836
rect 17438 -19300 17472 -18932
rect 18878 -19300 18912 -18932
rect 17534 -19396 18816 -19362
rect 17438 -20426 17472 -19458
rect 18878 -20426 18912 -19458
rect 17534 -20522 18816 -20488
rect 19134 -18870 20416 -18836
rect 19038 -19300 19072 -18932
rect 20478 -19300 20512 -18932
rect 19134 -19396 20416 -19362
rect 19038 -20426 19072 -19458
rect 20478 -20426 20512 -19458
rect 19134 -20522 20416 -20488
rect 20734 -18870 22016 -18836
rect 20638 -19300 20672 -18932
rect 22078 -19300 22112 -18932
rect 20734 -19396 22016 -19362
rect 20638 -20426 20672 -19458
rect 22078 -20426 22112 -19458
rect 20734 -20522 22016 -20488
rect 22334 -18870 23616 -18836
rect 22238 -19300 22272 -18932
rect 23678 -19300 23712 -18932
rect 22334 -19396 23616 -19362
rect 22238 -20426 22272 -19458
rect 23678 -20426 23712 -19458
rect 22334 -20522 23616 -20488
rect 23934 -18870 25216 -18836
rect 23838 -19300 23872 -18932
rect 25278 -19300 25312 -18932
rect 23934 -19396 25216 -19362
rect 23838 -20426 23872 -19458
rect 25278 -20426 25312 -19458
rect 23934 -20522 25216 -20488
rect 25534 -18870 26816 -18836
rect 25438 -19300 25472 -18932
rect 26878 -19300 26912 -18932
rect 25534 -19396 26816 -19362
rect 25438 -20426 25472 -19458
rect 26878 -20426 26912 -19458
rect 25534 -20522 26816 -20488
rect 27134 -18870 28416 -18836
rect 27038 -19300 27072 -18932
rect 28478 -19300 28512 -18932
rect 27134 -19396 28416 -19362
rect 27038 -20426 27072 -19458
rect 28478 -20426 28512 -19458
rect 27134 -20522 28416 -20488
rect 28734 -18870 30016 -18836
rect 28638 -19300 28672 -18932
rect 30078 -19300 30112 -18932
rect 28734 -19396 30016 -19362
rect 28638 -20426 28672 -19458
rect 30078 -20426 30112 -19458
rect 28734 -20522 30016 -20488
rect 30334 -18870 31616 -18836
rect 30238 -19300 30272 -18932
rect 31678 -19300 31712 -18932
rect 30334 -19396 31616 -19362
rect 30238 -20426 30272 -19458
rect 31678 -20426 31712 -19458
rect 30334 -20522 31616 -20488
rect 31934 -18870 33216 -18836
rect 31838 -19300 31872 -18932
rect 33278 -19300 33312 -18932
rect 31934 -19396 33216 -19362
rect 31838 -20426 31872 -19458
rect 33278 -20426 33312 -19458
rect 31934 -20522 33216 -20488
rect 33534 -18870 34816 -18836
rect 33438 -19300 33472 -18932
rect 34878 -19300 34912 -18932
rect 33534 -19396 34816 -19362
rect 33438 -20426 33472 -19458
rect 34878 -20426 34912 -19458
rect 33534 -20522 34816 -20488
rect 35134 -18870 36416 -18836
rect 35038 -19300 35072 -18932
rect 36478 -19300 36512 -18932
rect 35134 -19396 36416 -19362
rect 35038 -20426 35072 -19458
rect 36478 -20426 36512 -19458
rect 35134 -20522 36416 -20488
rect 36734 -18870 38016 -18836
rect 36638 -19300 36672 -18932
rect 38078 -19300 38112 -18932
rect 36734 -19396 38016 -19362
rect 36638 -20426 36672 -19458
rect 38078 -20426 38112 -19458
rect 36734 -20522 38016 -20488
rect -66 -20670 1216 -20636
rect -162 -21100 -128 -20732
rect 1278 -21100 1312 -20732
rect -66 -21196 1216 -21162
rect -162 -22226 -128 -21258
rect 1278 -22226 1312 -21258
rect -66 -22322 1216 -22288
rect 1534 -20670 2816 -20636
rect 1438 -21100 1472 -20732
rect 2878 -21100 2912 -20732
rect 1534 -21196 2816 -21162
rect 1438 -22226 1472 -21258
rect 2878 -22226 2912 -21258
rect 1534 -22322 2816 -22288
rect 3134 -20670 4416 -20636
rect 3038 -21100 3072 -20732
rect 4478 -21100 4512 -20732
rect 3134 -21196 4416 -21162
rect 3038 -22226 3072 -21258
rect 4478 -22226 4512 -21258
rect 3134 -22322 4416 -22288
rect 4734 -20670 6016 -20636
rect 4638 -21100 4672 -20732
rect 6078 -21100 6112 -20732
rect 4734 -21196 6016 -21162
rect 4638 -22226 4672 -21258
rect 6078 -22226 6112 -21258
rect 4734 -22322 6016 -22288
rect 6334 -20670 7616 -20636
rect 6238 -21100 6272 -20732
rect 7678 -21100 7712 -20732
rect 6334 -21196 7616 -21162
rect 6238 -22226 6272 -21258
rect 7678 -22226 7712 -21258
rect 6334 -22322 7616 -22288
rect 7934 -20670 9216 -20636
rect 7838 -21100 7872 -20732
rect 9278 -21100 9312 -20732
rect 7934 -21196 9216 -21162
rect 7838 -22226 7872 -21258
rect 9278 -22226 9312 -21258
rect 7934 -22322 9216 -22288
rect 9534 -20670 10816 -20636
rect 9438 -21100 9472 -20732
rect 10878 -21100 10912 -20732
rect 9534 -21196 10816 -21162
rect 9438 -22226 9472 -21258
rect 10878 -22226 10912 -21258
rect 9534 -22322 10816 -22288
rect 11134 -20670 12416 -20636
rect 11038 -21100 11072 -20732
rect 12478 -21100 12512 -20732
rect 11134 -21196 12416 -21162
rect 11038 -22226 11072 -21258
rect 12478 -22226 12512 -21258
rect 11134 -22322 12416 -22288
rect 12734 -20670 14016 -20636
rect 12638 -21100 12672 -20732
rect 14078 -21100 14112 -20732
rect 12734 -21196 14016 -21162
rect 12638 -22226 12672 -21258
rect 14078 -22226 14112 -21258
rect 12734 -22322 14016 -22288
rect 14334 -20670 15616 -20636
rect 14238 -21100 14272 -20732
rect 15678 -21100 15712 -20732
rect 14334 -21196 15616 -21162
rect 14238 -22226 14272 -21258
rect 15678 -22226 15712 -21258
rect 14334 -22322 15616 -22288
rect 15934 -20670 17216 -20636
rect 15838 -21100 15872 -20732
rect 17278 -21100 17312 -20732
rect 15934 -21196 17216 -21162
rect 15838 -22226 15872 -21258
rect 17278 -22226 17312 -21258
rect 15934 -22322 17216 -22288
rect 17534 -20670 18816 -20636
rect 17438 -21100 17472 -20732
rect 18878 -21100 18912 -20732
rect 17534 -21196 18816 -21162
rect 17438 -22226 17472 -21258
rect 18878 -22226 18912 -21258
rect 17534 -22322 18816 -22288
rect 19134 -20670 20416 -20636
rect 19038 -21100 19072 -20732
rect 20478 -21100 20512 -20732
rect 19134 -21196 20416 -21162
rect 19038 -22226 19072 -21258
rect 20478 -22226 20512 -21258
rect 19134 -22322 20416 -22288
rect 20734 -20670 22016 -20636
rect 20638 -21100 20672 -20732
rect 22078 -21100 22112 -20732
rect 20734 -21196 22016 -21162
rect 20638 -22226 20672 -21258
rect 22078 -22226 22112 -21258
rect 20734 -22322 22016 -22288
rect 22334 -20670 23616 -20636
rect 22238 -21100 22272 -20732
rect 23678 -21100 23712 -20732
rect 22334 -21196 23616 -21162
rect 22238 -22226 22272 -21258
rect 23678 -22226 23712 -21258
rect 22334 -22322 23616 -22288
rect 23934 -20670 25216 -20636
rect 23838 -21100 23872 -20732
rect 25278 -21100 25312 -20732
rect 23934 -21196 25216 -21162
rect 23838 -22226 23872 -21258
rect 25278 -22226 25312 -21258
rect 23934 -22322 25216 -22288
rect 25534 -20670 26816 -20636
rect 25438 -21100 25472 -20732
rect 26878 -21100 26912 -20732
rect 25534 -21196 26816 -21162
rect 25438 -22226 25472 -21258
rect 26878 -22226 26912 -21258
rect 25534 -22322 26816 -22288
rect 27134 -20670 28416 -20636
rect 27038 -21100 27072 -20732
rect 28478 -21100 28512 -20732
rect 27134 -21196 28416 -21162
rect 27038 -22226 27072 -21258
rect 28478 -22226 28512 -21258
rect 27134 -22322 28416 -22288
rect 28734 -20670 30016 -20636
rect 28638 -21100 28672 -20732
rect 30078 -21100 30112 -20732
rect 28734 -21196 30016 -21162
rect 28638 -22226 28672 -21258
rect 30078 -22226 30112 -21258
rect 28734 -22322 30016 -22288
rect 30334 -20670 31616 -20636
rect 30238 -21100 30272 -20732
rect 31678 -21100 31712 -20732
rect 30334 -21196 31616 -21162
rect 30238 -22226 30272 -21258
rect 31678 -22226 31712 -21258
rect 30334 -22322 31616 -22288
rect 31934 -20670 33216 -20636
rect 31838 -21100 31872 -20732
rect 33278 -21100 33312 -20732
rect 31934 -21196 33216 -21162
rect 31838 -22226 31872 -21258
rect 33278 -22226 33312 -21258
rect 31934 -22322 33216 -22288
rect 33534 -20670 34816 -20636
rect 33438 -21100 33472 -20732
rect 34878 -21100 34912 -20732
rect 33534 -21196 34816 -21162
rect 33438 -22226 33472 -21258
rect 34878 -22226 34912 -21258
rect 33534 -22322 34816 -22288
rect 35134 -20670 36416 -20636
rect 35038 -21100 35072 -20732
rect 36478 -21100 36512 -20732
rect 35134 -21196 36416 -21162
rect 35038 -22226 35072 -21258
rect 36478 -22226 36512 -21258
rect 35134 -22322 36416 -22288
rect 36734 -20670 38016 -20636
rect 36638 -21100 36672 -20732
rect 38078 -21100 38112 -20732
rect 36734 -21196 38016 -21162
rect 36638 -22226 36672 -21258
rect 38078 -22226 38112 -21258
rect 36734 -22322 38016 -22288
rect 32594 -22438 33336 -22404
rect 28314 -22558 29056 -22524
rect 28218 -23596 28252 -22620
rect 29118 -23596 29152 -22620
rect 32498 -23146 32532 -22500
rect 33398 -23146 33432 -22500
rect 32594 -23242 33336 -23208
rect 33964 -22458 34390 -22424
rect 33868 -23166 33902 -22520
rect 34452 -23166 34486 -22520
rect 33964 -23262 34390 -23228
rect 28314 -23692 29056 -23658
rect 33132 -23580 34190 -23546
rect 144 -24206 1990 -24172
rect 48 -24736 82 -24268
rect 2052 -24736 2086 -24268
rect 144 -24832 1990 -24798
rect 2344 -24206 4190 -24172
rect 2248 -24736 2282 -24268
rect 4252 -24736 4286 -24268
rect 2344 -24832 4190 -24798
rect 4544 -24206 6390 -24172
rect 4448 -24736 4482 -24268
rect 6452 -24736 6486 -24268
rect 4544 -24832 6390 -24798
rect 6744 -24206 8590 -24172
rect 6648 -24736 6682 -24268
rect 8652 -24736 8686 -24268
rect 6744 -24832 8590 -24798
rect 8944 -24206 10790 -24172
rect 8848 -24736 8882 -24268
rect 10852 -24736 10886 -24268
rect 8944 -24832 10790 -24798
rect 11144 -24206 12990 -24172
rect 11048 -24736 11082 -24268
rect 13052 -24736 13086 -24268
rect 11144 -24832 12990 -24798
rect 13344 -24206 15190 -24172
rect 13248 -24736 13282 -24268
rect 15252 -24736 15286 -24268
rect 13344 -24832 15190 -24798
rect 15544 -24206 17390 -24172
rect 15448 -24736 15482 -24268
rect 17452 -24736 17486 -24268
rect 15544 -24832 17390 -24798
rect 17744 -24206 19590 -24172
rect 17648 -24736 17682 -24268
rect 19652 -24736 19686 -24268
rect 17744 -24832 19590 -24798
rect 19944 -24206 21790 -24172
rect 19848 -24736 19882 -24268
rect 21852 -24736 21886 -24268
rect 33036 -24288 33070 -23642
rect 34252 -24288 34286 -23642
rect 33132 -24384 34190 -24350
rect 34504 -23578 37142 -23544
rect 34408 -24286 34442 -23640
rect 37204 -24286 37238 -23640
rect 34504 -24382 37142 -24348
rect 19944 -24832 21790 -24798
rect 22292 -24548 26968 -24514
rect 144 -25006 1990 -24972
rect 48 -25536 82 -25068
rect 2052 -25536 2086 -25068
rect 144 -25632 1990 -25598
rect 2344 -25006 4190 -24972
rect 2248 -25536 2282 -25068
rect 4252 -25536 4286 -25068
rect 2344 -25632 4190 -25598
rect 4544 -25006 6390 -24972
rect 4448 -25536 4482 -25068
rect 6452 -25536 6486 -25068
rect 4544 -25632 6390 -25598
rect 6744 -25006 8590 -24972
rect 6648 -25536 6682 -25068
rect 8652 -25536 8686 -25068
rect 6744 -25632 8590 -25598
rect 8944 -25006 10790 -24972
rect 8848 -25536 8882 -25068
rect 10852 -25536 10886 -25068
rect 8944 -25632 10790 -25598
rect 11144 -25006 12990 -24972
rect 11048 -25536 11082 -25068
rect 13052 -25536 13086 -25068
rect 11144 -25632 12990 -25598
rect 13344 -25006 15190 -24972
rect 13248 -25536 13282 -25068
rect 15252 -25536 15286 -25068
rect 13344 -25632 15190 -25598
rect 15544 -25006 17390 -24972
rect 15448 -25536 15482 -25068
rect 17452 -25536 17486 -25068
rect 15544 -25632 17390 -25598
rect 17744 -25006 19590 -24972
rect 17648 -25536 17682 -25068
rect 19652 -25536 19686 -25068
rect 17744 -25632 19590 -25598
rect 19944 -25006 21790 -24972
rect 19848 -25536 19882 -25068
rect 21852 -25536 21886 -25068
rect 19944 -25632 21790 -25598
rect 144 -25806 1990 -25772
rect 48 -26336 82 -25868
rect 2052 -26336 2086 -25868
rect 144 -26432 1990 -26398
rect 2344 -25806 4190 -25772
rect 2248 -26336 2282 -25868
rect 4252 -26336 4286 -25868
rect 2344 -26432 4190 -26398
rect 4544 -25806 6390 -25772
rect 4448 -26336 4482 -25868
rect 6452 -26336 6486 -25868
rect 4544 -26432 6390 -26398
rect 6744 -25806 8590 -25772
rect 6648 -26336 6682 -25868
rect 8652 -26336 8686 -25868
rect 6744 -26432 8590 -26398
rect 8944 -25806 10790 -25772
rect 8848 -26336 8882 -25868
rect 10852 -26336 10886 -25868
rect 8944 -26432 10790 -26398
rect 11144 -25806 12990 -25772
rect 11048 -26336 11082 -25868
rect 13052 -26336 13086 -25868
rect 11144 -26432 12990 -26398
rect 13344 -25806 15190 -25772
rect 13248 -26336 13282 -25868
rect 15252 -26336 15286 -25868
rect 13344 -26432 15190 -26398
rect 15544 -25806 17390 -25772
rect 15448 -26336 15482 -25868
rect 17452 -26336 17486 -25868
rect 15544 -26432 17390 -26398
rect 17744 -25806 19590 -25772
rect 17648 -26336 17682 -25868
rect 19652 -26336 19686 -25868
rect 17744 -26432 19590 -26398
rect 19944 -25806 21790 -25772
rect 19848 -26336 19882 -25868
rect 21852 -26336 21886 -25868
rect 19944 -26432 21790 -26398
rect 144 -26606 1990 -26572
rect 48 -27136 82 -26668
rect 2052 -27136 2086 -26668
rect 144 -27232 1990 -27198
rect 2344 -26606 4190 -26572
rect 2248 -27136 2282 -26668
rect 4252 -27136 4286 -26668
rect 2344 -27232 4190 -27198
rect 4544 -26606 6390 -26572
rect 4448 -27136 4482 -26668
rect 6452 -27136 6486 -26668
rect 4544 -27232 6390 -27198
rect 6744 -26606 8590 -26572
rect 6648 -27136 6682 -26668
rect 8652 -27136 8686 -26668
rect 6744 -27232 8590 -27198
rect 8944 -26606 10790 -26572
rect 8848 -27136 8882 -26668
rect 10852 -27136 10886 -26668
rect 8944 -27232 10790 -27198
rect 11144 -26606 12990 -26572
rect 11048 -27136 11082 -26668
rect 13052 -27136 13086 -26668
rect 11144 -27232 12990 -27198
rect 13344 -26606 15190 -26572
rect 13248 -27136 13282 -26668
rect 15252 -27136 15286 -26668
rect 13344 -27232 15190 -27198
rect 15544 -26606 17390 -26572
rect 15448 -27136 15482 -26668
rect 17452 -27136 17486 -26668
rect 15544 -27232 17390 -27198
rect 17744 -26606 19590 -26572
rect 17648 -27136 17682 -26668
rect 19652 -27136 19686 -26668
rect 17744 -27232 19590 -27198
rect 19944 -26606 21790 -26572
rect 19848 -27136 19882 -26668
rect 21852 -27136 21886 -26668
rect 19944 -27232 21790 -27198
rect 144 -27406 1990 -27372
rect 48 -27936 82 -27468
rect 2052 -27936 2086 -27468
rect 144 -28032 1990 -27998
rect 2344 -27406 4190 -27372
rect 2248 -27936 2282 -27468
rect 4252 -27936 4286 -27468
rect 2344 -28032 4190 -27998
rect 4544 -27406 6390 -27372
rect 4448 -27936 4482 -27468
rect 6452 -27936 6486 -27468
rect 4544 -28032 6390 -27998
rect 6744 -27406 8590 -27372
rect 6648 -27936 6682 -27468
rect 8652 -27936 8686 -27468
rect 6744 -28032 8590 -27998
rect 8944 -27406 10790 -27372
rect 8848 -27936 8882 -27468
rect 10852 -27936 10886 -27468
rect 8944 -28032 10790 -27998
rect 11144 -27406 12990 -27372
rect 11048 -27936 11082 -27468
rect 13052 -27936 13086 -27468
rect 11144 -28032 12990 -27998
rect 13344 -27406 15190 -27372
rect 13248 -27936 13282 -27468
rect 15252 -27936 15286 -27468
rect 13344 -28032 15190 -27998
rect 15544 -27406 17390 -27372
rect 15448 -27936 15482 -27468
rect 17452 -27936 17486 -27468
rect 15544 -28032 17390 -27998
rect 17744 -27406 19590 -27372
rect 17648 -27936 17682 -27468
rect 19652 -27936 19686 -27468
rect 17744 -28032 19590 -27998
rect 19944 -27406 21790 -27372
rect 19848 -27936 19882 -27468
rect 21852 -27936 21886 -27468
rect 19944 -28032 21790 -27998
rect 144 -28206 1990 -28172
rect 48 -28736 82 -28268
rect 2052 -28736 2086 -28268
rect 144 -28832 1990 -28798
rect 2344 -28206 4190 -28172
rect 2248 -28736 2282 -28268
rect 4252 -28736 4286 -28268
rect 2344 -28832 4190 -28798
rect 4544 -28206 6390 -28172
rect 4448 -28736 4482 -28268
rect 6452 -28736 6486 -28268
rect 4544 -28832 6390 -28798
rect 6744 -28206 8590 -28172
rect 6648 -28736 6682 -28268
rect 8652 -28736 8686 -28268
rect 6744 -28832 8590 -28798
rect 8944 -28206 10790 -28172
rect 8848 -28736 8882 -28268
rect 10852 -28736 10886 -28268
rect 8944 -28832 10790 -28798
rect 11144 -28206 12990 -28172
rect 11048 -28736 11082 -28268
rect 13052 -28736 13086 -28268
rect 11144 -28832 12990 -28798
rect 13344 -28206 15190 -28172
rect 13248 -28736 13282 -28268
rect 15252 -28736 15286 -28268
rect 13344 -28832 15190 -28798
rect 15544 -28206 17390 -28172
rect 15448 -28736 15482 -28268
rect 17452 -28736 17486 -28268
rect 15544 -28832 17390 -28798
rect 17744 -28206 19590 -28172
rect 17648 -28736 17682 -28268
rect 19652 -28736 19686 -28268
rect 17744 -28832 19590 -28798
rect 19944 -28206 21790 -28172
rect 19848 -28736 19882 -28268
rect 21852 -28736 21886 -28268
rect 19944 -28832 21790 -28798
rect 144 -29006 1990 -28972
rect 48 -29536 82 -29068
rect 2052 -29536 2086 -29068
rect 144 -29632 1990 -29598
rect 2344 -29006 4190 -28972
rect 2248 -29536 2282 -29068
rect 4252 -29536 4286 -29068
rect 2344 -29632 4190 -29598
rect 4544 -29006 6390 -28972
rect 4448 -29536 4482 -29068
rect 6452 -29536 6486 -29068
rect 4544 -29632 6390 -29598
rect 6744 -29006 8590 -28972
rect 6648 -29536 6682 -29068
rect 8652 -29536 8686 -29068
rect 6744 -29632 8590 -29598
rect 8944 -29006 10790 -28972
rect 8848 -29536 8882 -29068
rect 10852 -29536 10886 -29068
rect 8944 -29632 10790 -29598
rect 11144 -29006 12990 -28972
rect 11048 -29536 11082 -29068
rect 13052 -29536 13086 -29068
rect 11144 -29632 12990 -29598
rect 13344 -29006 15190 -28972
rect 13248 -29536 13282 -29068
rect 15252 -29536 15286 -29068
rect 13344 -29632 15190 -29598
rect 15544 -29006 17390 -28972
rect 15448 -29536 15482 -29068
rect 17452 -29536 17486 -29068
rect 15544 -29632 17390 -29598
rect 17744 -29006 19590 -28972
rect 17648 -29536 17682 -29068
rect 19652 -29536 19686 -29068
rect 17744 -29632 19590 -29598
rect 19944 -29006 21790 -28972
rect 19848 -29536 19882 -29068
rect 21852 -29536 21886 -29068
rect 19944 -29632 21790 -29598
rect 144 -29806 1990 -29772
rect 48 -30336 82 -29868
rect 2052 -30336 2086 -29868
rect 144 -30432 1990 -30398
rect 2344 -29806 4190 -29772
rect 2248 -30336 2282 -29868
rect 4252 -30336 4286 -29868
rect 2344 -30432 4190 -30398
rect 4544 -29806 6390 -29772
rect 4448 -30336 4482 -29868
rect 6452 -30336 6486 -29868
rect 4544 -30432 6390 -30398
rect 6744 -29806 8590 -29772
rect 6648 -30336 6682 -29868
rect 8652 -30336 8686 -29868
rect 6744 -30432 8590 -30398
rect 8944 -29806 10790 -29772
rect 8848 -30336 8882 -29868
rect 10852 -30336 10886 -29868
rect 8944 -30432 10790 -30398
rect 11144 -29806 12990 -29772
rect 11048 -30336 11082 -29868
rect 13052 -30336 13086 -29868
rect 11144 -30432 12990 -30398
rect 13344 -29806 15190 -29772
rect 13248 -30336 13282 -29868
rect 15252 -30336 15286 -29868
rect 13344 -30432 15190 -30398
rect 15544 -29806 17390 -29772
rect 15448 -30336 15482 -29868
rect 17452 -30336 17486 -29868
rect 15544 -30432 17390 -30398
rect 17744 -29806 19590 -29772
rect 17648 -30336 17682 -29868
rect 19652 -30336 19686 -29868
rect 17744 -30432 19590 -30398
rect 19944 -29806 21790 -29772
rect 19848 -30336 19882 -29868
rect 21852 -30336 21886 -29868
rect 19944 -30432 21790 -30398
rect 144 -30606 1990 -30572
rect 48 -31136 82 -30668
rect 2052 -31136 2086 -30668
rect 144 -31232 1990 -31198
rect 2344 -30606 4190 -30572
rect 2248 -31136 2282 -30668
rect 4252 -31136 4286 -30668
rect 2344 -31232 4190 -31198
rect 4544 -30606 6390 -30572
rect 4448 -31136 4482 -30668
rect 6452 -31136 6486 -30668
rect 4544 -31232 6390 -31198
rect 6744 -30606 8590 -30572
rect 6648 -31136 6682 -30668
rect 8652 -31136 8686 -30668
rect 6744 -31232 8590 -31198
rect 8944 -30606 10790 -30572
rect 8848 -31136 8882 -30668
rect 10852 -31136 10886 -30668
rect 8944 -31232 10790 -31198
rect 11144 -30606 12990 -30572
rect 11048 -31136 11082 -30668
rect 13052 -31136 13086 -30668
rect 11144 -31232 12990 -31198
rect 13344 -30606 15190 -30572
rect 13248 -31136 13282 -30668
rect 15252 -31136 15286 -30668
rect 13344 -31232 15190 -31198
rect 15544 -30606 17390 -30572
rect 15448 -31136 15482 -30668
rect 17452 -31136 17486 -30668
rect 15544 -31232 17390 -31198
rect 17744 -30606 19590 -30572
rect 17648 -31136 17682 -30668
rect 19652 -31136 19686 -30668
rect 17744 -31232 19590 -31198
rect 19944 -30606 21790 -30572
rect 19848 -31136 19882 -30668
rect 21852 -31136 21886 -30668
rect 19944 -31232 21790 -31198
rect 144 -31406 1990 -31372
rect 48 -31936 82 -31468
rect 2052 -31936 2086 -31468
rect 144 -32032 1990 -31998
rect 2344 -31406 4190 -31372
rect 2248 -31936 2282 -31468
rect 4252 -31936 4286 -31468
rect 2344 -32032 4190 -31998
rect 4544 -31406 6390 -31372
rect 4448 -31936 4482 -31468
rect 6452 -31936 6486 -31468
rect 4544 -32032 6390 -31998
rect 6744 -31406 8590 -31372
rect 6648 -31936 6682 -31468
rect 8652 -31936 8686 -31468
rect 6744 -32032 8590 -31998
rect 8944 -31406 10790 -31372
rect 8848 -31936 8882 -31468
rect 10852 -31936 10886 -31468
rect 8944 -32032 10790 -31998
rect 11144 -31406 12990 -31372
rect 11048 -31936 11082 -31468
rect 13052 -31936 13086 -31468
rect 11144 -32032 12990 -31998
rect 13344 -31406 15190 -31372
rect 13248 -31936 13282 -31468
rect 15252 -31936 15286 -31468
rect 13344 -32032 15190 -31998
rect 15544 -31406 17390 -31372
rect 15448 -31936 15482 -31468
rect 17452 -31936 17486 -31468
rect 15544 -32032 17390 -31998
rect 17744 -31406 19590 -31372
rect 17648 -31936 17682 -31468
rect 19652 -31936 19686 -31468
rect 17744 -32032 19590 -31998
rect 19944 -31406 21790 -31372
rect 19848 -31936 19882 -31468
rect 21852 -31936 21886 -31468
rect 19944 -32032 21790 -31998
rect 22196 -31968 22230 -24610
rect 27030 -31968 27064 -24610
rect 34854 -24730 35900 -24696
rect 34758 -26966 34792 -24792
rect 35962 -26966 35996 -24792
rect 34854 -27062 35900 -27028
rect 36194 -24730 37240 -24696
rect 36098 -26966 36132 -24792
rect 37302 -26966 37336 -24792
rect 36194 -27062 37240 -27028
rect 31774 -28336 32042 -28302
rect 32214 -28336 32482 -28302
rect 32654 -28336 32922 -28302
rect 31678 -29044 31712 -28398
rect 32104 -29044 32138 -28398
rect 33974 -28336 34242 -28302
rect 34414 -28336 34682 -28302
rect 34854 -28336 35122 -28302
rect 33068 -28636 33636 -28602
rect 32972 -29044 33006 -28698
rect 33698 -29044 33732 -28698
rect 31774 -29140 32042 -29106
rect 32214 -29140 32482 -29106
rect 32654 -29140 32922 -29106
rect 33068 -29140 33636 -29106
rect 33878 -29044 33912 -28398
rect 34304 -29044 34338 -28398
rect 36174 -28336 36442 -28302
rect 36614 -28336 36882 -28302
rect 37054 -28336 37322 -28302
rect 35268 -28636 35836 -28602
rect 35172 -29044 35206 -28698
rect 35898 -29044 35932 -28698
rect 33974 -29140 34242 -29106
rect 34414 -29140 34682 -29106
rect 34854 -29140 35122 -29106
rect 35268 -29140 35836 -29106
rect 36078 -29044 36112 -28398
rect 36504 -29044 36538 -28398
rect 37468 -28636 38036 -28602
rect 37372 -29044 37406 -28698
rect 38098 -29044 38132 -28698
rect 36174 -29140 36442 -29106
rect 36614 -29140 36882 -29106
rect 37054 -29140 37322 -29106
rect 37468 -29140 38036 -29106
rect 31786 -30918 32354 -30884
rect 32500 -30918 32768 -30884
rect 32940 -30918 33208 -30884
rect 33380 -30918 33648 -30884
rect 31690 -31326 31724 -30980
rect 32416 -31326 32450 -30980
rect 31786 -31422 32354 -31388
rect 33284 -31626 33318 -30980
rect 33710 -31626 33744 -30980
rect 33986 -30918 34554 -30884
rect 34700 -30918 34968 -30884
rect 35140 -30918 35408 -30884
rect 35580 -30918 35848 -30884
rect 33890 -31326 33924 -30980
rect 34616 -31326 34650 -30980
rect 33986 -31422 34554 -31388
rect 32500 -31722 32768 -31688
rect 32940 -31722 33208 -31688
rect 33380 -31722 33648 -31688
rect 35484 -31626 35518 -30980
rect 35910 -31626 35944 -30980
rect 36186 -30918 36754 -30884
rect 36900 -30918 37168 -30884
rect 37340 -30918 37608 -30884
rect 37780 -30918 38048 -30884
rect 36090 -31326 36124 -30980
rect 36816 -31326 36850 -30980
rect 36186 -31422 36754 -31388
rect 34700 -31722 34968 -31688
rect 35140 -31722 35408 -31688
rect 35580 -31722 35848 -31688
rect 37684 -31626 37718 -30980
rect 38110 -31626 38144 -30980
rect 36900 -31722 37168 -31688
rect 37340 -31722 37608 -31688
rect 37780 -31722 38048 -31688
rect 22292 -32064 26968 -32030
<< poly >>
rect 171 11713 259 11729
rect 171 11445 187 11713
rect 221 11445 259 11713
rect 171 11429 259 11445
rect 1859 11713 1947 11729
rect 1859 11445 1897 11713
rect 1931 11445 1947 11713
rect 1859 11429 1947 11445
rect 2371 11713 2459 11729
rect 2371 11445 2387 11713
rect 2421 11445 2459 11713
rect 2371 11429 2459 11445
rect 4059 11713 4147 11729
rect 4059 11445 4097 11713
rect 4131 11445 4147 11713
rect 4059 11429 4147 11445
rect 4571 11713 4659 11729
rect 4571 11445 4587 11713
rect 4621 11445 4659 11713
rect 4571 11429 4659 11445
rect 6259 11713 6347 11729
rect 6259 11445 6297 11713
rect 6331 11445 6347 11713
rect 6259 11429 6347 11445
rect 6771 11713 6859 11729
rect 6771 11445 6787 11713
rect 6821 11445 6859 11713
rect 6771 11429 6859 11445
rect 8459 11713 8547 11729
rect 8459 11445 8497 11713
rect 8531 11445 8547 11713
rect 8459 11429 8547 11445
rect 8971 11713 9059 11729
rect 8971 11445 8987 11713
rect 9021 11445 9059 11713
rect 8971 11429 9059 11445
rect 10659 11713 10747 11729
rect 10659 11445 10697 11713
rect 10731 11445 10747 11713
rect 10659 11429 10747 11445
rect 11171 11713 11259 11729
rect 11171 11445 11187 11713
rect 11221 11445 11259 11713
rect 11171 11429 11259 11445
rect 12859 11713 12947 11729
rect 12859 11445 12897 11713
rect 12931 11445 12947 11713
rect 12859 11429 12947 11445
rect 13371 11713 13459 11729
rect 13371 11445 13387 11713
rect 13421 11445 13459 11713
rect 13371 11429 13459 11445
rect 15059 11713 15147 11729
rect 15059 11445 15097 11713
rect 15131 11445 15147 11713
rect 15059 11429 15147 11445
rect 15571 11713 15659 11729
rect 15571 11445 15587 11713
rect 15621 11445 15659 11713
rect 15571 11429 15659 11445
rect 17259 11713 17347 11729
rect 17259 11445 17297 11713
rect 17331 11445 17347 11713
rect 17259 11429 17347 11445
rect 17771 11713 17859 11729
rect 17771 11445 17787 11713
rect 17821 11445 17859 11713
rect 17771 11429 17859 11445
rect 19459 11713 19547 11729
rect 19459 11445 19497 11713
rect 19531 11445 19547 11713
rect 19459 11429 19547 11445
rect 19971 11713 20059 11729
rect 19971 11445 19987 11713
rect 20021 11445 20059 11713
rect 19971 11429 20059 11445
rect 21659 11713 21747 11729
rect 21659 11445 21697 11713
rect 21731 11445 21747 11713
rect 21659 11429 21747 11445
rect 171 10913 259 10929
rect 171 10645 187 10913
rect 221 10645 259 10913
rect 171 10629 259 10645
rect 1859 10913 1947 10929
rect 1859 10645 1897 10913
rect 1931 10645 1947 10913
rect 1859 10629 1947 10645
rect 2370 10912 2458 10928
rect 2370 10644 2386 10912
rect 2420 10644 2458 10912
rect 2370 10628 2458 10644
rect 4058 10912 4146 10928
rect 4058 10644 4096 10912
rect 4130 10644 4146 10912
rect 4058 10628 4146 10644
rect 4570 10912 4658 10928
rect 4570 10644 4586 10912
rect 4620 10644 4658 10912
rect 4570 10628 4658 10644
rect 6258 10912 6346 10928
rect 6258 10644 6296 10912
rect 6330 10644 6346 10912
rect 6258 10628 6346 10644
rect 6770 10912 6858 10928
rect 6770 10644 6786 10912
rect 6820 10644 6858 10912
rect 6770 10628 6858 10644
rect 8458 10912 8546 10928
rect 8458 10644 8496 10912
rect 8530 10644 8546 10912
rect 8458 10628 8546 10644
rect 8970 10912 9058 10928
rect 8970 10644 8986 10912
rect 9020 10644 9058 10912
rect 8970 10628 9058 10644
rect 10658 10912 10746 10928
rect 10658 10644 10696 10912
rect 10730 10644 10746 10912
rect 10658 10628 10746 10644
rect 11170 10912 11258 10928
rect 11170 10644 11186 10912
rect 11220 10644 11258 10912
rect 11170 10628 11258 10644
rect 12858 10912 12946 10928
rect 12858 10644 12896 10912
rect 12930 10644 12946 10912
rect 12858 10628 12946 10644
rect 13370 10912 13458 10928
rect 13370 10644 13386 10912
rect 13420 10644 13458 10912
rect 13370 10628 13458 10644
rect 15058 10912 15146 10928
rect 15058 10644 15096 10912
rect 15130 10644 15146 10912
rect 15058 10628 15146 10644
rect 15570 10912 15658 10928
rect 15570 10644 15586 10912
rect 15620 10644 15658 10912
rect 15570 10628 15658 10644
rect 17258 10912 17346 10928
rect 17258 10644 17296 10912
rect 17330 10644 17346 10912
rect 17258 10628 17346 10644
rect 17770 10912 17858 10928
rect 17770 10644 17786 10912
rect 17820 10644 17858 10912
rect 17770 10628 17858 10644
rect 19458 10912 19546 10928
rect 19458 10644 19496 10912
rect 19530 10644 19546 10912
rect 19458 10628 19546 10644
rect 19971 10913 20059 10929
rect 19971 10645 19987 10913
rect 20021 10645 20059 10913
rect 19971 10629 20059 10645
rect 21659 10913 21747 10929
rect 21659 10645 21697 10913
rect 21731 10645 21747 10913
rect 21659 10629 21747 10645
rect 171 10113 259 10129
rect 171 9845 187 10113
rect 221 9845 259 10113
rect 171 9829 259 9845
rect 1859 10113 1947 10129
rect 1859 9845 1897 10113
rect 1931 9845 1947 10113
rect 1859 9829 1947 9845
rect 2370 10112 2458 10128
rect 2370 9844 2386 10112
rect 2420 9844 2458 10112
rect 2370 9828 2458 9844
rect 4058 10112 4146 10128
rect 4058 9844 4096 10112
rect 4130 9844 4146 10112
rect 4058 9828 4146 9844
rect 4570 10112 4658 10128
rect 4570 9844 4586 10112
rect 4620 9844 4658 10112
rect 4570 9828 4658 9844
rect 6258 10112 6346 10128
rect 6258 9844 6296 10112
rect 6330 9844 6346 10112
rect 6258 9828 6346 9844
rect 6770 10112 6858 10128
rect 6770 9844 6786 10112
rect 6820 9844 6858 10112
rect 6770 9828 6858 9844
rect 8458 10112 8546 10128
rect 8458 9844 8496 10112
rect 8530 9844 8546 10112
rect 8458 9828 8546 9844
rect 8970 10112 9058 10128
rect 8970 9844 8986 10112
rect 9020 9844 9058 10112
rect 8970 9828 9058 9844
rect 10658 10112 10746 10128
rect 10658 9844 10696 10112
rect 10730 9844 10746 10112
rect 10658 9828 10746 9844
rect 11170 10112 11258 10128
rect 11170 9844 11186 10112
rect 11220 9844 11258 10112
rect 11170 9828 11258 9844
rect 12858 10112 12946 10128
rect 12858 9844 12896 10112
rect 12930 9844 12946 10112
rect 12858 9828 12946 9844
rect 13370 10112 13458 10128
rect 13370 9844 13386 10112
rect 13420 9844 13458 10112
rect 13370 9828 13458 9844
rect 15058 10112 15146 10128
rect 15058 9844 15096 10112
rect 15130 9844 15146 10112
rect 15058 9828 15146 9844
rect 15570 10112 15658 10128
rect 15570 9844 15586 10112
rect 15620 9844 15658 10112
rect 15570 9828 15658 9844
rect 17258 10112 17346 10128
rect 17258 9844 17296 10112
rect 17330 9844 17346 10112
rect 17258 9828 17346 9844
rect 17770 10112 17858 10128
rect 17770 9844 17786 10112
rect 17820 9844 17858 10112
rect 17770 9828 17858 9844
rect 19458 10112 19546 10128
rect 19458 9844 19496 10112
rect 19530 9844 19546 10112
rect 19458 9828 19546 9844
rect 19971 10113 20059 10129
rect 19971 9845 19987 10113
rect 20021 9845 20059 10113
rect 19971 9829 20059 9845
rect 21659 10113 21747 10129
rect 21659 9845 21697 10113
rect 21731 9845 21747 10113
rect 21659 9829 21747 9845
rect 171 9313 259 9329
rect 171 9045 187 9313
rect 221 9045 259 9313
rect 171 9029 259 9045
rect 1859 9313 1947 9329
rect 1859 9045 1897 9313
rect 1931 9045 1947 9313
rect 1859 9029 1947 9045
rect 2370 9312 2458 9328
rect 2370 9044 2386 9312
rect 2420 9044 2458 9312
rect 2370 9028 2458 9044
rect 4058 9312 4146 9328
rect 4058 9044 4096 9312
rect 4130 9044 4146 9312
rect 4058 9028 4146 9044
rect 4570 9312 4658 9328
rect 4570 9044 4586 9312
rect 4620 9044 4658 9312
rect 4570 9028 4658 9044
rect 6258 9312 6346 9328
rect 6258 9044 6296 9312
rect 6330 9044 6346 9312
rect 6258 9028 6346 9044
rect 6770 9312 6858 9328
rect 6770 9044 6786 9312
rect 6820 9044 6858 9312
rect 6770 9028 6858 9044
rect 8458 9312 8546 9328
rect 8458 9044 8496 9312
rect 8530 9044 8546 9312
rect 8458 9028 8546 9044
rect 8970 9312 9058 9328
rect 8970 9044 8986 9312
rect 9020 9044 9058 9312
rect 8970 9028 9058 9044
rect 10658 9312 10746 9328
rect 10658 9044 10696 9312
rect 10730 9044 10746 9312
rect 10658 9028 10746 9044
rect 11170 9312 11258 9328
rect 11170 9044 11186 9312
rect 11220 9044 11258 9312
rect 11170 9028 11258 9044
rect 12858 9312 12946 9328
rect 12858 9044 12896 9312
rect 12930 9044 12946 9312
rect 12858 9028 12946 9044
rect 13370 9312 13458 9328
rect 13370 9044 13386 9312
rect 13420 9044 13458 9312
rect 13370 9028 13458 9044
rect 15058 9312 15146 9328
rect 15058 9044 15096 9312
rect 15130 9044 15146 9312
rect 15058 9028 15146 9044
rect 15570 9312 15658 9328
rect 15570 9044 15586 9312
rect 15620 9044 15658 9312
rect 15570 9028 15658 9044
rect 17258 9312 17346 9328
rect 17258 9044 17296 9312
rect 17330 9044 17346 9312
rect 17258 9028 17346 9044
rect 17770 9312 17858 9328
rect 17770 9044 17786 9312
rect 17820 9044 17858 9312
rect 17770 9028 17858 9044
rect 19458 9312 19546 9328
rect 19458 9044 19496 9312
rect 19530 9044 19546 9312
rect 19458 9028 19546 9044
rect 19971 9313 20059 9329
rect 19971 9045 19987 9313
rect 20021 9045 20059 9313
rect 19971 9029 20059 9045
rect 21659 9313 21747 9329
rect 21659 9045 21697 9313
rect 21731 9045 21747 9313
rect 21659 9029 21747 9045
rect 171 8513 259 8529
rect 171 8245 187 8513
rect 221 8245 259 8513
rect 171 8229 259 8245
rect 1859 8513 1947 8529
rect 1859 8245 1897 8513
rect 1931 8245 1947 8513
rect 1859 8229 1947 8245
rect 2370 8512 2458 8528
rect 2370 8244 2386 8512
rect 2420 8244 2458 8512
rect 2370 8228 2458 8244
rect 4058 8512 4146 8528
rect 4058 8244 4096 8512
rect 4130 8244 4146 8512
rect 4058 8228 4146 8244
rect 4570 8512 4658 8528
rect 4570 8244 4586 8512
rect 4620 8244 4658 8512
rect 4570 8228 4658 8244
rect 6258 8512 6346 8528
rect 6258 8244 6296 8512
rect 6330 8244 6346 8512
rect 6258 8228 6346 8244
rect 6770 8512 6858 8528
rect 6770 8244 6786 8512
rect 6820 8244 6858 8512
rect 6770 8228 6858 8244
rect 8458 8512 8546 8528
rect 8458 8244 8496 8512
rect 8530 8244 8546 8512
rect 8458 8228 8546 8244
rect 8970 8512 9058 8528
rect 8970 8244 8986 8512
rect 9020 8244 9058 8512
rect 8970 8228 9058 8244
rect 10658 8512 10746 8528
rect 10658 8244 10696 8512
rect 10730 8244 10746 8512
rect 10658 8228 10746 8244
rect 11170 8512 11258 8528
rect 11170 8244 11186 8512
rect 11220 8244 11258 8512
rect 11170 8228 11258 8244
rect 12858 8512 12946 8528
rect 12858 8244 12896 8512
rect 12930 8244 12946 8512
rect 12858 8228 12946 8244
rect 13370 8512 13458 8528
rect 13370 8244 13386 8512
rect 13420 8244 13458 8512
rect 13370 8228 13458 8244
rect 15058 8512 15146 8528
rect 15058 8244 15096 8512
rect 15130 8244 15146 8512
rect 15058 8228 15146 8244
rect 15570 8512 15658 8528
rect 15570 8244 15586 8512
rect 15620 8244 15658 8512
rect 15570 8228 15658 8244
rect 17258 8512 17346 8528
rect 17258 8244 17296 8512
rect 17330 8244 17346 8512
rect 17258 8228 17346 8244
rect 17770 8512 17858 8528
rect 17770 8244 17786 8512
rect 17820 8244 17858 8512
rect 17770 8228 17858 8244
rect 19458 8512 19546 8528
rect 19458 8244 19496 8512
rect 19530 8244 19546 8512
rect 19458 8228 19546 8244
rect 19971 8513 20059 8529
rect 19971 8245 19987 8513
rect 20021 8245 20059 8513
rect 19971 8229 20059 8245
rect 21659 8513 21747 8529
rect 21659 8245 21697 8513
rect 21731 8245 21747 8513
rect 21659 8229 21747 8245
rect 171 7713 259 7729
rect 171 7445 187 7713
rect 221 7445 259 7713
rect 171 7429 259 7445
rect 1859 7713 1947 7729
rect 1859 7445 1897 7713
rect 1931 7445 1947 7713
rect 1859 7429 1947 7445
rect 2370 7712 2458 7728
rect 2370 7444 2386 7712
rect 2420 7444 2458 7712
rect 2370 7428 2458 7444
rect 4058 7712 4146 7728
rect 4058 7444 4096 7712
rect 4130 7444 4146 7712
rect 4058 7428 4146 7444
rect 4570 7712 4658 7728
rect 4570 7444 4586 7712
rect 4620 7444 4658 7712
rect 4570 7428 4658 7444
rect 6258 7712 6346 7728
rect 6258 7444 6296 7712
rect 6330 7444 6346 7712
rect 6258 7428 6346 7444
rect 6770 7712 6858 7728
rect 6770 7444 6786 7712
rect 6820 7444 6858 7712
rect 6770 7428 6858 7444
rect 8458 7712 8546 7728
rect 8458 7444 8496 7712
rect 8530 7444 8546 7712
rect 8458 7428 8546 7444
rect 8970 7712 9058 7728
rect 8970 7444 8986 7712
rect 9020 7444 9058 7712
rect 8970 7428 9058 7444
rect 10658 7712 10746 7728
rect 10658 7444 10696 7712
rect 10730 7444 10746 7712
rect 10658 7428 10746 7444
rect 11170 7712 11258 7728
rect 11170 7444 11186 7712
rect 11220 7444 11258 7712
rect 11170 7428 11258 7444
rect 12858 7712 12946 7728
rect 12858 7444 12896 7712
rect 12930 7444 12946 7712
rect 12858 7428 12946 7444
rect 13370 7712 13458 7728
rect 13370 7444 13386 7712
rect 13420 7444 13458 7712
rect 13370 7428 13458 7444
rect 15058 7712 15146 7728
rect 15058 7444 15096 7712
rect 15130 7444 15146 7712
rect 15058 7428 15146 7444
rect 15570 7712 15658 7728
rect 15570 7444 15586 7712
rect 15620 7444 15658 7712
rect 15570 7428 15658 7444
rect 17258 7712 17346 7728
rect 17258 7444 17296 7712
rect 17330 7444 17346 7712
rect 17258 7428 17346 7444
rect 17770 7712 17858 7728
rect 17770 7444 17786 7712
rect 17820 7444 17858 7712
rect 17770 7428 17858 7444
rect 19458 7712 19546 7728
rect 19458 7444 19496 7712
rect 19530 7444 19546 7712
rect 19458 7428 19546 7444
rect 19971 7713 20059 7729
rect 19971 7445 19987 7713
rect 20021 7445 20059 7713
rect 19971 7429 20059 7445
rect 21659 7713 21747 7729
rect 21659 7445 21697 7713
rect 21731 7445 21747 7713
rect 21659 7429 21747 7445
rect 171 6913 259 6929
rect 171 6645 187 6913
rect 221 6645 259 6913
rect 171 6629 259 6645
rect 1859 6913 1947 6929
rect 1859 6645 1897 6913
rect 1931 6645 1947 6913
rect 1859 6629 1947 6645
rect 2370 6912 2458 6928
rect 2370 6644 2386 6912
rect 2420 6644 2458 6912
rect 2370 6628 2458 6644
rect 4058 6912 4146 6928
rect 4058 6644 4096 6912
rect 4130 6644 4146 6912
rect 4058 6628 4146 6644
rect 4570 6912 4658 6928
rect 4570 6644 4586 6912
rect 4620 6644 4658 6912
rect 4570 6628 4658 6644
rect 6258 6912 6346 6928
rect 6258 6644 6296 6912
rect 6330 6644 6346 6912
rect 6258 6628 6346 6644
rect 6770 6912 6858 6928
rect 6770 6644 6786 6912
rect 6820 6644 6858 6912
rect 6770 6628 6858 6644
rect 8458 6912 8546 6928
rect 8458 6644 8496 6912
rect 8530 6644 8546 6912
rect 8458 6628 8546 6644
rect 8970 6912 9058 6928
rect 8970 6644 8986 6912
rect 9020 6644 9058 6912
rect 8970 6628 9058 6644
rect 10658 6912 10746 6928
rect 10658 6644 10696 6912
rect 10730 6644 10746 6912
rect 10658 6628 10746 6644
rect 11170 6912 11258 6928
rect 11170 6644 11186 6912
rect 11220 6644 11258 6912
rect 11170 6628 11258 6644
rect 12858 6912 12946 6928
rect 12858 6644 12896 6912
rect 12930 6644 12946 6912
rect 12858 6628 12946 6644
rect 13370 6912 13458 6928
rect 13370 6644 13386 6912
rect 13420 6644 13458 6912
rect 13370 6628 13458 6644
rect 15058 6912 15146 6928
rect 15058 6644 15096 6912
rect 15130 6644 15146 6912
rect 15058 6628 15146 6644
rect 15570 6912 15658 6928
rect 15570 6644 15586 6912
rect 15620 6644 15658 6912
rect 15570 6628 15658 6644
rect 17258 6912 17346 6928
rect 17258 6644 17296 6912
rect 17330 6644 17346 6912
rect 17258 6628 17346 6644
rect 17770 6912 17858 6928
rect 17770 6644 17786 6912
rect 17820 6644 17858 6912
rect 17770 6628 17858 6644
rect 19458 6912 19546 6928
rect 19458 6644 19496 6912
rect 19530 6644 19546 6912
rect 19458 6628 19546 6644
rect 19971 6913 20059 6929
rect 19971 6645 19987 6913
rect 20021 6645 20059 6913
rect 19971 6629 20059 6645
rect 21659 6913 21747 6929
rect 21659 6645 21697 6913
rect 21731 6645 21747 6913
rect 21659 6629 21747 6645
rect 171 6113 259 6129
rect 171 5845 187 6113
rect 221 5845 259 6113
rect 171 5829 259 5845
rect 1859 6113 1947 6129
rect 1859 5845 1897 6113
rect 1931 5845 1947 6113
rect 1859 5829 1947 5845
rect 2370 6112 2458 6128
rect 2370 5844 2386 6112
rect 2420 5844 2458 6112
rect 2370 5828 2458 5844
rect 4058 6112 4146 6128
rect 4058 5844 4096 6112
rect 4130 5844 4146 6112
rect 4058 5828 4146 5844
rect 4570 6112 4658 6128
rect 4570 5844 4586 6112
rect 4620 5844 4658 6112
rect 4570 5828 4658 5844
rect 6258 6112 6346 6128
rect 6258 5844 6296 6112
rect 6330 5844 6346 6112
rect 6258 5828 6346 5844
rect 6770 6112 6858 6128
rect 6770 5844 6786 6112
rect 6820 5844 6858 6112
rect 6770 5828 6858 5844
rect 8458 6112 8546 6128
rect 8458 5844 8496 6112
rect 8530 5844 8546 6112
rect 8458 5828 8546 5844
rect 8970 6112 9058 6128
rect 8970 5844 8986 6112
rect 9020 5844 9058 6112
rect 8970 5828 9058 5844
rect 10658 6112 10746 6128
rect 10658 5844 10696 6112
rect 10730 5844 10746 6112
rect 10658 5828 10746 5844
rect 11170 6112 11258 6128
rect 11170 5844 11186 6112
rect 11220 5844 11258 6112
rect 11170 5828 11258 5844
rect 12858 6112 12946 6128
rect 12858 5844 12896 6112
rect 12930 5844 12946 6112
rect 12858 5828 12946 5844
rect 13370 6112 13458 6128
rect 13370 5844 13386 6112
rect 13420 5844 13458 6112
rect 13370 5828 13458 5844
rect 15058 6112 15146 6128
rect 15058 5844 15096 6112
rect 15130 5844 15146 6112
rect 15058 5828 15146 5844
rect 15570 6112 15658 6128
rect 15570 5844 15586 6112
rect 15620 5844 15658 6112
rect 15570 5828 15658 5844
rect 17258 6112 17346 6128
rect 17258 5844 17296 6112
rect 17330 5844 17346 6112
rect 17258 5828 17346 5844
rect 17770 6112 17858 6128
rect 17770 5844 17786 6112
rect 17820 5844 17858 6112
rect 17770 5828 17858 5844
rect 19458 6112 19546 6128
rect 19458 5844 19496 6112
rect 19530 5844 19546 6112
rect 19458 5828 19546 5844
rect 19971 6113 20059 6129
rect 19971 5845 19987 6113
rect 20021 5845 20059 6113
rect 19971 5829 20059 5845
rect 21659 6113 21747 6129
rect 21659 5845 21697 6113
rect 21731 5845 21747 6113
rect 21659 5829 21747 5845
rect 171 5313 259 5329
rect 171 5045 187 5313
rect 221 5045 259 5313
rect 171 5029 259 5045
rect 1859 5313 1947 5329
rect 1859 5045 1897 5313
rect 1931 5045 1947 5313
rect 1859 5029 1947 5045
rect 2370 5312 2458 5328
rect 2370 5044 2386 5312
rect 2420 5044 2458 5312
rect 2370 5028 2458 5044
rect 4058 5312 4146 5328
rect 4058 5044 4096 5312
rect 4130 5044 4146 5312
rect 4058 5028 4146 5044
rect 4570 5312 4658 5328
rect 4570 5044 4586 5312
rect 4620 5044 4658 5312
rect 4570 5028 4658 5044
rect 6258 5312 6346 5328
rect 6258 5044 6296 5312
rect 6330 5044 6346 5312
rect 6258 5028 6346 5044
rect 6770 5312 6858 5328
rect 6770 5044 6786 5312
rect 6820 5044 6858 5312
rect 6770 5028 6858 5044
rect 8458 5312 8546 5328
rect 8458 5044 8496 5312
rect 8530 5044 8546 5312
rect 8458 5028 8546 5044
rect 8970 5312 9058 5328
rect 8970 5044 8986 5312
rect 9020 5044 9058 5312
rect 8970 5028 9058 5044
rect 10658 5312 10746 5328
rect 10658 5044 10696 5312
rect 10730 5044 10746 5312
rect 10658 5028 10746 5044
rect 11170 5312 11258 5328
rect 11170 5044 11186 5312
rect 11220 5044 11258 5312
rect 11170 5028 11258 5044
rect 12858 5312 12946 5328
rect 12858 5044 12896 5312
rect 12930 5044 12946 5312
rect 12858 5028 12946 5044
rect 13370 5312 13458 5328
rect 13370 5044 13386 5312
rect 13420 5044 13458 5312
rect 13370 5028 13458 5044
rect 15058 5312 15146 5328
rect 15058 5044 15096 5312
rect 15130 5044 15146 5312
rect 15058 5028 15146 5044
rect 15570 5312 15658 5328
rect 15570 5044 15586 5312
rect 15620 5044 15658 5312
rect 15570 5028 15658 5044
rect 17258 5312 17346 5328
rect 17258 5044 17296 5312
rect 17330 5044 17346 5312
rect 17258 5028 17346 5044
rect 17770 5312 17858 5328
rect 17770 5044 17786 5312
rect 17820 5044 17858 5312
rect 17770 5028 17858 5044
rect 19458 5312 19546 5328
rect 19458 5044 19496 5312
rect 19530 5044 19546 5312
rect 19458 5028 19546 5044
rect 19971 5313 20059 5329
rect 19971 5045 19987 5313
rect 20021 5045 20059 5313
rect 19971 5029 20059 5045
rect 21659 5313 21747 5329
rect 21659 5045 21697 5313
rect 21731 5045 21747 5313
rect 21659 5029 21747 5045
rect 171 4513 259 4529
rect 171 4245 187 4513
rect 221 4245 259 4513
rect 171 4229 259 4245
rect 1859 4513 1947 4529
rect 1859 4245 1897 4513
rect 1931 4245 1947 4513
rect 1859 4229 1947 4245
rect 2371 4513 2459 4529
rect 2371 4245 2387 4513
rect 2421 4245 2459 4513
rect 2371 4229 2459 4245
rect 4059 4513 4147 4529
rect 4059 4245 4097 4513
rect 4131 4245 4147 4513
rect 4059 4229 4147 4245
rect 4571 4513 4659 4529
rect 4571 4245 4587 4513
rect 4621 4245 4659 4513
rect 4571 4229 4659 4245
rect 6259 4513 6347 4529
rect 6259 4245 6297 4513
rect 6331 4245 6347 4513
rect 6259 4229 6347 4245
rect 6771 4513 6859 4529
rect 6771 4245 6787 4513
rect 6821 4245 6859 4513
rect 6771 4229 6859 4245
rect 8459 4513 8547 4529
rect 8459 4245 8497 4513
rect 8531 4245 8547 4513
rect 8459 4229 8547 4245
rect 8972 4514 9060 4530
rect 8972 4246 8988 4514
rect 9022 4246 9060 4514
rect 8972 4230 9060 4246
rect 10660 4514 10748 4530
rect 10660 4246 10698 4514
rect 10732 4246 10748 4514
rect 10660 4230 10748 4246
rect 11172 4514 11260 4530
rect 11172 4246 11188 4514
rect 11222 4246 11260 4514
rect 11172 4230 11260 4246
rect 12860 4514 12948 4530
rect 12860 4246 12898 4514
rect 12932 4246 12948 4514
rect 12860 4230 12948 4246
rect 13371 4513 13459 4529
rect 13371 4245 13387 4513
rect 13421 4245 13459 4513
rect 13371 4229 13459 4245
rect 15059 4513 15147 4529
rect 15059 4245 15097 4513
rect 15131 4245 15147 4513
rect 15059 4229 15147 4245
rect 15571 4513 15659 4529
rect 15571 4245 15587 4513
rect 15621 4245 15659 4513
rect 15571 4229 15659 4245
rect 17259 4513 17347 4529
rect 17259 4245 17297 4513
rect 17331 4245 17347 4513
rect 17259 4229 17347 4245
rect 17771 4513 17859 4529
rect 17771 4245 17787 4513
rect 17821 4245 17859 4513
rect 17771 4229 17859 4245
rect 19459 4513 19547 4529
rect 19459 4245 19497 4513
rect 19531 4245 19547 4513
rect 19459 4229 19547 4245
rect 19971 4513 20059 4529
rect 19971 4245 19987 4513
rect 20021 4245 20059 4513
rect 19971 4229 20059 4245
rect 21659 4513 21747 4529
rect 21659 4245 21697 4513
rect 21731 4245 21747 4513
rect 21659 4229 21747 4245
rect 27900 11312 27926 11412
rect 28726 11396 28823 11412
rect 28726 11328 28773 11396
rect 28807 11328 28823 11396
rect 28726 11312 28823 11328
rect 27900 11154 27926 11254
rect 28726 11238 28823 11254
rect 28726 11170 28773 11238
rect 28807 11170 28823 11238
rect 28726 11154 28823 11170
rect 27900 10996 27926 11096
rect 28726 11080 28823 11096
rect 28726 11012 28773 11080
rect 28807 11012 28823 11080
rect 28726 10996 28823 11012
rect 27900 10838 27926 10938
rect 28726 10922 28823 10938
rect 28726 10854 28773 10922
rect 28807 10854 28823 10922
rect 28726 10838 28823 10854
rect 30148 11799 30248 11815
rect 30148 11765 30164 11799
rect 30232 11765 30248 11799
rect 30148 11727 30248 11765
rect 30306 11799 30406 11815
rect 30306 11765 30322 11799
rect 30390 11765 30406 11799
rect 30306 11727 30406 11765
rect 30464 11799 30564 11815
rect 30464 11765 30480 11799
rect 30548 11765 30564 11799
rect 30464 11727 30564 11765
rect 30148 11489 30248 11527
rect 30148 11455 30164 11489
rect 30232 11455 30248 11489
rect 30148 11439 30248 11455
rect 30306 11489 30406 11527
rect 30306 11455 30322 11489
rect 30390 11455 30406 11489
rect 30306 11439 30406 11455
rect 30464 11489 30564 11527
rect 30464 11455 30480 11489
rect 30548 11455 30564 11489
rect 30464 11439 30564 11455
rect 30903 11799 31003 11815
rect 30903 11765 30919 11799
rect 30987 11765 31003 11799
rect 30903 11727 31003 11765
rect 30903 11489 31003 11527
rect 30903 11455 30919 11489
rect 30987 11455 31003 11489
rect 30903 11439 31003 11455
rect 31343 11799 31443 11815
rect 31343 11765 31359 11799
rect 31427 11765 31443 11799
rect 31343 11727 31443 11765
rect 31343 11489 31443 11527
rect 31343 11455 31359 11489
rect 31427 11455 31443 11489
rect 31343 11439 31443 11455
rect 31783 11799 31883 11815
rect 31783 11765 31799 11799
rect 31867 11765 31883 11799
rect 31783 11727 31883 11765
rect 31783 11489 31883 11527
rect 31783 11455 31799 11489
rect 31867 11455 31883 11489
rect 31783 11439 31883 11455
rect 32348 11799 32448 11815
rect 32348 11765 32364 11799
rect 32432 11765 32448 11799
rect 32348 11727 32448 11765
rect 32506 11799 32606 11815
rect 32506 11765 32522 11799
rect 32590 11765 32606 11799
rect 32506 11727 32606 11765
rect 32664 11799 32764 11815
rect 32664 11765 32680 11799
rect 32748 11765 32764 11799
rect 32664 11727 32764 11765
rect 32348 11489 32448 11527
rect 32348 11455 32364 11489
rect 32432 11455 32448 11489
rect 32348 11439 32448 11455
rect 32506 11489 32606 11527
rect 32506 11455 32522 11489
rect 32590 11455 32606 11489
rect 32506 11439 32606 11455
rect 32664 11489 32764 11527
rect 32664 11455 32680 11489
rect 32748 11455 32764 11489
rect 32664 11439 32764 11455
rect 33103 11799 33203 11815
rect 33103 11765 33119 11799
rect 33187 11765 33203 11799
rect 33103 11727 33203 11765
rect 33103 11489 33203 11527
rect 33103 11455 33119 11489
rect 33187 11455 33203 11489
rect 33103 11439 33203 11455
rect 33543 11799 33643 11815
rect 33543 11765 33559 11799
rect 33627 11765 33643 11799
rect 33543 11727 33643 11765
rect 33543 11489 33643 11527
rect 33543 11455 33559 11489
rect 33627 11455 33643 11489
rect 33543 11439 33643 11455
rect 33983 11799 34083 11815
rect 33983 11765 33999 11799
rect 34067 11765 34083 11799
rect 33983 11727 34083 11765
rect 33983 11489 34083 11527
rect 33983 11455 33999 11489
rect 34067 11455 34083 11489
rect 33983 11439 34083 11455
rect 34548 11799 34648 11815
rect 34548 11765 34564 11799
rect 34632 11765 34648 11799
rect 34548 11727 34648 11765
rect 34706 11799 34806 11815
rect 34706 11765 34722 11799
rect 34790 11765 34806 11799
rect 34706 11727 34806 11765
rect 34864 11799 34964 11815
rect 34864 11765 34880 11799
rect 34948 11765 34964 11799
rect 34864 11727 34964 11765
rect 34548 11489 34648 11527
rect 34548 11455 34564 11489
rect 34632 11455 34648 11489
rect 34548 11439 34648 11455
rect 34706 11489 34806 11527
rect 34706 11455 34722 11489
rect 34790 11455 34806 11489
rect 34706 11439 34806 11455
rect 34864 11489 34964 11527
rect 34864 11455 34880 11489
rect 34948 11455 34964 11489
rect 34864 11439 34964 11455
rect 35303 11799 35403 11815
rect 35303 11765 35319 11799
rect 35387 11765 35403 11799
rect 35303 11727 35403 11765
rect 35303 11489 35403 11527
rect 35303 11455 35319 11489
rect 35387 11455 35403 11489
rect 35303 11439 35403 11455
rect 35743 11799 35843 11815
rect 35743 11765 35759 11799
rect 35827 11765 35843 11799
rect 35743 11727 35843 11765
rect 35743 11489 35843 11527
rect 35743 11455 35759 11489
rect 35827 11455 35843 11489
rect 35743 11439 35843 11455
rect 36183 11799 36283 11815
rect 36183 11765 36199 11799
rect 36267 11765 36283 11799
rect 36183 11727 36283 11765
rect 36183 11489 36283 11527
rect 36183 11455 36199 11489
rect 36267 11455 36283 11489
rect 36183 11439 36283 11455
rect 30190 10988 30590 11004
rect 30190 10954 30206 10988
rect 30574 10954 30590 10988
rect 30190 10907 30590 10954
rect 30190 10760 30590 10807
rect 30190 10726 30206 10760
rect 30574 10726 30590 10760
rect 30190 10710 30590 10726
rect 30904 10988 31004 11004
rect 30904 10954 30920 10988
rect 30988 10954 31004 10988
rect 30904 10907 31004 10954
rect 27900 10272 27926 10372
rect 28726 10356 28823 10372
rect 28726 10288 28773 10356
rect 28807 10288 28823 10356
rect 28726 10272 28823 10288
rect 27900 10114 27926 10214
rect 28726 10198 28823 10214
rect 28726 10130 28773 10198
rect 28807 10130 28823 10198
rect 28726 10114 28823 10130
rect 27900 9956 27926 10056
rect 28726 10040 28823 10056
rect 28726 9972 28773 10040
rect 28807 9972 28823 10040
rect 28726 9956 28823 9972
rect 27900 9798 27926 9898
rect 28726 9882 28823 9898
rect 28726 9814 28773 9882
rect 28807 9814 28823 9882
rect 28726 9798 28823 9814
rect 30904 10460 31004 10507
rect 30904 10426 30920 10460
rect 30988 10426 31004 10460
rect 30904 10410 31004 10426
rect 31344 10988 31444 11004
rect 31344 10954 31360 10988
rect 31428 10954 31444 10988
rect 31344 10907 31444 10954
rect 31344 10460 31444 10507
rect 31344 10426 31360 10460
rect 31428 10426 31444 10460
rect 31344 10410 31444 10426
rect 31784 10988 31884 11004
rect 31784 10954 31800 10988
rect 31868 10954 31884 10988
rect 31784 10907 31884 10954
rect 31784 10460 31884 10507
rect 31784 10426 31800 10460
rect 31868 10426 31884 10460
rect 31784 10410 31884 10426
rect 32390 10988 32790 11004
rect 32390 10954 32406 10988
rect 32774 10954 32790 10988
rect 32390 10907 32790 10954
rect 32390 10760 32790 10807
rect 32390 10726 32406 10760
rect 32774 10726 32790 10760
rect 32390 10710 32790 10726
rect 33104 10988 33204 11004
rect 33104 10954 33120 10988
rect 33188 10954 33204 10988
rect 33104 10907 33204 10954
rect 33104 10460 33204 10507
rect 33104 10426 33120 10460
rect 33188 10426 33204 10460
rect 33104 10410 33204 10426
rect 33544 10988 33644 11004
rect 33544 10954 33560 10988
rect 33628 10954 33644 10988
rect 33544 10907 33644 10954
rect 33544 10460 33644 10507
rect 33544 10426 33560 10460
rect 33628 10426 33644 10460
rect 33544 10410 33644 10426
rect 33984 10988 34084 11004
rect 33984 10954 34000 10988
rect 34068 10954 34084 10988
rect 33984 10907 34084 10954
rect 33984 10460 34084 10507
rect 33984 10426 34000 10460
rect 34068 10426 34084 10460
rect 33984 10410 34084 10426
rect 34590 10988 34990 11004
rect 34590 10954 34606 10988
rect 34974 10954 34990 10988
rect 34590 10907 34990 10954
rect 34590 10760 34990 10807
rect 34590 10726 34606 10760
rect 34974 10726 34990 10760
rect 34590 10710 34990 10726
rect 35304 10988 35404 11004
rect 35304 10954 35320 10988
rect 35388 10954 35404 10988
rect 35304 10907 35404 10954
rect 35304 10460 35404 10507
rect 35304 10426 35320 10460
rect 35388 10426 35404 10460
rect 35304 10410 35404 10426
rect 35744 10988 35844 11004
rect 35744 10954 35760 10988
rect 35828 10954 35844 10988
rect 35744 10907 35844 10954
rect 35744 10460 35844 10507
rect 35744 10426 35760 10460
rect 35828 10426 35844 10460
rect 35744 10410 35844 10426
rect 36184 10988 36284 11004
rect 36184 10954 36200 10988
rect 36268 10954 36284 10988
rect 36184 10907 36284 10954
rect 36184 10460 36284 10507
rect 36184 10426 36200 10460
rect 36268 10426 36284 10460
rect 36184 10410 36284 10426
rect 27900 9232 27926 9332
rect 28726 9316 28823 9332
rect 28726 9248 28773 9316
rect 28807 9248 28823 9316
rect 28726 9232 28823 9248
rect 27900 9074 27926 9174
rect 28726 9158 28823 9174
rect 28726 9090 28773 9158
rect 28807 9090 28823 9158
rect 28726 9074 28823 9090
rect 27900 8916 27926 9016
rect 28726 9000 28823 9016
rect 28726 8932 28773 9000
rect 28807 8932 28823 9000
rect 28726 8916 28823 8932
rect 27900 8758 27926 8858
rect 28726 8842 28823 8858
rect 28726 8774 28773 8842
rect 28807 8774 28823 8842
rect 28726 8758 28823 8774
rect 29778 9678 30578 9694
rect 29778 9644 29794 9678
rect 30562 9644 30578 9678
rect 29778 9597 30578 9644
rect 30636 9678 31436 9694
rect 30636 9644 30652 9678
rect 31420 9644 31436 9678
rect 30636 9597 31436 9644
rect 29778 9150 30578 9197
rect 29778 9116 29794 9150
rect 30562 9116 30578 9150
rect 29778 9100 30578 9116
rect 30636 9150 31436 9197
rect 30636 9116 30652 9150
rect 31420 9116 31436 9150
rect 30636 9100 31436 9116
rect 27900 8192 27926 8292
rect 28726 8276 28823 8292
rect 28726 8208 28773 8276
rect 28807 8208 28823 8276
rect 28726 8192 28823 8208
rect 27900 8034 27926 8134
rect 28726 8118 28823 8134
rect 28726 8050 28773 8118
rect 28807 8050 28823 8118
rect 28726 8034 28823 8050
rect 27900 7876 27926 7976
rect 28726 7960 28823 7976
rect 28726 7892 28773 7960
rect 28807 7892 28823 7960
rect 28726 7876 28823 7892
rect 27900 7718 27926 7818
rect 28726 7802 28823 7818
rect 28726 7734 28773 7802
rect 28807 7734 28823 7802
rect 28726 7718 28823 7734
rect 27900 7152 27926 7252
rect 28726 7236 28823 7252
rect 28726 7168 28773 7236
rect 28807 7168 28823 7236
rect 28726 7152 28823 7168
rect 27900 6994 27926 7094
rect 28726 7078 28823 7094
rect 28726 7010 28773 7078
rect 28807 7010 28823 7078
rect 28726 6994 28823 7010
rect 27900 6836 27926 6936
rect 28726 6920 28823 6936
rect 28726 6852 28773 6920
rect 28807 6852 28823 6920
rect 28726 6836 28823 6852
rect 27900 6678 27926 6778
rect 28726 6762 28823 6778
rect 28726 6694 28773 6762
rect 28807 6694 28823 6762
rect 28726 6678 28823 6694
rect 29778 8674 30578 8690
rect 29778 8640 29794 8674
rect 30562 8640 30578 8674
rect 29778 8593 30578 8640
rect 30636 8674 31436 8690
rect 30636 8640 30652 8674
rect 31420 8640 31436 8674
rect 30636 8593 31436 8640
rect 29778 8146 30578 8193
rect 29778 8112 29794 8146
rect 30562 8112 30578 8146
rect 29778 8096 30578 8112
rect 30636 8146 31436 8193
rect 30636 8112 30652 8146
rect 31420 8112 31436 8146
rect 30636 8096 31436 8112
rect 29778 8038 30578 8054
rect 29778 8004 29794 8038
rect 30562 8004 30578 8038
rect 29778 7957 30578 8004
rect 30636 8038 31436 8054
rect 30636 8004 30652 8038
rect 31420 8004 31436 8038
rect 30636 7957 31436 8004
rect 29778 7510 30578 7557
rect 29778 7476 29794 7510
rect 30562 7476 30578 7510
rect 29778 7460 30578 7476
rect 30636 7510 31436 7557
rect 30636 7476 30652 7510
rect 31420 7476 31436 7510
rect 30636 7460 31436 7476
rect 32956 8940 33156 8956
rect 32956 8906 32972 8940
rect 33140 8906 33156 8940
rect 32956 8859 33156 8906
rect 33214 8940 33414 8956
rect 33214 8906 33230 8940
rect 33398 8906 33414 8940
rect 33214 8859 33414 8906
rect 32956 8012 33156 8059
rect 32956 7978 32972 8012
rect 33140 7978 33156 8012
rect 32956 7962 33156 7978
rect 33214 8012 33414 8059
rect 33214 7978 33230 8012
rect 33398 7978 33414 8012
rect 33214 7962 33414 7978
rect 33796 8940 33996 8956
rect 33796 8906 33812 8940
rect 33980 8906 33996 8940
rect 33796 8859 33996 8906
rect 34054 8940 34254 8956
rect 34054 8906 34070 8940
rect 34238 8906 34254 8940
rect 34054 8859 34254 8906
rect 33796 8012 33996 8059
rect 33796 7978 33812 8012
rect 33980 7978 33996 8012
rect 33796 7962 33996 7978
rect 34054 8012 34254 8059
rect 34054 7978 34070 8012
rect 34238 7978 34254 8012
rect 34054 7962 34254 7978
rect 34618 8720 34684 8736
rect 34618 8686 34634 8720
rect 34668 8686 34684 8720
rect 34618 8670 34684 8686
rect 34636 8639 34666 8670
rect 34636 8208 34666 8239
rect 34618 8192 34684 8208
rect 34618 8158 34634 8192
rect 34668 8158 34684 8192
rect 34618 8142 34684 8158
rect 35038 8720 35104 8736
rect 35038 8686 35054 8720
rect 35088 8686 35104 8720
rect 35038 8670 35104 8686
rect 35056 8639 35086 8670
rect 35056 8208 35086 8239
rect 35038 8192 35104 8208
rect 35038 8158 35054 8192
rect 35088 8158 35104 8192
rect 35038 8142 35104 8158
rect 35458 8720 35524 8736
rect 35458 8686 35474 8720
rect 35508 8686 35524 8720
rect 35458 8670 35524 8686
rect 35476 8639 35506 8670
rect 35476 8208 35506 8239
rect 35458 8192 35524 8208
rect 35458 8158 35474 8192
rect 35508 8158 35524 8192
rect 35458 8142 35524 8158
rect 29660 7002 29757 7018
rect 29660 6834 29676 7002
rect 29710 6834 29757 7002
rect 29660 6818 29757 6834
rect 30557 7002 30654 7018
rect 30557 6834 30604 7002
rect 30638 6834 30654 7002
rect 30557 6818 30654 6834
rect 31000 7002 31097 7018
rect 31000 6834 31016 7002
rect 31050 6834 31097 7002
rect 31000 6818 31097 6834
rect 31897 7002 31994 7018
rect 31897 6834 31944 7002
rect 31978 6834 31994 7002
rect 31897 6818 31994 6834
rect 33518 7510 33618 7526
rect 33518 7476 33534 7510
rect 33602 7476 33618 7510
rect 33518 7438 33618 7476
rect 33676 7510 33776 7526
rect 33676 7476 33692 7510
rect 33760 7476 33776 7510
rect 33676 7438 33776 7476
rect 33834 7510 33934 7526
rect 33834 7476 33850 7510
rect 33918 7476 33934 7510
rect 33834 7438 33934 7476
rect 33992 7510 34092 7526
rect 33992 7476 34008 7510
rect 34076 7476 34092 7510
rect 33992 7438 34092 7476
rect 33518 7000 33618 7038
rect 33518 6966 33534 7000
rect 33602 6966 33618 7000
rect 33518 6950 33618 6966
rect 33676 7000 33776 7038
rect 33676 6966 33692 7000
rect 33760 6966 33776 7000
rect 33676 6950 33776 6966
rect 33834 7000 33934 7038
rect 33834 6966 33850 7000
rect 33918 6966 33934 7000
rect 33834 6950 33934 6966
rect 33992 7000 34092 7038
rect 33992 6966 34008 7000
rect 34076 6966 34092 7000
rect 33992 6950 34092 6966
rect 34618 7402 34684 7418
rect 34618 7368 34634 7402
rect 34668 7368 34684 7402
rect 34618 7352 34684 7368
rect 34636 7330 34666 7352
rect 34636 7108 34666 7130
rect 34618 7092 34684 7108
rect 34618 7058 34634 7092
rect 34668 7058 34684 7092
rect 34618 7042 34684 7058
rect 35038 7402 35104 7418
rect 35038 7368 35054 7402
rect 35088 7368 35104 7402
rect 35038 7352 35104 7368
rect 35056 7330 35086 7352
rect 35056 7108 35086 7130
rect 35038 7092 35104 7108
rect 35038 7058 35054 7092
rect 35088 7058 35104 7092
rect 35038 7042 35104 7058
rect 35458 7402 35524 7418
rect 35458 7368 35474 7402
rect 35508 7368 35524 7402
rect 35458 7352 35524 7368
rect 35476 7330 35506 7352
rect 35476 7108 35506 7130
rect 35458 7092 35524 7108
rect 35458 7058 35474 7092
rect 35508 7058 35524 7092
rect 35458 7042 35524 7058
rect 27900 6112 27926 6212
rect 28726 6196 28823 6212
rect 28726 6128 28773 6196
rect 28807 6128 28823 6196
rect 28726 6112 28823 6128
rect 27900 5954 27926 6054
rect 28726 6038 28823 6054
rect 28726 5970 28773 6038
rect 28807 5970 28823 6038
rect 28726 5954 28823 5970
rect 27900 5796 27926 5896
rect 28726 5880 28823 5896
rect 28726 5812 28773 5880
rect 28807 5812 28823 5880
rect 28726 5796 28823 5812
rect 27900 5638 27926 5738
rect 28726 5722 28823 5738
rect 28726 5654 28773 5722
rect 28807 5654 28823 5722
rect 28726 5638 28823 5654
rect 29670 6172 29758 6188
rect 29670 6004 29686 6172
rect 29720 6004 29758 6172
rect 29670 5988 29758 6004
rect 30558 6172 30646 6188
rect 30558 6004 30596 6172
rect 30630 6004 30646 6172
rect 30558 5988 30646 6004
rect 31010 6172 31098 6188
rect 31010 6004 31026 6172
rect 31060 6004 31098 6172
rect 31010 5988 31098 6004
rect 31898 6172 31986 6188
rect 31898 6004 31936 6172
rect 31970 6004 31986 6172
rect 31898 5988 31986 6004
rect 27958 5238 28758 5254
rect 27958 5204 27974 5238
rect 28742 5204 28758 5238
rect 27958 5157 28758 5204
rect 27958 4310 28758 4357
rect 27958 4276 27974 4310
rect 28742 4276 28758 4310
rect 27958 4260 28758 4276
rect 29968 5580 30368 5596
rect 29968 5546 29984 5580
rect 30352 5546 30368 5580
rect 29968 5508 30368 5546
rect 29968 5370 30368 5408
rect 29968 5336 29984 5370
rect 30352 5336 30368 5370
rect 29968 5320 30368 5336
rect 31278 5580 31678 5596
rect 31278 5546 31294 5580
rect 31662 5546 31678 5580
rect 31278 5508 31678 5546
rect 31278 5370 31678 5408
rect 31278 5336 31294 5370
rect 31662 5336 31678 5370
rect 31278 5320 31678 5336
rect 29670 4912 29758 4928
rect 29670 4744 29686 4912
rect 29720 4744 29758 4912
rect 29670 4728 29758 4744
rect 30558 4912 30646 4928
rect 30558 4744 30596 4912
rect 30630 4744 30646 4912
rect 30558 4728 30646 4744
rect 31010 4912 31098 4928
rect 31010 4744 31026 4912
rect 31060 4744 31098 4912
rect 31010 4728 31098 4744
rect 31898 4912 31986 4928
rect 31898 4744 31936 4912
rect 31970 4744 31986 4912
rect 31898 4728 31986 4744
rect 17148 3388 17248 3404
rect 17148 3354 17164 3388
rect 17232 3354 17248 3388
rect 17148 3316 17248 3354
rect 17306 3388 17406 3404
rect 17306 3354 17322 3388
rect 17390 3354 17406 3388
rect 17306 3316 17406 3354
rect 17464 3388 17564 3404
rect 17464 3354 17480 3388
rect 17548 3354 17564 3388
rect 17464 3316 17564 3354
rect 17622 3388 17722 3404
rect 17622 3354 17638 3388
rect 17706 3354 17722 3388
rect 17622 3316 17722 3354
rect 17148 2490 17248 2516
rect 17306 2490 17406 2516
rect 17464 2490 17564 2516
rect 17622 2490 17722 2516
rect 32768 4030 32868 4046
rect 32768 3996 32784 4030
rect 32852 3996 32868 4030
rect 32768 3958 32868 3996
rect 32926 4030 33026 4046
rect 32926 3996 32942 4030
rect 33010 3996 33026 4030
rect 32926 3958 33026 3996
rect 33084 4030 33184 4046
rect 33084 3996 33100 4030
rect 33168 3996 33184 4030
rect 33084 3958 33184 3996
rect 33242 4030 33342 4046
rect 33242 3996 33258 4030
rect 33326 3996 33342 4030
rect 33242 3958 33342 3996
rect 33400 4030 33500 4046
rect 33400 3996 33416 4030
rect 33484 3996 33500 4030
rect 33400 3958 33500 3996
rect 33558 4030 33658 4046
rect 33558 3996 33574 4030
rect 33642 3996 33658 4030
rect 33558 3958 33658 3996
rect 33716 4030 33816 4046
rect 33716 3996 33732 4030
rect 33800 3996 33816 4030
rect 33716 3958 33816 3996
rect 33874 4030 33974 4046
rect 33874 3996 33890 4030
rect 33958 3996 33974 4030
rect 33874 3958 33974 3996
rect 32768 3520 32868 3558
rect 32768 3486 32784 3520
rect 32852 3486 32868 3520
rect 32768 3470 32868 3486
rect 32926 3520 33026 3558
rect 32926 3486 32942 3520
rect 33010 3486 33026 3520
rect 32926 3470 33026 3486
rect 33084 3520 33184 3558
rect 33084 3486 33100 3520
rect 33168 3486 33184 3520
rect 33084 3470 33184 3486
rect 33242 3520 33342 3558
rect 33242 3486 33258 3520
rect 33326 3486 33342 3520
rect 33242 3470 33342 3486
rect 33400 3520 33500 3558
rect 33400 3486 33416 3520
rect 33484 3486 33500 3520
rect 33400 3470 33500 3486
rect 33558 3520 33658 3558
rect 33558 3486 33574 3520
rect 33642 3486 33658 3520
rect 33558 3470 33658 3486
rect 33716 3520 33816 3558
rect 33716 3486 33732 3520
rect 33800 3486 33816 3520
rect 33716 3470 33816 3486
rect 33874 3520 33974 3558
rect 33874 3486 33890 3520
rect 33958 3486 33974 3520
rect 33874 3470 33974 3486
rect 34958 4030 35058 4046
rect 34958 3996 34974 4030
rect 35042 3996 35058 4030
rect 34958 3958 35058 3996
rect 35116 4030 35216 4046
rect 35116 3996 35132 4030
rect 35200 3996 35216 4030
rect 35116 3958 35216 3996
rect 35274 4030 35374 4046
rect 35274 3996 35290 4030
rect 35358 3996 35374 4030
rect 35274 3958 35374 3996
rect 34958 3520 35058 3558
rect 34958 3486 34974 3520
rect 35042 3486 35058 3520
rect 34958 3470 35058 3486
rect 35116 3520 35216 3558
rect 35116 3486 35132 3520
rect 35200 3486 35216 3520
rect 35116 3470 35216 3486
rect 35274 3520 35374 3558
rect 35274 3486 35290 3520
rect 35358 3486 35374 3520
rect 35274 3470 35374 3486
rect 36360 5938 36448 5954
rect 36360 5770 36376 5938
rect 36410 5770 36448 5938
rect 36360 5754 36448 5770
rect 36848 5938 36936 5954
rect 36848 5770 36886 5938
rect 36920 5770 36936 5938
rect 36848 5754 36936 5770
rect 36360 5680 36448 5696
rect 36360 5512 36376 5680
rect 36410 5512 36448 5680
rect 36360 5496 36448 5512
rect 36848 5680 36936 5696
rect 36848 5512 36886 5680
rect 36920 5512 36936 5680
rect 36848 5496 36936 5512
rect 36360 5422 36448 5438
rect 36360 5254 36376 5422
rect 36410 5254 36448 5422
rect 36360 5238 36448 5254
rect 36848 5422 36936 5438
rect 36848 5254 36886 5422
rect 36920 5254 36936 5422
rect 36848 5238 36936 5254
rect 36360 5164 36448 5180
rect 36360 4996 36376 5164
rect 36410 4996 36448 5164
rect 36360 4980 36448 4996
rect 36848 5164 36936 5180
rect 36848 4996 36886 5164
rect 36920 4996 36936 5164
rect 36848 4980 36936 4996
rect 36360 4906 36448 4922
rect 36360 4738 36376 4906
rect 36410 4738 36448 4906
rect 36360 4722 36448 4738
rect 36848 4906 36936 4922
rect 36848 4738 36886 4906
rect 36920 4738 36936 4906
rect 36848 4722 36936 4738
rect 36360 4648 36448 4664
rect 36360 4480 36376 4648
rect 36410 4480 36448 4648
rect 36360 4464 36448 4480
rect 36848 4648 36936 4664
rect 36848 4480 36886 4648
rect 36920 4480 36936 4648
rect 36848 4464 36936 4480
rect 36360 4390 36448 4406
rect 36360 4222 36376 4390
rect 36410 4222 36448 4390
rect 36360 4206 36448 4222
rect 36848 4390 36936 4406
rect 36848 4222 36886 4390
rect 36920 4222 36936 4390
rect 36848 4206 36936 4222
rect 36360 4132 36448 4148
rect 36360 3964 36376 4132
rect 36410 3964 36448 4132
rect 36360 3948 36448 3964
rect 36848 4132 36936 4148
rect 36848 3964 36886 4132
rect 36920 3964 36936 4132
rect 36848 3948 36936 3964
rect 37146 5938 37234 5954
rect 37146 5770 37162 5938
rect 37196 5770 37234 5938
rect 37146 5754 37234 5770
rect 37634 5938 37722 5954
rect 37634 5770 37672 5938
rect 37706 5770 37722 5938
rect 37634 5754 37722 5770
rect 37146 5680 37234 5696
rect 37146 5512 37162 5680
rect 37196 5512 37234 5680
rect 37146 5496 37234 5512
rect 37634 5680 37722 5696
rect 37634 5512 37672 5680
rect 37706 5512 37722 5680
rect 37634 5496 37722 5512
rect 37146 5422 37234 5438
rect 37146 5254 37162 5422
rect 37196 5254 37234 5422
rect 37146 5238 37234 5254
rect 37634 5422 37722 5438
rect 37634 5254 37672 5422
rect 37706 5254 37722 5422
rect 37634 5238 37722 5254
rect 37146 5164 37234 5180
rect 37146 4996 37162 5164
rect 37196 4996 37234 5164
rect 37146 4980 37234 4996
rect 37634 5164 37722 5180
rect 37634 4996 37672 5164
rect 37706 4996 37722 5164
rect 37634 4980 37722 4996
rect 37146 4906 37234 4922
rect 37146 4738 37162 4906
rect 37196 4738 37234 4906
rect 37146 4722 37234 4738
rect 37634 4906 37722 4922
rect 37634 4738 37672 4906
rect 37706 4738 37722 4906
rect 37634 4722 37722 4738
rect 37146 4648 37234 4664
rect 37146 4480 37162 4648
rect 37196 4480 37234 4648
rect 37146 4464 37234 4480
rect 37634 4648 37722 4664
rect 37634 4480 37672 4648
rect 37706 4480 37722 4648
rect 37634 4464 37722 4480
rect 37146 4390 37234 4406
rect 37146 4222 37162 4390
rect 37196 4222 37234 4390
rect 37146 4206 37234 4222
rect 37634 4390 37722 4406
rect 37634 4222 37672 4390
rect 37706 4222 37722 4390
rect 37634 4206 37722 4222
rect 37146 4132 37234 4148
rect 37146 3964 37162 4132
rect 37196 3964 37234 4132
rect 37146 3948 37234 3964
rect 37634 4132 37722 4148
rect 37634 3964 37672 4132
rect 37706 3964 37722 4132
rect 37634 3948 37722 3964
rect 32438 3100 32538 3116
rect 32438 3066 32454 3100
rect 32522 3066 32538 3100
rect 32438 3028 32538 3066
rect 32596 3100 32696 3116
rect 32596 3066 32612 3100
rect 32680 3066 32696 3100
rect 32596 3028 32696 3066
rect 32438 2590 32538 2628
rect 32438 2556 32454 2590
rect 32522 2556 32538 2590
rect 32438 2540 32538 2556
rect 32596 2590 32696 2628
rect 32596 2556 32612 2590
rect 32680 2556 32696 2590
rect 32596 2540 32696 2556
rect 34038 3100 34138 3116
rect 34038 3066 34054 3100
rect 34122 3066 34138 3100
rect 34038 3028 34138 3066
rect 34196 3100 34296 3116
rect 34196 3066 34212 3100
rect 34280 3066 34296 3100
rect 34196 3028 34296 3066
rect 34038 2590 34138 2628
rect 34038 2556 34054 2590
rect 34122 2556 34138 2590
rect 34038 2540 34138 2556
rect 34196 2590 34296 2628
rect 34196 2556 34212 2590
rect 34280 2556 34296 2590
rect 34196 2540 34296 2556
rect 35638 3100 35738 3116
rect 35638 3066 35654 3100
rect 35722 3066 35738 3100
rect 35638 3028 35738 3066
rect 35796 3100 35896 3116
rect 35796 3066 35812 3100
rect 35880 3066 35896 3100
rect 35796 3028 35896 3066
rect 35638 2590 35738 2628
rect 35638 2556 35654 2590
rect 35722 2556 35738 2590
rect 35638 2540 35738 2556
rect 35796 2590 35896 2628
rect 35796 2556 35812 2590
rect 35880 2556 35896 2590
rect 35796 2540 35896 2556
rect -29 2033 59 2049
rect -29 1265 -13 2033
rect 21 1265 59 2033
rect -29 1249 59 1265
rect 459 2033 547 2049
rect 459 1265 497 2033
rect 531 1265 547 2033
rect 459 1249 547 1265
rect 589 2033 677 2049
rect 589 1265 605 2033
rect 639 1265 677 2033
rect 589 1249 677 1265
rect 1077 2033 1165 2049
rect 1077 1265 1115 2033
rect 1149 1265 1165 2033
rect 1077 1249 1165 1265
rect -29 887 59 903
rect -29 719 -13 887
rect 21 719 59 887
rect -29 703 59 719
rect 459 887 547 903
rect 459 719 497 887
rect 531 719 547 887
rect 459 703 547 719
rect 589 887 677 903
rect 589 719 605 887
rect 639 719 677 887
rect 589 703 677 719
rect 1077 887 1165 903
rect 1077 719 1115 887
rect 1149 719 1165 887
rect 1077 703 1165 719
rect 1571 2033 1659 2049
rect 1571 1265 1587 2033
rect 1621 1265 1659 2033
rect 1571 1249 1659 1265
rect 2059 2033 2147 2049
rect 2059 1265 2097 2033
rect 2131 1265 2147 2033
rect 2059 1249 2147 1265
rect 2189 2033 2277 2049
rect 2189 1265 2205 2033
rect 2239 1265 2277 2033
rect 2189 1249 2277 1265
rect 2677 2033 2765 2049
rect 2677 1265 2715 2033
rect 2749 1265 2765 2033
rect 2677 1249 2765 1265
rect 1571 887 1659 903
rect 1571 719 1587 887
rect 1621 719 1659 887
rect 1571 703 1659 719
rect 2059 887 2147 903
rect 2059 719 2097 887
rect 2131 719 2147 887
rect 2059 703 2147 719
rect 2189 887 2277 903
rect 2189 719 2205 887
rect 2239 719 2277 887
rect 2189 703 2277 719
rect 2677 887 2765 903
rect 2677 719 2715 887
rect 2749 719 2765 887
rect 2677 703 2765 719
rect 3171 2033 3259 2049
rect 3171 1265 3187 2033
rect 3221 1265 3259 2033
rect 3171 1249 3259 1265
rect 3659 2033 3747 2049
rect 3659 1265 3697 2033
rect 3731 1265 3747 2033
rect 3659 1249 3747 1265
rect 3789 2033 3877 2049
rect 3789 1265 3805 2033
rect 3839 1265 3877 2033
rect 3789 1249 3877 1265
rect 4277 2033 4365 2049
rect 4277 1265 4315 2033
rect 4349 1265 4365 2033
rect 4277 1249 4365 1265
rect 3171 887 3259 903
rect 3171 719 3187 887
rect 3221 719 3259 887
rect 3171 703 3259 719
rect 3659 887 3747 903
rect 3659 719 3697 887
rect 3731 719 3747 887
rect 3659 703 3747 719
rect 3789 887 3877 903
rect 3789 719 3805 887
rect 3839 719 3877 887
rect 3789 703 3877 719
rect 4277 887 4365 903
rect 4277 719 4315 887
rect 4349 719 4365 887
rect 4277 703 4365 719
rect 4771 2033 4859 2049
rect 4771 1265 4787 2033
rect 4821 1265 4859 2033
rect 4771 1249 4859 1265
rect 5259 2033 5347 2049
rect 5259 1265 5297 2033
rect 5331 1265 5347 2033
rect 5259 1249 5347 1265
rect 5389 2033 5477 2049
rect 5389 1265 5405 2033
rect 5439 1265 5477 2033
rect 5389 1249 5477 1265
rect 5877 2033 5965 2049
rect 5877 1265 5915 2033
rect 5949 1265 5965 2033
rect 5877 1249 5965 1265
rect 4771 887 4859 903
rect 4771 719 4787 887
rect 4821 719 4859 887
rect 4771 703 4859 719
rect 5259 887 5347 903
rect 5259 719 5297 887
rect 5331 719 5347 887
rect 5259 703 5347 719
rect 5389 887 5477 903
rect 5389 719 5405 887
rect 5439 719 5477 887
rect 5389 703 5477 719
rect 5877 887 5965 903
rect 5877 719 5915 887
rect 5949 719 5965 887
rect 5877 703 5965 719
rect 6371 2033 6459 2049
rect 6371 1265 6387 2033
rect 6421 1265 6459 2033
rect 6371 1249 6459 1265
rect 6859 2033 6947 2049
rect 6859 1265 6897 2033
rect 6931 1265 6947 2033
rect 6859 1249 6947 1265
rect 6989 2033 7077 2049
rect 6989 1265 7005 2033
rect 7039 1265 7077 2033
rect 6989 1249 7077 1265
rect 7477 2033 7565 2049
rect 7477 1265 7515 2033
rect 7549 1265 7565 2033
rect 7477 1249 7565 1265
rect 6371 887 6459 903
rect 6371 719 6387 887
rect 6421 719 6459 887
rect 6371 703 6459 719
rect 6859 887 6947 903
rect 6859 719 6897 887
rect 6931 719 6947 887
rect 6859 703 6947 719
rect 6989 887 7077 903
rect 6989 719 7005 887
rect 7039 719 7077 887
rect 6989 703 7077 719
rect 7477 887 7565 903
rect 7477 719 7515 887
rect 7549 719 7565 887
rect 7477 703 7565 719
rect 7971 2033 8059 2049
rect 7971 1265 7987 2033
rect 8021 1265 8059 2033
rect 7971 1249 8059 1265
rect 8459 2033 8547 2049
rect 8459 1265 8497 2033
rect 8531 1265 8547 2033
rect 8459 1249 8547 1265
rect 8589 2033 8677 2049
rect 8589 1265 8605 2033
rect 8639 1265 8677 2033
rect 8589 1249 8677 1265
rect 9077 2033 9165 2049
rect 9077 1265 9115 2033
rect 9149 1265 9165 2033
rect 9077 1249 9165 1265
rect 7971 887 8059 903
rect 7971 719 7987 887
rect 8021 719 8059 887
rect 7971 703 8059 719
rect 8459 887 8547 903
rect 8459 719 8497 887
rect 8531 719 8547 887
rect 8459 703 8547 719
rect 8589 887 8677 903
rect 8589 719 8605 887
rect 8639 719 8677 887
rect 8589 703 8677 719
rect 9077 887 9165 903
rect 9077 719 9115 887
rect 9149 719 9165 887
rect 9077 703 9165 719
rect 9571 2033 9659 2049
rect 9571 1265 9587 2033
rect 9621 1265 9659 2033
rect 9571 1249 9659 1265
rect 10059 2033 10147 2049
rect 10059 1265 10097 2033
rect 10131 1265 10147 2033
rect 10059 1249 10147 1265
rect 10189 2033 10277 2049
rect 10189 1265 10205 2033
rect 10239 1265 10277 2033
rect 10189 1249 10277 1265
rect 10677 2033 10765 2049
rect 10677 1265 10715 2033
rect 10749 1265 10765 2033
rect 10677 1249 10765 1265
rect 9571 887 9659 903
rect 9571 719 9587 887
rect 9621 719 9659 887
rect 9571 703 9659 719
rect 10059 887 10147 903
rect 10059 719 10097 887
rect 10131 719 10147 887
rect 10059 703 10147 719
rect 10189 887 10277 903
rect 10189 719 10205 887
rect 10239 719 10277 887
rect 10189 703 10277 719
rect 10677 887 10765 903
rect 10677 719 10715 887
rect 10749 719 10765 887
rect 10677 703 10765 719
rect 11171 2033 11259 2049
rect 11171 1265 11187 2033
rect 11221 1265 11259 2033
rect 11171 1249 11259 1265
rect 11659 2033 11747 2049
rect 11659 1265 11697 2033
rect 11731 1265 11747 2033
rect 11659 1249 11747 1265
rect 11789 2033 11877 2049
rect 11789 1265 11805 2033
rect 11839 1265 11877 2033
rect 11789 1249 11877 1265
rect 12277 2033 12365 2049
rect 12277 1265 12315 2033
rect 12349 1265 12365 2033
rect 12277 1249 12365 1265
rect 11171 887 11259 903
rect 11171 719 11187 887
rect 11221 719 11259 887
rect 11171 703 11259 719
rect 11659 887 11747 903
rect 11659 719 11697 887
rect 11731 719 11747 887
rect 11659 703 11747 719
rect 11789 887 11877 903
rect 11789 719 11805 887
rect 11839 719 11877 887
rect 11789 703 11877 719
rect 12277 887 12365 903
rect 12277 719 12315 887
rect 12349 719 12365 887
rect 12277 703 12365 719
rect 12771 2033 12859 2049
rect 12771 1265 12787 2033
rect 12821 1265 12859 2033
rect 12771 1249 12859 1265
rect 13259 2033 13347 2049
rect 13259 1265 13297 2033
rect 13331 1265 13347 2033
rect 13259 1249 13347 1265
rect 13389 2033 13477 2049
rect 13389 1265 13405 2033
rect 13439 1265 13477 2033
rect 13389 1249 13477 1265
rect 13877 2033 13965 2049
rect 13877 1265 13915 2033
rect 13949 1265 13965 2033
rect 13877 1249 13965 1265
rect 12771 887 12859 903
rect 12771 719 12787 887
rect 12821 719 12859 887
rect 12771 703 12859 719
rect 13259 887 13347 903
rect 13259 719 13297 887
rect 13331 719 13347 887
rect 13259 703 13347 719
rect 13389 887 13477 903
rect 13389 719 13405 887
rect 13439 719 13477 887
rect 13389 703 13477 719
rect 13877 887 13965 903
rect 13877 719 13915 887
rect 13949 719 13965 887
rect 13877 703 13965 719
rect 14371 2033 14459 2049
rect 14371 1265 14387 2033
rect 14421 1265 14459 2033
rect 14371 1249 14459 1265
rect 14859 2033 14947 2049
rect 14859 1265 14897 2033
rect 14931 1265 14947 2033
rect 14859 1249 14947 1265
rect 14989 2033 15077 2049
rect 14989 1265 15005 2033
rect 15039 1265 15077 2033
rect 14989 1249 15077 1265
rect 15477 2033 15565 2049
rect 15477 1265 15515 2033
rect 15549 1265 15565 2033
rect 15477 1249 15565 1265
rect 14371 887 14459 903
rect 14371 719 14387 887
rect 14421 719 14459 887
rect 14371 703 14459 719
rect 14859 887 14947 903
rect 14859 719 14897 887
rect 14931 719 14947 887
rect 14859 703 14947 719
rect 14989 887 15077 903
rect 14989 719 15005 887
rect 15039 719 15077 887
rect 14989 703 15077 719
rect 15477 887 15565 903
rect 15477 719 15515 887
rect 15549 719 15565 887
rect 15477 703 15565 719
rect 15971 2033 16059 2049
rect 15971 1265 15987 2033
rect 16021 1265 16059 2033
rect 15971 1249 16059 1265
rect 16459 2033 16547 2049
rect 16459 1265 16497 2033
rect 16531 1265 16547 2033
rect 16459 1249 16547 1265
rect 16589 2033 16677 2049
rect 16589 1265 16605 2033
rect 16639 1265 16677 2033
rect 16589 1249 16677 1265
rect 17077 2033 17165 2049
rect 17077 1265 17115 2033
rect 17149 1265 17165 2033
rect 17077 1249 17165 1265
rect 15971 887 16059 903
rect 15971 719 15987 887
rect 16021 719 16059 887
rect 15971 703 16059 719
rect 16459 887 16547 903
rect 16459 719 16497 887
rect 16531 719 16547 887
rect 16459 703 16547 719
rect 16589 887 16677 903
rect 16589 719 16605 887
rect 16639 719 16677 887
rect 16589 703 16677 719
rect 17077 887 17165 903
rect 17077 719 17115 887
rect 17149 719 17165 887
rect 17077 703 17165 719
rect 17571 2033 17659 2049
rect 17571 1265 17587 2033
rect 17621 1265 17659 2033
rect 17571 1249 17659 1265
rect 18059 2033 18147 2049
rect 18059 1265 18097 2033
rect 18131 1265 18147 2033
rect 18059 1249 18147 1265
rect 18189 2033 18277 2049
rect 18189 1265 18205 2033
rect 18239 1265 18277 2033
rect 18189 1249 18277 1265
rect 18677 2033 18765 2049
rect 18677 1265 18715 2033
rect 18749 1265 18765 2033
rect 18677 1249 18765 1265
rect 17571 887 17659 903
rect 17571 719 17587 887
rect 17621 719 17659 887
rect 17571 703 17659 719
rect 18059 887 18147 903
rect 18059 719 18097 887
rect 18131 719 18147 887
rect 18059 703 18147 719
rect 18189 887 18277 903
rect 18189 719 18205 887
rect 18239 719 18277 887
rect 18189 703 18277 719
rect 18677 887 18765 903
rect 18677 719 18715 887
rect 18749 719 18765 887
rect 18677 703 18765 719
rect 19171 2033 19259 2049
rect 19171 1265 19187 2033
rect 19221 1265 19259 2033
rect 19171 1249 19259 1265
rect 19659 2033 19747 2049
rect 19659 1265 19697 2033
rect 19731 1265 19747 2033
rect 19659 1249 19747 1265
rect 19789 2033 19877 2049
rect 19789 1265 19805 2033
rect 19839 1265 19877 2033
rect 19789 1249 19877 1265
rect 20277 2033 20365 2049
rect 20277 1265 20315 2033
rect 20349 1265 20365 2033
rect 20277 1249 20365 1265
rect 19171 887 19259 903
rect 19171 719 19187 887
rect 19221 719 19259 887
rect 19171 703 19259 719
rect 19659 887 19747 903
rect 19659 719 19697 887
rect 19731 719 19747 887
rect 19659 703 19747 719
rect 19789 887 19877 903
rect 19789 719 19805 887
rect 19839 719 19877 887
rect 19789 703 19877 719
rect 20277 887 20365 903
rect 20277 719 20315 887
rect 20349 719 20365 887
rect 20277 703 20365 719
rect 20771 2033 20859 2049
rect 20771 1265 20787 2033
rect 20821 1265 20859 2033
rect 20771 1249 20859 1265
rect 21259 2033 21347 2049
rect 21259 1265 21297 2033
rect 21331 1265 21347 2033
rect 21259 1249 21347 1265
rect 21389 2033 21477 2049
rect 21389 1265 21405 2033
rect 21439 1265 21477 2033
rect 21389 1249 21477 1265
rect 21877 2033 21965 2049
rect 21877 1265 21915 2033
rect 21949 1265 21965 2033
rect 21877 1249 21965 1265
rect 20771 887 20859 903
rect 20771 719 20787 887
rect 20821 719 20859 887
rect 20771 703 20859 719
rect 21259 887 21347 903
rect 21259 719 21297 887
rect 21331 719 21347 887
rect 21259 703 21347 719
rect 21389 887 21477 903
rect 21389 719 21405 887
rect 21439 719 21477 887
rect 21389 703 21477 719
rect 21877 887 21965 903
rect 21877 719 21915 887
rect 21949 719 21965 887
rect 21877 703 21965 719
rect 22371 2033 22459 2049
rect 22371 1265 22387 2033
rect 22421 1265 22459 2033
rect 22371 1249 22459 1265
rect 22859 2033 22947 2049
rect 22859 1265 22897 2033
rect 22931 1265 22947 2033
rect 22859 1249 22947 1265
rect 22989 2033 23077 2049
rect 22989 1265 23005 2033
rect 23039 1265 23077 2033
rect 22989 1249 23077 1265
rect 23477 2033 23565 2049
rect 23477 1265 23515 2033
rect 23549 1265 23565 2033
rect 23477 1249 23565 1265
rect 22371 887 22459 903
rect 22371 719 22387 887
rect 22421 719 22459 887
rect 22371 703 22459 719
rect 22859 887 22947 903
rect 22859 719 22897 887
rect 22931 719 22947 887
rect 22859 703 22947 719
rect 22989 887 23077 903
rect 22989 719 23005 887
rect 23039 719 23077 887
rect 22989 703 23077 719
rect 23477 887 23565 903
rect 23477 719 23515 887
rect 23549 719 23565 887
rect 23477 703 23565 719
rect 23971 2033 24059 2049
rect 23971 1265 23987 2033
rect 24021 1265 24059 2033
rect 23971 1249 24059 1265
rect 24459 2033 24547 2049
rect 24459 1265 24497 2033
rect 24531 1265 24547 2033
rect 24459 1249 24547 1265
rect 24589 2033 24677 2049
rect 24589 1265 24605 2033
rect 24639 1265 24677 2033
rect 24589 1249 24677 1265
rect 25077 2033 25165 2049
rect 25077 1265 25115 2033
rect 25149 1265 25165 2033
rect 25077 1249 25165 1265
rect 23971 887 24059 903
rect 23971 719 23987 887
rect 24021 719 24059 887
rect 23971 703 24059 719
rect 24459 887 24547 903
rect 24459 719 24497 887
rect 24531 719 24547 887
rect 24459 703 24547 719
rect 24589 887 24677 903
rect 24589 719 24605 887
rect 24639 719 24677 887
rect 24589 703 24677 719
rect 25077 887 25165 903
rect 25077 719 25115 887
rect 25149 719 25165 887
rect 25077 703 25165 719
rect 25571 2033 25659 2049
rect 25571 1265 25587 2033
rect 25621 1265 25659 2033
rect 25571 1249 25659 1265
rect 26059 2033 26147 2049
rect 26059 1265 26097 2033
rect 26131 1265 26147 2033
rect 26059 1249 26147 1265
rect 26189 2033 26277 2049
rect 26189 1265 26205 2033
rect 26239 1265 26277 2033
rect 26189 1249 26277 1265
rect 26677 2033 26765 2049
rect 26677 1265 26715 2033
rect 26749 1265 26765 2033
rect 26677 1249 26765 1265
rect 25571 887 25659 903
rect 25571 719 25587 887
rect 25621 719 25659 887
rect 25571 703 25659 719
rect 26059 887 26147 903
rect 26059 719 26097 887
rect 26131 719 26147 887
rect 26059 703 26147 719
rect 26189 887 26277 903
rect 26189 719 26205 887
rect 26239 719 26277 887
rect 26189 703 26277 719
rect 26677 887 26765 903
rect 26677 719 26715 887
rect 26749 719 26765 887
rect 26677 703 26765 719
rect 27171 2033 27259 2049
rect 27171 1265 27187 2033
rect 27221 1265 27259 2033
rect 27171 1249 27259 1265
rect 27659 2033 27747 2049
rect 27659 1265 27697 2033
rect 27731 1265 27747 2033
rect 27659 1249 27747 1265
rect 27789 2033 27877 2049
rect 27789 1265 27805 2033
rect 27839 1265 27877 2033
rect 27789 1249 27877 1265
rect 28277 2033 28365 2049
rect 28277 1265 28315 2033
rect 28349 1265 28365 2033
rect 28277 1249 28365 1265
rect 27171 887 27259 903
rect 27171 719 27187 887
rect 27221 719 27259 887
rect 27171 703 27259 719
rect 27659 887 27747 903
rect 27659 719 27697 887
rect 27731 719 27747 887
rect 27659 703 27747 719
rect 27789 887 27877 903
rect 27789 719 27805 887
rect 27839 719 27877 887
rect 27789 703 27877 719
rect 28277 887 28365 903
rect 28277 719 28315 887
rect 28349 719 28365 887
rect 28277 703 28365 719
rect 28771 2033 28859 2049
rect 28771 1265 28787 2033
rect 28821 1265 28859 2033
rect 28771 1249 28859 1265
rect 29259 2033 29347 2049
rect 29259 1265 29297 2033
rect 29331 1265 29347 2033
rect 29259 1249 29347 1265
rect 29389 2033 29477 2049
rect 29389 1265 29405 2033
rect 29439 1265 29477 2033
rect 29389 1249 29477 1265
rect 29877 2033 29965 2049
rect 29877 1265 29915 2033
rect 29949 1265 29965 2033
rect 29877 1249 29965 1265
rect 28771 887 28859 903
rect 28771 719 28787 887
rect 28821 719 28859 887
rect 28771 703 28859 719
rect 29259 887 29347 903
rect 29259 719 29297 887
rect 29331 719 29347 887
rect 29259 703 29347 719
rect 29389 887 29477 903
rect 29389 719 29405 887
rect 29439 719 29477 887
rect 29389 703 29477 719
rect 29877 887 29965 903
rect 29877 719 29915 887
rect 29949 719 29965 887
rect 29877 703 29965 719
rect 30371 2033 30459 2049
rect 30371 1265 30387 2033
rect 30421 1265 30459 2033
rect 30371 1249 30459 1265
rect 30859 2033 30947 2049
rect 30859 1265 30897 2033
rect 30931 1265 30947 2033
rect 30859 1249 30947 1265
rect 30989 2033 31077 2049
rect 30989 1265 31005 2033
rect 31039 1265 31077 2033
rect 30989 1249 31077 1265
rect 31477 2033 31565 2049
rect 31477 1265 31515 2033
rect 31549 1265 31565 2033
rect 31477 1249 31565 1265
rect 30371 887 30459 903
rect 30371 719 30387 887
rect 30421 719 30459 887
rect 30371 703 30459 719
rect 30859 887 30947 903
rect 30859 719 30897 887
rect 30931 719 30947 887
rect 30859 703 30947 719
rect 30989 887 31077 903
rect 30989 719 31005 887
rect 31039 719 31077 887
rect 30989 703 31077 719
rect 31477 887 31565 903
rect 31477 719 31515 887
rect 31549 719 31565 887
rect 31477 703 31565 719
rect 31971 2033 32059 2049
rect 31971 1265 31987 2033
rect 32021 1265 32059 2033
rect 31971 1249 32059 1265
rect 32459 2033 32547 2049
rect 32459 1265 32497 2033
rect 32531 1265 32547 2033
rect 32459 1249 32547 1265
rect 32589 2033 32677 2049
rect 32589 1265 32605 2033
rect 32639 1265 32677 2033
rect 32589 1249 32677 1265
rect 33077 2033 33165 2049
rect 33077 1265 33115 2033
rect 33149 1265 33165 2033
rect 33077 1249 33165 1265
rect 31971 887 32059 903
rect 31971 719 31987 887
rect 32021 719 32059 887
rect 31971 703 32059 719
rect 32459 887 32547 903
rect 32459 719 32497 887
rect 32531 719 32547 887
rect 32459 703 32547 719
rect 32589 887 32677 903
rect 32589 719 32605 887
rect 32639 719 32677 887
rect 32589 703 32677 719
rect 33077 887 33165 903
rect 33077 719 33115 887
rect 33149 719 33165 887
rect 33077 703 33165 719
rect 33571 2033 33659 2049
rect 33571 1265 33587 2033
rect 33621 1265 33659 2033
rect 33571 1249 33659 1265
rect 34059 2033 34147 2049
rect 34059 1265 34097 2033
rect 34131 1265 34147 2033
rect 34059 1249 34147 1265
rect 34189 2033 34277 2049
rect 34189 1265 34205 2033
rect 34239 1265 34277 2033
rect 34189 1249 34277 1265
rect 34677 2033 34765 2049
rect 34677 1265 34715 2033
rect 34749 1265 34765 2033
rect 34677 1249 34765 1265
rect 33571 887 33659 903
rect 33571 719 33587 887
rect 33621 719 33659 887
rect 33571 703 33659 719
rect 34059 887 34147 903
rect 34059 719 34097 887
rect 34131 719 34147 887
rect 34059 703 34147 719
rect 34189 887 34277 903
rect 34189 719 34205 887
rect 34239 719 34277 887
rect 34189 703 34277 719
rect 34677 887 34765 903
rect 34677 719 34715 887
rect 34749 719 34765 887
rect 34677 703 34765 719
rect 35171 2033 35259 2049
rect 35171 1265 35187 2033
rect 35221 1265 35259 2033
rect 35171 1249 35259 1265
rect 35659 2033 35747 2049
rect 35659 1265 35697 2033
rect 35731 1265 35747 2033
rect 35659 1249 35747 1265
rect 35789 2033 35877 2049
rect 35789 1265 35805 2033
rect 35839 1265 35877 2033
rect 35789 1249 35877 1265
rect 36277 2033 36365 2049
rect 36277 1265 36315 2033
rect 36349 1265 36365 2033
rect 36277 1249 36365 1265
rect 35171 887 35259 903
rect 35171 719 35187 887
rect 35221 719 35259 887
rect 35171 703 35259 719
rect 35659 887 35747 903
rect 35659 719 35697 887
rect 35731 719 35747 887
rect 35659 703 35747 719
rect 35789 887 35877 903
rect 35789 719 35805 887
rect 35839 719 35877 887
rect 35789 703 35877 719
rect 36277 887 36365 903
rect 36277 719 36315 887
rect 36349 719 36365 887
rect 36277 703 36365 719
rect 36771 2033 36859 2049
rect 36771 1265 36787 2033
rect 36821 1265 36859 2033
rect 36771 1249 36859 1265
rect 37259 2033 37347 2049
rect 37259 1265 37297 2033
rect 37331 1265 37347 2033
rect 37259 1249 37347 1265
rect 37389 2033 37477 2049
rect 37389 1265 37405 2033
rect 37439 1265 37477 2033
rect 37389 1249 37477 1265
rect 37877 2033 37965 2049
rect 37877 1265 37915 2033
rect 37949 1265 37965 2033
rect 37877 1249 37965 1265
rect 36771 887 36859 903
rect 36771 719 36787 887
rect 36821 719 36859 887
rect 36771 703 36859 719
rect 37259 887 37347 903
rect 37259 719 37297 887
rect 37331 719 37347 887
rect 37259 703 37347 719
rect 37389 887 37477 903
rect 37389 719 37405 887
rect 37439 719 37477 887
rect 37389 703 37477 719
rect 37877 887 37965 903
rect 37877 719 37915 887
rect 37949 719 37965 887
rect 37877 703 37965 719
rect -29 233 59 249
rect -29 -535 -13 233
rect 21 -535 59 233
rect -29 -551 59 -535
rect 459 233 547 249
rect 459 -535 497 233
rect 531 -535 547 233
rect 459 -551 547 -535
rect 589 233 677 249
rect 589 -535 605 233
rect 639 -535 677 233
rect 589 -551 677 -535
rect 1077 233 1165 249
rect 1077 -535 1115 233
rect 1149 -535 1165 233
rect 1077 -551 1165 -535
rect -29 -913 59 -897
rect -29 -1081 -13 -913
rect 21 -1081 59 -913
rect -29 -1097 59 -1081
rect 459 -913 547 -897
rect 459 -1081 497 -913
rect 531 -1081 547 -913
rect 459 -1097 547 -1081
rect 589 -913 677 -897
rect 589 -1081 605 -913
rect 639 -1081 677 -913
rect 589 -1097 677 -1081
rect 1077 -913 1165 -897
rect 1077 -1081 1115 -913
rect 1149 -1081 1165 -913
rect 1077 -1097 1165 -1081
rect 1571 233 1659 249
rect 1571 -535 1587 233
rect 1621 -535 1659 233
rect 1571 -551 1659 -535
rect 2059 233 2147 249
rect 2059 -535 2097 233
rect 2131 -535 2147 233
rect 2059 -551 2147 -535
rect 2189 233 2277 249
rect 2189 -535 2205 233
rect 2239 -535 2277 233
rect 2189 -551 2277 -535
rect 2677 233 2765 249
rect 2677 -535 2715 233
rect 2749 -535 2765 233
rect 2677 -551 2765 -535
rect 1571 -913 1659 -897
rect 1571 -1081 1587 -913
rect 1621 -1081 1659 -913
rect 1571 -1097 1659 -1081
rect 2059 -913 2147 -897
rect 2059 -1081 2097 -913
rect 2131 -1081 2147 -913
rect 2059 -1097 2147 -1081
rect 2189 -913 2277 -897
rect 2189 -1081 2205 -913
rect 2239 -1081 2277 -913
rect 2189 -1097 2277 -1081
rect 2677 -913 2765 -897
rect 2677 -1081 2715 -913
rect 2749 -1081 2765 -913
rect 2677 -1097 2765 -1081
rect 3171 233 3259 249
rect 3171 -535 3187 233
rect 3221 -535 3259 233
rect 3171 -551 3259 -535
rect 3659 233 3747 249
rect 3659 -535 3697 233
rect 3731 -535 3747 233
rect 3659 -551 3747 -535
rect 3789 233 3877 249
rect 3789 -535 3805 233
rect 3839 -535 3877 233
rect 3789 -551 3877 -535
rect 4277 233 4365 249
rect 4277 -535 4315 233
rect 4349 -535 4365 233
rect 4277 -551 4365 -535
rect 3171 -913 3259 -897
rect 3171 -1081 3187 -913
rect 3221 -1081 3259 -913
rect 3171 -1097 3259 -1081
rect 3659 -913 3747 -897
rect 3659 -1081 3697 -913
rect 3731 -1081 3747 -913
rect 3659 -1097 3747 -1081
rect 3789 -913 3877 -897
rect 3789 -1081 3805 -913
rect 3839 -1081 3877 -913
rect 3789 -1097 3877 -1081
rect 4277 -913 4365 -897
rect 4277 -1081 4315 -913
rect 4349 -1081 4365 -913
rect 4277 -1097 4365 -1081
rect 4771 233 4859 249
rect 4771 -535 4787 233
rect 4821 -535 4859 233
rect 4771 -551 4859 -535
rect 5259 233 5347 249
rect 5259 -535 5297 233
rect 5331 -535 5347 233
rect 5259 -551 5347 -535
rect 5389 233 5477 249
rect 5389 -535 5405 233
rect 5439 -535 5477 233
rect 5389 -551 5477 -535
rect 5877 233 5965 249
rect 5877 -535 5915 233
rect 5949 -535 5965 233
rect 5877 -551 5965 -535
rect 4771 -913 4859 -897
rect 4771 -1081 4787 -913
rect 4821 -1081 4859 -913
rect 4771 -1097 4859 -1081
rect 5259 -913 5347 -897
rect 5259 -1081 5297 -913
rect 5331 -1081 5347 -913
rect 5259 -1097 5347 -1081
rect 5389 -913 5477 -897
rect 5389 -1081 5405 -913
rect 5439 -1081 5477 -913
rect 5389 -1097 5477 -1081
rect 5877 -913 5965 -897
rect 5877 -1081 5915 -913
rect 5949 -1081 5965 -913
rect 5877 -1097 5965 -1081
rect 6371 233 6459 249
rect 6371 -535 6387 233
rect 6421 -535 6459 233
rect 6371 -551 6459 -535
rect 6859 233 6947 249
rect 6859 -535 6897 233
rect 6931 -535 6947 233
rect 6859 -551 6947 -535
rect 6989 233 7077 249
rect 6989 -535 7005 233
rect 7039 -535 7077 233
rect 6989 -551 7077 -535
rect 7477 233 7565 249
rect 7477 -535 7515 233
rect 7549 -535 7565 233
rect 7477 -551 7565 -535
rect 6371 -913 6459 -897
rect 6371 -1081 6387 -913
rect 6421 -1081 6459 -913
rect 6371 -1097 6459 -1081
rect 6859 -913 6947 -897
rect 6859 -1081 6897 -913
rect 6931 -1081 6947 -913
rect 6859 -1097 6947 -1081
rect 6989 -913 7077 -897
rect 6989 -1081 7005 -913
rect 7039 -1081 7077 -913
rect 6989 -1097 7077 -1081
rect 7477 -913 7565 -897
rect 7477 -1081 7515 -913
rect 7549 -1081 7565 -913
rect 7477 -1097 7565 -1081
rect 7971 233 8059 249
rect 7971 -535 7987 233
rect 8021 -535 8059 233
rect 7971 -551 8059 -535
rect 8459 233 8547 249
rect 8459 -535 8497 233
rect 8531 -535 8547 233
rect 8459 -551 8547 -535
rect 8589 233 8677 249
rect 8589 -535 8605 233
rect 8639 -535 8677 233
rect 8589 -551 8677 -535
rect 9077 233 9165 249
rect 9077 -535 9115 233
rect 9149 -535 9165 233
rect 9077 -551 9165 -535
rect 7971 -913 8059 -897
rect 7971 -1081 7987 -913
rect 8021 -1081 8059 -913
rect 7971 -1097 8059 -1081
rect 8459 -913 8547 -897
rect 8459 -1081 8497 -913
rect 8531 -1081 8547 -913
rect 8459 -1097 8547 -1081
rect 8589 -913 8677 -897
rect 8589 -1081 8605 -913
rect 8639 -1081 8677 -913
rect 8589 -1097 8677 -1081
rect 9077 -913 9165 -897
rect 9077 -1081 9115 -913
rect 9149 -1081 9165 -913
rect 9077 -1097 9165 -1081
rect 9571 233 9659 249
rect 9571 -535 9587 233
rect 9621 -535 9659 233
rect 9571 -551 9659 -535
rect 10059 233 10147 249
rect 10059 -535 10097 233
rect 10131 -535 10147 233
rect 10059 -551 10147 -535
rect 10189 233 10277 249
rect 10189 -535 10205 233
rect 10239 -535 10277 233
rect 10189 -551 10277 -535
rect 10677 233 10765 249
rect 10677 -535 10715 233
rect 10749 -535 10765 233
rect 10677 -551 10765 -535
rect 9571 -913 9659 -897
rect 9571 -1081 9587 -913
rect 9621 -1081 9659 -913
rect 9571 -1097 9659 -1081
rect 10059 -913 10147 -897
rect 10059 -1081 10097 -913
rect 10131 -1081 10147 -913
rect 10059 -1097 10147 -1081
rect 10189 -913 10277 -897
rect 10189 -1081 10205 -913
rect 10239 -1081 10277 -913
rect 10189 -1097 10277 -1081
rect 10677 -913 10765 -897
rect 10677 -1081 10715 -913
rect 10749 -1081 10765 -913
rect 10677 -1097 10765 -1081
rect 11171 233 11259 249
rect 11171 -535 11187 233
rect 11221 -535 11259 233
rect 11171 -551 11259 -535
rect 11659 233 11747 249
rect 11659 -535 11697 233
rect 11731 -535 11747 233
rect 11659 -551 11747 -535
rect 11789 233 11877 249
rect 11789 -535 11805 233
rect 11839 -535 11877 233
rect 11789 -551 11877 -535
rect 12277 233 12365 249
rect 12277 -535 12315 233
rect 12349 -535 12365 233
rect 12277 -551 12365 -535
rect 11171 -913 11259 -897
rect 11171 -1081 11187 -913
rect 11221 -1081 11259 -913
rect 11171 -1097 11259 -1081
rect 11659 -913 11747 -897
rect 11659 -1081 11697 -913
rect 11731 -1081 11747 -913
rect 11659 -1097 11747 -1081
rect 11789 -913 11877 -897
rect 11789 -1081 11805 -913
rect 11839 -1081 11877 -913
rect 11789 -1097 11877 -1081
rect 12277 -913 12365 -897
rect 12277 -1081 12315 -913
rect 12349 -1081 12365 -913
rect 12277 -1097 12365 -1081
rect 12771 233 12859 249
rect 12771 -535 12787 233
rect 12821 -535 12859 233
rect 12771 -551 12859 -535
rect 13259 233 13347 249
rect 13259 -535 13297 233
rect 13331 -535 13347 233
rect 13259 -551 13347 -535
rect 13389 233 13477 249
rect 13389 -535 13405 233
rect 13439 -535 13477 233
rect 13389 -551 13477 -535
rect 13877 233 13965 249
rect 13877 -535 13915 233
rect 13949 -535 13965 233
rect 13877 -551 13965 -535
rect 12771 -913 12859 -897
rect 12771 -1081 12787 -913
rect 12821 -1081 12859 -913
rect 12771 -1097 12859 -1081
rect 13259 -913 13347 -897
rect 13259 -1081 13297 -913
rect 13331 -1081 13347 -913
rect 13259 -1097 13347 -1081
rect 13389 -913 13477 -897
rect 13389 -1081 13405 -913
rect 13439 -1081 13477 -913
rect 13389 -1097 13477 -1081
rect 13877 -913 13965 -897
rect 13877 -1081 13915 -913
rect 13949 -1081 13965 -913
rect 13877 -1097 13965 -1081
rect 14371 233 14459 249
rect 14371 -535 14387 233
rect 14421 -535 14459 233
rect 14371 -551 14459 -535
rect 14859 233 14947 249
rect 14859 -535 14897 233
rect 14931 -535 14947 233
rect 14859 -551 14947 -535
rect 14989 233 15077 249
rect 14989 -535 15005 233
rect 15039 -535 15077 233
rect 14989 -551 15077 -535
rect 15477 233 15565 249
rect 15477 -535 15515 233
rect 15549 -535 15565 233
rect 15477 -551 15565 -535
rect 14371 -913 14459 -897
rect 14371 -1081 14387 -913
rect 14421 -1081 14459 -913
rect 14371 -1097 14459 -1081
rect 14859 -913 14947 -897
rect 14859 -1081 14897 -913
rect 14931 -1081 14947 -913
rect 14859 -1097 14947 -1081
rect 14989 -913 15077 -897
rect 14989 -1081 15005 -913
rect 15039 -1081 15077 -913
rect 14989 -1097 15077 -1081
rect 15477 -913 15565 -897
rect 15477 -1081 15515 -913
rect 15549 -1081 15565 -913
rect 15477 -1097 15565 -1081
rect 15971 233 16059 249
rect 15971 -535 15987 233
rect 16021 -535 16059 233
rect 15971 -551 16059 -535
rect 16459 233 16547 249
rect 16459 -535 16497 233
rect 16531 -535 16547 233
rect 16459 -551 16547 -535
rect 16589 233 16677 249
rect 16589 -535 16605 233
rect 16639 -535 16677 233
rect 16589 -551 16677 -535
rect 17077 233 17165 249
rect 17077 -535 17115 233
rect 17149 -535 17165 233
rect 17077 -551 17165 -535
rect 15971 -913 16059 -897
rect 15971 -1081 15987 -913
rect 16021 -1081 16059 -913
rect 15971 -1097 16059 -1081
rect 16459 -913 16547 -897
rect 16459 -1081 16497 -913
rect 16531 -1081 16547 -913
rect 16459 -1097 16547 -1081
rect 16589 -913 16677 -897
rect 16589 -1081 16605 -913
rect 16639 -1081 16677 -913
rect 16589 -1097 16677 -1081
rect 17077 -913 17165 -897
rect 17077 -1081 17115 -913
rect 17149 -1081 17165 -913
rect 17077 -1097 17165 -1081
rect 17571 233 17659 249
rect 17571 -535 17587 233
rect 17621 -535 17659 233
rect 17571 -551 17659 -535
rect 18059 233 18147 249
rect 18059 -535 18097 233
rect 18131 -535 18147 233
rect 18059 -551 18147 -535
rect 18189 233 18277 249
rect 18189 -535 18205 233
rect 18239 -535 18277 233
rect 18189 -551 18277 -535
rect 18677 233 18765 249
rect 18677 -535 18715 233
rect 18749 -535 18765 233
rect 18677 -551 18765 -535
rect 17571 -913 17659 -897
rect 17571 -1081 17587 -913
rect 17621 -1081 17659 -913
rect 17571 -1097 17659 -1081
rect 18059 -913 18147 -897
rect 18059 -1081 18097 -913
rect 18131 -1081 18147 -913
rect 18059 -1097 18147 -1081
rect 18189 -913 18277 -897
rect 18189 -1081 18205 -913
rect 18239 -1081 18277 -913
rect 18189 -1097 18277 -1081
rect 18677 -913 18765 -897
rect 18677 -1081 18715 -913
rect 18749 -1081 18765 -913
rect 18677 -1097 18765 -1081
rect 19171 233 19259 249
rect 19171 -535 19187 233
rect 19221 -535 19259 233
rect 19171 -551 19259 -535
rect 19659 233 19747 249
rect 19659 -535 19697 233
rect 19731 -535 19747 233
rect 19659 -551 19747 -535
rect 19789 233 19877 249
rect 19789 -535 19805 233
rect 19839 -535 19877 233
rect 19789 -551 19877 -535
rect 20277 233 20365 249
rect 20277 -535 20315 233
rect 20349 -535 20365 233
rect 20277 -551 20365 -535
rect 19171 -913 19259 -897
rect 19171 -1081 19187 -913
rect 19221 -1081 19259 -913
rect 19171 -1097 19259 -1081
rect 19659 -913 19747 -897
rect 19659 -1081 19697 -913
rect 19731 -1081 19747 -913
rect 19659 -1097 19747 -1081
rect 19789 -913 19877 -897
rect 19789 -1081 19805 -913
rect 19839 -1081 19877 -913
rect 19789 -1097 19877 -1081
rect 20277 -913 20365 -897
rect 20277 -1081 20315 -913
rect 20349 -1081 20365 -913
rect 20277 -1097 20365 -1081
rect 20771 233 20859 249
rect 20771 -535 20787 233
rect 20821 -535 20859 233
rect 20771 -551 20859 -535
rect 21259 233 21347 249
rect 21259 -535 21297 233
rect 21331 -535 21347 233
rect 21259 -551 21347 -535
rect 21389 233 21477 249
rect 21389 -535 21405 233
rect 21439 -535 21477 233
rect 21389 -551 21477 -535
rect 21877 233 21965 249
rect 21877 -535 21915 233
rect 21949 -535 21965 233
rect 21877 -551 21965 -535
rect 20771 -913 20859 -897
rect 20771 -1081 20787 -913
rect 20821 -1081 20859 -913
rect 20771 -1097 20859 -1081
rect 21259 -913 21347 -897
rect 21259 -1081 21297 -913
rect 21331 -1081 21347 -913
rect 21259 -1097 21347 -1081
rect 21389 -913 21477 -897
rect 21389 -1081 21405 -913
rect 21439 -1081 21477 -913
rect 21389 -1097 21477 -1081
rect 21877 -913 21965 -897
rect 21877 -1081 21915 -913
rect 21949 -1081 21965 -913
rect 21877 -1097 21965 -1081
rect 22371 233 22459 249
rect 22371 -535 22387 233
rect 22421 -535 22459 233
rect 22371 -551 22459 -535
rect 22859 233 22947 249
rect 22859 -535 22897 233
rect 22931 -535 22947 233
rect 22859 -551 22947 -535
rect 22989 233 23077 249
rect 22989 -535 23005 233
rect 23039 -535 23077 233
rect 22989 -551 23077 -535
rect 23477 233 23565 249
rect 23477 -535 23515 233
rect 23549 -535 23565 233
rect 23477 -551 23565 -535
rect 22371 -913 22459 -897
rect 22371 -1081 22387 -913
rect 22421 -1081 22459 -913
rect 22371 -1097 22459 -1081
rect 22859 -913 22947 -897
rect 22859 -1081 22897 -913
rect 22931 -1081 22947 -913
rect 22859 -1097 22947 -1081
rect 22989 -913 23077 -897
rect 22989 -1081 23005 -913
rect 23039 -1081 23077 -913
rect 22989 -1097 23077 -1081
rect 23477 -913 23565 -897
rect 23477 -1081 23515 -913
rect 23549 -1081 23565 -913
rect 23477 -1097 23565 -1081
rect 23971 233 24059 249
rect 23971 -535 23987 233
rect 24021 -535 24059 233
rect 23971 -551 24059 -535
rect 24459 233 24547 249
rect 24459 -535 24497 233
rect 24531 -535 24547 233
rect 24459 -551 24547 -535
rect 24589 233 24677 249
rect 24589 -535 24605 233
rect 24639 -535 24677 233
rect 24589 -551 24677 -535
rect 25077 233 25165 249
rect 25077 -535 25115 233
rect 25149 -535 25165 233
rect 25077 -551 25165 -535
rect 23971 -913 24059 -897
rect 23971 -1081 23987 -913
rect 24021 -1081 24059 -913
rect 23971 -1097 24059 -1081
rect 24459 -913 24547 -897
rect 24459 -1081 24497 -913
rect 24531 -1081 24547 -913
rect 24459 -1097 24547 -1081
rect 24589 -913 24677 -897
rect 24589 -1081 24605 -913
rect 24639 -1081 24677 -913
rect 24589 -1097 24677 -1081
rect 25077 -913 25165 -897
rect 25077 -1081 25115 -913
rect 25149 -1081 25165 -913
rect 25077 -1097 25165 -1081
rect 25571 233 25659 249
rect 25571 -535 25587 233
rect 25621 -535 25659 233
rect 25571 -551 25659 -535
rect 26059 233 26147 249
rect 26059 -535 26097 233
rect 26131 -535 26147 233
rect 26059 -551 26147 -535
rect 26189 233 26277 249
rect 26189 -535 26205 233
rect 26239 -535 26277 233
rect 26189 -551 26277 -535
rect 26677 233 26765 249
rect 26677 -535 26715 233
rect 26749 -535 26765 233
rect 26677 -551 26765 -535
rect 25571 -913 25659 -897
rect 25571 -1081 25587 -913
rect 25621 -1081 25659 -913
rect 25571 -1097 25659 -1081
rect 26059 -913 26147 -897
rect 26059 -1081 26097 -913
rect 26131 -1081 26147 -913
rect 26059 -1097 26147 -1081
rect 26189 -913 26277 -897
rect 26189 -1081 26205 -913
rect 26239 -1081 26277 -913
rect 26189 -1097 26277 -1081
rect 26677 -913 26765 -897
rect 26677 -1081 26715 -913
rect 26749 -1081 26765 -913
rect 26677 -1097 26765 -1081
rect 27171 233 27259 249
rect 27171 -535 27187 233
rect 27221 -535 27259 233
rect 27171 -551 27259 -535
rect 27659 233 27747 249
rect 27659 -535 27697 233
rect 27731 -535 27747 233
rect 27659 -551 27747 -535
rect 27789 233 27877 249
rect 27789 -535 27805 233
rect 27839 -535 27877 233
rect 27789 -551 27877 -535
rect 28277 233 28365 249
rect 28277 -535 28315 233
rect 28349 -535 28365 233
rect 28277 -551 28365 -535
rect 27171 -913 27259 -897
rect 27171 -1081 27187 -913
rect 27221 -1081 27259 -913
rect 27171 -1097 27259 -1081
rect 27659 -913 27747 -897
rect 27659 -1081 27697 -913
rect 27731 -1081 27747 -913
rect 27659 -1097 27747 -1081
rect 27789 -913 27877 -897
rect 27789 -1081 27805 -913
rect 27839 -1081 27877 -913
rect 27789 -1097 27877 -1081
rect 28277 -913 28365 -897
rect 28277 -1081 28315 -913
rect 28349 -1081 28365 -913
rect 28277 -1097 28365 -1081
rect 28771 233 28859 249
rect 28771 -535 28787 233
rect 28821 -535 28859 233
rect 28771 -551 28859 -535
rect 29259 233 29347 249
rect 29259 -535 29297 233
rect 29331 -535 29347 233
rect 29259 -551 29347 -535
rect 29389 233 29477 249
rect 29389 -535 29405 233
rect 29439 -535 29477 233
rect 29389 -551 29477 -535
rect 29877 233 29965 249
rect 29877 -535 29915 233
rect 29949 -535 29965 233
rect 29877 -551 29965 -535
rect 28771 -913 28859 -897
rect 28771 -1081 28787 -913
rect 28821 -1081 28859 -913
rect 28771 -1097 28859 -1081
rect 29259 -913 29347 -897
rect 29259 -1081 29297 -913
rect 29331 -1081 29347 -913
rect 29259 -1097 29347 -1081
rect 29389 -913 29477 -897
rect 29389 -1081 29405 -913
rect 29439 -1081 29477 -913
rect 29389 -1097 29477 -1081
rect 29877 -913 29965 -897
rect 29877 -1081 29915 -913
rect 29949 -1081 29965 -913
rect 29877 -1097 29965 -1081
rect 30371 233 30459 249
rect 30371 -535 30387 233
rect 30421 -535 30459 233
rect 30371 -551 30459 -535
rect 30859 233 30947 249
rect 30859 -535 30897 233
rect 30931 -535 30947 233
rect 30859 -551 30947 -535
rect 30989 233 31077 249
rect 30989 -535 31005 233
rect 31039 -535 31077 233
rect 30989 -551 31077 -535
rect 31477 233 31565 249
rect 31477 -535 31515 233
rect 31549 -535 31565 233
rect 31477 -551 31565 -535
rect 30371 -913 30459 -897
rect 30371 -1081 30387 -913
rect 30421 -1081 30459 -913
rect 30371 -1097 30459 -1081
rect 30859 -913 30947 -897
rect 30859 -1081 30897 -913
rect 30931 -1081 30947 -913
rect 30859 -1097 30947 -1081
rect 30989 -913 31077 -897
rect 30989 -1081 31005 -913
rect 31039 -1081 31077 -913
rect 30989 -1097 31077 -1081
rect 31477 -913 31565 -897
rect 31477 -1081 31515 -913
rect 31549 -1081 31565 -913
rect 31477 -1097 31565 -1081
rect 31971 233 32059 249
rect 31971 -535 31987 233
rect 32021 -535 32059 233
rect 31971 -551 32059 -535
rect 32459 233 32547 249
rect 32459 -535 32497 233
rect 32531 -535 32547 233
rect 32459 -551 32547 -535
rect 32589 233 32677 249
rect 32589 -535 32605 233
rect 32639 -535 32677 233
rect 32589 -551 32677 -535
rect 33077 233 33165 249
rect 33077 -535 33115 233
rect 33149 -535 33165 233
rect 33077 -551 33165 -535
rect 31971 -913 32059 -897
rect 31971 -1081 31987 -913
rect 32021 -1081 32059 -913
rect 31971 -1097 32059 -1081
rect 32459 -913 32547 -897
rect 32459 -1081 32497 -913
rect 32531 -1081 32547 -913
rect 32459 -1097 32547 -1081
rect 32589 -913 32677 -897
rect 32589 -1081 32605 -913
rect 32639 -1081 32677 -913
rect 32589 -1097 32677 -1081
rect 33077 -913 33165 -897
rect 33077 -1081 33115 -913
rect 33149 -1081 33165 -913
rect 33077 -1097 33165 -1081
rect 33571 233 33659 249
rect 33571 -535 33587 233
rect 33621 -535 33659 233
rect 33571 -551 33659 -535
rect 34059 233 34147 249
rect 34059 -535 34097 233
rect 34131 -535 34147 233
rect 34059 -551 34147 -535
rect 34189 233 34277 249
rect 34189 -535 34205 233
rect 34239 -535 34277 233
rect 34189 -551 34277 -535
rect 34677 233 34765 249
rect 34677 -535 34715 233
rect 34749 -535 34765 233
rect 34677 -551 34765 -535
rect 33571 -913 33659 -897
rect 33571 -1081 33587 -913
rect 33621 -1081 33659 -913
rect 33571 -1097 33659 -1081
rect 34059 -913 34147 -897
rect 34059 -1081 34097 -913
rect 34131 -1081 34147 -913
rect 34059 -1097 34147 -1081
rect 34189 -913 34277 -897
rect 34189 -1081 34205 -913
rect 34239 -1081 34277 -913
rect 34189 -1097 34277 -1081
rect 34677 -913 34765 -897
rect 34677 -1081 34715 -913
rect 34749 -1081 34765 -913
rect 34677 -1097 34765 -1081
rect 35171 233 35259 249
rect 35171 -535 35187 233
rect 35221 -535 35259 233
rect 35171 -551 35259 -535
rect 35659 233 35747 249
rect 35659 -535 35697 233
rect 35731 -535 35747 233
rect 35659 -551 35747 -535
rect 35789 233 35877 249
rect 35789 -535 35805 233
rect 35839 -535 35877 233
rect 35789 -551 35877 -535
rect 36277 233 36365 249
rect 36277 -535 36315 233
rect 36349 -535 36365 233
rect 36277 -551 36365 -535
rect 35171 -913 35259 -897
rect 35171 -1081 35187 -913
rect 35221 -1081 35259 -913
rect 35171 -1097 35259 -1081
rect 35659 -913 35747 -897
rect 35659 -1081 35697 -913
rect 35731 -1081 35747 -913
rect 35659 -1097 35747 -1081
rect 35789 -913 35877 -897
rect 35789 -1081 35805 -913
rect 35839 -1081 35877 -913
rect 35789 -1097 35877 -1081
rect 36277 -913 36365 -897
rect 36277 -1081 36315 -913
rect 36349 -1081 36365 -913
rect 36277 -1097 36365 -1081
rect 36771 233 36859 249
rect 36771 -535 36787 233
rect 36821 -535 36859 233
rect 36771 -551 36859 -535
rect 37259 233 37347 249
rect 37259 -535 37297 233
rect 37331 -535 37347 233
rect 37259 -551 37347 -535
rect 37389 233 37477 249
rect 37389 -535 37405 233
rect 37439 -535 37477 233
rect 37389 -551 37477 -535
rect 37877 233 37965 249
rect 37877 -535 37915 233
rect 37949 -535 37965 233
rect 37877 -551 37965 -535
rect 36771 -913 36859 -897
rect 36771 -1081 36787 -913
rect 36821 -1081 36859 -913
rect 36771 -1097 36859 -1081
rect 37259 -913 37347 -897
rect 37259 -1081 37297 -913
rect 37331 -1081 37347 -913
rect 37259 -1097 37347 -1081
rect 37389 -913 37477 -897
rect 37389 -1081 37405 -913
rect 37439 -1081 37477 -913
rect 37389 -1097 37477 -1081
rect 37877 -913 37965 -897
rect 37877 -1081 37915 -913
rect 37949 -1081 37965 -913
rect 37877 -1097 37965 -1081
rect -29 -1567 59 -1551
rect -29 -2335 -13 -1567
rect 21 -2335 59 -1567
rect -29 -2351 59 -2335
rect 459 -1567 547 -1551
rect 459 -2335 497 -1567
rect 531 -2335 547 -1567
rect 459 -2351 547 -2335
rect 589 -1567 677 -1551
rect 589 -2335 605 -1567
rect 639 -2335 677 -1567
rect 589 -2351 677 -2335
rect 1077 -1567 1165 -1551
rect 1077 -2335 1115 -1567
rect 1149 -2335 1165 -1567
rect 1077 -2351 1165 -2335
rect -29 -2713 59 -2697
rect -29 -2881 -13 -2713
rect 21 -2881 59 -2713
rect -29 -2897 59 -2881
rect 459 -2713 547 -2697
rect 459 -2881 497 -2713
rect 531 -2881 547 -2713
rect 459 -2897 547 -2881
rect 589 -2713 677 -2697
rect 589 -2881 605 -2713
rect 639 -2881 677 -2713
rect 589 -2897 677 -2881
rect 1077 -2713 1165 -2697
rect 1077 -2881 1115 -2713
rect 1149 -2881 1165 -2713
rect 1077 -2897 1165 -2881
rect 1571 -1567 1659 -1551
rect 1571 -2335 1587 -1567
rect 1621 -2335 1659 -1567
rect 1571 -2351 1659 -2335
rect 2059 -1567 2147 -1551
rect 2059 -2335 2097 -1567
rect 2131 -2335 2147 -1567
rect 2059 -2351 2147 -2335
rect 2189 -1567 2277 -1551
rect 2189 -2335 2205 -1567
rect 2239 -2335 2277 -1567
rect 2189 -2351 2277 -2335
rect 2677 -1567 2765 -1551
rect 2677 -2335 2715 -1567
rect 2749 -2335 2765 -1567
rect 2677 -2351 2765 -2335
rect 1571 -2713 1659 -2697
rect 1571 -2881 1587 -2713
rect 1621 -2881 1659 -2713
rect 1571 -2897 1659 -2881
rect 2059 -2713 2147 -2697
rect 2059 -2881 2097 -2713
rect 2131 -2881 2147 -2713
rect 2059 -2897 2147 -2881
rect 2189 -2713 2277 -2697
rect 2189 -2881 2205 -2713
rect 2239 -2881 2277 -2713
rect 2189 -2897 2277 -2881
rect 2677 -2713 2765 -2697
rect 2677 -2881 2715 -2713
rect 2749 -2881 2765 -2713
rect 2677 -2897 2765 -2881
rect 3171 -1567 3259 -1551
rect 3171 -2335 3187 -1567
rect 3221 -2335 3259 -1567
rect 3171 -2351 3259 -2335
rect 3659 -1567 3747 -1551
rect 3659 -2335 3697 -1567
rect 3731 -2335 3747 -1567
rect 3659 -2351 3747 -2335
rect 3789 -1567 3877 -1551
rect 3789 -2335 3805 -1567
rect 3839 -2335 3877 -1567
rect 3789 -2351 3877 -2335
rect 4277 -1567 4365 -1551
rect 4277 -2335 4315 -1567
rect 4349 -2335 4365 -1567
rect 4277 -2351 4365 -2335
rect 3171 -2713 3259 -2697
rect 3171 -2881 3187 -2713
rect 3221 -2881 3259 -2713
rect 3171 -2897 3259 -2881
rect 3659 -2713 3747 -2697
rect 3659 -2881 3697 -2713
rect 3731 -2881 3747 -2713
rect 3659 -2897 3747 -2881
rect 3789 -2713 3877 -2697
rect 3789 -2881 3805 -2713
rect 3839 -2881 3877 -2713
rect 3789 -2897 3877 -2881
rect 4277 -2713 4365 -2697
rect 4277 -2881 4315 -2713
rect 4349 -2881 4365 -2713
rect 4277 -2897 4365 -2881
rect 4771 -1567 4859 -1551
rect 4771 -2335 4787 -1567
rect 4821 -2335 4859 -1567
rect 4771 -2351 4859 -2335
rect 5259 -1567 5347 -1551
rect 5259 -2335 5297 -1567
rect 5331 -2335 5347 -1567
rect 5259 -2351 5347 -2335
rect 5389 -1567 5477 -1551
rect 5389 -2335 5405 -1567
rect 5439 -2335 5477 -1567
rect 5389 -2351 5477 -2335
rect 5877 -1567 5965 -1551
rect 5877 -2335 5915 -1567
rect 5949 -2335 5965 -1567
rect 5877 -2351 5965 -2335
rect 4771 -2713 4859 -2697
rect 4771 -2881 4787 -2713
rect 4821 -2881 4859 -2713
rect 4771 -2897 4859 -2881
rect 5259 -2713 5347 -2697
rect 5259 -2881 5297 -2713
rect 5331 -2881 5347 -2713
rect 5259 -2897 5347 -2881
rect 5389 -2713 5477 -2697
rect 5389 -2881 5405 -2713
rect 5439 -2881 5477 -2713
rect 5389 -2897 5477 -2881
rect 5877 -2713 5965 -2697
rect 5877 -2881 5915 -2713
rect 5949 -2881 5965 -2713
rect 5877 -2897 5965 -2881
rect 6371 -1567 6459 -1551
rect 6371 -2335 6387 -1567
rect 6421 -2335 6459 -1567
rect 6371 -2351 6459 -2335
rect 6859 -1567 6947 -1551
rect 6859 -2335 6897 -1567
rect 6931 -2335 6947 -1567
rect 6859 -2351 6947 -2335
rect 6989 -1567 7077 -1551
rect 6989 -2335 7005 -1567
rect 7039 -2335 7077 -1567
rect 6989 -2351 7077 -2335
rect 7477 -1567 7565 -1551
rect 7477 -2335 7515 -1567
rect 7549 -2335 7565 -1567
rect 7477 -2351 7565 -2335
rect 6371 -2713 6459 -2697
rect 6371 -2881 6387 -2713
rect 6421 -2881 6459 -2713
rect 6371 -2897 6459 -2881
rect 6859 -2713 6947 -2697
rect 6859 -2881 6897 -2713
rect 6931 -2881 6947 -2713
rect 6859 -2897 6947 -2881
rect 6989 -2713 7077 -2697
rect 6989 -2881 7005 -2713
rect 7039 -2881 7077 -2713
rect 6989 -2897 7077 -2881
rect 7477 -2713 7565 -2697
rect 7477 -2881 7515 -2713
rect 7549 -2881 7565 -2713
rect 7477 -2897 7565 -2881
rect 7971 -1567 8059 -1551
rect 7971 -2335 7987 -1567
rect 8021 -2335 8059 -1567
rect 7971 -2351 8059 -2335
rect 8459 -1567 8547 -1551
rect 8459 -2335 8497 -1567
rect 8531 -2335 8547 -1567
rect 8459 -2351 8547 -2335
rect 8589 -1567 8677 -1551
rect 8589 -2335 8605 -1567
rect 8639 -2335 8677 -1567
rect 8589 -2351 8677 -2335
rect 9077 -1567 9165 -1551
rect 9077 -2335 9115 -1567
rect 9149 -2335 9165 -1567
rect 9077 -2351 9165 -2335
rect 7971 -2713 8059 -2697
rect 7971 -2881 7987 -2713
rect 8021 -2881 8059 -2713
rect 7971 -2897 8059 -2881
rect 8459 -2713 8547 -2697
rect 8459 -2881 8497 -2713
rect 8531 -2881 8547 -2713
rect 8459 -2897 8547 -2881
rect 8589 -2713 8677 -2697
rect 8589 -2881 8605 -2713
rect 8639 -2881 8677 -2713
rect 8589 -2897 8677 -2881
rect 9077 -2713 9165 -2697
rect 9077 -2881 9115 -2713
rect 9149 -2881 9165 -2713
rect 9077 -2897 9165 -2881
rect 9571 -1567 9659 -1551
rect 9571 -2335 9587 -1567
rect 9621 -2335 9659 -1567
rect 9571 -2351 9659 -2335
rect 10059 -1567 10147 -1551
rect 10059 -2335 10097 -1567
rect 10131 -2335 10147 -1567
rect 10059 -2351 10147 -2335
rect 10189 -1567 10277 -1551
rect 10189 -2335 10205 -1567
rect 10239 -2335 10277 -1567
rect 10189 -2351 10277 -2335
rect 10677 -1567 10765 -1551
rect 10677 -2335 10715 -1567
rect 10749 -2335 10765 -1567
rect 10677 -2351 10765 -2335
rect 9571 -2713 9659 -2697
rect 9571 -2881 9587 -2713
rect 9621 -2881 9659 -2713
rect 9571 -2897 9659 -2881
rect 10059 -2713 10147 -2697
rect 10059 -2881 10097 -2713
rect 10131 -2881 10147 -2713
rect 10059 -2897 10147 -2881
rect 10189 -2713 10277 -2697
rect 10189 -2881 10205 -2713
rect 10239 -2881 10277 -2713
rect 10189 -2897 10277 -2881
rect 10677 -2713 10765 -2697
rect 10677 -2881 10715 -2713
rect 10749 -2881 10765 -2713
rect 10677 -2897 10765 -2881
rect 11171 -1567 11259 -1551
rect 11171 -2335 11187 -1567
rect 11221 -2335 11259 -1567
rect 11171 -2351 11259 -2335
rect 11659 -1567 11747 -1551
rect 11659 -2335 11697 -1567
rect 11731 -2335 11747 -1567
rect 11659 -2351 11747 -2335
rect 11789 -1567 11877 -1551
rect 11789 -2335 11805 -1567
rect 11839 -2335 11877 -1567
rect 11789 -2351 11877 -2335
rect 12277 -1567 12365 -1551
rect 12277 -2335 12315 -1567
rect 12349 -2335 12365 -1567
rect 12277 -2351 12365 -2335
rect 11171 -2713 11259 -2697
rect 11171 -2881 11187 -2713
rect 11221 -2881 11259 -2713
rect 11171 -2897 11259 -2881
rect 11659 -2713 11747 -2697
rect 11659 -2881 11697 -2713
rect 11731 -2881 11747 -2713
rect 11659 -2897 11747 -2881
rect 11789 -2713 11877 -2697
rect 11789 -2881 11805 -2713
rect 11839 -2881 11877 -2713
rect 11789 -2897 11877 -2881
rect 12277 -2713 12365 -2697
rect 12277 -2881 12315 -2713
rect 12349 -2881 12365 -2713
rect 12277 -2897 12365 -2881
rect 12771 -1567 12859 -1551
rect 12771 -2335 12787 -1567
rect 12821 -2335 12859 -1567
rect 12771 -2351 12859 -2335
rect 13259 -1567 13347 -1551
rect 13259 -2335 13297 -1567
rect 13331 -2335 13347 -1567
rect 13259 -2351 13347 -2335
rect 13389 -1567 13477 -1551
rect 13389 -2335 13405 -1567
rect 13439 -2335 13477 -1567
rect 13389 -2351 13477 -2335
rect 13877 -1567 13965 -1551
rect 13877 -2335 13915 -1567
rect 13949 -2335 13965 -1567
rect 13877 -2351 13965 -2335
rect 12771 -2713 12859 -2697
rect 12771 -2881 12787 -2713
rect 12821 -2881 12859 -2713
rect 12771 -2897 12859 -2881
rect 13259 -2713 13347 -2697
rect 13259 -2881 13297 -2713
rect 13331 -2881 13347 -2713
rect 13259 -2897 13347 -2881
rect 13389 -2713 13477 -2697
rect 13389 -2881 13405 -2713
rect 13439 -2881 13477 -2713
rect 13389 -2897 13477 -2881
rect 13877 -2713 13965 -2697
rect 13877 -2881 13915 -2713
rect 13949 -2881 13965 -2713
rect 13877 -2897 13965 -2881
rect 14371 -1567 14459 -1551
rect 14371 -2335 14387 -1567
rect 14421 -2335 14459 -1567
rect 14371 -2351 14459 -2335
rect 14859 -1567 14947 -1551
rect 14859 -2335 14897 -1567
rect 14931 -2335 14947 -1567
rect 14859 -2351 14947 -2335
rect 14989 -1567 15077 -1551
rect 14989 -2335 15005 -1567
rect 15039 -2335 15077 -1567
rect 14989 -2351 15077 -2335
rect 15477 -1567 15565 -1551
rect 15477 -2335 15515 -1567
rect 15549 -2335 15565 -1567
rect 15477 -2351 15565 -2335
rect 14371 -2713 14459 -2697
rect 14371 -2881 14387 -2713
rect 14421 -2881 14459 -2713
rect 14371 -2897 14459 -2881
rect 14859 -2713 14947 -2697
rect 14859 -2881 14897 -2713
rect 14931 -2881 14947 -2713
rect 14859 -2897 14947 -2881
rect 14989 -2713 15077 -2697
rect 14989 -2881 15005 -2713
rect 15039 -2881 15077 -2713
rect 14989 -2897 15077 -2881
rect 15477 -2713 15565 -2697
rect 15477 -2881 15515 -2713
rect 15549 -2881 15565 -2713
rect 15477 -2897 15565 -2881
rect 15971 -1567 16059 -1551
rect 15971 -2335 15987 -1567
rect 16021 -2335 16059 -1567
rect 15971 -2351 16059 -2335
rect 16459 -1567 16547 -1551
rect 16459 -2335 16497 -1567
rect 16531 -2335 16547 -1567
rect 16459 -2351 16547 -2335
rect 16589 -1567 16677 -1551
rect 16589 -2335 16605 -1567
rect 16639 -2335 16677 -1567
rect 16589 -2351 16677 -2335
rect 17077 -1567 17165 -1551
rect 17077 -2335 17115 -1567
rect 17149 -2335 17165 -1567
rect 17077 -2351 17165 -2335
rect 15971 -2713 16059 -2697
rect 15971 -2881 15987 -2713
rect 16021 -2881 16059 -2713
rect 15971 -2897 16059 -2881
rect 16459 -2713 16547 -2697
rect 16459 -2881 16497 -2713
rect 16531 -2881 16547 -2713
rect 16459 -2897 16547 -2881
rect 16589 -2713 16677 -2697
rect 16589 -2881 16605 -2713
rect 16639 -2881 16677 -2713
rect 16589 -2897 16677 -2881
rect 17077 -2713 17165 -2697
rect 17077 -2881 17115 -2713
rect 17149 -2881 17165 -2713
rect 17077 -2897 17165 -2881
rect 17571 -1567 17659 -1551
rect 17571 -2335 17587 -1567
rect 17621 -2335 17659 -1567
rect 17571 -2351 17659 -2335
rect 18059 -1567 18147 -1551
rect 18059 -2335 18097 -1567
rect 18131 -2335 18147 -1567
rect 18059 -2351 18147 -2335
rect 18189 -1567 18277 -1551
rect 18189 -2335 18205 -1567
rect 18239 -2335 18277 -1567
rect 18189 -2351 18277 -2335
rect 18677 -1567 18765 -1551
rect 18677 -2335 18715 -1567
rect 18749 -2335 18765 -1567
rect 18677 -2351 18765 -2335
rect 17571 -2713 17659 -2697
rect 17571 -2881 17587 -2713
rect 17621 -2881 17659 -2713
rect 17571 -2897 17659 -2881
rect 18059 -2713 18147 -2697
rect 18059 -2881 18097 -2713
rect 18131 -2881 18147 -2713
rect 18059 -2897 18147 -2881
rect 18189 -2713 18277 -2697
rect 18189 -2881 18205 -2713
rect 18239 -2881 18277 -2713
rect 18189 -2897 18277 -2881
rect 18677 -2713 18765 -2697
rect 18677 -2881 18715 -2713
rect 18749 -2881 18765 -2713
rect 18677 -2897 18765 -2881
rect 19171 -1567 19259 -1551
rect 19171 -2335 19187 -1567
rect 19221 -2335 19259 -1567
rect 19171 -2351 19259 -2335
rect 19659 -1567 19747 -1551
rect 19659 -2335 19697 -1567
rect 19731 -2335 19747 -1567
rect 19659 -2351 19747 -2335
rect 19789 -1567 19877 -1551
rect 19789 -2335 19805 -1567
rect 19839 -2335 19877 -1567
rect 19789 -2351 19877 -2335
rect 20277 -1567 20365 -1551
rect 20277 -2335 20315 -1567
rect 20349 -2335 20365 -1567
rect 20277 -2351 20365 -2335
rect 19171 -2713 19259 -2697
rect 19171 -2881 19187 -2713
rect 19221 -2881 19259 -2713
rect 19171 -2897 19259 -2881
rect 19659 -2713 19747 -2697
rect 19659 -2881 19697 -2713
rect 19731 -2881 19747 -2713
rect 19659 -2897 19747 -2881
rect 19789 -2713 19877 -2697
rect 19789 -2881 19805 -2713
rect 19839 -2881 19877 -2713
rect 19789 -2897 19877 -2881
rect 20277 -2713 20365 -2697
rect 20277 -2881 20315 -2713
rect 20349 -2881 20365 -2713
rect 20277 -2897 20365 -2881
rect 20771 -1567 20859 -1551
rect 20771 -2335 20787 -1567
rect 20821 -2335 20859 -1567
rect 20771 -2351 20859 -2335
rect 21259 -1567 21347 -1551
rect 21259 -2335 21297 -1567
rect 21331 -2335 21347 -1567
rect 21259 -2351 21347 -2335
rect 21389 -1567 21477 -1551
rect 21389 -2335 21405 -1567
rect 21439 -2335 21477 -1567
rect 21389 -2351 21477 -2335
rect 21877 -1567 21965 -1551
rect 21877 -2335 21915 -1567
rect 21949 -2335 21965 -1567
rect 21877 -2351 21965 -2335
rect 20771 -2713 20859 -2697
rect 20771 -2881 20787 -2713
rect 20821 -2881 20859 -2713
rect 20771 -2897 20859 -2881
rect 21259 -2713 21347 -2697
rect 21259 -2881 21297 -2713
rect 21331 -2881 21347 -2713
rect 21259 -2897 21347 -2881
rect 21389 -2713 21477 -2697
rect 21389 -2881 21405 -2713
rect 21439 -2881 21477 -2713
rect 21389 -2897 21477 -2881
rect 21877 -2713 21965 -2697
rect 21877 -2881 21915 -2713
rect 21949 -2881 21965 -2713
rect 21877 -2897 21965 -2881
rect 22371 -1567 22459 -1551
rect 22371 -2335 22387 -1567
rect 22421 -2335 22459 -1567
rect 22371 -2351 22459 -2335
rect 22859 -1567 22947 -1551
rect 22859 -2335 22897 -1567
rect 22931 -2335 22947 -1567
rect 22859 -2351 22947 -2335
rect 22989 -1567 23077 -1551
rect 22989 -2335 23005 -1567
rect 23039 -2335 23077 -1567
rect 22989 -2351 23077 -2335
rect 23477 -1567 23565 -1551
rect 23477 -2335 23515 -1567
rect 23549 -2335 23565 -1567
rect 23477 -2351 23565 -2335
rect 22371 -2713 22459 -2697
rect 22371 -2881 22387 -2713
rect 22421 -2881 22459 -2713
rect 22371 -2897 22459 -2881
rect 22859 -2713 22947 -2697
rect 22859 -2881 22897 -2713
rect 22931 -2881 22947 -2713
rect 22859 -2897 22947 -2881
rect 22989 -2713 23077 -2697
rect 22989 -2881 23005 -2713
rect 23039 -2881 23077 -2713
rect 22989 -2897 23077 -2881
rect 23477 -2713 23565 -2697
rect 23477 -2881 23515 -2713
rect 23549 -2881 23565 -2713
rect 23477 -2897 23565 -2881
rect 23971 -1567 24059 -1551
rect 23971 -2335 23987 -1567
rect 24021 -2335 24059 -1567
rect 23971 -2351 24059 -2335
rect 24459 -1567 24547 -1551
rect 24459 -2335 24497 -1567
rect 24531 -2335 24547 -1567
rect 24459 -2351 24547 -2335
rect 24589 -1567 24677 -1551
rect 24589 -2335 24605 -1567
rect 24639 -2335 24677 -1567
rect 24589 -2351 24677 -2335
rect 25077 -1567 25165 -1551
rect 25077 -2335 25115 -1567
rect 25149 -2335 25165 -1567
rect 25077 -2351 25165 -2335
rect 23971 -2713 24059 -2697
rect 23971 -2881 23987 -2713
rect 24021 -2881 24059 -2713
rect 23971 -2897 24059 -2881
rect 24459 -2713 24547 -2697
rect 24459 -2881 24497 -2713
rect 24531 -2881 24547 -2713
rect 24459 -2897 24547 -2881
rect 24589 -2713 24677 -2697
rect 24589 -2881 24605 -2713
rect 24639 -2881 24677 -2713
rect 24589 -2897 24677 -2881
rect 25077 -2713 25165 -2697
rect 25077 -2881 25115 -2713
rect 25149 -2881 25165 -2713
rect 25077 -2897 25165 -2881
rect 25571 -1567 25659 -1551
rect 25571 -2335 25587 -1567
rect 25621 -2335 25659 -1567
rect 25571 -2351 25659 -2335
rect 26059 -1567 26147 -1551
rect 26059 -2335 26097 -1567
rect 26131 -2335 26147 -1567
rect 26059 -2351 26147 -2335
rect 26189 -1567 26277 -1551
rect 26189 -2335 26205 -1567
rect 26239 -2335 26277 -1567
rect 26189 -2351 26277 -2335
rect 26677 -1567 26765 -1551
rect 26677 -2335 26715 -1567
rect 26749 -2335 26765 -1567
rect 26677 -2351 26765 -2335
rect 25571 -2713 25659 -2697
rect 25571 -2881 25587 -2713
rect 25621 -2881 25659 -2713
rect 25571 -2897 25659 -2881
rect 26059 -2713 26147 -2697
rect 26059 -2881 26097 -2713
rect 26131 -2881 26147 -2713
rect 26059 -2897 26147 -2881
rect 26189 -2713 26277 -2697
rect 26189 -2881 26205 -2713
rect 26239 -2881 26277 -2713
rect 26189 -2897 26277 -2881
rect 26677 -2713 26765 -2697
rect 26677 -2881 26715 -2713
rect 26749 -2881 26765 -2713
rect 26677 -2897 26765 -2881
rect 27171 -1567 27259 -1551
rect 27171 -2335 27187 -1567
rect 27221 -2335 27259 -1567
rect 27171 -2351 27259 -2335
rect 27659 -1567 27747 -1551
rect 27659 -2335 27697 -1567
rect 27731 -2335 27747 -1567
rect 27659 -2351 27747 -2335
rect 27789 -1567 27877 -1551
rect 27789 -2335 27805 -1567
rect 27839 -2335 27877 -1567
rect 27789 -2351 27877 -2335
rect 28277 -1567 28365 -1551
rect 28277 -2335 28315 -1567
rect 28349 -2335 28365 -1567
rect 28277 -2351 28365 -2335
rect 27171 -2713 27259 -2697
rect 27171 -2881 27187 -2713
rect 27221 -2881 27259 -2713
rect 27171 -2897 27259 -2881
rect 27659 -2713 27747 -2697
rect 27659 -2881 27697 -2713
rect 27731 -2881 27747 -2713
rect 27659 -2897 27747 -2881
rect 27789 -2713 27877 -2697
rect 27789 -2881 27805 -2713
rect 27839 -2881 27877 -2713
rect 27789 -2897 27877 -2881
rect 28277 -2713 28365 -2697
rect 28277 -2881 28315 -2713
rect 28349 -2881 28365 -2713
rect 28277 -2897 28365 -2881
rect 28771 -1567 28859 -1551
rect 28771 -2335 28787 -1567
rect 28821 -2335 28859 -1567
rect 28771 -2351 28859 -2335
rect 29259 -1567 29347 -1551
rect 29259 -2335 29297 -1567
rect 29331 -2335 29347 -1567
rect 29259 -2351 29347 -2335
rect 29389 -1567 29477 -1551
rect 29389 -2335 29405 -1567
rect 29439 -2335 29477 -1567
rect 29389 -2351 29477 -2335
rect 29877 -1567 29965 -1551
rect 29877 -2335 29915 -1567
rect 29949 -2335 29965 -1567
rect 29877 -2351 29965 -2335
rect 28771 -2713 28859 -2697
rect 28771 -2881 28787 -2713
rect 28821 -2881 28859 -2713
rect 28771 -2897 28859 -2881
rect 29259 -2713 29347 -2697
rect 29259 -2881 29297 -2713
rect 29331 -2881 29347 -2713
rect 29259 -2897 29347 -2881
rect 29389 -2713 29477 -2697
rect 29389 -2881 29405 -2713
rect 29439 -2881 29477 -2713
rect 29389 -2897 29477 -2881
rect 29877 -2713 29965 -2697
rect 29877 -2881 29915 -2713
rect 29949 -2881 29965 -2713
rect 29877 -2897 29965 -2881
rect 30371 -1567 30459 -1551
rect 30371 -2335 30387 -1567
rect 30421 -2335 30459 -1567
rect 30371 -2351 30459 -2335
rect 30859 -1567 30947 -1551
rect 30859 -2335 30897 -1567
rect 30931 -2335 30947 -1567
rect 30859 -2351 30947 -2335
rect 30989 -1567 31077 -1551
rect 30989 -2335 31005 -1567
rect 31039 -2335 31077 -1567
rect 30989 -2351 31077 -2335
rect 31477 -1567 31565 -1551
rect 31477 -2335 31515 -1567
rect 31549 -2335 31565 -1567
rect 31477 -2351 31565 -2335
rect 30371 -2713 30459 -2697
rect 30371 -2881 30387 -2713
rect 30421 -2881 30459 -2713
rect 30371 -2897 30459 -2881
rect 30859 -2713 30947 -2697
rect 30859 -2881 30897 -2713
rect 30931 -2881 30947 -2713
rect 30859 -2897 30947 -2881
rect 30989 -2713 31077 -2697
rect 30989 -2881 31005 -2713
rect 31039 -2881 31077 -2713
rect 30989 -2897 31077 -2881
rect 31477 -2713 31565 -2697
rect 31477 -2881 31515 -2713
rect 31549 -2881 31565 -2713
rect 31477 -2897 31565 -2881
rect 31971 -1567 32059 -1551
rect 31971 -2335 31987 -1567
rect 32021 -2335 32059 -1567
rect 31971 -2351 32059 -2335
rect 32459 -1567 32547 -1551
rect 32459 -2335 32497 -1567
rect 32531 -2335 32547 -1567
rect 32459 -2351 32547 -2335
rect 32589 -1567 32677 -1551
rect 32589 -2335 32605 -1567
rect 32639 -2335 32677 -1567
rect 32589 -2351 32677 -2335
rect 33077 -1567 33165 -1551
rect 33077 -2335 33115 -1567
rect 33149 -2335 33165 -1567
rect 33077 -2351 33165 -2335
rect 31971 -2713 32059 -2697
rect 31971 -2881 31987 -2713
rect 32021 -2881 32059 -2713
rect 31971 -2897 32059 -2881
rect 32459 -2713 32547 -2697
rect 32459 -2881 32497 -2713
rect 32531 -2881 32547 -2713
rect 32459 -2897 32547 -2881
rect 32589 -2713 32677 -2697
rect 32589 -2881 32605 -2713
rect 32639 -2881 32677 -2713
rect 32589 -2897 32677 -2881
rect 33077 -2713 33165 -2697
rect 33077 -2881 33115 -2713
rect 33149 -2881 33165 -2713
rect 33077 -2897 33165 -2881
rect 33571 -1567 33659 -1551
rect 33571 -2335 33587 -1567
rect 33621 -2335 33659 -1567
rect 33571 -2351 33659 -2335
rect 34059 -1567 34147 -1551
rect 34059 -2335 34097 -1567
rect 34131 -2335 34147 -1567
rect 34059 -2351 34147 -2335
rect 34189 -1567 34277 -1551
rect 34189 -2335 34205 -1567
rect 34239 -2335 34277 -1567
rect 34189 -2351 34277 -2335
rect 34677 -1567 34765 -1551
rect 34677 -2335 34715 -1567
rect 34749 -2335 34765 -1567
rect 34677 -2351 34765 -2335
rect 33571 -2713 33659 -2697
rect 33571 -2881 33587 -2713
rect 33621 -2881 33659 -2713
rect 33571 -2897 33659 -2881
rect 34059 -2713 34147 -2697
rect 34059 -2881 34097 -2713
rect 34131 -2881 34147 -2713
rect 34059 -2897 34147 -2881
rect 34189 -2713 34277 -2697
rect 34189 -2881 34205 -2713
rect 34239 -2881 34277 -2713
rect 34189 -2897 34277 -2881
rect 34677 -2713 34765 -2697
rect 34677 -2881 34715 -2713
rect 34749 -2881 34765 -2713
rect 34677 -2897 34765 -2881
rect 35171 -1567 35259 -1551
rect 35171 -2335 35187 -1567
rect 35221 -2335 35259 -1567
rect 35171 -2351 35259 -2335
rect 35659 -1567 35747 -1551
rect 35659 -2335 35697 -1567
rect 35731 -2335 35747 -1567
rect 35659 -2351 35747 -2335
rect 35789 -1567 35877 -1551
rect 35789 -2335 35805 -1567
rect 35839 -2335 35877 -1567
rect 35789 -2351 35877 -2335
rect 36277 -1567 36365 -1551
rect 36277 -2335 36315 -1567
rect 36349 -2335 36365 -1567
rect 36277 -2351 36365 -2335
rect 35171 -2713 35259 -2697
rect 35171 -2881 35187 -2713
rect 35221 -2881 35259 -2713
rect 35171 -2897 35259 -2881
rect 35659 -2713 35747 -2697
rect 35659 -2881 35697 -2713
rect 35731 -2881 35747 -2713
rect 35659 -2897 35747 -2881
rect 35789 -2713 35877 -2697
rect 35789 -2881 35805 -2713
rect 35839 -2881 35877 -2713
rect 35789 -2897 35877 -2881
rect 36277 -2713 36365 -2697
rect 36277 -2881 36315 -2713
rect 36349 -2881 36365 -2713
rect 36277 -2897 36365 -2881
rect 36771 -1567 36859 -1551
rect 36771 -2335 36787 -1567
rect 36821 -2335 36859 -1567
rect 36771 -2351 36859 -2335
rect 37259 -1567 37347 -1551
rect 37259 -2335 37297 -1567
rect 37331 -2335 37347 -1567
rect 37259 -2351 37347 -2335
rect 37389 -1567 37477 -1551
rect 37389 -2335 37405 -1567
rect 37439 -2335 37477 -1567
rect 37389 -2351 37477 -2335
rect 37877 -1567 37965 -1551
rect 37877 -2335 37915 -1567
rect 37949 -2335 37965 -1567
rect 37877 -2351 37965 -2335
rect 36771 -2713 36859 -2697
rect 36771 -2881 36787 -2713
rect 36821 -2881 36859 -2713
rect 36771 -2897 36859 -2881
rect 37259 -2713 37347 -2697
rect 37259 -2881 37297 -2713
rect 37331 -2881 37347 -2713
rect 37259 -2897 37347 -2881
rect 37389 -2713 37477 -2697
rect 37389 -2881 37405 -2713
rect 37439 -2881 37477 -2713
rect 37389 -2897 37477 -2881
rect 37877 -2713 37965 -2697
rect 37877 -2881 37915 -2713
rect 37949 -2881 37965 -2713
rect 37877 -2897 37965 -2881
rect -29 -3367 59 -3351
rect -29 -4135 -13 -3367
rect 21 -4135 59 -3367
rect -29 -4151 59 -4135
rect 459 -3367 547 -3351
rect 459 -4135 497 -3367
rect 531 -4135 547 -3367
rect 459 -4151 547 -4135
rect 589 -3367 677 -3351
rect 589 -4135 605 -3367
rect 639 -4135 677 -3367
rect 589 -4151 677 -4135
rect 1077 -3367 1165 -3351
rect 1077 -4135 1115 -3367
rect 1149 -4135 1165 -3367
rect 1077 -4151 1165 -4135
rect -29 -4513 59 -4497
rect -29 -4681 -13 -4513
rect 21 -4681 59 -4513
rect -29 -4697 59 -4681
rect 459 -4513 547 -4497
rect 459 -4681 497 -4513
rect 531 -4681 547 -4513
rect 459 -4697 547 -4681
rect 589 -4513 677 -4497
rect 589 -4681 605 -4513
rect 639 -4681 677 -4513
rect 589 -4697 677 -4681
rect 1077 -4513 1165 -4497
rect 1077 -4681 1115 -4513
rect 1149 -4681 1165 -4513
rect 1077 -4697 1165 -4681
rect 1571 -3367 1659 -3351
rect 1571 -4135 1587 -3367
rect 1621 -4135 1659 -3367
rect 1571 -4151 1659 -4135
rect 2059 -3367 2147 -3351
rect 2059 -4135 2097 -3367
rect 2131 -4135 2147 -3367
rect 2059 -4151 2147 -4135
rect 2189 -3367 2277 -3351
rect 2189 -4135 2205 -3367
rect 2239 -4135 2277 -3367
rect 2189 -4151 2277 -4135
rect 2677 -3367 2765 -3351
rect 2677 -4135 2715 -3367
rect 2749 -4135 2765 -3367
rect 2677 -4151 2765 -4135
rect 1571 -4513 1659 -4497
rect 1571 -4681 1587 -4513
rect 1621 -4681 1659 -4513
rect 1571 -4697 1659 -4681
rect 2059 -4513 2147 -4497
rect 2059 -4681 2097 -4513
rect 2131 -4681 2147 -4513
rect 2059 -4697 2147 -4681
rect 2189 -4513 2277 -4497
rect 2189 -4681 2205 -4513
rect 2239 -4681 2277 -4513
rect 2189 -4697 2277 -4681
rect 2677 -4513 2765 -4497
rect 2677 -4681 2715 -4513
rect 2749 -4681 2765 -4513
rect 2677 -4697 2765 -4681
rect 3171 -3367 3259 -3351
rect 3171 -4135 3187 -3367
rect 3221 -4135 3259 -3367
rect 3171 -4151 3259 -4135
rect 3659 -3367 3747 -3351
rect 3659 -4135 3697 -3367
rect 3731 -4135 3747 -3367
rect 3659 -4151 3747 -4135
rect 3789 -3367 3877 -3351
rect 3789 -4135 3805 -3367
rect 3839 -4135 3877 -3367
rect 3789 -4151 3877 -4135
rect 4277 -3367 4365 -3351
rect 4277 -4135 4315 -3367
rect 4349 -4135 4365 -3367
rect 4277 -4151 4365 -4135
rect 3171 -4513 3259 -4497
rect 3171 -4681 3187 -4513
rect 3221 -4681 3259 -4513
rect 3171 -4697 3259 -4681
rect 3659 -4513 3747 -4497
rect 3659 -4681 3697 -4513
rect 3731 -4681 3747 -4513
rect 3659 -4697 3747 -4681
rect 3789 -4513 3877 -4497
rect 3789 -4681 3805 -4513
rect 3839 -4681 3877 -4513
rect 3789 -4697 3877 -4681
rect 4277 -4513 4365 -4497
rect 4277 -4681 4315 -4513
rect 4349 -4681 4365 -4513
rect 4277 -4697 4365 -4681
rect 4771 -3367 4859 -3351
rect 4771 -4135 4787 -3367
rect 4821 -4135 4859 -3367
rect 4771 -4151 4859 -4135
rect 5259 -3367 5347 -3351
rect 5259 -4135 5297 -3367
rect 5331 -4135 5347 -3367
rect 5259 -4151 5347 -4135
rect 5389 -3367 5477 -3351
rect 5389 -4135 5405 -3367
rect 5439 -4135 5477 -3367
rect 5389 -4151 5477 -4135
rect 5877 -3367 5965 -3351
rect 5877 -4135 5915 -3367
rect 5949 -4135 5965 -3367
rect 5877 -4151 5965 -4135
rect 4771 -4513 4859 -4497
rect 4771 -4681 4787 -4513
rect 4821 -4681 4859 -4513
rect 4771 -4697 4859 -4681
rect 5259 -4513 5347 -4497
rect 5259 -4681 5297 -4513
rect 5331 -4681 5347 -4513
rect 5259 -4697 5347 -4681
rect 5389 -4513 5477 -4497
rect 5389 -4681 5405 -4513
rect 5439 -4681 5477 -4513
rect 5389 -4697 5477 -4681
rect 5877 -4513 5965 -4497
rect 5877 -4681 5915 -4513
rect 5949 -4681 5965 -4513
rect 5877 -4697 5965 -4681
rect 6371 -3367 6459 -3351
rect 6371 -4135 6387 -3367
rect 6421 -4135 6459 -3367
rect 6371 -4151 6459 -4135
rect 6859 -3367 6947 -3351
rect 6859 -4135 6897 -3367
rect 6931 -4135 6947 -3367
rect 6859 -4151 6947 -4135
rect 6989 -3367 7077 -3351
rect 6989 -4135 7005 -3367
rect 7039 -4135 7077 -3367
rect 6989 -4151 7077 -4135
rect 7477 -3367 7565 -3351
rect 7477 -4135 7515 -3367
rect 7549 -4135 7565 -3367
rect 7477 -4151 7565 -4135
rect 6371 -4513 6459 -4497
rect 6371 -4681 6387 -4513
rect 6421 -4681 6459 -4513
rect 6371 -4697 6459 -4681
rect 6859 -4513 6947 -4497
rect 6859 -4681 6897 -4513
rect 6931 -4681 6947 -4513
rect 6859 -4697 6947 -4681
rect 6989 -4513 7077 -4497
rect 6989 -4681 7005 -4513
rect 7039 -4681 7077 -4513
rect 6989 -4697 7077 -4681
rect 7477 -4513 7565 -4497
rect 7477 -4681 7515 -4513
rect 7549 -4681 7565 -4513
rect 7477 -4697 7565 -4681
rect 7971 -3367 8059 -3351
rect 7971 -4135 7987 -3367
rect 8021 -4135 8059 -3367
rect 7971 -4151 8059 -4135
rect 8459 -3367 8547 -3351
rect 8459 -4135 8497 -3367
rect 8531 -4135 8547 -3367
rect 8459 -4151 8547 -4135
rect 8589 -3367 8677 -3351
rect 8589 -4135 8605 -3367
rect 8639 -4135 8677 -3367
rect 8589 -4151 8677 -4135
rect 9077 -3367 9165 -3351
rect 9077 -4135 9115 -3367
rect 9149 -4135 9165 -3367
rect 9077 -4151 9165 -4135
rect 7971 -4513 8059 -4497
rect 7971 -4681 7987 -4513
rect 8021 -4681 8059 -4513
rect 7971 -4697 8059 -4681
rect 8459 -4513 8547 -4497
rect 8459 -4681 8497 -4513
rect 8531 -4681 8547 -4513
rect 8459 -4697 8547 -4681
rect 8589 -4513 8677 -4497
rect 8589 -4681 8605 -4513
rect 8639 -4681 8677 -4513
rect 8589 -4697 8677 -4681
rect 9077 -4513 9165 -4497
rect 9077 -4681 9115 -4513
rect 9149 -4681 9165 -4513
rect 9077 -4697 9165 -4681
rect 9571 -3367 9659 -3351
rect 9571 -4135 9587 -3367
rect 9621 -4135 9659 -3367
rect 9571 -4151 9659 -4135
rect 10059 -3367 10147 -3351
rect 10059 -4135 10097 -3367
rect 10131 -4135 10147 -3367
rect 10059 -4151 10147 -4135
rect 10189 -3367 10277 -3351
rect 10189 -4135 10205 -3367
rect 10239 -4135 10277 -3367
rect 10189 -4151 10277 -4135
rect 10677 -3367 10765 -3351
rect 10677 -4135 10715 -3367
rect 10749 -4135 10765 -3367
rect 10677 -4151 10765 -4135
rect 9571 -4513 9659 -4497
rect 9571 -4681 9587 -4513
rect 9621 -4681 9659 -4513
rect 9571 -4697 9659 -4681
rect 10059 -4513 10147 -4497
rect 10059 -4681 10097 -4513
rect 10131 -4681 10147 -4513
rect 10059 -4697 10147 -4681
rect 10189 -4513 10277 -4497
rect 10189 -4681 10205 -4513
rect 10239 -4681 10277 -4513
rect 10189 -4697 10277 -4681
rect 10677 -4513 10765 -4497
rect 10677 -4681 10715 -4513
rect 10749 -4681 10765 -4513
rect 10677 -4697 10765 -4681
rect 11171 -3367 11259 -3351
rect 11171 -4135 11187 -3367
rect 11221 -4135 11259 -3367
rect 11171 -4151 11259 -4135
rect 11659 -3367 11747 -3351
rect 11659 -4135 11697 -3367
rect 11731 -4135 11747 -3367
rect 11659 -4151 11747 -4135
rect 11789 -3367 11877 -3351
rect 11789 -4135 11805 -3367
rect 11839 -4135 11877 -3367
rect 11789 -4151 11877 -4135
rect 12277 -3367 12365 -3351
rect 12277 -4135 12315 -3367
rect 12349 -4135 12365 -3367
rect 12277 -4151 12365 -4135
rect 11171 -4513 11259 -4497
rect 11171 -4681 11187 -4513
rect 11221 -4681 11259 -4513
rect 11171 -4697 11259 -4681
rect 11659 -4513 11747 -4497
rect 11659 -4681 11697 -4513
rect 11731 -4681 11747 -4513
rect 11659 -4697 11747 -4681
rect 11789 -4513 11877 -4497
rect 11789 -4681 11805 -4513
rect 11839 -4681 11877 -4513
rect 11789 -4697 11877 -4681
rect 12277 -4513 12365 -4497
rect 12277 -4681 12315 -4513
rect 12349 -4681 12365 -4513
rect 12277 -4697 12365 -4681
rect 12771 -3367 12859 -3351
rect 12771 -4135 12787 -3367
rect 12821 -4135 12859 -3367
rect 12771 -4151 12859 -4135
rect 13259 -3367 13347 -3351
rect 13259 -4135 13297 -3367
rect 13331 -4135 13347 -3367
rect 13259 -4151 13347 -4135
rect 13389 -3367 13477 -3351
rect 13389 -4135 13405 -3367
rect 13439 -4135 13477 -3367
rect 13389 -4151 13477 -4135
rect 13877 -3367 13965 -3351
rect 13877 -4135 13915 -3367
rect 13949 -4135 13965 -3367
rect 13877 -4151 13965 -4135
rect 12771 -4513 12859 -4497
rect 12771 -4681 12787 -4513
rect 12821 -4681 12859 -4513
rect 12771 -4697 12859 -4681
rect 13259 -4513 13347 -4497
rect 13259 -4681 13297 -4513
rect 13331 -4681 13347 -4513
rect 13259 -4697 13347 -4681
rect 13389 -4513 13477 -4497
rect 13389 -4681 13405 -4513
rect 13439 -4681 13477 -4513
rect 13389 -4697 13477 -4681
rect 13877 -4513 13965 -4497
rect 13877 -4681 13915 -4513
rect 13949 -4681 13965 -4513
rect 13877 -4697 13965 -4681
rect 14371 -3367 14459 -3351
rect 14371 -4135 14387 -3367
rect 14421 -4135 14459 -3367
rect 14371 -4151 14459 -4135
rect 14859 -3367 14947 -3351
rect 14859 -4135 14897 -3367
rect 14931 -4135 14947 -3367
rect 14859 -4151 14947 -4135
rect 14989 -3367 15077 -3351
rect 14989 -4135 15005 -3367
rect 15039 -4135 15077 -3367
rect 14989 -4151 15077 -4135
rect 15477 -3367 15565 -3351
rect 15477 -4135 15515 -3367
rect 15549 -4135 15565 -3367
rect 15477 -4151 15565 -4135
rect 14371 -4513 14459 -4497
rect 14371 -4681 14387 -4513
rect 14421 -4681 14459 -4513
rect 14371 -4697 14459 -4681
rect 14859 -4513 14947 -4497
rect 14859 -4681 14897 -4513
rect 14931 -4681 14947 -4513
rect 14859 -4697 14947 -4681
rect 14989 -4513 15077 -4497
rect 14989 -4681 15005 -4513
rect 15039 -4681 15077 -4513
rect 14989 -4697 15077 -4681
rect 15477 -4513 15565 -4497
rect 15477 -4681 15515 -4513
rect 15549 -4681 15565 -4513
rect 15477 -4697 15565 -4681
rect 15971 -3367 16059 -3351
rect 15971 -4135 15987 -3367
rect 16021 -4135 16059 -3367
rect 15971 -4151 16059 -4135
rect 16459 -3367 16547 -3351
rect 16459 -4135 16497 -3367
rect 16531 -4135 16547 -3367
rect 16459 -4151 16547 -4135
rect 16589 -3367 16677 -3351
rect 16589 -4135 16605 -3367
rect 16639 -4135 16677 -3367
rect 16589 -4151 16677 -4135
rect 17077 -3367 17165 -3351
rect 17077 -4135 17115 -3367
rect 17149 -4135 17165 -3367
rect 17077 -4151 17165 -4135
rect 15971 -4513 16059 -4497
rect 15971 -4681 15987 -4513
rect 16021 -4681 16059 -4513
rect 15971 -4697 16059 -4681
rect 16459 -4513 16547 -4497
rect 16459 -4681 16497 -4513
rect 16531 -4681 16547 -4513
rect 16459 -4697 16547 -4681
rect 16589 -4513 16677 -4497
rect 16589 -4681 16605 -4513
rect 16639 -4681 16677 -4513
rect 16589 -4697 16677 -4681
rect 17077 -4513 17165 -4497
rect 17077 -4681 17115 -4513
rect 17149 -4681 17165 -4513
rect 17077 -4697 17165 -4681
rect 17571 -3367 17659 -3351
rect 17571 -4135 17587 -3367
rect 17621 -4135 17659 -3367
rect 17571 -4151 17659 -4135
rect 18059 -3367 18147 -3351
rect 18059 -4135 18097 -3367
rect 18131 -4135 18147 -3367
rect 18059 -4151 18147 -4135
rect 18189 -3367 18277 -3351
rect 18189 -4135 18205 -3367
rect 18239 -4135 18277 -3367
rect 18189 -4151 18277 -4135
rect 18677 -3367 18765 -3351
rect 18677 -4135 18715 -3367
rect 18749 -4135 18765 -3367
rect 18677 -4151 18765 -4135
rect 17571 -4513 17659 -4497
rect 17571 -4681 17587 -4513
rect 17621 -4681 17659 -4513
rect 17571 -4697 17659 -4681
rect 18059 -4513 18147 -4497
rect 18059 -4681 18097 -4513
rect 18131 -4681 18147 -4513
rect 18059 -4697 18147 -4681
rect 18189 -4513 18277 -4497
rect 18189 -4681 18205 -4513
rect 18239 -4681 18277 -4513
rect 18189 -4697 18277 -4681
rect 18677 -4513 18765 -4497
rect 18677 -4681 18715 -4513
rect 18749 -4681 18765 -4513
rect 18677 -4697 18765 -4681
rect 19171 -3367 19259 -3351
rect 19171 -4135 19187 -3367
rect 19221 -4135 19259 -3367
rect 19171 -4151 19259 -4135
rect 19659 -3367 19747 -3351
rect 19659 -4135 19697 -3367
rect 19731 -4135 19747 -3367
rect 19659 -4151 19747 -4135
rect 19789 -3367 19877 -3351
rect 19789 -4135 19805 -3367
rect 19839 -4135 19877 -3367
rect 19789 -4151 19877 -4135
rect 20277 -3367 20365 -3351
rect 20277 -4135 20315 -3367
rect 20349 -4135 20365 -3367
rect 20277 -4151 20365 -4135
rect 19171 -4513 19259 -4497
rect 19171 -4681 19187 -4513
rect 19221 -4681 19259 -4513
rect 19171 -4697 19259 -4681
rect 19659 -4513 19747 -4497
rect 19659 -4681 19697 -4513
rect 19731 -4681 19747 -4513
rect 19659 -4697 19747 -4681
rect 19789 -4513 19877 -4497
rect 19789 -4681 19805 -4513
rect 19839 -4681 19877 -4513
rect 19789 -4697 19877 -4681
rect 20277 -4513 20365 -4497
rect 20277 -4681 20315 -4513
rect 20349 -4681 20365 -4513
rect 20277 -4697 20365 -4681
rect 20771 -3367 20859 -3351
rect 20771 -4135 20787 -3367
rect 20821 -4135 20859 -3367
rect 20771 -4151 20859 -4135
rect 21259 -3367 21347 -3351
rect 21259 -4135 21297 -3367
rect 21331 -4135 21347 -3367
rect 21259 -4151 21347 -4135
rect 21389 -3367 21477 -3351
rect 21389 -4135 21405 -3367
rect 21439 -4135 21477 -3367
rect 21389 -4151 21477 -4135
rect 21877 -3367 21965 -3351
rect 21877 -4135 21915 -3367
rect 21949 -4135 21965 -3367
rect 21877 -4151 21965 -4135
rect 20771 -4513 20859 -4497
rect 20771 -4681 20787 -4513
rect 20821 -4681 20859 -4513
rect 20771 -4697 20859 -4681
rect 21259 -4513 21347 -4497
rect 21259 -4681 21297 -4513
rect 21331 -4681 21347 -4513
rect 21259 -4697 21347 -4681
rect 21389 -4513 21477 -4497
rect 21389 -4681 21405 -4513
rect 21439 -4681 21477 -4513
rect 21389 -4697 21477 -4681
rect 21877 -4513 21965 -4497
rect 21877 -4681 21915 -4513
rect 21949 -4681 21965 -4513
rect 21877 -4697 21965 -4681
rect 22371 -3367 22459 -3351
rect 22371 -4135 22387 -3367
rect 22421 -4135 22459 -3367
rect 22371 -4151 22459 -4135
rect 22859 -3367 22947 -3351
rect 22859 -4135 22897 -3367
rect 22931 -4135 22947 -3367
rect 22859 -4151 22947 -4135
rect 22989 -3367 23077 -3351
rect 22989 -4135 23005 -3367
rect 23039 -4135 23077 -3367
rect 22989 -4151 23077 -4135
rect 23477 -3367 23565 -3351
rect 23477 -4135 23515 -3367
rect 23549 -4135 23565 -3367
rect 23477 -4151 23565 -4135
rect 22371 -4513 22459 -4497
rect 22371 -4681 22387 -4513
rect 22421 -4681 22459 -4513
rect 22371 -4697 22459 -4681
rect 22859 -4513 22947 -4497
rect 22859 -4681 22897 -4513
rect 22931 -4681 22947 -4513
rect 22859 -4697 22947 -4681
rect 22989 -4513 23077 -4497
rect 22989 -4681 23005 -4513
rect 23039 -4681 23077 -4513
rect 22989 -4697 23077 -4681
rect 23477 -4513 23565 -4497
rect 23477 -4681 23515 -4513
rect 23549 -4681 23565 -4513
rect 23477 -4697 23565 -4681
rect 23971 -3367 24059 -3351
rect 23971 -4135 23987 -3367
rect 24021 -4135 24059 -3367
rect 23971 -4151 24059 -4135
rect 24459 -3367 24547 -3351
rect 24459 -4135 24497 -3367
rect 24531 -4135 24547 -3367
rect 24459 -4151 24547 -4135
rect 24589 -3367 24677 -3351
rect 24589 -4135 24605 -3367
rect 24639 -4135 24677 -3367
rect 24589 -4151 24677 -4135
rect 25077 -3367 25165 -3351
rect 25077 -4135 25115 -3367
rect 25149 -4135 25165 -3367
rect 25077 -4151 25165 -4135
rect 23971 -4513 24059 -4497
rect 23971 -4681 23987 -4513
rect 24021 -4681 24059 -4513
rect 23971 -4697 24059 -4681
rect 24459 -4513 24547 -4497
rect 24459 -4681 24497 -4513
rect 24531 -4681 24547 -4513
rect 24459 -4697 24547 -4681
rect 24589 -4513 24677 -4497
rect 24589 -4681 24605 -4513
rect 24639 -4681 24677 -4513
rect 24589 -4697 24677 -4681
rect 25077 -4513 25165 -4497
rect 25077 -4681 25115 -4513
rect 25149 -4681 25165 -4513
rect 25077 -4697 25165 -4681
rect 25571 -3367 25659 -3351
rect 25571 -4135 25587 -3367
rect 25621 -4135 25659 -3367
rect 25571 -4151 25659 -4135
rect 26059 -3367 26147 -3351
rect 26059 -4135 26097 -3367
rect 26131 -4135 26147 -3367
rect 26059 -4151 26147 -4135
rect 26189 -3367 26277 -3351
rect 26189 -4135 26205 -3367
rect 26239 -4135 26277 -3367
rect 26189 -4151 26277 -4135
rect 26677 -3367 26765 -3351
rect 26677 -4135 26715 -3367
rect 26749 -4135 26765 -3367
rect 26677 -4151 26765 -4135
rect 25571 -4513 25659 -4497
rect 25571 -4681 25587 -4513
rect 25621 -4681 25659 -4513
rect 25571 -4697 25659 -4681
rect 26059 -4513 26147 -4497
rect 26059 -4681 26097 -4513
rect 26131 -4681 26147 -4513
rect 26059 -4697 26147 -4681
rect 26189 -4513 26277 -4497
rect 26189 -4681 26205 -4513
rect 26239 -4681 26277 -4513
rect 26189 -4697 26277 -4681
rect 26677 -4513 26765 -4497
rect 26677 -4681 26715 -4513
rect 26749 -4681 26765 -4513
rect 26677 -4697 26765 -4681
rect 27171 -3367 27259 -3351
rect 27171 -4135 27187 -3367
rect 27221 -4135 27259 -3367
rect 27171 -4151 27259 -4135
rect 27659 -3367 27747 -3351
rect 27659 -4135 27697 -3367
rect 27731 -4135 27747 -3367
rect 27659 -4151 27747 -4135
rect 27789 -3367 27877 -3351
rect 27789 -4135 27805 -3367
rect 27839 -4135 27877 -3367
rect 27789 -4151 27877 -4135
rect 28277 -3367 28365 -3351
rect 28277 -4135 28315 -3367
rect 28349 -4135 28365 -3367
rect 28277 -4151 28365 -4135
rect 27171 -4513 27259 -4497
rect 27171 -4681 27187 -4513
rect 27221 -4681 27259 -4513
rect 27171 -4697 27259 -4681
rect 27659 -4513 27747 -4497
rect 27659 -4681 27697 -4513
rect 27731 -4681 27747 -4513
rect 27659 -4697 27747 -4681
rect 27789 -4513 27877 -4497
rect 27789 -4681 27805 -4513
rect 27839 -4681 27877 -4513
rect 27789 -4697 27877 -4681
rect 28277 -4513 28365 -4497
rect 28277 -4681 28315 -4513
rect 28349 -4681 28365 -4513
rect 28277 -4697 28365 -4681
rect 28771 -3367 28859 -3351
rect 28771 -4135 28787 -3367
rect 28821 -4135 28859 -3367
rect 28771 -4151 28859 -4135
rect 29259 -3367 29347 -3351
rect 29259 -4135 29297 -3367
rect 29331 -4135 29347 -3367
rect 29259 -4151 29347 -4135
rect 29389 -3367 29477 -3351
rect 29389 -4135 29405 -3367
rect 29439 -4135 29477 -3367
rect 29389 -4151 29477 -4135
rect 29877 -3367 29965 -3351
rect 29877 -4135 29915 -3367
rect 29949 -4135 29965 -3367
rect 29877 -4151 29965 -4135
rect 28771 -4513 28859 -4497
rect 28771 -4681 28787 -4513
rect 28821 -4681 28859 -4513
rect 28771 -4697 28859 -4681
rect 29259 -4513 29347 -4497
rect 29259 -4681 29297 -4513
rect 29331 -4681 29347 -4513
rect 29259 -4697 29347 -4681
rect 29389 -4513 29477 -4497
rect 29389 -4681 29405 -4513
rect 29439 -4681 29477 -4513
rect 29389 -4697 29477 -4681
rect 29877 -4513 29965 -4497
rect 29877 -4681 29915 -4513
rect 29949 -4681 29965 -4513
rect 29877 -4697 29965 -4681
rect 30371 -3367 30459 -3351
rect 30371 -4135 30387 -3367
rect 30421 -4135 30459 -3367
rect 30371 -4151 30459 -4135
rect 30859 -3367 30947 -3351
rect 30859 -4135 30897 -3367
rect 30931 -4135 30947 -3367
rect 30859 -4151 30947 -4135
rect 30989 -3367 31077 -3351
rect 30989 -4135 31005 -3367
rect 31039 -4135 31077 -3367
rect 30989 -4151 31077 -4135
rect 31477 -3367 31565 -3351
rect 31477 -4135 31515 -3367
rect 31549 -4135 31565 -3367
rect 31477 -4151 31565 -4135
rect 30371 -4513 30459 -4497
rect 30371 -4681 30387 -4513
rect 30421 -4681 30459 -4513
rect 30371 -4697 30459 -4681
rect 30859 -4513 30947 -4497
rect 30859 -4681 30897 -4513
rect 30931 -4681 30947 -4513
rect 30859 -4697 30947 -4681
rect 30989 -4513 31077 -4497
rect 30989 -4681 31005 -4513
rect 31039 -4681 31077 -4513
rect 30989 -4697 31077 -4681
rect 31477 -4513 31565 -4497
rect 31477 -4681 31515 -4513
rect 31549 -4681 31565 -4513
rect 31477 -4697 31565 -4681
rect 31971 -3367 32059 -3351
rect 31971 -4135 31987 -3367
rect 32021 -4135 32059 -3367
rect 31971 -4151 32059 -4135
rect 32459 -3367 32547 -3351
rect 32459 -4135 32497 -3367
rect 32531 -4135 32547 -3367
rect 32459 -4151 32547 -4135
rect 32589 -3367 32677 -3351
rect 32589 -4135 32605 -3367
rect 32639 -4135 32677 -3367
rect 32589 -4151 32677 -4135
rect 33077 -3367 33165 -3351
rect 33077 -4135 33115 -3367
rect 33149 -4135 33165 -3367
rect 33077 -4151 33165 -4135
rect 31971 -4513 32059 -4497
rect 31971 -4681 31987 -4513
rect 32021 -4681 32059 -4513
rect 31971 -4697 32059 -4681
rect 32459 -4513 32547 -4497
rect 32459 -4681 32497 -4513
rect 32531 -4681 32547 -4513
rect 32459 -4697 32547 -4681
rect 32589 -4513 32677 -4497
rect 32589 -4681 32605 -4513
rect 32639 -4681 32677 -4513
rect 32589 -4697 32677 -4681
rect 33077 -4513 33165 -4497
rect 33077 -4681 33115 -4513
rect 33149 -4681 33165 -4513
rect 33077 -4697 33165 -4681
rect 33571 -3367 33659 -3351
rect 33571 -4135 33587 -3367
rect 33621 -4135 33659 -3367
rect 33571 -4151 33659 -4135
rect 34059 -3367 34147 -3351
rect 34059 -4135 34097 -3367
rect 34131 -4135 34147 -3367
rect 34059 -4151 34147 -4135
rect 34189 -3367 34277 -3351
rect 34189 -4135 34205 -3367
rect 34239 -4135 34277 -3367
rect 34189 -4151 34277 -4135
rect 34677 -3367 34765 -3351
rect 34677 -4135 34715 -3367
rect 34749 -4135 34765 -3367
rect 34677 -4151 34765 -4135
rect 33571 -4513 33659 -4497
rect 33571 -4681 33587 -4513
rect 33621 -4681 33659 -4513
rect 33571 -4697 33659 -4681
rect 34059 -4513 34147 -4497
rect 34059 -4681 34097 -4513
rect 34131 -4681 34147 -4513
rect 34059 -4697 34147 -4681
rect 34189 -4513 34277 -4497
rect 34189 -4681 34205 -4513
rect 34239 -4681 34277 -4513
rect 34189 -4697 34277 -4681
rect 34677 -4513 34765 -4497
rect 34677 -4681 34715 -4513
rect 34749 -4681 34765 -4513
rect 34677 -4697 34765 -4681
rect 35171 -3367 35259 -3351
rect 35171 -4135 35187 -3367
rect 35221 -4135 35259 -3367
rect 35171 -4151 35259 -4135
rect 35659 -3367 35747 -3351
rect 35659 -4135 35697 -3367
rect 35731 -4135 35747 -3367
rect 35659 -4151 35747 -4135
rect 35789 -3367 35877 -3351
rect 35789 -4135 35805 -3367
rect 35839 -4135 35877 -3367
rect 35789 -4151 35877 -4135
rect 36277 -3367 36365 -3351
rect 36277 -4135 36315 -3367
rect 36349 -4135 36365 -3367
rect 36277 -4151 36365 -4135
rect 35171 -4513 35259 -4497
rect 35171 -4681 35187 -4513
rect 35221 -4681 35259 -4513
rect 35171 -4697 35259 -4681
rect 35659 -4513 35747 -4497
rect 35659 -4681 35697 -4513
rect 35731 -4681 35747 -4513
rect 35659 -4697 35747 -4681
rect 35789 -4513 35877 -4497
rect 35789 -4681 35805 -4513
rect 35839 -4681 35877 -4513
rect 35789 -4697 35877 -4681
rect 36277 -4513 36365 -4497
rect 36277 -4681 36315 -4513
rect 36349 -4681 36365 -4513
rect 36277 -4697 36365 -4681
rect 36771 -3367 36859 -3351
rect 36771 -4135 36787 -3367
rect 36821 -4135 36859 -3367
rect 36771 -4151 36859 -4135
rect 37259 -3367 37347 -3351
rect 37259 -4135 37297 -3367
rect 37331 -4135 37347 -3367
rect 37259 -4151 37347 -4135
rect 37389 -3367 37477 -3351
rect 37389 -4135 37405 -3367
rect 37439 -4135 37477 -3367
rect 37389 -4151 37477 -4135
rect 37877 -3367 37965 -3351
rect 37877 -4135 37915 -3367
rect 37949 -4135 37965 -3367
rect 37877 -4151 37965 -4135
rect 36771 -4513 36859 -4497
rect 36771 -4681 36787 -4513
rect 36821 -4681 36859 -4513
rect 36771 -4697 36859 -4681
rect 37259 -4513 37347 -4497
rect 37259 -4681 37297 -4513
rect 37331 -4681 37347 -4513
rect 37259 -4697 37347 -4681
rect 37389 -4513 37477 -4497
rect 37389 -4681 37405 -4513
rect 37439 -4681 37477 -4513
rect 37389 -4697 37477 -4681
rect 37877 -4513 37965 -4497
rect 37877 -4681 37915 -4513
rect 37949 -4681 37965 -4513
rect 37877 -4697 37965 -4681
rect -40 -8232 57 -8216
rect -40 -8400 -24 -8232
rect 10 -8400 57 -8232
rect -40 -8416 57 -8400
rect 457 -8232 554 -8216
rect 457 -8400 504 -8232
rect 538 -8400 554 -8232
rect 457 -8416 554 -8400
rect 596 -8232 693 -8216
rect 596 -8400 612 -8232
rect 646 -8400 693 -8232
rect 596 -8416 693 -8400
rect 1093 -8232 1190 -8216
rect 1093 -8400 1140 -8232
rect 1174 -8400 1190 -8232
rect 1093 -8416 1190 -8400
rect -40 -8758 57 -8742
rect -40 -9526 -24 -8758
rect 10 -9526 57 -8758
rect -40 -9542 57 -9526
rect 457 -8758 554 -8742
rect 457 -9526 504 -8758
rect 538 -9526 554 -8758
rect 457 -9542 554 -9526
rect 596 -8758 693 -8742
rect 596 -9526 612 -8758
rect 646 -9526 693 -8758
rect 596 -9542 693 -9526
rect 1093 -8758 1190 -8742
rect 1093 -9526 1140 -8758
rect 1174 -9526 1190 -8758
rect 1093 -9542 1190 -9526
rect 1560 -8232 1657 -8216
rect 1560 -8400 1576 -8232
rect 1610 -8400 1657 -8232
rect 1560 -8416 1657 -8400
rect 2057 -8232 2154 -8216
rect 2057 -8400 2104 -8232
rect 2138 -8400 2154 -8232
rect 2057 -8416 2154 -8400
rect 2196 -8232 2293 -8216
rect 2196 -8400 2212 -8232
rect 2246 -8400 2293 -8232
rect 2196 -8416 2293 -8400
rect 2693 -8232 2790 -8216
rect 2693 -8400 2740 -8232
rect 2774 -8400 2790 -8232
rect 2693 -8416 2790 -8400
rect 1560 -8758 1657 -8742
rect 1560 -9526 1576 -8758
rect 1610 -9526 1657 -8758
rect 1560 -9542 1657 -9526
rect 2057 -8758 2154 -8742
rect 2057 -9526 2104 -8758
rect 2138 -9526 2154 -8758
rect 2057 -9542 2154 -9526
rect 2196 -8758 2293 -8742
rect 2196 -9526 2212 -8758
rect 2246 -9526 2293 -8758
rect 2196 -9542 2293 -9526
rect 2693 -8758 2790 -8742
rect 2693 -9526 2740 -8758
rect 2774 -9526 2790 -8758
rect 2693 -9542 2790 -9526
rect 3160 -8232 3257 -8216
rect 3160 -8400 3176 -8232
rect 3210 -8400 3257 -8232
rect 3160 -8416 3257 -8400
rect 3657 -8232 3754 -8216
rect 3657 -8400 3704 -8232
rect 3738 -8400 3754 -8232
rect 3657 -8416 3754 -8400
rect 3796 -8232 3893 -8216
rect 3796 -8400 3812 -8232
rect 3846 -8400 3893 -8232
rect 3796 -8416 3893 -8400
rect 4293 -8232 4390 -8216
rect 4293 -8400 4340 -8232
rect 4374 -8400 4390 -8232
rect 4293 -8416 4390 -8400
rect 3160 -8758 3257 -8742
rect 3160 -9526 3176 -8758
rect 3210 -9526 3257 -8758
rect 3160 -9542 3257 -9526
rect 3657 -8758 3754 -8742
rect 3657 -9526 3704 -8758
rect 3738 -9526 3754 -8758
rect 3657 -9542 3754 -9526
rect 3796 -8758 3893 -8742
rect 3796 -9526 3812 -8758
rect 3846 -9526 3893 -8758
rect 3796 -9542 3893 -9526
rect 4293 -8758 4390 -8742
rect 4293 -9526 4340 -8758
rect 4374 -9526 4390 -8758
rect 4293 -9542 4390 -9526
rect 4760 -8232 4857 -8216
rect 4760 -8400 4776 -8232
rect 4810 -8400 4857 -8232
rect 4760 -8416 4857 -8400
rect 5257 -8232 5354 -8216
rect 5257 -8400 5304 -8232
rect 5338 -8400 5354 -8232
rect 5257 -8416 5354 -8400
rect 5396 -8232 5493 -8216
rect 5396 -8400 5412 -8232
rect 5446 -8400 5493 -8232
rect 5396 -8416 5493 -8400
rect 5893 -8232 5990 -8216
rect 5893 -8400 5940 -8232
rect 5974 -8400 5990 -8232
rect 5893 -8416 5990 -8400
rect 4760 -8758 4857 -8742
rect 4760 -9526 4776 -8758
rect 4810 -9526 4857 -8758
rect 4760 -9542 4857 -9526
rect 5257 -8758 5354 -8742
rect 5257 -9526 5304 -8758
rect 5338 -9526 5354 -8758
rect 5257 -9542 5354 -9526
rect 5396 -8758 5493 -8742
rect 5396 -9526 5412 -8758
rect 5446 -9526 5493 -8758
rect 5396 -9542 5493 -9526
rect 5893 -8758 5990 -8742
rect 5893 -9526 5940 -8758
rect 5974 -9526 5990 -8758
rect 5893 -9542 5990 -9526
rect 6360 -8232 6457 -8216
rect 6360 -8400 6376 -8232
rect 6410 -8400 6457 -8232
rect 6360 -8416 6457 -8400
rect 6857 -8232 6954 -8216
rect 6857 -8400 6904 -8232
rect 6938 -8400 6954 -8232
rect 6857 -8416 6954 -8400
rect 6996 -8232 7093 -8216
rect 6996 -8400 7012 -8232
rect 7046 -8400 7093 -8232
rect 6996 -8416 7093 -8400
rect 7493 -8232 7590 -8216
rect 7493 -8400 7540 -8232
rect 7574 -8400 7590 -8232
rect 7493 -8416 7590 -8400
rect 6360 -8758 6457 -8742
rect 6360 -9526 6376 -8758
rect 6410 -9526 6457 -8758
rect 6360 -9542 6457 -9526
rect 6857 -8758 6954 -8742
rect 6857 -9526 6904 -8758
rect 6938 -9526 6954 -8758
rect 6857 -9542 6954 -9526
rect 6996 -8758 7093 -8742
rect 6996 -9526 7012 -8758
rect 7046 -9526 7093 -8758
rect 6996 -9542 7093 -9526
rect 7493 -8758 7590 -8742
rect 7493 -9526 7540 -8758
rect 7574 -9526 7590 -8758
rect 7493 -9542 7590 -9526
rect 7960 -8232 8057 -8216
rect 7960 -8400 7976 -8232
rect 8010 -8400 8057 -8232
rect 7960 -8416 8057 -8400
rect 8457 -8232 8554 -8216
rect 8457 -8400 8504 -8232
rect 8538 -8400 8554 -8232
rect 8457 -8416 8554 -8400
rect 8596 -8232 8693 -8216
rect 8596 -8400 8612 -8232
rect 8646 -8400 8693 -8232
rect 8596 -8416 8693 -8400
rect 9093 -8232 9190 -8216
rect 9093 -8400 9140 -8232
rect 9174 -8400 9190 -8232
rect 9093 -8416 9190 -8400
rect 7960 -8758 8057 -8742
rect 7960 -9526 7976 -8758
rect 8010 -9526 8057 -8758
rect 7960 -9542 8057 -9526
rect 8457 -8758 8554 -8742
rect 8457 -9526 8504 -8758
rect 8538 -9526 8554 -8758
rect 8457 -9542 8554 -9526
rect 8596 -8758 8693 -8742
rect 8596 -9526 8612 -8758
rect 8646 -9526 8693 -8758
rect 8596 -9542 8693 -9526
rect 9093 -8758 9190 -8742
rect 9093 -9526 9140 -8758
rect 9174 -9526 9190 -8758
rect 9093 -9542 9190 -9526
rect 9560 -8232 9657 -8216
rect 9560 -8400 9576 -8232
rect 9610 -8400 9657 -8232
rect 9560 -8416 9657 -8400
rect 10057 -8232 10154 -8216
rect 10057 -8400 10104 -8232
rect 10138 -8400 10154 -8232
rect 10057 -8416 10154 -8400
rect 10196 -8232 10293 -8216
rect 10196 -8400 10212 -8232
rect 10246 -8400 10293 -8232
rect 10196 -8416 10293 -8400
rect 10693 -8232 10790 -8216
rect 10693 -8400 10740 -8232
rect 10774 -8400 10790 -8232
rect 10693 -8416 10790 -8400
rect 9560 -8758 9657 -8742
rect 9560 -9526 9576 -8758
rect 9610 -9526 9657 -8758
rect 9560 -9542 9657 -9526
rect 10057 -8758 10154 -8742
rect 10057 -9526 10104 -8758
rect 10138 -9526 10154 -8758
rect 10057 -9542 10154 -9526
rect 10196 -8758 10293 -8742
rect 10196 -9526 10212 -8758
rect 10246 -9526 10293 -8758
rect 10196 -9542 10293 -9526
rect 10693 -8758 10790 -8742
rect 10693 -9526 10740 -8758
rect 10774 -9526 10790 -8758
rect 10693 -9542 10790 -9526
rect 11160 -8232 11257 -8216
rect 11160 -8400 11176 -8232
rect 11210 -8400 11257 -8232
rect 11160 -8416 11257 -8400
rect 11657 -8232 11754 -8216
rect 11657 -8400 11704 -8232
rect 11738 -8400 11754 -8232
rect 11657 -8416 11754 -8400
rect 11796 -8232 11893 -8216
rect 11796 -8400 11812 -8232
rect 11846 -8400 11893 -8232
rect 11796 -8416 11893 -8400
rect 12293 -8232 12390 -8216
rect 12293 -8400 12340 -8232
rect 12374 -8400 12390 -8232
rect 12293 -8416 12390 -8400
rect 11160 -8758 11257 -8742
rect 11160 -9526 11176 -8758
rect 11210 -9526 11257 -8758
rect 11160 -9542 11257 -9526
rect 11657 -8758 11754 -8742
rect 11657 -9526 11704 -8758
rect 11738 -9526 11754 -8758
rect 11657 -9542 11754 -9526
rect 11796 -8758 11893 -8742
rect 11796 -9526 11812 -8758
rect 11846 -9526 11893 -8758
rect 11796 -9542 11893 -9526
rect 12293 -8758 12390 -8742
rect 12293 -9526 12340 -8758
rect 12374 -9526 12390 -8758
rect 12293 -9542 12390 -9526
rect 12760 -8232 12857 -8216
rect 12760 -8400 12776 -8232
rect 12810 -8400 12857 -8232
rect 12760 -8416 12857 -8400
rect 13257 -8232 13354 -8216
rect 13257 -8400 13304 -8232
rect 13338 -8400 13354 -8232
rect 13257 -8416 13354 -8400
rect 13396 -8232 13493 -8216
rect 13396 -8400 13412 -8232
rect 13446 -8400 13493 -8232
rect 13396 -8416 13493 -8400
rect 13893 -8232 13990 -8216
rect 13893 -8400 13940 -8232
rect 13974 -8400 13990 -8232
rect 13893 -8416 13990 -8400
rect 12760 -8758 12857 -8742
rect 12760 -9526 12776 -8758
rect 12810 -9526 12857 -8758
rect 12760 -9542 12857 -9526
rect 13257 -8758 13354 -8742
rect 13257 -9526 13304 -8758
rect 13338 -9526 13354 -8758
rect 13257 -9542 13354 -9526
rect 13396 -8758 13493 -8742
rect 13396 -9526 13412 -8758
rect 13446 -9526 13493 -8758
rect 13396 -9542 13493 -9526
rect 13893 -8758 13990 -8742
rect 13893 -9526 13940 -8758
rect 13974 -9526 13990 -8758
rect 13893 -9542 13990 -9526
rect 14360 -8232 14457 -8216
rect 14360 -8400 14376 -8232
rect 14410 -8400 14457 -8232
rect 14360 -8416 14457 -8400
rect 14857 -8232 14954 -8216
rect 14857 -8400 14904 -8232
rect 14938 -8400 14954 -8232
rect 14857 -8416 14954 -8400
rect 14996 -8232 15093 -8216
rect 14996 -8400 15012 -8232
rect 15046 -8400 15093 -8232
rect 14996 -8416 15093 -8400
rect 15493 -8232 15590 -8216
rect 15493 -8400 15540 -8232
rect 15574 -8400 15590 -8232
rect 15493 -8416 15590 -8400
rect 14360 -8758 14457 -8742
rect 14360 -9526 14376 -8758
rect 14410 -9526 14457 -8758
rect 14360 -9542 14457 -9526
rect 14857 -8758 14954 -8742
rect 14857 -9526 14904 -8758
rect 14938 -9526 14954 -8758
rect 14857 -9542 14954 -9526
rect 14996 -8758 15093 -8742
rect 14996 -9526 15012 -8758
rect 15046 -9526 15093 -8758
rect 14996 -9542 15093 -9526
rect 15493 -8758 15590 -8742
rect 15493 -9526 15540 -8758
rect 15574 -9526 15590 -8758
rect 15493 -9542 15590 -9526
rect 15960 -8232 16057 -8216
rect 15960 -8400 15976 -8232
rect 16010 -8400 16057 -8232
rect 15960 -8416 16057 -8400
rect 16457 -8232 16554 -8216
rect 16457 -8400 16504 -8232
rect 16538 -8400 16554 -8232
rect 16457 -8416 16554 -8400
rect 16596 -8232 16693 -8216
rect 16596 -8400 16612 -8232
rect 16646 -8400 16693 -8232
rect 16596 -8416 16693 -8400
rect 17093 -8232 17190 -8216
rect 17093 -8400 17140 -8232
rect 17174 -8400 17190 -8232
rect 17093 -8416 17190 -8400
rect 15960 -8758 16057 -8742
rect 15960 -9526 15976 -8758
rect 16010 -9526 16057 -8758
rect 15960 -9542 16057 -9526
rect 16457 -8758 16554 -8742
rect 16457 -9526 16504 -8758
rect 16538 -9526 16554 -8758
rect 16457 -9542 16554 -9526
rect 16596 -8758 16693 -8742
rect 16596 -9526 16612 -8758
rect 16646 -9526 16693 -8758
rect 16596 -9542 16693 -9526
rect 17093 -8758 17190 -8742
rect 17093 -9526 17140 -8758
rect 17174 -9526 17190 -8758
rect 17093 -9542 17190 -9526
rect 17560 -8232 17657 -8216
rect 17560 -8400 17576 -8232
rect 17610 -8400 17657 -8232
rect 17560 -8416 17657 -8400
rect 18057 -8232 18154 -8216
rect 18057 -8400 18104 -8232
rect 18138 -8400 18154 -8232
rect 18057 -8416 18154 -8400
rect 18196 -8232 18293 -8216
rect 18196 -8400 18212 -8232
rect 18246 -8400 18293 -8232
rect 18196 -8416 18293 -8400
rect 18693 -8232 18790 -8216
rect 18693 -8400 18740 -8232
rect 18774 -8400 18790 -8232
rect 18693 -8416 18790 -8400
rect 17560 -8758 17657 -8742
rect 17560 -9526 17576 -8758
rect 17610 -9526 17657 -8758
rect 17560 -9542 17657 -9526
rect 18057 -8758 18154 -8742
rect 18057 -9526 18104 -8758
rect 18138 -9526 18154 -8758
rect 18057 -9542 18154 -9526
rect 18196 -8758 18293 -8742
rect 18196 -9526 18212 -8758
rect 18246 -9526 18293 -8758
rect 18196 -9542 18293 -9526
rect 18693 -8758 18790 -8742
rect 18693 -9526 18740 -8758
rect 18774 -9526 18790 -8758
rect 18693 -9542 18790 -9526
rect 19160 -8232 19257 -8216
rect 19160 -8400 19176 -8232
rect 19210 -8400 19257 -8232
rect 19160 -8416 19257 -8400
rect 19657 -8232 19754 -8216
rect 19657 -8400 19704 -8232
rect 19738 -8400 19754 -8232
rect 19657 -8416 19754 -8400
rect 19796 -8232 19893 -8216
rect 19796 -8400 19812 -8232
rect 19846 -8400 19893 -8232
rect 19796 -8416 19893 -8400
rect 20293 -8232 20390 -8216
rect 20293 -8400 20340 -8232
rect 20374 -8400 20390 -8232
rect 20293 -8416 20390 -8400
rect 19160 -8758 19257 -8742
rect 19160 -9526 19176 -8758
rect 19210 -9526 19257 -8758
rect 19160 -9542 19257 -9526
rect 19657 -8758 19754 -8742
rect 19657 -9526 19704 -8758
rect 19738 -9526 19754 -8758
rect 19657 -9542 19754 -9526
rect 19796 -8758 19893 -8742
rect 19796 -9526 19812 -8758
rect 19846 -9526 19893 -8758
rect 19796 -9542 19893 -9526
rect 20293 -8758 20390 -8742
rect 20293 -9526 20340 -8758
rect 20374 -9526 20390 -8758
rect 20293 -9542 20390 -9526
rect 20760 -8232 20857 -8216
rect 20760 -8400 20776 -8232
rect 20810 -8400 20857 -8232
rect 20760 -8416 20857 -8400
rect 21257 -8232 21354 -8216
rect 21257 -8400 21304 -8232
rect 21338 -8400 21354 -8232
rect 21257 -8416 21354 -8400
rect 21396 -8232 21493 -8216
rect 21396 -8400 21412 -8232
rect 21446 -8400 21493 -8232
rect 21396 -8416 21493 -8400
rect 21893 -8232 21990 -8216
rect 21893 -8400 21940 -8232
rect 21974 -8400 21990 -8232
rect 21893 -8416 21990 -8400
rect 20760 -8758 20857 -8742
rect 20760 -9526 20776 -8758
rect 20810 -9526 20857 -8758
rect 20760 -9542 20857 -9526
rect 21257 -8758 21354 -8742
rect 21257 -9526 21304 -8758
rect 21338 -9526 21354 -8758
rect 21257 -9542 21354 -9526
rect 21396 -8758 21493 -8742
rect 21396 -9526 21412 -8758
rect 21446 -9526 21493 -8758
rect 21396 -9542 21493 -9526
rect 21893 -8758 21990 -8742
rect 21893 -9526 21940 -8758
rect 21974 -9526 21990 -8758
rect 21893 -9542 21990 -9526
rect 22360 -8232 22457 -8216
rect 22360 -8400 22376 -8232
rect 22410 -8400 22457 -8232
rect 22360 -8416 22457 -8400
rect 22857 -8232 22954 -8216
rect 22857 -8400 22904 -8232
rect 22938 -8400 22954 -8232
rect 22857 -8416 22954 -8400
rect 22996 -8232 23093 -8216
rect 22996 -8400 23012 -8232
rect 23046 -8400 23093 -8232
rect 22996 -8416 23093 -8400
rect 23493 -8232 23590 -8216
rect 23493 -8400 23540 -8232
rect 23574 -8400 23590 -8232
rect 23493 -8416 23590 -8400
rect 22360 -8758 22457 -8742
rect 22360 -9526 22376 -8758
rect 22410 -9526 22457 -8758
rect 22360 -9542 22457 -9526
rect 22857 -8758 22954 -8742
rect 22857 -9526 22904 -8758
rect 22938 -9526 22954 -8758
rect 22857 -9542 22954 -9526
rect 22996 -8758 23093 -8742
rect 22996 -9526 23012 -8758
rect 23046 -9526 23093 -8758
rect 22996 -9542 23093 -9526
rect 23493 -8758 23590 -8742
rect 23493 -9526 23540 -8758
rect 23574 -9526 23590 -8758
rect 23493 -9542 23590 -9526
rect 23960 -8232 24057 -8216
rect 23960 -8400 23976 -8232
rect 24010 -8400 24057 -8232
rect 23960 -8416 24057 -8400
rect 24457 -8232 24554 -8216
rect 24457 -8400 24504 -8232
rect 24538 -8400 24554 -8232
rect 24457 -8416 24554 -8400
rect 24596 -8232 24693 -8216
rect 24596 -8400 24612 -8232
rect 24646 -8400 24693 -8232
rect 24596 -8416 24693 -8400
rect 25093 -8232 25190 -8216
rect 25093 -8400 25140 -8232
rect 25174 -8400 25190 -8232
rect 25093 -8416 25190 -8400
rect 23960 -8758 24057 -8742
rect 23960 -9526 23976 -8758
rect 24010 -9526 24057 -8758
rect 23960 -9542 24057 -9526
rect 24457 -8758 24554 -8742
rect 24457 -9526 24504 -8758
rect 24538 -9526 24554 -8758
rect 24457 -9542 24554 -9526
rect 24596 -8758 24693 -8742
rect 24596 -9526 24612 -8758
rect 24646 -9526 24693 -8758
rect 24596 -9542 24693 -9526
rect 25093 -8758 25190 -8742
rect 25093 -9526 25140 -8758
rect 25174 -9526 25190 -8758
rect 25093 -9542 25190 -9526
rect 25560 -8232 25657 -8216
rect 25560 -8400 25576 -8232
rect 25610 -8400 25657 -8232
rect 25560 -8416 25657 -8400
rect 26057 -8232 26154 -8216
rect 26057 -8400 26104 -8232
rect 26138 -8400 26154 -8232
rect 26057 -8416 26154 -8400
rect 26196 -8232 26293 -8216
rect 26196 -8400 26212 -8232
rect 26246 -8400 26293 -8232
rect 26196 -8416 26293 -8400
rect 26693 -8232 26790 -8216
rect 26693 -8400 26740 -8232
rect 26774 -8400 26790 -8232
rect 26693 -8416 26790 -8400
rect 25560 -8758 25657 -8742
rect 25560 -9526 25576 -8758
rect 25610 -9526 25657 -8758
rect 25560 -9542 25657 -9526
rect 26057 -8758 26154 -8742
rect 26057 -9526 26104 -8758
rect 26138 -9526 26154 -8758
rect 26057 -9542 26154 -9526
rect 26196 -8758 26293 -8742
rect 26196 -9526 26212 -8758
rect 26246 -9526 26293 -8758
rect 26196 -9542 26293 -9526
rect 26693 -8758 26790 -8742
rect 26693 -9526 26740 -8758
rect 26774 -9526 26790 -8758
rect 26693 -9542 26790 -9526
rect 27160 -8232 27257 -8216
rect 27160 -8400 27176 -8232
rect 27210 -8400 27257 -8232
rect 27160 -8416 27257 -8400
rect 27657 -8232 27754 -8216
rect 27657 -8400 27704 -8232
rect 27738 -8400 27754 -8232
rect 27657 -8416 27754 -8400
rect 27796 -8232 27893 -8216
rect 27796 -8400 27812 -8232
rect 27846 -8400 27893 -8232
rect 27796 -8416 27893 -8400
rect 28293 -8232 28390 -8216
rect 28293 -8400 28340 -8232
rect 28374 -8400 28390 -8232
rect 28293 -8416 28390 -8400
rect 27160 -8758 27257 -8742
rect 27160 -9526 27176 -8758
rect 27210 -9526 27257 -8758
rect 27160 -9542 27257 -9526
rect 27657 -8758 27754 -8742
rect 27657 -9526 27704 -8758
rect 27738 -9526 27754 -8758
rect 27657 -9542 27754 -9526
rect 27796 -8758 27893 -8742
rect 27796 -9526 27812 -8758
rect 27846 -9526 27893 -8758
rect 27796 -9542 27893 -9526
rect 28293 -8758 28390 -8742
rect 28293 -9526 28340 -8758
rect 28374 -9526 28390 -8758
rect 28293 -9542 28390 -9526
rect 28760 -8232 28857 -8216
rect 28760 -8400 28776 -8232
rect 28810 -8400 28857 -8232
rect 28760 -8416 28857 -8400
rect 29257 -8232 29354 -8216
rect 29257 -8400 29304 -8232
rect 29338 -8400 29354 -8232
rect 29257 -8416 29354 -8400
rect 29396 -8232 29493 -8216
rect 29396 -8400 29412 -8232
rect 29446 -8400 29493 -8232
rect 29396 -8416 29493 -8400
rect 29893 -8232 29990 -8216
rect 29893 -8400 29940 -8232
rect 29974 -8400 29990 -8232
rect 29893 -8416 29990 -8400
rect 28760 -8758 28857 -8742
rect 28760 -9526 28776 -8758
rect 28810 -9526 28857 -8758
rect 28760 -9542 28857 -9526
rect 29257 -8758 29354 -8742
rect 29257 -9526 29304 -8758
rect 29338 -9526 29354 -8758
rect 29257 -9542 29354 -9526
rect 29396 -8758 29493 -8742
rect 29396 -9526 29412 -8758
rect 29446 -9526 29493 -8758
rect 29396 -9542 29493 -9526
rect 29893 -8758 29990 -8742
rect 29893 -9526 29940 -8758
rect 29974 -9526 29990 -8758
rect 29893 -9542 29990 -9526
rect 30360 -8232 30457 -8216
rect 30360 -8400 30376 -8232
rect 30410 -8400 30457 -8232
rect 30360 -8416 30457 -8400
rect 30857 -8232 30954 -8216
rect 30857 -8400 30904 -8232
rect 30938 -8400 30954 -8232
rect 30857 -8416 30954 -8400
rect 30996 -8232 31093 -8216
rect 30996 -8400 31012 -8232
rect 31046 -8400 31093 -8232
rect 30996 -8416 31093 -8400
rect 31493 -8232 31590 -8216
rect 31493 -8400 31540 -8232
rect 31574 -8400 31590 -8232
rect 31493 -8416 31590 -8400
rect 30360 -8758 30457 -8742
rect 30360 -9526 30376 -8758
rect 30410 -9526 30457 -8758
rect 30360 -9542 30457 -9526
rect 30857 -8758 30954 -8742
rect 30857 -9526 30904 -8758
rect 30938 -9526 30954 -8758
rect 30857 -9542 30954 -9526
rect 30996 -8758 31093 -8742
rect 30996 -9526 31012 -8758
rect 31046 -9526 31093 -8758
rect 30996 -9542 31093 -9526
rect 31493 -8758 31590 -8742
rect 31493 -9526 31540 -8758
rect 31574 -9526 31590 -8758
rect 31493 -9542 31590 -9526
rect 31960 -8232 32057 -8216
rect 31960 -8400 31976 -8232
rect 32010 -8400 32057 -8232
rect 31960 -8416 32057 -8400
rect 32457 -8232 32554 -8216
rect 32457 -8400 32504 -8232
rect 32538 -8400 32554 -8232
rect 32457 -8416 32554 -8400
rect 32596 -8232 32693 -8216
rect 32596 -8400 32612 -8232
rect 32646 -8400 32693 -8232
rect 32596 -8416 32693 -8400
rect 33093 -8232 33190 -8216
rect 33093 -8400 33140 -8232
rect 33174 -8400 33190 -8232
rect 33093 -8416 33190 -8400
rect 31960 -8758 32057 -8742
rect 31960 -9526 31976 -8758
rect 32010 -9526 32057 -8758
rect 31960 -9542 32057 -9526
rect 32457 -8758 32554 -8742
rect 32457 -9526 32504 -8758
rect 32538 -9526 32554 -8758
rect 32457 -9542 32554 -9526
rect 32596 -8758 32693 -8742
rect 32596 -9526 32612 -8758
rect 32646 -9526 32693 -8758
rect 32596 -9542 32693 -9526
rect 33093 -8758 33190 -8742
rect 33093 -9526 33140 -8758
rect 33174 -9526 33190 -8758
rect 33093 -9542 33190 -9526
rect 33560 -8232 33657 -8216
rect 33560 -8400 33576 -8232
rect 33610 -8400 33657 -8232
rect 33560 -8416 33657 -8400
rect 34057 -8232 34154 -8216
rect 34057 -8400 34104 -8232
rect 34138 -8400 34154 -8232
rect 34057 -8416 34154 -8400
rect 34196 -8232 34293 -8216
rect 34196 -8400 34212 -8232
rect 34246 -8400 34293 -8232
rect 34196 -8416 34293 -8400
rect 34693 -8232 34790 -8216
rect 34693 -8400 34740 -8232
rect 34774 -8400 34790 -8232
rect 34693 -8416 34790 -8400
rect 33560 -8758 33657 -8742
rect 33560 -9526 33576 -8758
rect 33610 -9526 33657 -8758
rect 33560 -9542 33657 -9526
rect 34057 -8758 34154 -8742
rect 34057 -9526 34104 -8758
rect 34138 -9526 34154 -8758
rect 34057 -9542 34154 -9526
rect 34196 -8758 34293 -8742
rect 34196 -9526 34212 -8758
rect 34246 -9526 34293 -8758
rect 34196 -9542 34293 -9526
rect 34693 -8758 34790 -8742
rect 34693 -9526 34740 -8758
rect 34774 -9526 34790 -8758
rect 34693 -9542 34790 -9526
rect 35160 -8232 35257 -8216
rect 35160 -8400 35176 -8232
rect 35210 -8400 35257 -8232
rect 35160 -8416 35257 -8400
rect 35657 -8232 35754 -8216
rect 35657 -8400 35704 -8232
rect 35738 -8400 35754 -8232
rect 35657 -8416 35754 -8400
rect 35796 -8232 35893 -8216
rect 35796 -8400 35812 -8232
rect 35846 -8400 35893 -8232
rect 35796 -8416 35893 -8400
rect 36293 -8232 36390 -8216
rect 36293 -8400 36340 -8232
rect 36374 -8400 36390 -8232
rect 36293 -8416 36390 -8400
rect 35160 -8758 35257 -8742
rect 35160 -9526 35176 -8758
rect 35210 -9526 35257 -8758
rect 35160 -9542 35257 -9526
rect 35657 -8758 35754 -8742
rect 35657 -9526 35704 -8758
rect 35738 -9526 35754 -8758
rect 35657 -9542 35754 -9526
rect 35796 -8758 35893 -8742
rect 35796 -9526 35812 -8758
rect 35846 -9526 35893 -8758
rect 35796 -9542 35893 -9526
rect 36293 -8758 36390 -8742
rect 36293 -9526 36340 -8758
rect 36374 -9526 36390 -8758
rect 36293 -9542 36390 -9526
rect 36760 -8232 36857 -8216
rect 36760 -8400 36776 -8232
rect 36810 -8400 36857 -8232
rect 36760 -8416 36857 -8400
rect 37257 -8232 37354 -8216
rect 37257 -8400 37304 -8232
rect 37338 -8400 37354 -8232
rect 37257 -8416 37354 -8400
rect 37396 -8232 37493 -8216
rect 37396 -8400 37412 -8232
rect 37446 -8400 37493 -8232
rect 37396 -8416 37493 -8400
rect 37893 -8232 37990 -8216
rect 37893 -8400 37940 -8232
rect 37974 -8400 37990 -8232
rect 37893 -8416 37990 -8400
rect 36760 -8758 36857 -8742
rect 36760 -9526 36776 -8758
rect 36810 -9526 36857 -8758
rect 36760 -9542 36857 -9526
rect 37257 -8758 37354 -8742
rect 37257 -9526 37304 -8758
rect 37338 -9526 37354 -8758
rect 37257 -9542 37354 -9526
rect 37396 -8758 37493 -8742
rect 37396 -9526 37412 -8758
rect 37446 -9526 37493 -8758
rect 37396 -9542 37493 -9526
rect 37893 -8758 37990 -8742
rect 37893 -9526 37940 -8758
rect 37974 -9526 37990 -8758
rect 37893 -9542 37990 -9526
rect -40 -10032 57 -10016
rect -40 -10200 -24 -10032
rect 10 -10200 57 -10032
rect -40 -10216 57 -10200
rect 457 -10032 554 -10016
rect 457 -10200 504 -10032
rect 538 -10200 554 -10032
rect 457 -10216 554 -10200
rect 596 -10032 693 -10016
rect 596 -10200 612 -10032
rect 646 -10200 693 -10032
rect 596 -10216 693 -10200
rect 1093 -10032 1190 -10016
rect 1093 -10200 1140 -10032
rect 1174 -10200 1190 -10032
rect 1093 -10216 1190 -10200
rect -40 -10558 57 -10542
rect -40 -11326 -24 -10558
rect 10 -11326 57 -10558
rect -40 -11342 57 -11326
rect 457 -10558 554 -10542
rect 457 -11326 504 -10558
rect 538 -11326 554 -10558
rect 457 -11342 554 -11326
rect 596 -10558 693 -10542
rect 596 -11326 612 -10558
rect 646 -11326 693 -10558
rect 596 -11342 693 -11326
rect 1093 -10558 1190 -10542
rect 1093 -11326 1140 -10558
rect 1174 -11326 1190 -10558
rect 1093 -11342 1190 -11326
rect 1560 -10032 1657 -10016
rect 1560 -10200 1576 -10032
rect 1610 -10200 1657 -10032
rect 1560 -10216 1657 -10200
rect 2057 -10032 2154 -10016
rect 2057 -10200 2104 -10032
rect 2138 -10200 2154 -10032
rect 2057 -10216 2154 -10200
rect 2196 -10032 2293 -10016
rect 2196 -10200 2212 -10032
rect 2246 -10200 2293 -10032
rect 2196 -10216 2293 -10200
rect 2693 -10032 2790 -10016
rect 2693 -10200 2740 -10032
rect 2774 -10200 2790 -10032
rect 2693 -10216 2790 -10200
rect 1560 -10558 1657 -10542
rect 1560 -11326 1576 -10558
rect 1610 -11326 1657 -10558
rect 1560 -11342 1657 -11326
rect 2057 -10558 2154 -10542
rect 2057 -11326 2104 -10558
rect 2138 -11326 2154 -10558
rect 2057 -11342 2154 -11326
rect 2196 -10558 2293 -10542
rect 2196 -11326 2212 -10558
rect 2246 -11326 2293 -10558
rect 2196 -11342 2293 -11326
rect 2693 -10558 2790 -10542
rect 2693 -11326 2740 -10558
rect 2774 -11326 2790 -10558
rect 2693 -11342 2790 -11326
rect 3160 -10032 3257 -10016
rect 3160 -10200 3176 -10032
rect 3210 -10200 3257 -10032
rect 3160 -10216 3257 -10200
rect 3657 -10032 3754 -10016
rect 3657 -10200 3704 -10032
rect 3738 -10200 3754 -10032
rect 3657 -10216 3754 -10200
rect 3796 -10032 3893 -10016
rect 3796 -10200 3812 -10032
rect 3846 -10200 3893 -10032
rect 3796 -10216 3893 -10200
rect 4293 -10032 4390 -10016
rect 4293 -10200 4340 -10032
rect 4374 -10200 4390 -10032
rect 4293 -10216 4390 -10200
rect 3160 -10558 3257 -10542
rect 3160 -11326 3176 -10558
rect 3210 -11326 3257 -10558
rect 3160 -11342 3257 -11326
rect 3657 -10558 3754 -10542
rect 3657 -11326 3704 -10558
rect 3738 -11326 3754 -10558
rect 3657 -11342 3754 -11326
rect 3796 -10558 3893 -10542
rect 3796 -11326 3812 -10558
rect 3846 -11326 3893 -10558
rect 3796 -11342 3893 -11326
rect 4293 -10558 4390 -10542
rect 4293 -11326 4340 -10558
rect 4374 -11326 4390 -10558
rect 4293 -11342 4390 -11326
rect 4760 -10032 4857 -10016
rect 4760 -10200 4776 -10032
rect 4810 -10200 4857 -10032
rect 4760 -10216 4857 -10200
rect 5257 -10032 5354 -10016
rect 5257 -10200 5304 -10032
rect 5338 -10200 5354 -10032
rect 5257 -10216 5354 -10200
rect 5396 -10032 5493 -10016
rect 5396 -10200 5412 -10032
rect 5446 -10200 5493 -10032
rect 5396 -10216 5493 -10200
rect 5893 -10032 5990 -10016
rect 5893 -10200 5940 -10032
rect 5974 -10200 5990 -10032
rect 5893 -10216 5990 -10200
rect 4760 -10558 4857 -10542
rect 4760 -11326 4776 -10558
rect 4810 -11326 4857 -10558
rect 4760 -11342 4857 -11326
rect 5257 -10558 5354 -10542
rect 5257 -11326 5304 -10558
rect 5338 -11326 5354 -10558
rect 5257 -11342 5354 -11326
rect 5396 -10558 5493 -10542
rect 5396 -11326 5412 -10558
rect 5446 -11326 5493 -10558
rect 5396 -11342 5493 -11326
rect 5893 -10558 5990 -10542
rect 5893 -11326 5940 -10558
rect 5974 -11326 5990 -10558
rect 5893 -11342 5990 -11326
rect 6360 -10032 6457 -10016
rect 6360 -10200 6376 -10032
rect 6410 -10200 6457 -10032
rect 6360 -10216 6457 -10200
rect 6857 -10032 6954 -10016
rect 6857 -10200 6904 -10032
rect 6938 -10200 6954 -10032
rect 6857 -10216 6954 -10200
rect 6996 -10032 7093 -10016
rect 6996 -10200 7012 -10032
rect 7046 -10200 7093 -10032
rect 6996 -10216 7093 -10200
rect 7493 -10032 7590 -10016
rect 7493 -10200 7540 -10032
rect 7574 -10200 7590 -10032
rect 7493 -10216 7590 -10200
rect 6360 -10558 6457 -10542
rect 6360 -11326 6376 -10558
rect 6410 -11326 6457 -10558
rect 6360 -11342 6457 -11326
rect 6857 -10558 6954 -10542
rect 6857 -11326 6904 -10558
rect 6938 -11326 6954 -10558
rect 6857 -11342 6954 -11326
rect 6996 -10558 7093 -10542
rect 6996 -11326 7012 -10558
rect 7046 -11326 7093 -10558
rect 6996 -11342 7093 -11326
rect 7493 -10558 7590 -10542
rect 7493 -11326 7540 -10558
rect 7574 -11326 7590 -10558
rect 7493 -11342 7590 -11326
rect 7960 -10032 8057 -10016
rect 7960 -10200 7976 -10032
rect 8010 -10200 8057 -10032
rect 7960 -10216 8057 -10200
rect 8457 -10032 8554 -10016
rect 8457 -10200 8504 -10032
rect 8538 -10200 8554 -10032
rect 8457 -10216 8554 -10200
rect 8596 -10032 8693 -10016
rect 8596 -10200 8612 -10032
rect 8646 -10200 8693 -10032
rect 8596 -10216 8693 -10200
rect 9093 -10032 9190 -10016
rect 9093 -10200 9140 -10032
rect 9174 -10200 9190 -10032
rect 9093 -10216 9190 -10200
rect 7960 -10558 8057 -10542
rect 7960 -11326 7976 -10558
rect 8010 -11326 8057 -10558
rect 7960 -11342 8057 -11326
rect 8457 -10558 8554 -10542
rect 8457 -11326 8504 -10558
rect 8538 -11326 8554 -10558
rect 8457 -11342 8554 -11326
rect 8596 -10558 8693 -10542
rect 8596 -11326 8612 -10558
rect 8646 -11326 8693 -10558
rect 8596 -11342 8693 -11326
rect 9093 -10558 9190 -10542
rect 9093 -11326 9140 -10558
rect 9174 -11326 9190 -10558
rect 9093 -11342 9190 -11326
rect 9560 -10032 9657 -10016
rect 9560 -10200 9576 -10032
rect 9610 -10200 9657 -10032
rect 9560 -10216 9657 -10200
rect 10057 -10032 10154 -10016
rect 10057 -10200 10104 -10032
rect 10138 -10200 10154 -10032
rect 10057 -10216 10154 -10200
rect 10196 -10032 10293 -10016
rect 10196 -10200 10212 -10032
rect 10246 -10200 10293 -10032
rect 10196 -10216 10293 -10200
rect 10693 -10032 10790 -10016
rect 10693 -10200 10740 -10032
rect 10774 -10200 10790 -10032
rect 10693 -10216 10790 -10200
rect 9560 -10558 9657 -10542
rect 9560 -11326 9576 -10558
rect 9610 -11326 9657 -10558
rect 9560 -11342 9657 -11326
rect 10057 -10558 10154 -10542
rect 10057 -11326 10104 -10558
rect 10138 -11326 10154 -10558
rect 10057 -11342 10154 -11326
rect 10196 -10558 10293 -10542
rect 10196 -11326 10212 -10558
rect 10246 -11326 10293 -10558
rect 10196 -11342 10293 -11326
rect 10693 -10558 10790 -10542
rect 10693 -11326 10740 -10558
rect 10774 -11326 10790 -10558
rect 10693 -11342 10790 -11326
rect 11160 -10032 11257 -10016
rect 11160 -10200 11176 -10032
rect 11210 -10200 11257 -10032
rect 11160 -10216 11257 -10200
rect 11657 -10032 11754 -10016
rect 11657 -10200 11704 -10032
rect 11738 -10200 11754 -10032
rect 11657 -10216 11754 -10200
rect 11796 -10032 11893 -10016
rect 11796 -10200 11812 -10032
rect 11846 -10200 11893 -10032
rect 11796 -10216 11893 -10200
rect 12293 -10032 12390 -10016
rect 12293 -10200 12340 -10032
rect 12374 -10200 12390 -10032
rect 12293 -10216 12390 -10200
rect 11160 -10558 11257 -10542
rect 11160 -11326 11176 -10558
rect 11210 -11326 11257 -10558
rect 11160 -11342 11257 -11326
rect 11657 -10558 11754 -10542
rect 11657 -11326 11704 -10558
rect 11738 -11326 11754 -10558
rect 11657 -11342 11754 -11326
rect 11796 -10558 11893 -10542
rect 11796 -11326 11812 -10558
rect 11846 -11326 11893 -10558
rect 11796 -11342 11893 -11326
rect 12293 -10558 12390 -10542
rect 12293 -11326 12340 -10558
rect 12374 -11326 12390 -10558
rect 12293 -11342 12390 -11326
rect 12760 -10032 12857 -10016
rect 12760 -10200 12776 -10032
rect 12810 -10200 12857 -10032
rect 12760 -10216 12857 -10200
rect 13257 -10032 13354 -10016
rect 13257 -10200 13304 -10032
rect 13338 -10200 13354 -10032
rect 13257 -10216 13354 -10200
rect 13396 -10032 13493 -10016
rect 13396 -10200 13412 -10032
rect 13446 -10200 13493 -10032
rect 13396 -10216 13493 -10200
rect 13893 -10032 13990 -10016
rect 13893 -10200 13940 -10032
rect 13974 -10200 13990 -10032
rect 13893 -10216 13990 -10200
rect 12760 -10558 12857 -10542
rect 12760 -11326 12776 -10558
rect 12810 -11326 12857 -10558
rect 12760 -11342 12857 -11326
rect 13257 -10558 13354 -10542
rect 13257 -11326 13304 -10558
rect 13338 -11326 13354 -10558
rect 13257 -11342 13354 -11326
rect 13396 -10558 13493 -10542
rect 13396 -11326 13412 -10558
rect 13446 -11326 13493 -10558
rect 13396 -11342 13493 -11326
rect 13893 -10558 13990 -10542
rect 13893 -11326 13940 -10558
rect 13974 -11326 13990 -10558
rect 13893 -11342 13990 -11326
rect 14360 -10032 14457 -10016
rect 14360 -10200 14376 -10032
rect 14410 -10200 14457 -10032
rect 14360 -10216 14457 -10200
rect 14857 -10032 14954 -10016
rect 14857 -10200 14904 -10032
rect 14938 -10200 14954 -10032
rect 14857 -10216 14954 -10200
rect 14996 -10032 15093 -10016
rect 14996 -10200 15012 -10032
rect 15046 -10200 15093 -10032
rect 14996 -10216 15093 -10200
rect 15493 -10032 15590 -10016
rect 15493 -10200 15540 -10032
rect 15574 -10200 15590 -10032
rect 15493 -10216 15590 -10200
rect 14360 -10558 14457 -10542
rect 14360 -11326 14376 -10558
rect 14410 -11326 14457 -10558
rect 14360 -11342 14457 -11326
rect 14857 -10558 14954 -10542
rect 14857 -11326 14904 -10558
rect 14938 -11326 14954 -10558
rect 14857 -11342 14954 -11326
rect 14996 -10558 15093 -10542
rect 14996 -11326 15012 -10558
rect 15046 -11326 15093 -10558
rect 14996 -11342 15093 -11326
rect 15493 -10558 15590 -10542
rect 15493 -11326 15540 -10558
rect 15574 -11326 15590 -10558
rect 15493 -11342 15590 -11326
rect 15960 -10032 16057 -10016
rect 15960 -10200 15976 -10032
rect 16010 -10200 16057 -10032
rect 15960 -10216 16057 -10200
rect 16457 -10032 16554 -10016
rect 16457 -10200 16504 -10032
rect 16538 -10200 16554 -10032
rect 16457 -10216 16554 -10200
rect 16596 -10032 16693 -10016
rect 16596 -10200 16612 -10032
rect 16646 -10200 16693 -10032
rect 16596 -10216 16693 -10200
rect 17093 -10032 17190 -10016
rect 17093 -10200 17140 -10032
rect 17174 -10200 17190 -10032
rect 17093 -10216 17190 -10200
rect 15960 -10558 16057 -10542
rect 15960 -11326 15976 -10558
rect 16010 -11326 16057 -10558
rect 15960 -11342 16057 -11326
rect 16457 -10558 16554 -10542
rect 16457 -11326 16504 -10558
rect 16538 -11326 16554 -10558
rect 16457 -11342 16554 -11326
rect 16596 -10558 16693 -10542
rect 16596 -11326 16612 -10558
rect 16646 -11326 16693 -10558
rect 16596 -11342 16693 -11326
rect 17093 -10558 17190 -10542
rect 17093 -11326 17140 -10558
rect 17174 -11326 17190 -10558
rect 17093 -11342 17190 -11326
rect 17560 -10032 17657 -10016
rect 17560 -10200 17576 -10032
rect 17610 -10200 17657 -10032
rect 17560 -10216 17657 -10200
rect 18057 -10032 18154 -10016
rect 18057 -10200 18104 -10032
rect 18138 -10200 18154 -10032
rect 18057 -10216 18154 -10200
rect 18196 -10032 18293 -10016
rect 18196 -10200 18212 -10032
rect 18246 -10200 18293 -10032
rect 18196 -10216 18293 -10200
rect 18693 -10032 18790 -10016
rect 18693 -10200 18740 -10032
rect 18774 -10200 18790 -10032
rect 18693 -10216 18790 -10200
rect 17560 -10558 17657 -10542
rect 17560 -11326 17576 -10558
rect 17610 -11326 17657 -10558
rect 17560 -11342 17657 -11326
rect 18057 -10558 18154 -10542
rect 18057 -11326 18104 -10558
rect 18138 -11326 18154 -10558
rect 18057 -11342 18154 -11326
rect 18196 -10558 18293 -10542
rect 18196 -11326 18212 -10558
rect 18246 -11326 18293 -10558
rect 18196 -11342 18293 -11326
rect 18693 -10558 18790 -10542
rect 18693 -11326 18740 -10558
rect 18774 -11326 18790 -10558
rect 18693 -11342 18790 -11326
rect 19160 -10032 19257 -10016
rect 19160 -10200 19176 -10032
rect 19210 -10200 19257 -10032
rect 19160 -10216 19257 -10200
rect 19657 -10032 19754 -10016
rect 19657 -10200 19704 -10032
rect 19738 -10200 19754 -10032
rect 19657 -10216 19754 -10200
rect 19796 -10032 19893 -10016
rect 19796 -10200 19812 -10032
rect 19846 -10200 19893 -10032
rect 19796 -10216 19893 -10200
rect 20293 -10032 20390 -10016
rect 20293 -10200 20340 -10032
rect 20374 -10200 20390 -10032
rect 20293 -10216 20390 -10200
rect 19160 -10558 19257 -10542
rect 19160 -11326 19176 -10558
rect 19210 -11326 19257 -10558
rect 19160 -11342 19257 -11326
rect 19657 -10558 19754 -10542
rect 19657 -11326 19704 -10558
rect 19738 -11326 19754 -10558
rect 19657 -11342 19754 -11326
rect 19796 -10558 19893 -10542
rect 19796 -11326 19812 -10558
rect 19846 -11326 19893 -10558
rect 19796 -11342 19893 -11326
rect 20293 -10558 20390 -10542
rect 20293 -11326 20340 -10558
rect 20374 -11326 20390 -10558
rect 20293 -11342 20390 -11326
rect 20760 -10032 20857 -10016
rect 20760 -10200 20776 -10032
rect 20810 -10200 20857 -10032
rect 20760 -10216 20857 -10200
rect 21257 -10032 21354 -10016
rect 21257 -10200 21304 -10032
rect 21338 -10200 21354 -10032
rect 21257 -10216 21354 -10200
rect 21396 -10032 21493 -10016
rect 21396 -10200 21412 -10032
rect 21446 -10200 21493 -10032
rect 21396 -10216 21493 -10200
rect 21893 -10032 21990 -10016
rect 21893 -10200 21940 -10032
rect 21974 -10200 21990 -10032
rect 21893 -10216 21990 -10200
rect 20760 -10558 20857 -10542
rect 20760 -11326 20776 -10558
rect 20810 -11326 20857 -10558
rect 20760 -11342 20857 -11326
rect 21257 -10558 21354 -10542
rect 21257 -11326 21304 -10558
rect 21338 -11326 21354 -10558
rect 21257 -11342 21354 -11326
rect 21396 -10558 21493 -10542
rect 21396 -11326 21412 -10558
rect 21446 -11326 21493 -10558
rect 21396 -11342 21493 -11326
rect 21893 -10558 21990 -10542
rect 21893 -11326 21940 -10558
rect 21974 -11326 21990 -10558
rect 21893 -11342 21990 -11326
rect 22360 -10032 22457 -10016
rect 22360 -10200 22376 -10032
rect 22410 -10200 22457 -10032
rect 22360 -10216 22457 -10200
rect 22857 -10032 22954 -10016
rect 22857 -10200 22904 -10032
rect 22938 -10200 22954 -10032
rect 22857 -10216 22954 -10200
rect 22996 -10032 23093 -10016
rect 22996 -10200 23012 -10032
rect 23046 -10200 23093 -10032
rect 22996 -10216 23093 -10200
rect 23493 -10032 23590 -10016
rect 23493 -10200 23540 -10032
rect 23574 -10200 23590 -10032
rect 23493 -10216 23590 -10200
rect 22360 -10558 22457 -10542
rect 22360 -11326 22376 -10558
rect 22410 -11326 22457 -10558
rect 22360 -11342 22457 -11326
rect 22857 -10558 22954 -10542
rect 22857 -11326 22904 -10558
rect 22938 -11326 22954 -10558
rect 22857 -11342 22954 -11326
rect 22996 -10558 23093 -10542
rect 22996 -11326 23012 -10558
rect 23046 -11326 23093 -10558
rect 22996 -11342 23093 -11326
rect 23493 -10558 23590 -10542
rect 23493 -11326 23540 -10558
rect 23574 -11326 23590 -10558
rect 23493 -11342 23590 -11326
rect 23960 -10032 24057 -10016
rect 23960 -10200 23976 -10032
rect 24010 -10200 24057 -10032
rect 23960 -10216 24057 -10200
rect 24457 -10032 24554 -10016
rect 24457 -10200 24504 -10032
rect 24538 -10200 24554 -10032
rect 24457 -10216 24554 -10200
rect 24596 -10032 24693 -10016
rect 24596 -10200 24612 -10032
rect 24646 -10200 24693 -10032
rect 24596 -10216 24693 -10200
rect 25093 -10032 25190 -10016
rect 25093 -10200 25140 -10032
rect 25174 -10200 25190 -10032
rect 25093 -10216 25190 -10200
rect 23960 -10558 24057 -10542
rect 23960 -11326 23976 -10558
rect 24010 -11326 24057 -10558
rect 23960 -11342 24057 -11326
rect 24457 -10558 24554 -10542
rect 24457 -11326 24504 -10558
rect 24538 -11326 24554 -10558
rect 24457 -11342 24554 -11326
rect 24596 -10558 24693 -10542
rect 24596 -11326 24612 -10558
rect 24646 -11326 24693 -10558
rect 24596 -11342 24693 -11326
rect 25093 -10558 25190 -10542
rect 25093 -11326 25140 -10558
rect 25174 -11326 25190 -10558
rect 25093 -11342 25190 -11326
rect 25560 -10032 25657 -10016
rect 25560 -10200 25576 -10032
rect 25610 -10200 25657 -10032
rect 25560 -10216 25657 -10200
rect 26057 -10032 26154 -10016
rect 26057 -10200 26104 -10032
rect 26138 -10200 26154 -10032
rect 26057 -10216 26154 -10200
rect 26196 -10032 26293 -10016
rect 26196 -10200 26212 -10032
rect 26246 -10200 26293 -10032
rect 26196 -10216 26293 -10200
rect 26693 -10032 26790 -10016
rect 26693 -10200 26740 -10032
rect 26774 -10200 26790 -10032
rect 26693 -10216 26790 -10200
rect 25560 -10558 25657 -10542
rect 25560 -11326 25576 -10558
rect 25610 -11326 25657 -10558
rect 25560 -11342 25657 -11326
rect 26057 -10558 26154 -10542
rect 26057 -11326 26104 -10558
rect 26138 -11326 26154 -10558
rect 26057 -11342 26154 -11326
rect 26196 -10558 26293 -10542
rect 26196 -11326 26212 -10558
rect 26246 -11326 26293 -10558
rect 26196 -11342 26293 -11326
rect 26693 -10558 26790 -10542
rect 26693 -11326 26740 -10558
rect 26774 -11326 26790 -10558
rect 26693 -11342 26790 -11326
rect 27160 -10032 27257 -10016
rect 27160 -10200 27176 -10032
rect 27210 -10200 27257 -10032
rect 27160 -10216 27257 -10200
rect 27657 -10032 27754 -10016
rect 27657 -10200 27704 -10032
rect 27738 -10200 27754 -10032
rect 27657 -10216 27754 -10200
rect 27796 -10032 27893 -10016
rect 27796 -10200 27812 -10032
rect 27846 -10200 27893 -10032
rect 27796 -10216 27893 -10200
rect 28293 -10032 28390 -10016
rect 28293 -10200 28340 -10032
rect 28374 -10200 28390 -10032
rect 28293 -10216 28390 -10200
rect 27160 -10558 27257 -10542
rect 27160 -11326 27176 -10558
rect 27210 -11326 27257 -10558
rect 27160 -11342 27257 -11326
rect 27657 -10558 27754 -10542
rect 27657 -11326 27704 -10558
rect 27738 -11326 27754 -10558
rect 27657 -11342 27754 -11326
rect 27796 -10558 27893 -10542
rect 27796 -11326 27812 -10558
rect 27846 -11326 27893 -10558
rect 27796 -11342 27893 -11326
rect 28293 -10558 28390 -10542
rect 28293 -11326 28340 -10558
rect 28374 -11326 28390 -10558
rect 28293 -11342 28390 -11326
rect 28760 -10032 28857 -10016
rect 28760 -10200 28776 -10032
rect 28810 -10200 28857 -10032
rect 28760 -10216 28857 -10200
rect 29257 -10032 29354 -10016
rect 29257 -10200 29304 -10032
rect 29338 -10200 29354 -10032
rect 29257 -10216 29354 -10200
rect 29396 -10032 29493 -10016
rect 29396 -10200 29412 -10032
rect 29446 -10200 29493 -10032
rect 29396 -10216 29493 -10200
rect 29893 -10032 29990 -10016
rect 29893 -10200 29940 -10032
rect 29974 -10200 29990 -10032
rect 29893 -10216 29990 -10200
rect 28760 -10558 28857 -10542
rect 28760 -11326 28776 -10558
rect 28810 -11326 28857 -10558
rect 28760 -11342 28857 -11326
rect 29257 -10558 29354 -10542
rect 29257 -11326 29304 -10558
rect 29338 -11326 29354 -10558
rect 29257 -11342 29354 -11326
rect 29396 -10558 29493 -10542
rect 29396 -11326 29412 -10558
rect 29446 -11326 29493 -10558
rect 29396 -11342 29493 -11326
rect 29893 -10558 29990 -10542
rect 29893 -11326 29940 -10558
rect 29974 -11326 29990 -10558
rect 29893 -11342 29990 -11326
rect 30360 -10032 30457 -10016
rect 30360 -10200 30376 -10032
rect 30410 -10200 30457 -10032
rect 30360 -10216 30457 -10200
rect 30857 -10032 30954 -10016
rect 30857 -10200 30904 -10032
rect 30938 -10200 30954 -10032
rect 30857 -10216 30954 -10200
rect 30996 -10032 31093 -10016
rect 30996 -10200 31012 -10032
rect 31046 -10200 31093 -10032
rect 30996 -10216 31093 -10200
rect 31493 -10032 31590 -10016
rect 31493 -10200 31540 -10032
rect 31574 -10200 31590 -10032
rect 31493 -10216 31590 -10200
rect 30360 -10558 30457 -10542
rect 30360 -11326 30376 -10558
rect 30410 -11326 30457 -10558
rect 30360 -11342 30457 -11326
rect 30857 -10558 30954 -10542
rect 30857 -11326 30904 -10558
rect 30938 -11326 30954 -10558
rect 30857 -11342 30954 -11326
rect 30996 -10558 31093 -10542
rect 30996 -11326 31012 -10558
rect 31046 -11326 31093 -10558
rect 30996 -11342 31093 -11326
rect 31493 -10558 31590 -10542
rect 31493 -11326 31540 -10558
rect 31574 -11326 31590 -10558
rect 31493 -11342 31590 -11326
rect 31960 -10032 32057 -10016
rect 31960 -10200 31976 -10032
rect 32010 -10200 32057 -10032
rect 31960 -10216 32057 -10200
rect 32457 -10032 32554 -10016
rect 32457 -10200 32504 -10032
rect 32538 -10200 32554 -10032
rect 32457 -10216 32554 -10200
rect 32596 -10032 32693 -10016
rect 32596 -10200 32612 -10032
rect 32646 -10200 32693 -10032
rect 32596 -10216 32693 -10200
rect 33093 -10032 33190 -10016
rect 33093 -10200 33140 -10032
rect 33174 -10200 33190 -10032
rect 33093 -10216 33190 -10200
rect 31960 -10558 32057 -10542
rect 31960 -11326 31976 -10558
rect 32010 -11326 32057 -10558
rect 31960 -11342 32057 -11326
rect 32457 -10558 32554 -10542
rect 32457 -11326 32504 -10558
rect 32538 -11326 32554 -10558
rect 32457 -11342 32554 -11326
rect 32596 -10558 32693 -10542
rect 32596 -11326 32612 -10558
rect 32646 -11326 32693 -10558
rect 32596 -11342 32693 -11326
rect 33093 -10558 33190 -10542
rect 33093 -11326 33140 -10558
rect 33174 -11326 33190 -10558
rect 33093 -11342 33190 -11326
rect 33560 -10032 33657 -10016
rect 33560 -10200 33576 -10032
rect 33610 -10200 33657 -10032
rect 33560 -10216 33657 -10200
rect 34057 -10032 34154 -10016
rect 34057 -10200 34104 -10032
rect 34138 -10200 34154 -10032
rect 34057 -10216 34154 -10200
rect 34196 -10032 34293 -10016
rect 34196 -10200 34212 -10032
rect 34246 -10200 34293 -10032
rect 34196 -10216 34293 -10200
rect 34693 -10032 34790 -10016
rect 34693 -10200 34740 -10032
rect 34774 -10200 34790 -10032
rect 34693 -10216 34790 -10200
rect 33560 -10558 33657 -10542
rect 33560 -11326 33576 -10558
rect 33610 -11326 33657 -10558
rect 33560 -11342 33657 -11326
rect 34057 -10558 34154 -10542
rect 34057 -11326 34104 -10558
rect 34138 -11326 34154 -10558
rect 34057 -11342 34154 -11326
rect 34196 -10558 34293 -10542
rect 34196 -11326 34212 -10558
rect 34246 -11326 34293 -10558
rect 34196 -11342 34293 -11326
rect 34693 -10558 34790 -10542
rect 34693 -11326 34740 -10558
rect 34774 -11326 34790 -10558
rect 34693 -11342 34790 -11326
rect 35160 -10032 35257 -10016
rect 35160 -10200 35176 -10032
rect 35210 -10200 35257 -10032
rect 35160 -10216 35257 -10200
rect 35657 -10032 35754 -10016
rect 35657 -10200 35704 -10032
rect 35738 -10200 35754 -10032
rect 35657 -10216 35754 -10200
rect 35796 -10032 35893 -10016
rect 35796 -10200 35812 -10032
rect 35846 -10200 35893 -10032
rect 35796 -10216 35893 -10200
rect 36293 -10032 36390 -10016
rect 36293 -10200 36340 -10032
rect 36374 -10200 36390 -10032
rect 36293 -10216 36390 -10200
rect 35160 -10558 35257 -10542
rect 35160 -11326 35176 -10558
rect 35210 -11326 35257 -10558
rect 35160 -11342 35257 -11326
rect 35657 -10558 35754 -10542
rect 35657 -11326 35704 -10558
rect 35738 -11326 35754 -10558
rect 35657 -11342 35754 -11326
rect 35796 -10558 35893 -10542
rect 35796 -11326 35812 -10558
rect 35846 -11326 35893 -10558
rect 35796 -11342 35893 -11326
rect 36293 -10558 36390 -10542
rect 36293 -11326 36340 -10558
rect 36374 -11326 36390 -10558
rect 36293 -11342 36390 -11326
rect 36760 -10032 36857 -10016
rect 36760 -10200 36776 -10032
rect 36810 -10200 36857 -10032
rect 36760 -10216 36857 -10200
rect 37257 -10032 37354 -10016
rect 37257 -10200 37304 -10032
rect 37338 -10200 37354 -10032
rect 37257 -10216 37354 -10200
rect 37396 -10032 37493 -10016
rect 37396 -10200 37412 -10032
rect 37446 -10200 37493 -10032
rect 37396 -10216 37493 -10200
rect 37893 -10032 37990 -10016
rect 37893 -10200 37940 -10032
rect 37974 -10200 37990 -10032
rect 37893 -10216 37990 -10200
rect 36760 -10558 36857 -10542
rect 36760 -11326 36776 -10558
rect 36810 -11326 36857 -10558
rect 36760 -11342 36857 -11326
rect 37257 -10558 37354 -10542
rect 37257 -11326 37304 -10558
rect 37338 -11326 37354 -10558
rect 37257 -11342 37354 -11326
rect 37396 -10558 37493 -10542
rect 37396 -11326 37412 -10558
rect 37446 -11326 37493 -10558
rect 37396 -11342 37493 -11326
rect 37893 -10558 37990 -10542
rect 37893 -11326 37940 -10558
rect 37974 -11326 37990 -10558
rect 37893 -11342 37990 -11326
rect -40 -11832 57 -11816
rect -40 -12000 -24 -11832
rect 10 -12000 57 -11832
rect -40 -12016 57 -12000
rect 457 -11832 554 -11816
rect 457 -12000 504 -11832
rect 538 -12000 554 -11832
rect 457 -12016 554 -12000
rect 596 -11832 693 -11816
rect 596 -12000 612 -11832
rect 646 -12000 693 -11832
rect 596 -12016 693 -12000
rect 1093 -11832 1190 -11816
rect 1093 -12000 1140 -11832
rect 1174 -12000 1190 -11832
rect 1093 -12016 1190 -12000
rect -40 -12358 57 -12342
rect -40 -13126 -24 -12358
rect 10 -13126 57 -12358
rect -40 -13142 57 -13126
rect 457 -12358 554 -12342
rect 457 -13126 504 -12358
rect 538 -13126 554 -12358
rect 457 -13142 554 -13126
rect 596 -12358 693 -12342
rect 596 -13126 612 -12358
rect 646 -13126 693 -12358
rect 596 -13142 693 -13126
rect 1093 -12358 1190 -12342
rect 1093 -13126 1140 -12358
rect 1174 -13126 1190 -12358
rect 1093 -13142 1190 -13126
rect 1560 -11832 1657 -11816
rect 1560 -12000 1576 -11832
rect 1610 -12000 1657 -11832
rect 1560 -12016 1657 -12000
rect 2057 -11832 2154 -11816
rect 2057 -12000 2104 -11832
rect 2138 -12000 2154 -11832
rect 2057 -12016 2154 -12000
rect 2196 -11832 2293 -11816
rect 2196 -12000 2212 -11832
rect 2246 -12000 2293 -11832
rect 2196 -12016 2293 -12000
rect 2693 -11832 2790 -11816
rect 2693 -12000 2740 -11832
rect 2774 -12000 2790 -11832
rect 2693 -12016 2790 -12000
rect 1560 -12358 1657 -12342
rect 1560 -13126 1576 -12358
rect 1610 -13126 1657 -12358
rect 1560 -13142 1657 -13126
rect 2057 -12358 2154 -12342
rect 2057 -13126 2104 -12358
rect 2138 -13126 2154 -12358
rect 2057 -13142 2154 -13126
rect 2196 -12358 2293 -12342
rect 2196 -13126 2212 -12358
rect 2246 -13126 2293 -12358
rect 2196 -13142 2293 -13126
rect 2693 -12358 2790 -12342
rect 2693 -13126 2740 -12358
rect 2774 -13126 2790 -12358
rect 2693 -13142 2790 -13126
rect 3160 -11832 3257 -11816
rect 3160 -12000 3176 -11832
rect 3210 -12000 3257 -11832
rect 3160 -12016 3257 -12000
rect 3657 -11832 3754 -11816
rect 3657 -12000 3704 -11832
rect 3738 -12000 3754 -11832
rect 3657 -12016 3754 -12000
rect 3796 -11832 3893 -11816
rect 3796 -12000 3812 -11832
rect 3846 -12000 3893 -11832
rect 3796 -12016 3893 -12000
rect 4293 -11832 4390 -11816
rect 4293 -12000 4340 -11832
rect 4374 -12000 4390 -11832
rect 4293 -12016 4390 -12000
rect 3160 -12358 3257 -12342
rect 3160 -13126 3176 -12358
rect 3210 -13126 3257 -12358
rect 3160 -13142 3257 -13126
rect 3657 -12358 3754 -12342
rect 3657 -13126 3704 -12358
rect 3738 -13126 3754 -12358
rect 3657 -13142 3754 -13126
rect 3796 -12358 3893 -12342
rect 3796 -13126 3812 -12358
rect 3846 -13126 3893 -12358
rect 3796 -13142 3893 -13126
rect 4293 -12358 4390 -12342
rect 4293 -13126 4340 -12358
rect 4374 -13126 4390 -12358
rect 4293 -13142 4390 -13126
rect 4760 -11832 4857 -11816
rect 4760 -12000 4776 -11832
rect 4810 -12000 4857 -11832
rect 4760 -12016 4857 -12000
rect 5257 -11832 5354 -11816
rect 5257 -12000 5304 -11832
rect 5338 -12000 5354 -11832
rect 5257 -12016 5354 -12000
rect 5396 -11832 5493 -11816
rect 5396 -12000 5412 -11832
rect 5446 -12000 5493 -11832
rect 5396 -12016 5493 -12000
rect 5893 -11832 5990 -11816
rect 5893 -12000 5940 -11832
rect 5974 -12000 5990 -11832
rect 5893 -12016 5990 -12000
rect 4760 -12358 4857 -12342
rect 4760 -13126 4776 -12358
rect 4810 -13126 4857 -12358
rect 4760 -13142 4857 -13126
rect 5257 -12358 5354 -12342
rect 5257 -13126 5304 -12358
rect 5338 -13126 5354 -12358
rect 5257 -13142 5354 -13126
rect 5396 -12358 5493 -12342
rect 5396 -13126 5412 -12358
rect 5446 -13126 5493 -12358
rect 5396 -13142 5493 -13126
rect 5893 -12358 5990 -12342
rect 5893 -13126 5940 -12358
rect 5974 -13126 5990 -12358
rect 5893 -13142 5990 -13126
rect 6360 -11832 6457 -11816
rect 6360 -12000 6376 -11832
rect 6410 -12000 6457 -11832
rect 6360 -12016 6457 -12000
rect 6857 -11832 6954 -11816
rect 6857 -12000 6904 -11832
rect 6938 -12000 6954 -11832
rect 6857 -12016 6954 -12000
rect 6996 -11832 7093 -11816
rect 6996 -12000 7012 -11832
rect 7046 -12000 7093 -11832
rect 6996 -12016 7093 -12000
rect 7493 -11832 7590 -11816
rect 7493 -12000 7540 -11832
rect 7574 -12000 7590 -11832
rect 7493 -12016 7590 -12000
rect 6360 -12358 6457 -12342
rect 6360 -13126 6376 -12358
rect 6410 -13126 6457 -12358
rect 6360 -13142 6457 -13126
rect 6857 -12358 6954 -12342
rect 6857 -13126 6904 -12358
rect 6938 -13126 6954 -12358
rect 6857 -13142 6954 -13126
rect 6996 -12358 7093 -12342
rect 6996 -13126 7012 -12358
rect 7046 -13126 7093 -12358
rect 6996 -13142 7093 -13126
rect 7493 -12358 7590 -12342
rect 7493 -13126 7540 -12358
rect 7574 -13126 7590 -12358
rect 7493 -13142 7590 -13126
rect 7960 -11832 8057 -11816
rect 7960 -12000 7976 -11832
rect 8010 -12000 8057 -11832
rect 7960 -12016 8057 -12000
rect 8457 -11832 8554 -11816
rect 8457 -12000 8504 -11832
rect 8538 -12000 8554 -11832
rect 8457 -12016 8554 -12000
rect 8596 -11832 8693 -11816
rect 8596 -12000 8612 -11832
rect 8646 -12000 8693 -11832
rect 8596 -12016 8693 -12000
rect 9093 -11832 9190 -11816
rect 9093 -12000 9140 -11832
rect 9174 -12000 9190 -11832
rect 9093 -12016 9190 -12000
rect 7960 -12358 8057 -12342
rect 7960 -13126 7976 -12358
rect 8010 -13126 8057 -12358
rect 7960 -13142 8057 -13126
rect 8457 -12358 8554 -12342
rect 8457 -13126 8504 -12358
rect 8538 -13126 8554 -12358
rect 8457 -13142 8554 -13126
rect 8596 -12358 8693 -12342
rect 8596 -13126 8612 -12358
rect 8646 -13126 8693 -12358
rect 8596 -13142 8693 -13126
rect 9093 -12358 9190 -12342
rect 9093 -13126 9140 -12358
rect 9174 -13126 9190 -12358
rect 9093 -13142 9190 -13126
rect 9560 -11832 9657 -11816
rect 9560 -12000 9576 -11832
rect 9610 -12000 9657 -11832
rect 9560 -12016 9657 -12000
rect 10057 -11832 10154 -11816
rect 10057 -12000 10104 -11832
rect 10138 -12000 10154 -11832
rect 10057 -12016 10154 -12000
rect 10196 -11832 10293 -11816
rect 10196 -12000 10212 -11832
rect 10246 -12000 10293 -11832
rect 10196 -12016 10293 -12000
rect 10693 -11832 10790 -11816
rect 10693 -12000 10740 -11832
rect 10774 -12000 10790 -11832
rect 10693 -12016 10790 -12000
rect 9560 -12358 9657 -12342
rect 9560 -13126 9576 -12358
rect 9610 -13126 9657 -12358
rect 9560 -13142 9657 -13126
rect 10057 -12358 10154 -12342
rect 10057 -13126 10104 -12358
rect 10138 -13126 10154 -12358
rect 10057 -13142 10154 -13126
rect 10196 -12358 10293 -12342
rect 10196 -13126 10212 -12358
rect 10246 -13126 10293 -12358
rect 10196 -13142 10293 -13126
rect 10693 -12358 10790 -12342
rect 10693 -13126 10740 -12358
rect 10774 -13126 10790 -12358
rect 10693 -13142 10790 -13126
rect 11160 -11832 11257 -11816
rect 11160 -12000 11176 -11832
rect 11210 -12000 11257 -11832
rect 11160 -12016 11257 -12000
rect 11657 -11832 11754 -11816
rect 11657 -12000 11704 -11832
rect 11738 -12000 11754 -11832
rect 11657 -12016 11754 -12000
rect 11796 -11832 11893 -11816
rect 11796 -12000 11812 -11832
rect 11846 -12000 11893 -11832
rect 11796 -12016 11893 -12000
rect 12293 -11832 12390 -11816
rect 12293 -12000 12340 -11832
rect 12374 -12000 12390 -11832
rect 12293 -12016 12390 -12000
rect 11160 -12358 11257 -12342
rect 11160 -13126 11176 -12358
rect 11210 -13126 11257 -12358
rect 11160 -13142 11257 -13126
rect 11657 -12358 11754 -12342
rect 11657 -13126 11704 -12358
rect 11738 -13126 11754 -12358
rect 11657 -13142 11754 -13126
rect 11796 -12358 11893 -12342
rect 11796 -13126 11812 -12358
rect 11846 -13126 11893 -12358
rect 11796 -13142 11893 -13126
rect 12293 -12358 12390 -12342
rect 12293 -13126 12340 -12358
rect 12374 -13126 12390 -12358
rect 12293 -13142 12390 -13126
rect 12760 -11832 12857 -11816
rect 12760 -12000 12776 -11832
rect 12810 -12000 12857 -11832
rect 12760 -12016 12857 -12000
rect 13257 -11832 13354 -11816
rect 13257 -12000 13304 -11832
rect 13338 -12000 13354 -11832
rect 13257 -12016 13354 -12000
rect 13396 -11832 13493 -11816
rect 13396 -12000 13412 -11832
rect 13446 -12000 13493 -11832
rect 13396 -12016 13493 -12000
rect 13893 -11832 13990 -11816
rect 13893 -12000 13940 -11832
rect 13974 -12000 13990 -11832
rect 13893 -12016 13990 -12000
rect 12760 -12358 12857 -12342
rect 12760 -13126 12776 -12358
rect 12810 -13126 12857 -12358
rect 12760 -13142 12857 -13126
rect 13257 -12358 13354 -12342
rect 13257 -13126 13304 -12358
rect 13338 -13126 13354 -12358
rect 13257 -13142 13354 -13126
rect 13396 -12358 13493 -12342
rect 13396 -13126 13412 -12358
rect 13446 -13126 13493 -12358
rect 13396 -13142 13493 -13126
rect 13893 -12358 13990 -12342
rect 13893 -13126 13940 -12358
rect 13974 -13126 13990 -12358
rect 13893 -13142 13990 -13126
rect 14360 -11832 14457 -11816
rect 14360 -12000 14376 -11832
rect 14410 -12000 14457 -11832
rect 14360 -12016 14457 -12000
rect 14857 -11832 14954 -11816
rect 14857 -12000 14904 -11832
rect 14938 -12000 14954 -11832
rect 14857 -12016 14954 -12000
rect 14996 -11832 15093 -11816
rect 14996 -12000 15012 -11832
rect 15046 -12000 15093 -11832
rect 14996 -12016 15093 -12000
rect 15493 -11832 15590 -11816
rect 15493 -12000 15540 -11832
rect 15574 -12000 15590 -11832
rect 15493 -12016 15590 -12000
rect 14360 -12358 14457 -12342
rect 14360 -13126 14376 -12358
rect 14410 -13126 14457 -12358
rect 14360 -13142 14457 -13126
rect 14857 -12358 14954 -12342
rect 14857 -13126 14904 -12358
rect 14938 -13126 14954 -12358
rect 14857 -13142 14954 -13126
rect 14996 -12358 15093 -12342
rect 14996 -13126 15012 -12358
rect 15046 -13126 15093 -12358
rect 14996 -13142 15093 -13126
rect 15493 -12358 15590 -12342
rect 15493 -13126 15540 -12358
rect 15574 -13126 15590 -12358
rect 15493 -13142 15590 -13126
rect 15960 -11832 16057 -11816
rect 15960 -12000 15976 -11832
rect 16010 -12000 16057 -11832
rect 15960 -12016 16057 -12000
rect 16457 -11832 16554 -11816
rect 16457 -12000 16504 -11832
rect 16538 -12000 16554 -11832
rect 16457 -12016 16554 -12000
rect 16596 -11832 16693 -11816
rect 16596 -12000 16612 -11832
rect 16646 -12000 16693 -11832
rect 16596 -12016 16693 -12000
rect 17093 -11832 17190 -11816
rect 17093 -12000 17140 -11832
rect 17174 -12000 17190 -11832
rect 17093 -12016 17190 -12000
rect 15960 -12358 16057 -12342
rect 15960 -13126 15976 -12358
rect 16010 -13126 16057 -12358
rect 15960 -13142 16057 -13126
rect 16457 -12358 16554 -12342
rect 16457 -13126 16504 -12358
rect 16538 -13126 16554 -12358
rect 16457 -13142 16554 -13126
rect 16596 -12358 16693 -12342
rect 16596 -13126 16612 -12358
rect 16646 -13126 16693 -12358
rect 16596 -13142 16693 -13126
rect 17093 -12358 17190 -12342
rect 17093 -13126 17140 -12358
rect 17174 -13126 17190 -12358
rect 17093 -13142 17190 -13126
rect 17560 -11832 17657 -11816
rect 17560 -12000 17576 -11832
rect 17610 -12000 17657 -11832
rect 17560 -12016 17657 -12000
rect 18057 -11832 18154 -11816
rect 18057 -12000 18104 -11832
rect 18138 -12000 18154 -11832
rect 18057 -12016 18154 -12000
rect 18196 -11832 18293 -11816
rect 18196 -12000 18212 -11832
rect 18246 -12000 18293 -11832
rect 18196 -12016 18293 -12000
rect 18693 -11832 18790 -11816
rect 18693 -12000 18740 -11832
rect 18774 -12000 18790 -11832
rect 18693 -12016 18790 -12000
rect 17560 -12358 17657 -12342
rect 17560 -13126 17576 -12358
rect 17610 -13126 17657 -12358
rect 17560 -13142 17657 -13126
rect 18057 -12358 18154 -12342
rect 18057 -13126 18104 -12358
rect 18138 -13126 18154 -12358
rect 18057 -13142 18154 -13126
rect 18196 -12358 18293 -12342
rect 18196 -13126 18212 -12358
rect 18246 -13126 18293 -12358
rect 18196 -13142 18293 -13126
rect 18693 -12358 18790 -12342
rect 18693 -13126 18740 -12358
rect 18774 -13126 18790 -12358
rect 18693 -13142 18790 -13126
rect 19160 -11832 19257 -11816
rect 19160 -12000 19176 -11832
rect 19210 -12000 19257 -11832
rect 19160 -12016 19257 -12000
rect 19657 -11832 19754 -11816
rect 19657 -12000 19704 -11832
rect 19738 -12000 19754 -11832
rect 19657 -12016 19754 -12000
rect 19796 -11832 19893 -11816
rect 19796 -12000 19812 -11832
rect 19846 -12000 19893 -11832
rect 19796 -12016 19893 -12000
rect 20293 -11832 20390 -11816
rect 20293 -12000 20340 -11832
rect 20374 -12000 20390 -11832
rect 20293 -12016 20390 -12000
rect 19160 -12358 19257 -12342
rect 19160 -13126 19176 -12358
rect 19210 -13126 19257 -12358
rect 19160 -13142 19257 -13126
rect 19657 -12358 19754 -12342
rect 19657 -13126 19704 -12358
rect 19738 -13126 19754 -12358
rect 19657 -13142 19754 -13126
rect 19796 -12358 19893 -12342
rect 19796 -13126 19812 -12358
rect 19846 -13126 19893 -12358
rect 19796 -13142 19893 -13126
rect 20293 -12358 20390 -12342
rect 20293 -13126 20340 -12358
rect 20374 -13126 20390 -12358
rect 20293 -13142 20390 -13126
rect 20760 -11832 20857 -11816
rect 20760 -12000 20776 -11832
rect 20810 -12000 20857 -11832
rect 20760 -12016 20857 -12000
rect 21257 -11832 21354 -11816
rect 21257 -12000 21304 -11832
rect 21338 -12000 21354 -11832
rect 21257 -12016 21354 -12000
rect 21396 -11832 21493 -11816
rect 21396 -12000 21412 -11832
rect 21446 -12000 21493 -11832
rect 21396 -12016 21493 -12000
rect 21893 -11832 21990 -11816
rect 21893 -12000 21940 -11832
rect 21974 -12000 21990 -11832
rect 21893 -12016 21990 -12000
rect 20760 -12358 20857 -12342
rect 20760 -13126 20776 -12358
rect 20810 -13126 20857 -12358
rect 20760 -13142 20857 -13126
rect 21257 -12358 21354 -12342
rect 21257 -13126 21304 -12358
rect 21338 -13126 21354 -12358
rect 21257 -13142 21354 -13126
rect 21396 -12358 21493 -12342
rect 21396 -13126 21412 -12358
rect 21446 -13126 21493 -12358
rect 21396 -13142 21493 -13126
rect 21893 -12358 21990 -12342
rect 21893 -13126 21940 -12358
rect 21974 -13126 21990 -12358
rect 21893 -13142 21990 -13126
rect 22360 -11832 22457 -11816
rect 22360 -12000 22376 -11832
rect 22410 -12000 22457 -11832
rect 22360 -12016 22457 -12000
rect 22857 -11832 22954 -11816
rect 22857 -12000 22904 -11832
rect 22938 -12000 22954 -11832
rect 22857 -12016 22954 -12000
rect 22996 -11832 23093 -11816
rect 22996 -12000 23012 -11832
rect 23046 -12000 23093 -11832
rect 22996 -12016 23093 -12000
rect 23493 -11832 23590 -11816
rect 23493 -12000 23540 -11832
rect 23574 -12000 23590 -11832
rect 23493 -12016 23590 -12000
rect 22360 -12358 22457 -12342
rect 22360 -13126 22376 -12358
rect 22410 -13126 22457 -12358
rect 22360 -13142 22457 -13126
rect 22857 -12358 22954 -12342
rect 22857 -13126 22904 -12358
rect 22938 -13126 22954 -12358
rect 22857 -13142 22954 -13126
rect 22996 -12358 23093 -12342
rect 22996 -13126 23012 -12358
rect 23046 -13126 23093 -12358
rect 22996 -13142 23093 -13126
rect 23493 -12358 23590 -12342
rect 23493 -13126 23540 -12358
rect 23574 -13126 23590 -12358
rect 23493 -13142 23590 -13126
rect 23960 -11832 24057 -11816
rect 23960 -12000 23976 -11832
rect 24010 -12000 24057 -11832
rect 23960 -12016 24057 -12000
rect 24457 -11832 24554 -11816
rect 24457 -12000 24504 -11832
rect 24538 -12000 24554 -11832
rect 24457 -12016 24554 -12000
rect 24596 -11832 24693 -11816
rect 24596 -12000 24612 -11832
rect 24646 -12000 24693 -11832
rect 24596 -12016 24693 -12000
rect 25093 -11832 25190 -11816
rect 25093 -12000 25140 -11832
rect 25174 -12000 25190 -11832
rect 25093 -12016 25190 -12000
rect 23960 -12358 24057 -12342
rect 23960 -13126 23976 -12358
rect 24010 -13126 24057 -12358
rect 23960 -13142 24057 -13126
rect 24457 -12358 24554 -12342
rect 24457 -13126 24504 -12358
rect 24538 -13126 24554 -12358
rect 24457 -13142 24554 -13126
rect 24596 -12358 24693 -12342
rect 24596 -13126 24612 -12358
rect 24646 -13126 24693 -12358
rect 24596 -13142 24693 -13126
rect 25093 -12358 25190 -12342
rect 25093 -13126 25140 -12358
rect 25174 -13126 25190 -12358
rect 25093 -13142 25190 -13126
rect 25560 -11832 25657 -11816
rect 25560 -12000 25576 -11832
rect 25610 -12000 25657 -11832
rect 25560 -12016 25657 -12000
rect 26057 -11832 26154 -11816
rect 26057 -12000 26104 -11832
rect 26138 -12000 26154 -11832
rect 26057 -12016 26154 -12000
rect 26196 -11832 26293 -11816
rect 26196 -12000 26212 -11832
rect 26246 -12000 26293 -11832
rect 26196 -12016 26293 -12000
rect 26693 -11832 26790 -11816
rect 26693 -12000 26740 -11832
rect 26774 -12000 26790 -11832
rect 26693 -12016 26790 -12000
rect 25560 -12358 25657 -12342
rect 25560 -13126 25576 -12358
rect 25610 -13126 25657 -12358
rect 25560 -13142 25657 -13126
rect 26057 -12358 26154 -12342
rect 26057 -13126 26104 -12358
rect 26138 -13126 26154 -12358
rect 26057 -13142 26154 -13126
rect 26196 -12358 26293 -12342
rect 26196 -13126 26212 -12358
rect 26246 -13126 26293 -12358
rect 26196 -13142 26293 -13126
rect 26693 -12358 26790 -12342
rect 26693 -13126 26740 -12358
rect 26774 -13126 26790 -12358
rect 26693 -13142 26790 -13126
rect 27160 -11832 27257 -11816
rect 27160 -12000 27176 -11832
rect 27210 -12000 27257 -11832
rect 27160 -12016 27257 -12000
rect 27657 -11832 27754 -11816
rect 27657 -12000 27704 -11832
rect 27738 -12000 27754 -11832
rect 27657 -12016 27754 -12000
rect 27796 -11832 27893 -11816
rect 27796 -12000 27812 -11832
rect 27846 -12000 27893 -11832
rect 27796 -12016 27893 -12000
rect 28293 -11832 28390 -11816
rect 28293 -12000 28340 -11832
rect 28374 -12000 28390 -11832
rect 28293 -12016 28390 -12000
rect 27160 -12358 27257 -12342
rect 27160 -13126 27176 -12358
rect 27210 -13126 27257 -12358
rect 27160 -13142 27257 -13126
rect 27657 -12358 27754 -12342
rect 27657 -13126 27704 -12358
rect 27738 -13126 27754 -12358
rect 27657 -13142 27754 -13126
rect 27796 -12358 27893 -12342
rect 27796 -13126 27812 -12358
rect 27846 -13126 27893 -12358
rect 27796 -13142 27893 -13126
rect 28293 -12358 28390 -12342
rect 28293 -13126 28340 -12358
rect 28374 -13126 28390 -12358
rect 28293 -13142 28390 -13126
rect 28760 -11832 28857 -11816
rect 28760 -12000 28776 -11832
rect 28810 -12000 28857 -11832
rect 28760 -12016 28857 -12000
rect 29257 -11832 29354 -11816
rect 29257 -12000 29304 -11832
rect 29338 -12000 29354 -11832
rect 29257 -12016 29354 -12000
rect 29396 -11832 29493 -11816
rect 29396 -12000 29412 -11832
rect 29446 -12000 29493 -11832
rect 29396 -12016 29493 -12000
rect 29893 -11832 29990 -11816
rect 29893 -12000 29940 -11832
rect 29974 -12000 29990 -11832
rect 29893 -12016 29990 -12000
rect 28760 -12358 28857 -12342
rect 28760 -13126 28776 -12358
rect 28810 -13126 28857 -12358
rect 28760 -13142 28857 -13126
rect 29257 -12358 29354 -12342
rect 29257 -13126 29304 -12358
rect 29338 -13126 29354 -12358
rect 29257 -13142 29354 -13126
rect 29396 -12358 29493 -12342
rect 29396 -13126 29412 -12358
rect 29446 -13126 29493 -12358
rect 29396 -13142 29493 -13126
rect 29893 -12358 29990 -12342
rect 29893 -13126 29940 -12358
rect 29974 -13126 29990 -12358
rect 29893 -13142 29990 -13126
rect 30360 -11832 30457 -11816
rect 30360 -12000 30376 -11832
rect 30410 -12000 30457 -11832
rect 30360 -12016 30457 -12000
rect 30857 -11832 30954 -11816
rect 30857 -12000 30904 -11832
rect 30938 -12000 30954 -11832
rect 30857 -12016 30954 -12000
rect 30996 -11832 31093 -11816
rect 30996 -12000 31012 -11832
rect 31046 -12000 31093 -11832
rect 30996 -12016 31093 -12000
rect 31493 -11832 31590 -11816
rect 31493 -12000 31540 -11832
rect 31574 -12000 31590 -11832
rect 31493 -12016 31590 -12000
rect 30360 -12358 30457 -12342
rect 30360 -13126 30376 -12358
rect 30410 -13126 30457 -12358
rect 30360 -13142 30457 -13126
rect 30857 -12358 30954 -12342
rect 30857 -13126 30904 -12358
rect 30938 -13126 30954 -12358
rect 30857 -13142 30954 -13126
rect 30996 -12358 31093 -12342
rect 30996 -13126 31012 -12358
rect 31046 -13126 31093 -12358
rect 30996 -13142 31093 -13126
rect 31493 -12358 31590 -12342
rect 31493 -13126 31540 -12358
rect 31574 -13126 31590 -12358
rect 31493 -13142 31590 -13126
rect 31960 -11832 32057 -11816
rect 31960 -12000 31976 -11832
rect 32010 -12000 32057 -11832
rect 31960 -12016 32057 -12000
rect 32457 -11832 32554 -11816
rect 32457 -12000 32504 -11832
rect 32538 -12000 32554 -11832
rect 32457 -12016 32554 -12000
rect 32596 -11832 32693 -11816
rect 32596 -12000 32612 -11832
rect 32646 -12000 32693 -11832
rect 32596 -12016 32693 -12000
rect 33093 -11832 33190 -11816
rect 33093 -12000 33140 -11832
rect 33174 -12000 33190 -11832
rect 33093 -12016 33190 -12000
rect 31960 -12358 32057 -12342
rect 31960 -13126 31976 -12358
rect 32010 -13126 32057 -12358
rect 31960 -13142 32057 -13126
rect 32457 -12358 32554 -12342
rect 32457 -13126 32504 -12358
rect 32538 -13126 32554 -12358
rect 32457 -13142 32554 -13126
rect 32596 -12358 32693 -12342
rect 32596 -13126 32612 -12358
rect 32646 -13126 32693 -12358
rect 32596 -13142 32693 -13126
rect 33093 -12358 33190 -12342
rect 33093 -13126 33140 -12358
rect 33174 -13126 33190 -12358
rect 33093 -13142 33190 -13126
rect 33560 -11832 33657 -11816
rect 33560 -12000 33576 -11832
rect 33610 -12000 33657 -11832
rect 33560 -12016 33657 -12000
rect 34057 -11832 34154 -11816
rect 34057 -12000 34104 -11832
rect 34138 -12000 34154 -11832
rect 34057 -12016 34154 -12000
rect 34196 -11832 34293 -11816
rect 34196 -12000 34212 -11832
rect 34246 -12000 34293 -11832
rect 34196 -12016 34293 -12000
rect 34693 -11832 34790 -11816
rect 34693 -12000 34740 -11832
rect 34774 -12000 34790 -11832
rect 34693 -12016 34790 -12000
rect 33560 -12358 33657 -12342
rect 33560 -13126 33576 -12358
rect 33610 -13126 33657 -12358
rect 33560 -13142 33657 -13126
rect 34057 -12358 34154 -12342
rect 34057 -13126 34104 -12358
rect 34138 -13126 34154 -12358
rect 34057 -13142 34154 -13126
rect 34196 -12358 34293 -12342
rect 34196 -13126 34212 -12358
rect 34246 -13126 34293 -12358
rect 34196 -13142 34293 -13126
rect 34693 -12358 34790 -12342
rect 34693 -13126 34740 -12358
rect 34774 -13126 34790 -12358
rect 34693 -13142 34790 -13126
rect 35160 -11832 35257 -11816
rect 35160 -12000 35176 -11832
rect 35210 -12000 35257 -11832
rect 35160 -12016 35257 -12000
rect 35657 -11832 35754 -11816
rect 35657 -12000 35704 -11832
rect 35738 -12000 35754 -11832
rect 35657 -12016 35754 -12000
rect 35796 -11832 35893 -11816
rect 35796 -12000 35812 -11832
rect 35846 -12000 35893 -11832
rect 35796 -12016 35893 -12000
rect 36293 -11832 36390 -11816
rect 36293 -12000 36340 -11832
rect 36374 -12000 36390 -11832
rect 36293 -12016 36390 -12000
rect 35160 -12358 35257 -12342
rect 35160 -13126 35176 -12358
rect 35210 -13126 35257 -12358
rect 35160 -13142 35257 -13126
rect 35657 -12358 35754 -12342
rect 35657 -13126 35704 -12358
rect 35738 -13126 35754 -12358
rect 35657 -13142 35754 -13126
rect 35796 -12358 35893 -12342
rect 35796 -13126 35812 -12358
rect 35846 -13126 35893 -12358
rect 35796 -13142 35893 -13126
rect 36293 -12358 36390 -12342
rect 36293 -13126 36340 -12358
rect 36374 -13126 36390 -12358
rect 36293 -13142 36390 -13126
rect 36760 -11832 36857 -11816
rect 36760 -12000 36776 -11832
rect 36810 -12000 36857 -11832
rect 36760 -12016 36857 -12000
rect 37257 -11832 37354 -11816
rect 37257 -12000 37304 -11832
rect 37338 -12000 37354 -11832
rect 37257 -12016 37354 -12000
rect 37396 -11832 37493 -11816
rect 37396 -12000 37412 -11832
rect 37446 -12000 37493 -11832
rect 37396 -12016 37493 -12000
rect 37893 -11832 37990 -11816
rect 37893 -12000 37940 -11832
rect 37974 -12000 37990 -11832
rect 37893 -12016 37990 -12000
rect 36760 -12358 36857 -12342
rect 36760 -13126 36776 -12358
rect 36810 -13126 36857 -12358
rect 36760 -13142 36857 -13126
rect 37257 -12358 37354 -12342
rect 37257 -13126 37304 -12358
rect 37338 -13126 37354 -12358
rect 37257 -13142 37354 -13126
rect 37396 -12358 37493 -12342
rect 37396 -13126 37412 -12358
rect 37446 -13126 37493 -12358
rect 37396 -13142 37493 -13126
rect 37893 -12358 37990 -12342
rect 37893 -13126 37940 -12358
rect 37974 -13126 37990 -12358
rect 37893 -13142 37990 -13126
rect -40 -13632 57 -13616
rect -40 -13800 -24 -13632
rect 10 -13800 57 -13632
rect -40 -13816 57 -13800
rect 457 -13632 554 -13616
rect 457 -13800 504 -13632
rect 538 -13800 554 -13632
rect 457 -13816 554 -13800
rect 596 -13632 693 -13616
rect 596 -13800 612 -13632
rect 646 -13800 693 -13632
rect 596 -13816 693 -13800
rect 1093 -13632 1190 -13616
rect 1093 -13800 1140 -13632
rect 1174 -13800 1190 -13632
rect 1093 -13816 1190 -13800
rect -40 -14158 57 -14142
rect -40 -14926 -24 -14158
rect 10 -14926 57 -14158
rect -40 -14942 57 -14926
rect 457 -14158 554 -14142
rect 457 -14926 504 -14158
rect 538 -14926 554 -14158
rect 457 -14942 554 -14926
rect 596 -14158 693 -14142
rect 596 -14926 612 -14158
rect 646 -14926 693 -14158
rect 596 -14942 693 -14926
rect 1093 -14158 1190 -14142
rect 1093 -14926 1140 -14158
rect 1174 -14926 1190 -14158
rect 1093 -14942 1190 -14926
rect 1560 -13632 1657 -13616
rect 1560 -13800 1576 -13632
rect 1610 -13800 1657 -13632
rect 1560 -13816 1657 -13800
rect 2057 -13632 2154 -13616
rect 2057 -13800 2104 -13632
rect 2138 -13800 2154 -13632
rect 2057 -13816 2154 -13800
rect 2196 -13632 2293 -13616
rect 2196 -13800 2212 -13632
rect 2246 -13800 2293 -13632
rect 2196 -13816 2293 -13800
rect 2693 -13632 2790 -13616
rect 2693 -13800 2740 -13632
rect 2774 -13800 2790 -13632
rect 2693 -13816 2790 -13800
rect 1560 -14158 1657 -14142
rect 1560 -14926 1576 -14158
rect 1610 -14926 1657 -14158
rect 1560 -14942 1657 -14926
rect 2057 -14158 2154 -14142
rect 2057 -14926 2104 -14158
rect 2138 -14926 2154 -14158
rect 2057 -14942 2154 -14926
rect 2196 -14158 2293 -14142
rect 2196 -14926 2212 -14158
rect 2246 -14926 2293 -14158
rect 2196 -14942 2293 -14926
rect 2693 -14158 2790 -14142
rect 2693 -14926 2740 -14158
rect 2774 -14926 2790 -14158
rect 2693 -14942 2790 -14926
rect 3160 -13632 3257 -13616
rect 3160 -13800 3176 -13632
rect 3210 -13800 3257 -13632
rect 3160 -13816 3257 -13800
rect 3657 -13632 3754 -13616
rect 3657 -13800 3704 -13632
rect 3738 -13800 3754 -13632
rect 3657 -13816 3754 -13800
rect 3796 -13632 3893 -13616
rect 3796 -13800 3812 -13632
rect 3846 -13800 3893 -13632
rect 3796 -13816 3893 -13800
rect 4293 -13632 4390 -13616
rect 4293 -13800 4340 -13632
rect 4374 -13800 4390 -13632
rect 4293 -13816 4390 -13800
rect 3160 -14158 3257 -14142
rect 3160 -14926 3176 -14158
rect 3210 -14926 3257 -14158
rect 3160 -14942 3257 -14926
rect 3657 -14158 3754 -14142
rect 3657 -14926 3704 -14158
rect 3738 -14926 3754 -14158
rect 3657 -14942 3754 -14926
rect 3796 -14158 3893 -14142
rect 3796 -14926 3812 -14158
rect 3846 -14926 3893 -14158
rect 3796 -14942 3893 -14926
rect 4293 -14158 4390 -14142
rect 4293 -14926 4340 -14158
rect 4374 -14926 4390 -14158
rect 4293 -14942 4390 -14926
rect 4760 -13632 4857 -13616
rect 4760 -13800 4776 -13632
rect 4810 -13800 4857 -13632
rect 4760 -13816 4857 -13800
rect 5257 -13632 5354 -13616
rect 5257 -13800 5304 -13632
rect 5338 -13800 5354 -13632
rect 5257 -13816 5354 -13800
rect 5396 -13632 5493 -13616
rect 5396 -13800 5412 -13632
rect 5446 -13800 5493 -13632
rect 5396 -13816 5493 -13800
rect 5893 -13632 5990 -13616
rect 5893 -13800 5940 -13632
rect 5974 -13800 5990 -13632
rect 5893 -13816 5990 -13800
rect 4760 -14158 4857 -14142
rect 4760 -14926 4776 -14158
rect 4810 -14926 4857 -14158
rect 4760 -14942 4857 -14926
rect 5257 -14158 5354 -14142
rect 5257 -14926 5304 -14158
rect 5338 -14926 5354 -14158
rect 5257 -14942 5354 -14926
rect 5396 -14158 5493 -14142
rect 5396 -14926 5412 -14158
rect 5446 -14926 5493 -14158
rect 5396 -14942 5493 -14926
rect 5893 -14158 5990 -14142
rect 5893 -14926 5940 -14158
rect 5974 -14926 5990 -14158
rect 5893 -14942 5990 -14926
rect 6360 -13632 6457 -13616
rect 6360 -13800 6376 -13632
rect 6410 -13800 6457 -13632
rect 6360 -13816 6457 -13800
rect 6857 -13632 6954 -13616
rect 6857 -13800 6904 -13632
rect 6938 -13800 6954 -13632
rect 6857 -13816 6954 -13800
rect 6996 -13632 7093 -13616
rect 6996 -13800 7012 -13632
rect 7046 -13800 7093 -13632
rect 6996 -13816 7093 -13800
rect 7493 -13632 7590 -13616
rect 7493 -13800 7540 -13632
rect 7574 -13800 7590 -13632
rect 7493 -13816 7590 -13800
rect 6360 -14158 6457 -14142
rect 6360 -14926 6376 -14158
rect 6410 -14926 6457 -14158
rect 6360 -14942 6457 -14926
rect 6857 -14158 6954 -14142
rect 6857 -14926 6904 -14158
rect 6938 -14926 6954 -14158
rect 6857 -14942 6954 -14926
rect 6996 -14158 7093 -14142
rect 6996 -14926 7012 -14158
rect 7046 -14926 7093 -14158
rect 6996 -14942 7093 -14926
rect 7493 -14158 7590 -14142
rect 7493 -14926 7540 -14158
rect 7574 -14926 7590 -14158
rect 7493 -14942 7590 -14926
rect 7960 -13632 8057 -13616
rect 7960 -13800 7976 -13632
rect 8010 -13800 8057 -13632
rect 7960 -13816 8057 -13800
rect 8457 -13632 8554 -13616
rect 8457 -13800 8504 -13632
rect 8538 -13800 8554 -13632
rect 8457 -13816 8554 -13800
rect 8596 -13632 8693 -13616
rect 8596 -13800 8612 -13632
rect 8646 -13800 8693 -13632
rect 8596 -13816 8693 -13800
rect 9093 -13632 9190 -13616
rect 9093 -13800 9140 -13632
rect 9174 -13800 9190 -13632
rect 9093 -13816 9190 -13800
rect 7960 -14158 8057 -14142
rect 7960 -14926 7976 -14158
rect 8010 -14926 8057 -14158
rect 7960 -14942 8057 -14926
rect 8457 -14158 8554 -14142
rect 8457 -14926 8504 -14158
rect 8538 -14926 8554 -14158
rect 8457 -14942 8554 -14926
rect 8596 -14158 8693 -14142
rect 8596 -14926 8612 -14158
rect 8646 -14926 8693 -14158
rect 8596 -14942 8693 -14926
rect 9093 -14158 9190 -14142
rect 9093 -14926 9140 -14158
rect 9174 -14926 9190 -14158
rect 9093 -14942 9190 -14926
rect 9560 -13632 9657 -13616
rect 9560 -13800 9576 -13632
rect 9610 -13800 9657 -13632
rect 9560 -13816 9657 -13800
rect 10057 -13632 10154 -13616
rect 10057 -13800 10104 -13632
rect 10138 -13800 10154 -13632
rect 10057 -13816 10154 -13800
rect 10196 -13632 10293 -13616
rect 10196 -13800 10212 -13632
rect 10246 -13800 10293 -13632
rect 10196 -13816 10293 -13800
rect 10693 -13632 10790 -13616
rect 10693 -13800 10740 -13632
rect 10774 -13800 10790 -13632
rect 10693 -13816 10790 -13800
rect 9560 -14158 9657 -14142
rect 9560 -14926 9576 -14158
rect 9610 -14926 9657 -14158
rect 9560 -14942 9657 -14926
rect 10057 -14158 10154 -14142
rect 10057 -14926 10104 -14158
rect 10138 -14926 10154 -14158
rect 10057 -14942 10154 -14926
rect 10196 -14158 10293 -14142
rect 10196 -14926 10212 -14158
rect 10246 -14926 10293 -14158
rect 10196 -14942 10293 -14926
rect 10693 -14158 10790 -14142
rect 10693 -14926 10740 -14158
rect 10774 -14926 10790 -14158
rect 10693 -14942 10790 -14926
rect 11160 -13632 11257 -13616
rect 11160 -13800 11176 -13632
rect 11210 -13800 11257 -13632
rect 11160 -13816 11257 -13800
rect 11657 -13632 11754 -13616
rect 11657 -13800 11704 -13632
rect 11738 -13800 11754 -13632
rect 11657 -13816 11754 -13800
rect 11796 -13632 11893 -13616
rect 11796 -13800 11812 -13632
rect 11846 -13800 11893 -13632
rect 11796 -13816 11893 -13800
rect 12293 -13632 12390 -13616
rect 12293 -13800 12340 -13632
rect 12374 -13800 12390 -13632
rect 12293 -13816 12390 -13800
rect 11160 -14158 11257 -14142
rect 11160 -14926 11176 -14158
rect 11210 -14926 11257 -14158
rect 11160 -14942 11257 -14926
rect 11657 -14158 11754 -14142
rect 11657 -14926 11704 -14158
rect 11738 -14926 11754 -14158
rect 11657 -14942 11754 -14926
rect 11796 -14158 11893 -14142
rect 11796 -14926 11812 -14158
rect 11846 -14926 11893 -14158
rect 11796 -14942 11893 -14926
rect 12293 -14158 12390 -14142
rect 12293 -14926 12340 -14158
rect 12374 -14926 12390 -14158
rect 12293 -14942 12390 -14926
rect 12760 -13632 12857 -13616
rect 12760 -13800 12776 -13632
rect 12810 -13800 12857 -13632
rect 12760 -13816 12857 -13800
rect 13257 -13632 13354 -13616
rect 13257 -13800 13304 -13632
rect 13338 -13800 13354 -13632
rect 13257 -13816 13354 -13800
rect 13396 -13632 13493 -13616
rect 13396 -13800 13412 -13632
rect 13446 -13800 13493 -13632
rect 13396 -13816 13493 -13800
rect 13893 -13632 13990 -13616
rect 13893 -13800 13940 -13632
rect 13974 -13800 13990 -13632
rect 13893 -13816 13990 -13800
rect 12760 -14158 12857 -14142
rect 12760 -14926 12776 -14158
rect 12810 -14926 12857 -14158
rect 12760 -14942 12857 -14926
rect 13257 -14158 13354 -14142
rect 13257 -14926 13304 -14158
rect 13338 -14926 13354 -14158
rect 13257 -14942 13354 -14926
rect 13396 -14158 13493 -14142
rect 13396 -14926 13412 -14158
rect 13446 -14926 13493 -14158
rect 13396 -14942 13493 -14926
rect 13893 -14158 13990 -14142
rect 13893 -14926 13940 -14158
rect 13974 -14926 13990 -14158
rect 13893 -14942 13990 -14926
rect 14360 -13632 14457 -13616
rect 14360 -13800 14376 -13632
rect 14410 -13800 14457 -13632
rect 14360 -13816 14457 -13800
rect 14857 -13632 14954 -13616
rect 14857 -13800 14904 -13632
rect 14938 -13800 14954 -13632
rect 14857 -13816 14954 -13800
rect 14996 -13632 15093 -13616
rect 14996 -13800 15012 -13632
rect 15046 -13800 15093 -13632
rect 14996 -13816 15093 -13800
rect 15493 -13632 15590 -13616
rect 15493 -13800 15540 -13632
rect 15574 -13800 15590 -13632
rect 15493 -13816 15590 -13800
rect 14360 -14158 14457 -14142
rect 14360 -14926 14376 -14158
rect 14410 -14926 14457 -14158
rect 14360 -14942 14457 -14926
rect 14857 -14158 14954 -14142
rect 14857 -14926 14904 -14158
rect 14938 -14926 14954 -14158
rect 14857 -14942 14954 -14926
rect 14996 -14158 15093 -14142
rect 14996 -14926 15012 -14158
rect 15046 -14926 15093 -14158
rect 14996 -14942 15093 -14926
rect 15493 -14158 15590 -14142
rect 15493 -14926 15540 -14158
rect 15574 -14926 15590 -14158
rect 15493 -14942 15590 -14926
rect 15960 -13632 16057 -13616
rect 15960 -13800 15976 -13632
rect 16010 -13800 16057 -13632
rect 15960 -13816 16057 -13800
rect 16457 -13632 16554 -13616
rect 16457 -13800 16504 -13632
rect 16538 -13800 16554 -13632
rect 16457 -13816 16554 -13800
rect 16596 -13632 16693 -13616
rect 16596 -13800 16612 -13632
rect 16646 -13800 16693 -13632
rect 16596 -13816 16693 -13800
rect 17093 -13632 17190 -13616
rect 17093 -13800 17140 -13632
rect 17174 -13800 17190 -13632
rect 17093 -13816 17190 -13800
rect 15960 -14158 16057 -14142
rect 15960 -14926 15976 -14158
rect 16010 -14926 16057 -14158
rect 15960 -14942 16057 -14926
rect 16457 -14158 16554 -14142
rect 16457 -14926 16504 -14158
rect 16538 -14926 16554 -14158
rect 16457 -14942 16554 -14926
rect 16596 -14158 16693 -14142
rect 16596 -14926 16612 -14158
rect 16646 -14926 16693 -14158
rect 16596 -14942 16693 -14926
rect 17093 -14158 17190 -14142
rect 17093 -14926 17140 -14158
rect 17174 -14926 17190 -14158
rect 17093 -14942 17190 -14926
rect 17560 -13632 17657 -13616
rect 17560 -13800 17576 -13632
rect 17610 -13800 17657 -13632
rect 17560 -13816 17657 -13800
rect 18057 -13632 18154 -13616
rect 18057 -13800 18104 -13632
rect 18138 -13800 18154 -13632
rect 18057 -13816 18154 -13800
rect 18196 -13632 18293 -13616
rect 18196 -13800 18212 -13632
rect 18246 -13800 18293 -13632
rect 18196 -13816 18293 -13800
rect 18693 -13632 18790 -13616
rect 18693 -13800 18740 -13632
rect 18774 -13800 18790 -13632
rect 18693 -13816 18790 -13800
rect 17560 -14158 17657 -14142
rect 17560 -14926 17576 -14158
rect 17610 -14926 17657 -14158
rect 17560 -14942 17657 -14926
rect 18057 -14158 18154 -14142
rect 18057 -14926 18104 -14158
rect 18138 -14926 18154 -14158
rect 18057 -14942 18154 -14926
rect 18196 -14158 18293 -14142
rect 18196 -14926 18212 -14158
rect 18246 -14926 18293 -14158
rect 18196 -14942 18293 -14926
rect 18693 -14158 18790 -14142
rect 18693 -14926 18740 -14158
rect 18774 -14926 18790 -14158
rect 18693 -14942 18790 -14926
rect 19160 -13632 19257 -13616
rect 19160 -13800 19176 -13632
rect 19210 -13800 19257 -13632
rect 19160 -13816 19257 -13800
rect 19657 -13632 19754 -13616
rect 19657 -13800 19704 -13632
rect 19738 -13800 19754 -13632
rect 19657 -13816 19754 -13800
rect 19796 -13632 19893 -13616
rect 19796 -13800 19812 -13632
rect 19846 -13800 19893 -13632
rect 19796 -13816 19893 -13800
rect 20293 -13632 20390 -13616
rect 20293 -13800 20340 -13632
rect 20374 -13800 20390 -13632
rect 20293 -13816 20390 -13800
rect 19160 -14158 19257 -14142
rect 19160 -14926 19176 -14158
rect 19210 -14926 19257 -14158
rect 19160 -14942 19257 -14926
rect 19657 -14158 19754 -14142
rect 19657 -14926 19704 -14158
rect 19738 -14926 19754 -14158
rect 19657 -14942 19754 -14926
rect 19796 -14158 19893 -14142
rect 19796 -14926 19812 -14158
rect 19846 -14926 19893 -14158
rect 19796 -14942 19893 -14926
rect 20293 -14158 20390 -14142
rect 20293 -14926 20340 -14158
rect 20374 -14926 20390 -14158
rect 20293 -14942 20390 -14926
rect 20760 -13632 20857 -13616
rect 20760 -13800 20776 -13632
rect 20810 -13800 20857 -13632
rect 20760 -13816 20857 -13800
rect 21257 -13632 21354 -13616
rect 21257 -13800 21304 -13632
rect 21338 -13800 21354 -13632
rect 21257 -13816 21354 -13800
rect 21396 -13632 21493 -13616
rect 21396 -13800 21412 -13632
rect 21446 -13800 21493 -13632
rect 21396 -13816 21493 -13800
rect 21893 -13632 21990 -13616
rect 21893 -13800 21940 -13632
rect 21974 -13800 21990 -13632
rect 21893 -13816 21990 -13800
rect 20760 -14158 20857 -14142
rect 20760 -14926 20776 -14158
rect 20810 -14926 20857 -14158
rect 20760 -14942 20857 -14926
rect 21257 -14158 21354 -14142
rect 21257 -14926 21304 -14158
rect 21338 -14926 21354 -14158
rect 21257 -14942 21354 -14926
rect 21396 -14158 21493 -14142
rect 21396 -14926 21412 -14158
rect 21446 -14926 21493 -14158
rect 21396 -14942 21493 -14926
rect 21893 -14158 21990 -14142
rect 21893 -14926 21940 -14158
rect 21974 -14926 21990 -14158
rect 21893 -14942 21990 -14926
rect 22360 -13632 22457 -13616
rect 22360 -13800 22376 -13632
rect 22410 -13800 22457 -13632
rect 22360 -13816 22457 -13800
rect 22857 -13632 22954 -13616
rect 22857 -13800 22904 -13632
rect 22938 -13800 22954 -13632
rect 22857 -13816 22954 -13800
rect 22996 -13632 23093 -13616
rect 22996 -13800 23012 -13632
rect 23046 -13800 23093 -13632
rect 22996 -13816 23093 -13800
rect 23493 -13632 23590 -13616
rect 23493 -13800 23540 -13632
rect 23574 -13800 23590 -13632
rect 23493 -13816 23590 -13800
rect 22360 -14158 22457 -14142
rect 22360 -14926 22376 -14158
rect 22410 -14926 22457 -14158
rect 22360 -14942 22457 -14926
rect 22857 -14158 22954 -14142
rect 22857 -14926 22904 -14158
rect 22938 -14926 22954 -14158
rect 22857 -14942 22954 -14926
rect 22996 -14158 23093 -14142
rect 22996 -14926 23012 -14158
rect 23046 -14926 23093 -14158
rect 22996 -14942 23093 -14926
rect 23493 -14158 23590 -14142
rect 23493 -14926 23540 -14158
rect 23574 -14926 23590 -14158
rect 23493 -14942 23590 -14926
rect 23960 -13632 24057 -13616
rect 23960 -13800 23976 -13632
rect 24010 -13800 24057 -13632
rect 23960 -13816 24057 -13800
rect 24457 -13632 24554 -13616
rect 24457 -13800 24504 -13632
rect 24538 -13800 24554 -13632
rect 24457 -13816 24554 -13800
rect 24596 -13632 24693 -13616
rect 24596 -13800 24612 -13632
rect 24646 -13800 24693 -13632
rect 24596 -13816 24693 -13800
rect 25093 -13632 25190 -13616
rect 25093 -13800 25140 -13632
rect 25174 -13800 25190 -13632
rect 25093 -13816 25190 -13800
rect 23960 -14158 24057 -14142
rect 23960 -14926 23976 -14158
rect 24010 -14926 24057 -14158
rect 23960 -14942 24057 -14926
rect 24457 -14158 24554 -14142
rect 24457 -14926 24504 -14158
rect 24538 -14926 24554 -14158
rect 24457 -14942 24554 -14926
rect 24596 -14158 24693 -14142
rect 24596 -14926 24612 -14158
rect 24646 -14926 24693 -14158
rect 24596 -14942 24693 -14926
rect 25093 -14158 25190 -14142
rect 25093 -14926 25140 -14158
rect 25174 -14926 25190 -14158
rect 25093 -14942 25190 -14926
rect 25560 -13632 25657 -13616
rect 25560 -13800 25576 -13632
rect 25610 -13800 25657 -13632
rect 25560 -13816 25657 -13800
rect 26057 -13632 26154 -13616
rect 26057 -13800 26104 -13632
rect 26138 -13800 26154 -13632
rect 26057 -13816 26154 -13800
rect 26196 -13632 26293 -13616
rect 26196 -13800 26212 -13632
rect 26246 -13800 26293 -13632
rect 26196 -13816 26293 -13800
rect 26693 -13632 26790 -13616
rect 26693 -13800 26740 -13632
rect 26774 -13800 26790 -13632
rect 26693 -13816 26790 -13800
rect 25560 -14158 25657 -14142
rect 25560 -14926 25576 -14158
rect 25610 -14926 25657 -14158
rect 25560 -14942 25657 -14926
rect 26057 -14158 26154 -14142
rect 26057 -14926 26104 -14158
rect 26138 -14926 26154 -14158
rect 26057 -14942 26154 -14926
rect 26196 -14158 26293 -14142
rect 26196 -14926 26212 -14158
rect 26246 -14926 26293 -14158
rect 26196 -14942 26293 -14926
rect 26693 -14158 26790 -14142
rect 26693 -14926 26740 -14158
rect 26774 -14926 26790 -14158
rect 26693 -14942 26790 -14926
rect 27160 -13632 27257 -13616
rect 27160 -13800 27176 -13632
rect 27210 -13800 27257 -13632
rect 27160 -13816 27257 -13800
rect 27657 -13632 27754 -13616
rect 27657 -13800 27704 -13632
rect 27738 -13800 27754 -13632
rect 27657 -13816 27754 -13800
rect 27796 -13632 27893 -13616
rect 27796 -13800 27812 -13632
rect 27846 -13800 27893 -13632
rect 27796 -13816 27893 -13800
rect 28293 -13632 28390 -13616
rect 28293 -13800 28340 -13632
rect 28374 -13800 28390 -13632
rect 28293 -13816 28390 -13800
rect 27160 -14158 27257 -14142
rect 27160 -14926 27176 -14158
rect 27210 -14926 27257 -14158
rect 27160 -14942 27257 -14926
rect 27657 -14158 27754 -14142
rect 27657 -14926 27704 -14158
rect 27738 -14926 27754 -14158
rect 27657 -14942 27754 -14926
rect 27796 -14158 27893 -14142
rect 27796 -14926 27812 -14158
rect 27846 -14926 27893 -14158
rect 27796 -14942 27893 -14926
rect 28293 -14158 28390 -14142
rect 28293 -14926 28340 -14158
rect 28374 -14926 28390 -14158
rect 28293 -14942 28390 -14926
rect 28760 -13632 28857 -13616
rect 28760 -13800 28776 -13632
rect 28810 -13800 28857 -13632
rect 28760 -13816 28857 -13800
rect 29257 -13632 29354 -13616
rect 29257 -13800 29304 -13632
rect 29338 -13800 29354 -13632
rect 29257 -13816 29354 -13800
rect 29396 -13632 29493 -13616
rect 29396 -13800 29412 -13632
rect 29446 -13800 29493 -13632
rect 29396 -13816 29493 -13800
rect 29893 -13632 29990 -13616
rect 29893 -13800 29940 -13632
rect 29974 -13800 29990 -13632
rect 29893 -13816 29990 -13800
rect 28760 -14158 28857 -14142
rect 28760 -14926 28776 -14158
rect 28810 -14926 28857 -14158
rect 28760 -14942 28857 -14926
rect 29257 -14158 29354 -14142
rect 29257 -14926 29304 -14158
rect 29338 -14926 29354 -14158
rect 29257 -14942 29354 -14926
rect 29396 -14158 29493 -14142
rect 29396 -14926 29412 -14158
rect 29446 -14926 29493 -14158
rect 29396 -14942 29493 -14926
rect 29893 -14158 29990 -14142
rect 29893 -14926 29940 -14158
rect 29974 -14926 29990 -14158
rect 29893 -14942 29990 -14926
rect 30360 -13632 30457 -13616
rect 30360 -13800 30376 -13632
rect 30410 -13800 30457 -13632
rect 30360 -13816 30457 -13800
rect 30857 -13632 30954 -13616
rect 30857 -13800 30904 -13632
rect 30938 -13800 30954 -13632
rect 30857 -13816 30954 -13800
rect 30996 -13632 31093 -13616
rect 30996 -13800 31012 -13632
rect 31046 -13800 31093 -13632
rect 30996 -13816 31093 -13800
rect 31493 -13632 31590 -13616
rect 31493 -13800 31540 -13632
rect 31574 -13800 31590 -13632
rect 31493 -13816 31590 -13800
rect 30360 -14158 30457 -14142
rect 30360 -14926 30376 -14158
rect 30410 -14926 30457 -14158
rect 30360 -14942 30457 -14926
rect 30857 -14158 30954 -14142
rect 30857 -14926 30904 -14158
rect 30938 -14926 30954 -14158
rect 30857 -14942 30954 -14926
rect 30996 -14158 31093 -14142
rect 30996 -14926 31012 -14158
rect 31046 -14926 31093 -14158
rect 30996 -14942 31093 -14926
rect 31493 -14158 31590 -14142
rect 31493 -14926 31540 -14158
rect 31574 -14926 31590 -14158
rect 31493 -14942 31590 -14926
rect 31960 -13632 32057 -13616
rect 31960 -13800 31976 -13632
rect 32010 -13800 32057 -13632
rect 31960 -13816 32057 -13800
rect 32457 -13632 32554 -13616
rect 32457 -13800 32504 -13632
rect 32538 -13800 32554 -13632
rect 32457 -13816 32554 -13800
rect 32596 -13632 32693 -13616
rect 32596 -13800 32612 -13632
rect 32646 -13800 32693 -13632
rect 32596 -13816 32693 -13800
rect 33093 -13632 33190 -13616
rect 33093 -13800 33140 -13632
rect 33174 -13800 33190 -13632
rect 33093 -13816 33190 -13800
rect 31960 -14158 32057 -14142
rect 31960 -14926 31976 -14158
rect 32010 -14926 32057 -14158
rect 31960 -14942 32057 -14926
rect 32457 -14158 32554 -14142
rect 32457 -14926 32504 -14158
rect 32538 -14926 32554 -14158
rect 32457 -14942 32554 -14926
rect 32596 -14158 32693 -14142
rect 32596 -14926 32612 -14158
rect 32646 -14926 32693 -14158
rect 32596 -14942 32693 -14926
rect 33093 -14158 33190 -14142
rect 33093 -14926 33140 -14158
rect 33174 -14926 33190 -14158
rect 33093 -14942 33190 -14926
rect 33560 -13632 33657 -13616
rect 33560 -13800 33576 -13632
rect 33610 -13800 33657 -13632
rect 33560 -13816 33657 -13800
rect 34057 -13632 34154 -13616
rect 34057 -13800 34104 -13632
rect 34138 -13800 34154 -13632
rect 34057 -13816 34154 -13800
rect 34196 -13632 34293 -13616
rect 34196 -13800 34212 -13632
rect 34246 -13800 34293 -13632
rect 34196 -13816 34293 -13800
rect 34693 -13632 34790 -13616
rect 34693 -13800 34740 -13632
rect 34774 -13800 34790 -13632
rect 34693 -13816 34790 -13800
rect 33560 -14158 33657 -14142
rect 33560 -14926 33576 -14158
rect 33610 -14926 33657 -14158
rect 33560 -14942 33657 -14926
rect 34057 -14158 34154 -14142
rect 34057 -14926 34104 -14158
rect 34138 -14926 34154 -14158
rect 34057 -14942 34154 -14926
rect 34196 -14158 34293 -14142
rect 34196 -14926 34212 -14158
rect 34246 -14926 34293 -14158
rect 34196 -14942 34293 -14926
rect 34693 -14158 34790 -14142
rect 34693 -14926 34740 -14158
rect 34774 -14926 34790 -14158
rect 34693 -14942 34790 -14926
rect 35160 -13632 35257 -13616
rect 35160 -13800 35176 -13632
rect 35210 -13800 35257 -13632
rect 35160 -13816 35257 -13800
rect 35657 -13632 35754 -13616
rect 35657 -13800 35704 -13632
rect 35738 -13800 35754 -13632
rect 35657 -13816 35754 -13800
rect 35796 -13632 35893 -13616
rect 35796 -13800 35812 -13632
rect 35846 -13800 35893 -13632
rect 35796 -13816 35893 -13800
rect 36293 -13632 36390 -13616
rect 36293 -13800 36340 -13632
rect 36374 -13800 36390 -13632
rect 36293 -13816 36390 -13800
rect 35160 -14158 35257 -14142
rect 35160 -14926 35176 -14158
rect 35210 -14926 35257 -14158
rect 35160 -14942 35257 -14926
rect 35657 -14158 35754 -14142
rect 35657 -14926 35704 -14158
rect 35738 -14926 35754 -14158
rect 35657 -14942 35754 -14926
rect 35796 -14158 35893 -14142
rect 35796 -14926 35812 -14158
rect 35846 -14926 35893 -14158
rect 35796 -14942 35893 -14926
rect 36293 -14158 36390 -14142
rect 36293 -14926 36340 -14158
rect 36374 -14926 36390 -14158
rect 36293 -14942 36390 -14926
rect 36760 -13632 36857 -13616
rect 36760 -13800 36776 -13632
rect 36810 -13800 36857 -13632
rect 36760 -13816 36857 -13800
rect 37257 -13632 37354 -13616
rect 37257 -13800 37304 -13632
rect 37338 -13800 37354 -13632
rect 37257 -13816 37354 -13800
rect 37396 -13632 37493 -13616
rect 37396 -13800 37412 -13632
rect 37446 -13800 37493 -13632
rect 37396 -13816 37493 -13800
rect 37893 -13632 37990 -13616
rect 37893 -13800 37940 -13632
rect 37974 -13800 37990 -13632
rect 37893 -13816 37990 -13800
rect 36760 -14158 36857 -14142
rect 36760 -14926 36776 -14158
rect 36810 -14926 36857 -14158
rect 36760 -14942 36857 -14926
rect 37257 -14158 37354 -14142
rect 37257 -14926 37304 -14158
rect 37338 -14926 37354 -14158
rect 37257 -14942 37354 -14926
rect 37396 -14158 37493 -14142
rect 37396 -14926 37412 -14158
rect 37446 -14926 37493 -14158
rect 37396 -14942 37493 -14926
rect 37893 -14158 37990 -14142
rect 37893 -14926 37940 -14158
rect 37974 -14926 37990 -14158
rect 37893 -14942 37990 -14926
rect -40 -15432 57 -15416
rect -40 -15600 -24 -15432
rect 10 -15600 57 -15432
rect -40 -15616 57 -15600
rect 457 -15432 554 -15416
rect 457 -15600 504 -15432
rect 538 -15600 554 -15432
rect 457 -15616 554 -15600
rect 596 -15432 693 -15416
rect 596 -15600 612 -15432
rect 646 -15600 693 -15432
rect 596 -15616 693 -15600
rect 1093 -15432 1190 -15416
rect 1093 -15600 1140 -15432
rect 1174 -15600 1190 -15432
rect 1093 -15616 1190 -15600
rect -40 -15958 57 -15942
rect -40 -16726 -24 -15958
rect 10 -16726 57 -15958
rect -40 -16742 57 -16726
rect 457 -15958 554 -15942
rect 457 -16726 504 -15958
rect 538 -16726 554 -15958
rect 457 -16742 554 -16726
rect 596 -15958 693 -15942
rect 596 -16726 612 -15958
rect 646 -16726 693 -15958
rect 596 -16742 693 -16726
rect 1093 -15958 1190 -15942
rect 1093 -16726 1140 -15958
rect 1174 -16726 1190 -15958
rect 1093 -16742 1190 -16726
rect 1560 -15432 1657 -15416
rect 1560 -15600 1576 -15432
rect 1610 -15600 1657 -15432
rect 1560 -15616 1657 -15600
rect 2057 -15432 2154 -15416
rect 2057 -15600 2104 -15432
rect 2138 -15600 2154 -15432
rect 2057 -15616 2154 -15600
rect 2196 -15432 2293 -15416
rect 2196 -15600 2212 -15432
rect 2246 -15600 2293 -15432
rect 2196 -15616 2293 -15600
rect 2693 -15432 2790 -15416
rect 2693 -15600 2740 -15432
rect 2774 -15600 2790 -15432
rect 2693 -15616 2790 -15600
rect 1560 -15958 1657 -15942
rect 1560 -16726 1576 -15958
rect 1610 -16726 1657 -15958
rect 1560 -16742 1657 -16726
rect 2057 -15958 2154 -15942
rect 2057 -16726 2104 -15958
rect 2138 -16726 2154 -15958
rect 2057 -16742 2154 -16726
rect 2196 -15958 2293 -15942
rect 2196 -16726 2212 -15958
rect 2246 -16726 2293 -15958
rect 2196 -16742 2293 -16726
rect 2693 -15958 2790 -15942
rect 2693 -16726 2740 -15958
rect 2774 -16726 2790 -15958
rect 2693 -16742 2790 -16726
rect 3160 -15432 3257 -15416
rect 3160 -15600 3176 -15432
rect 3210 -15600 3257 -15432
rect 3160 -15616 3257 -15600
rect 3657 -15432 3754 -15416
rect 3657 -15600 3704 -15432
rect 3738 -15600 3754 -15432
rect 3657 -15616 3754 -15600
rect 3796 -15432 3893 -15416
rect 3796 -15600 3812 -15432
rect 3846 -15600 3893 -15432
rect 3796 -15616 3893 -15600
rect 4293 -15432 4390 -15416
rect 4293 -15600 4340 -15432
rect 4374 -15600 4390 -15432
rect 4293 -15616 4390 -15600
rect 3160 -15958 3257 -15942
rect 3160 -16726 3176 -15958
rect 3210 -16726 3257 -15958
rect 3160 -16742 3257 -16726
rect 3657 -15958 3754 -15942
rect 3657 -16726 3704 -15958
rect 3738 -16726 3754 -15958
rect 3657 -16742 3754 -16726
rect 3796 -15958 3893 -15942
rect 3796 -16726 3812 -15958
rect 3846 -16726 3893 -15958
rect 3796 -16742 3893 -16726
rect 4293 -15958 4390 -15942
rect 4293 -16726 4340 -15958
rect 4374 -16726 4390 -15958
rect 4293 -16742 4390 -16726
rect 4760 -15432 4857 -15416
rect 4760 -15600 4776 -15432
rect 4810 -15600 4857 -15432
rect 4760 -15616 4857 -15600
rect 5257 -15432 5354 -15416
rect 5257 -15600 5304 -15432
rect 5338 -15600 5354 -15432
rect 5257 -15616 5354 -15600
rect 5396 -15432 5493 -15416
rect 5396 -15600 5412 -15432
rect 5446 -15600 5493 -15432
rect 5396 -15616 5493 -15600
rect 5893 -15432 5990 -15416
rect 5893 -15600 5940 -15432
rect 5974 -15600 5990 -15432
rect 5893 -15616 5990 -15600
rect 4760 -15958 4857 -15942
rect 4760 -16726 4776 -15958
rect 4810 -16726 4857 -15958
rect 4760 -16742 4857 -16726
rect 5257 -15958 5354 -15942
rect 5257 -16726 5304 -15958
rect 5338 -16726 5354 -15958
rect 5257 -16742 5354 -16726
rect 5396 -15958 5493 -15942
rect 5396 -16726 5412 -15958
rect 5446 -16726 5493 -15958
rect 5396 -16742 5493 -16726
rect 5893 -15958 5990 -15942
rect 5893 -16726 5940 -15958
rect 5974 -16726 5990 -15958
rect 5893 -16742 5990 -16726
rect 6360 -15432 6457 -15416
rect 6360 -15600 6376 -15432
rect 6410 -15600 6457 -15432
rect 6360 -15616 6457 -15600
rect 6857 -15432 6954 -15416
rect 6857 -15600 6904 -15432
rect 6938 -15600 6954 -15432
rect 6857 -15616 6954 -15600
rect 6996 -15432 7093 -15416
rect 6996 -15600 7012 -15432
rect 7046 -15600 7093 -15432
rect 6996 -15616 7093 -15600
rect 7493 -15432 7590 -15416
rect 7493 -15600 7540 -15432
rect 7574 -15600 7590 -15432
rect 7493 -15616 7590 -15600
rect 6360 -15958 6457 -15942
rect 6360 -16726 6376 -15958
rect 6410 -16726 6457 -15958
rect 6360 -16742 6457 -16726
rect 6857 -15958 6954 -15942
rect 6857 -16726 6904 -15958
rect 6938 -16726 6954 -15958
rect 6857 -16742 6954 -16726
rect 6996 -15958 7093 -15942
rect 6996 -16726 7012 -15958
rect 7046 -16726 7093 -15958
rect 6996 -16742 7093 -16726
rect 7493 -15958 7590 -15942
rect 7493 -16726 7540 -15958
rect 7574 -16726 7590 -15958
rect 7493 -16742 7590 -16726
rect 7960 -15432 8057 -15416
rect 7960 -15600 7976 -15432
rect 8010 -15600 8057 -15432
rect 7960 -15616 8057 -15600
rect 8457 -15432 8554 -15416
rect 8457 -15600 8504 -15432
rect 8538 -15600 8554 -15432
rect 8457 -15616 8554 -15600
rect 8596 -15432 8693 -15416
rect 8596 -15600 8612 -15432
rect 8646 -15600 8693 -15432
rect 8596 -15616 8693 -15600
rect 9093 -15432 9190 -15416
rect 9093 -15600 9140 -15432
rect 9174 -15600 9190 -15432
rect 9093 -15616 9190 -15600
rect 7960 -15958 8057 -15942
rect 7960 -16726 7976 -15958
rect 8010 -16726 8057 -15958
rect 7960 -16742 8057 -16726
rect 8457 -15958 8554 -15942
rect 8457 -16726 8504 -15958
rect 8538 -16726 8554 -15958
rect 8457 -16742 8554 -16726
rect 8596 -15958 8693 -15942
rect 8596 -16726 8612 -15958
rect 8646 -16726 8693 -15958
rect 8596 -16742 8693 -16726
rect 9093 -15958 9190 -15942
rect 9093 -16726 9140 -15958
rect 9174 -16726 9190 -15958
rect 9093 -16742 9190 -16726
rect 9560 -15432 9657 -15416
rect 9560 -15600 9576 -15432
rect 9610 -15600 9657 -15432
rect 9560 -15616 9657 -15600
rect 10057 -15432 10154 -15416
rect 10057 -15600 10104 -15432
rect 10138 -15600 10154 -15432
rect 10057 -15616 10154 -15600
rect 10196 -15432 10293 -15416
rect 10196 -15600 10212 -15432
rect 10246 -15600 10293 -15432
rect 10196 -15616 10293 -15600
rect 10693 -15432 10790 -15416
rect 10693 -15600 10740 -15432
rect 10774 -15600 10790 -15432
rect 10693 -15616 10790 -15600
rect 9560 -15958 9657 -15942
rect 9560 -16726 9576 -15958
rect 9610 -16726 9657 -15958
rect 9560 -16742 9657 -16726
rect 10057 -15958 10154 -15942
rect 10057 -16726 10104 -15958
rect 10138 -16726 10154 -15958
rect 10057 -16742 10154 -16726
rect 10196 -15958 10293 -15942
rect 10196 -16726 10212 -15958
rect 10246 -16726 10293 -15958
rect 10196 -16742 10293 -16726
rect 10693 -15958 10790 -15942
rect 10693 -16726 10740 -15958
rect 10774 -16726 10790 -15958
rect 10693 -16742 10790 -16726
rect 11160 -15432 11257 -15416
rect 11160 -15600 11176 -15432
rect 11210 -15600 11257 -15432
rect 11160 -15616 11257 -15600
rect 11657 -15432 11754 -15416
rect 11657 -15600 11704 -15432
rect 11738 -15600 11754 -15432
rect 11657 -15616 11754 -15600
rect 11796 -15432 11893 -15416
rect 11796 -15600 11812 -15432
rect 11846 -15600 11893 -15432
rect 11796 -15616 11893 -15600
rect 12293 -15432 12390 -15416
rect 12293 -15600 12340 -15432
rect 12374 -15600 12390 -15432
rect 12293 -15616 12390 -15600
rect 11160 -15958 11257 -15942
rect 11160 -16726 11176 -15958
rect 11210 -16726 11257 -15958
rect 11160 -16742 11257 -16726
rect 11657 -15958 11754 -15942
rect 11657 -16726 11704 -15958
rect 11738 -16726 11754 -15958
rect 11657 -16742 11754 -16726
rect 11796 -15958 11893 -15942
rect 11796 -16726 11812 -15958
rect 11846 -16726 11893 -15958
rect 11796 -16742 11893 -16726
rect 12293 -15958 12390 -15942
rect 12293 -16726 12340 -15958
rect 12374 -16726 12390 -15958
rect 12293 -16742 12390 -16726
rect 12760 -15432 12857 -15416
rect 12760 -15600 12776 -15432
rect 12810 -15600 12857 -15432
rect 12760 -15616 12857 -15600
rect 13257 -15432 13354 -15416
rect 13257 -15600 13304 -15432
rect 13338 -15600 13354 -15432
rect 13257 -15616 13354 -15600
rect 13396 -15432 13493 -15416
rect 13396 -15600 13412 -15432
rect 13446 -15600 13493 -15432
rect 13396 -15616 13493 -15600
rect 13893 -15432 13990 -15416
rect 13893 -15600 13940 -15432
rect 13974 -15600 13990 -15432
rect 13893 -15616 13990 -15600
rect 12760 -15958 12857 -15942
rect 12760 -16726 12776 -15958
rect 12810 -16726 12857 -15958
rect 12760 -16742 12857 -16726
rect 13257 -15958 13354 -15942
rect 13257 -16726 13304 -15958
rect 13338 -16726 13354 -15958
rect 13257 -16742 13354 -16726
rect 13396 -15958 13493 -15942
rect 13396 -16726 13412 -15958
rect 13446 -16726 13493 -15958
rect 13396 -16742 13493 -16726
rect 13893 -15958 13990 -15942
rect 13893 -16726 13940 -15958
rect 13974 -16726 13990 -15958
rect 13893 -16742 13990 -16726
rect 14360 -15432 14457 -15416
rect 14360 -15600 14376 -15432
rect 14410 -15600 14457 -15432
rect 14360 -15616 14457 -15600
rect 14857 -15432 14954 -15416
rect 14857 -15600 14904 -15432
rect 14938 -15600 14954 -15432
rect 14857 -15616 14954 -15600
rect 14996 -15432 15093 -15416
rect 14996 -15600 15012 -15432
rect 15046 -15600 15093 -15432
rect 14996 -15616 15093 -15600
rect 15493 -15432 15590 -15416
rect 15493 -15600 15540 -15432
rect 15574 -15600 15590 -15432
rect 15493 -15616 15590 -15600
rect 14360 -15958 14457 -15942
rect 14360 -16726 14376 -15958
rect 14410 -16726 14457 -15958
rect 14360 -16742 14457 -16726
rect 14857 -15958 14954 -15942
rect 14857 -16726 14904 -15958
rect 14938 -16726 14954 -15958
rect 14857 -16742 14954 -16726
rect 14996 -15958 15093 -15942
rect 14996 -16726 15012 -15958
rect 15046 -16726 15093 -15958
rect 14996 -16742 15093 -16726
rect 15493 -15958 15590 -15942
rect 15493 -16726 15540 -15958
rect 15574 -16726 15590 -15958
rect 15493 -16742 15590 -16726
rect 15960 -15432 16057 -15416
rect 15960 -15600 15976 -15432
rect 16010 -15600 16057 -15432
rect 15960 -15616 16057 -15600
rect 16457 -15432 16554 -15416
rect 16457 -15600 16504 -15432
rect 16538 -15600 16554 -15432
rect 16457 -15616 16554 -15600
rect 16596 -15432 16693 -15416
rect 16596 -15600 16612 -15432
rect 16646 -15600 16693 -15432
rect 16596 -15616 16693 -15600
rect 17093 -15432 17190 -15416
rect 17093 -15600 17140 -15432
rect 17174 -15600 17190 -15432
rect 17093 -15616 17190 -15600
rect 15960 -15958 16057 -15942
rect 15960 -16726 15976 -15958
rect 16010 -16726 16057 -15958
rect 15960 -16742 16057 -16726
rect 16457 -15958 16554 -15942
rect 16457 -16726 16504 -15958
rect 16538 -16726 16554 -15958
rect 16457 -16742 16554 -16726
rect 16596 -15958 16693 -15942
rect 16596 -16726 16612 -15958
rect 16646 -16726 16693 -15958
rect 16596 -16742 16693 -16726
rect 17093 -15958 17190 -15942
rect 17093 -16726 17140 -15958
rect 17174 -16726 17190 -15958
rect 17093 -16742 17190 -16726
rect 17560 -15432 17657 -15416
rect 17560 -15600 17576 -15432
rect 17610 -15600 17657 -15432
rect 17560 -15616 17657 -15600
rect 18057 -15432 18154 -15416
rect 18057 -15600 18104 -15432
rect 18138 -15600 18154 -15432
rect 18057 -15616 18154 -15600
rect 18196 -15432 18293 -15416
rect 18196 -15600 18212 -15432
rect 18246 -15600 18293 -15432
rect 18196 -15616 18293 -15600
rect 18693 -15432 18790 -15416
rect 18693 -15600 18740 -15432
rect 18774 -15600 18790 -15432
rect 18693 -15616 18790 -15600
rect 17560 -15958 17657 -15942
rect 17560 -16726 17576 -15958
rect 17610 -16726 17657 -15958
rect 17560 -16742 17657 -16726
rect 18057 -15958 18154 -15942
rect 18057 -16726 18104 -15958
rect 18138 -16726 18154 -15958
rect 18057 -16742 18154 -16726
rect 18196 -15958 18293 -15942
rect 18196 -16726 18212 -15958
rect 18246 -16726 18293 -15958
rect 18196 -16742 18293 -16726
rect 18693 -15958 18790 -15942
rect 18693 -16726 18740 -15958
rect 18774 -16726 18790 -15958
rect 18693 -16742 18790 -16726
rect 19160 -15432 19257 -15416
rect 19160 -15600 19176 -15432
rect 19210 -15600 19257 -15432
rect 19160 -15616 19257 -15600
rect 19657 -15432 19754 -15416
rect 19657 -15600 19704 -15432
rect 19738 -15600 19754 -15432
rect 19657 -15616 19754 -15600
rect 19796 -15432 19893 -15416
rect 19796 -15600 19812 -15432
rect 19846 -15600 19893 -15432
rect 19796 -15616 19893 -15600
rect 20293 -15432 20390 -15416
rect 20293 -15600 20340 -15432
rect 20374 -15600 20390 -15432
rect 20293 -15616 20390 -15600
rect 19160 -15958 19257 -15942
rect 19160 -16726 19176 -15958
rect 19210 -16726 19257 -15958
rect 19160 -16742 19257 -16726
rect 19657 -15958 19754 -15942
rect 19657 -16726 19704 -15958
rect 19738 -16726 19754 -15958
rect 19657 -16742 19754 -16726
rect 19796 -15958 19893 -15942
rect 19796 -16726 19812 -15958
rect 19846 -16726 19893 -15958
rect 19796 -16742 19893 -16726
rect 20293 -15958 20390 -15942
rect 20293 -16726 20340 -15958
rect 20374 -16726 20390 -15958
rect 20293 -16742 20390 -16726
rect 20760 -15432 20857 -15416
rect 20760 -15600 20776 -15432
rect 20810 -15600 20857 -15432
rect 20760 -15616 20857 -15600
rect 21257 -15432 21354 -15416
rect 21257 -15600 21304 -15432
rect 21338 -15600 21354 -15432
rect 21257 -15616 21354 -15600
rect 21396 -15432 21493 -15416
rect 21396 -15600 21412 -15432
rect 21446 -15600 21493 -15432
rect 21396 -15616 21493 -15600
rect 21893 -15432 21990 -15416
rect 21893 -15600 21940 -15432
rect 21974 -15600 21990 -15432
rect 21893 -15616 21990 -15600
rect 20760 -15958 20857 -15942
rect 20760 -16726 20776 -15958
rect 20810 -16726 20857 -15958
rect 20760 -16742 20857 -16726
rect 21257 -15958 21354 -15942
rect 21257 -16726 21304 -15958
rect 21338 -16726 21354 -15958
rect 21257 -16742 21354 -16726
rect 21396 -15958 21493 -15942
rect 21396 -16726 21412 -15958
rect 21446 -16726 21493 -15958
rect 21396 -16742 21493 -16726
rect 21893 -15958 21990 -15942
rect 21893 -16726 21940 -15958
rect 21974 -16726 21990 -15958
rect 21893 -16742 21990 -16726
rect 22360 -15432 22457 -15416
rect 22360 -15600 22376 -15432
rect 22410 -15600 22457 -15432
rect 22360 -15616 22457 -15600
rect 22857 -15432 22954 -15416
rect 22857 -15600 22904 -15432
rect 22938 -15600 22954 -15432
rect 22857 -15616 22954 -15600
rect 22996 -15432 23093 -15416
rect 22996 -15600 23012 -15432
rect 23046 -15600 23093 -15432
rect 22996 -15616 23093 -15600
rect 23493 -15432 23590 -15416
rect 23493 -15600 23540 -15432
rect 23574 -15600 23590 -15432
rect 23493 -15616 23590 -15600
rect 22360 -15958 22457 -15942
rect 22360 -16726 22376 -15958
rect 22410 -16726 22457 -15958
rect 22360 -16742 22457 -16726
rect 22857 -15958 22954 -15942
rect 22857 -16726 22904 -15958
rect 22938 -16726 22954 -15958
rect 22857 -16742 22954 -16726
rect 22996 -15958 23093 -15942
rect 22996 -16726 23012 -15958
rect 23046 -16726 23093 -15958
rect 22996 -16742 23093 -16726
rect 23493 -15958 23590 -15942
rect 23493 -16726 23540 -15958
rect 23574 -16726 23590 -15958
rect 23493 -16742 23590 -16726
rect 23960 -15432 24057 -15416
rect 23960 -15600 23976 -15432
rect 24010 -15600 24057 -15432
rect 23960 -15616 24057 -15600
rect 24457 -15432 24554 -15416
rect 24457 -15600 24504 -15432
rect 24538 -15600 24554 -15432
rect 24457 -15616 24554 -15600
rect 24596 -15432 24693 -15416
rect 24596 -15600 24612 -15432
rect 24646 -15600 24693 -15432
rect 24596 -15616 24693 -15600
rect 25093 -15432 25190 -15416
rect 25093 -15600 25140 -15432
rect 25174 -15600 25190 -15432
rect 25093 -15616 25190 -15600
rect 23960 -15958 24057 -15942
rect 23960 -16726 23976 -15958
rect 24010 -16726 24057 -15958
rect 23960 -16742 24057 -16726
rect 24457 -15958 24554 -15942
rect 24457 -16726 24504 -15958
rect 24538 -16726 24554 -15958
rect 24457 -16742 24554 -16726
rect 24596 -15958 24693 -15942
rect 24596 -16726 24612 -15958
rect 24646 -16726 24693 -15958
rect 24596 -16742 24693 -16726
rect 25093 -15958 25190 -15942
rect 25093 -16726 25140 -15958
rect 25174 -16726 25190 -15958
rect 25093 -16742 25190 -16726
rect 25560 -15432 25657 -15416
rect 25560 -15600 25576 -15432
rect 25610 -15600 25657 -15432
rect 25560 -15616 25657 -15600
rect 26057 -15432 26154 -15416
rect 26057 -15600 26104 -15432
rect 26138 -15600 26154 -15432
rect 26057 -15616 26154 -15600
rect 26196 -15432 26293 -15416
rect 26196 -15600 26212 -15432
rect 26246 -15600 26293 -15432
rect 26196 -15616 26293 -15600
rect 26693 -15432 26790 -15416
rect 26693 -15600 26740 -15432
rect 26774 -15600 26790 -15432
rect 26693 -15616 26790 -15600
rect 25560 -15958 25657 -15942
rect 25560 -16726 25576 -15958
rect 25610 -16726 25657 -15958
rect 25560 -16742 25657 -16726
rect 26057 -15958 26154 -15942
rect 26057 -16726 26104 -15958
rect 26138 -16726 26154 -15958
rect 26057 -16742 26154 -16726
rect 26196 -15958 26293 -15942
rect 26196 -16726 26212 -15958
rect 26246 -16726 26293 -15958
rect 26196 -16742 26293 -16726
rect 26693 -15958 26790 -15942
rect 26693 -16726 26740 -15958
rect 26774 -16726 26790 -15958
rect 26693 -16742 26790 -16726
rect 27160 -15432 27257 -15416
rect 27160 -15600 27176 -15432
rect 27210 -15600 27257 -15432
rect 27160 -15616 27257 -15600
rect 27657 -15432 27754 -15416
rect 27657 -15600 27704 -15432
rect 27738 -15600 27754 -15432
rect 27657 -15616 27754 -15600
rect 27796 -15432 27893 -15416
rect 27796 -15600 27812 -15432
rect 27846 -15600 27893 -15432
rect 27796 -15616 27893 -15600
rect 28293 -15432 28390 -15416
rect 28293 -15600 28340 -15432
rect 28374 -15600 28390 -15432
rect 28293 -15616 28390 -15600
rect 27160 -15958 27257 -15942
rect 27160 -16726 27176 -15958
rect 27210 -16726 27257 -15958
rect 27160 -16742 27257 -16726
rect 27657 -15958 27754 -15942
rect 27657 -16726 27704 -15958
rect 27738 -16726 27754 -15958
rect 27657 -16742 27754 -16726
rect 27796 -15958 27893 -15942
rect 27796 -16726 27812 -15958
rect 27846 -16726 27893 -15958
rect 27796 -16742 27893 -16726
rect 28293 -15958 28390 -15942
rect 28293 -16726 28340 -15958
rect 28374 -16726 28390 -15958
rect 28293 -16742 28390 -16726
rect 28760 -15432 28857 -15416
rect 28760 -15600 28776 -15432
rect 28810 -15600 28857 -15432
rect 28760 -15616 28857 -15600
rect 29257 -15432 29354 -15416
rect 29257 -15600 29304 -15432
rect 29338 -15600 29354 -15432
rect 29257 -15616 29354 -15600
rect 29396 -15432 29493 -15416
rect 29396 -15600 29412 -15432
rect 29446 -15600 29493 -15432
rect 29396 -15616 29493 -15600
rect 29893 -15432 29990 -15416
rect 29893 -15600 29940 -15432
rect 29974 -15600 29990 -15432
rect 29893 -15616 29990 -15600
rect 28760 -15958 28857 -15942
rect 28760 -16726 28776 -15958
rect 28810 -16726 28857 -15958
rect 28760 -16742 28857 -16726
rect 29257 -15958 29354 -15942
rect 29257 -16726 29304 -15958
rect 29338 -16726 29354 -15958
rect 29257 -16742 29354 -16726
rect 29396 -15958 29493 -15942
rect 29396 -16726 29412 -15958
rect 29446 -16726 29493 -15958
rect 29396 -16742 29493 -16726
rect 29893 -15958 29990 -15942
rect 29893 -16726 29940 -15958
rect 29974 -16726 29990 -15958
rect 29893 -16742 29990 -16726
rect 30360 -15432 30457 -15416
rect 30360 -15600 30376 -15432
rect 30410 -15600 30457 -15432
rect 30360 -15616 30457 -15600
rect 30857 -15432 30954 -15416
rect 30857 -15600 30904 -15432
rect 30938 -15600 30954 -15432
rect 30857 -15616 30954 -15600
rect 30996 -15432 31093 -15416
rect 30996 -15600 31012 -15432
rect 31046 -15600 31093 -15432
rect 30996 -15616 31093 -15600
rect 31493 -15432 31590 -15416
rect 31493 -15600 31540 -15432
rect 31574 -15600 31590 -15432
rect 31493 -15616 31590 -15600
rect 30360 -15958 30457 -15942
rect 30360 -16726 30376 -15958
rect 30410 -16726 30457 -15958
rect 30360 -16742 30457 -16726
rect 30857 -15958 30954 -15942
rect 30857 -16726 30904 -15958
rect 30938 -16726 30954 -15958
rect 30857 -16742 30954 -16726
rect 30996 -15958 31093 -15942
rect 30996 -16726 31012 -15958
rect 31046 -16726 31093 -15958
rect 30996 -16742 31093 -16726
rect 31493 -15958 31590 -15942
rect 31493 -16726 31540 -15958
rect 31574 -16726 31590 -15958
rect 31493 -16742 31590 -16726
rect 31960 -15432 32057 -15416
rect 31960 -15600 31976 -15432
rect 32010 -15600 32057 -15432
rect 31960 -15616 32057 -15600
rect 32457 -15432 32554 -15416
rect 32457 -15600 32504 -15432
rect 32538 -15600 32554 -15432
rect 32457 -15616 32554 -15600
rect 32596 -15432 32693 -15416
rect 32596 -15600 32612 -15432
rect 32646 -15600 32693 -15432
rect 32596 -15616 32693 -15600
rect 33093 -15432 33190 -15416
rect 33093 -15600 33140 -15432
rect 33174 -15600 33190 -15432
rect 33093 -15616 33190 -15600
rect 31960 -15958 32057 -15942
rect 31960 -16726 31976 -15958
rect 32010 -16726 32057 -15958
rect 31960 -16742 32057 -16726
rect 32457 -15958 32554 -15942
rect 32457 -16726 32504 -15958
rect 32538 -16726 32554 -15958
rect 32457 -16742 32554 -16726
rect 32596 -15958 32693 -15942
rect 32596 -16726 32612 -15958
rect 32646 -16726 32693 -15958
rect 32596 -16742 32693 -16726
rect 33093 -15958 33190 -15942
rect 33093 -16726 33140 -15958
rect 33174 -16726 33190 -15958
rect 33093 -16742 33190 -16726
rect 33560 -15432 33657 -15416
rect 33560 -15600 33576 -15432
rect 33610 -15600 33657 -15432
rect 33560 -15616 33657 -15600
rect 34057 -15432 34154 -15416
rect 34057 -15600 34104 -15432
rect 34138 -15600 34154 -15432
rect 34057 -15616 34154 -15600
rect 34196 -15432 34293 -15416
rect 34196 -15600 34212 -15432
rect 34246 -15600 34293 -15432
rect 34196 -15616 34293 -15600
rect 34693 -15432 34790 -15416
rect 34693 -15600 34740 -15432
rect 34774 -15600 34790 -15432
rect 34693 -15616 34790 -15600
rect 33560 -15958 33657 -15942
rect 33560 -16726 33576 -15958
rect 33610 -16726 33657 -15958
rect 33560 -16742 33657 -16726
rect 34057 -15958 34154 -15942
rect 34057 -16726 34104 -15958
rect 34138 -16726 34154 -15958
rect 34057 -16742 34154 -16726
rect 34196 -15958 34293 -15942
rect 34196 -16726 34212 -15958
rect 34246 -16726 34293 -15958
rect 34196 -16742 34293 -16726
rect 34693 -15958 34790 -15942
rect 34693 -16726 34740 -15958
rect 34774 -16726 34790 -15958
rect 34693 -16742 34790 -16726
rect 35160 -15432 35257 -15416
rect 35160 -15600 35176 -15432
rect 35210 -15600 35257 -15432
rect 35160 -15616 35257 -15600
rect 35657 -15432 35754 -15416
rect 35657 -15600 35704 -15432
rect 35738 -15600 35754 -15432
rect 35657 -15616 35754 -15600
rect 35796 -15432 35893 -15416
rect 35796 -15600 35812 -15432
rect 35846 -15600 35893 -15432
rect 35796 -15616 35893 -15600
rect 36293 -15432 36390 -15416
rect 36293 -15600 36340 -15432
rect 36374 -15600 36390 -15432
rect 36293 -15616 36390 -15600
rect 35160 -15958 35257 -15942
rect 35160 -16726 35176 -15958
rect 35210 -16726 35257 -15958
rect 35160 -16742 35257 -16726
rect 35657 -15958 35754 -15942
rect 35657 -16726 35704 -15958
rect 35738 -16726 35754 -15958
rect 35657 -16742 35754 -16726
rect 35796 -15958 35893 -15942
rect 35796 -16726 35812 -15958
rect 35846 -16726 35893 -15958
rect 35796 -16742 35893 -16726
rect 36293 -15958 36390 -15942
rect 36293 -16726 36340 -15958
rect 36374 -16726 36390 -15958
rect 36293 -16742 36390 -16726
rect 36760 -15432 36857 -15416
rect 36760 -15600 36776 -15432
rect 36810 -15600 36857 -15432
rect 36760 -15616 36857 -15600
rect 37257 -15432 37354 -15416
rect 37257 -15600 37304 -15432
rect 37338 -15600 37354 -15432
rect 37257 -15616 37354 -15600
rect 37396 -15432 37493 -15416
rect 37396 -15600 37412 -15432
rect 37446 -15600 37493 -15432
rect 37396 -15616 37493 -15600
rect 37893 -15432 37990 -15416
rect 37893 -15600 37940 -15432
rect 37974 -15600 37990 -15432
rect 37893 -15616 37990 -15600
rect 36760 -15958 36857 -15942
rect 36760 -16726 36776 -15958
rect 36810 -16726 36857 -15958
rect 36760 -16742 36857 -16726
rect 37257 -15958 37354 -15942
rect 37257 -16726 37304 -15958
rect 37338 -16726 37354 -15958
rect 37257 -16742 37354 -16726
rect 37396 -15958 37493 -15942
rect 37396 -16726 37412 -15958
rect 37446 -16726 37493 -15958
rect 37396 -16742 37493 -16726
rect 37893 -15958 37990 -15942
rect 37893 -16726 37940 -15958
rect 37974 -16726 37990 -15958
rect 37893 -16742 37990 -16726
rect -40 -17232 57 -17216
rect -40 -17400 -24 -17232
rect 10 -17400 57 -17232
rect -40 -17416 57 -17400
rect 457 -17232 554 -17216
rect 457 -17400 504 -17232
rect 538 -17400 554 -17232
rect 457 -17416 554 -17400
rect 596 -17232 693 -17216
rect 596 -17400 612 -17232
rect 646 -17400 693 -17232
rect 596 -17416 693 -17400
rect 1093 -17232 1190 -17216
rect 1093 -17400 1140 -17232
rect 1174 -17400 1190 -17232
rect 1093 -17416 1190 -17400
rect -40 -17758 57 -17742
rect -40 -18526 -24 -17758
rect 10 -18526 57 -17758
rect -40 -18542 57 -18526
rect 457 -17758 554 -17742
rect 457 -18526 504 -17758
rect 538 -18526 554 -17758
rect 457 -18542 554 -18526
rect 596 -17758 693 -17742
rect 596 -18526 612 -17758
rect 646 -18526 693 -17758
rect 596 -18542 693 -18526
rect 1093 -17758 1190 -17742
rect 1093 -18526 1140 -17758
rect 1174 -18526 1190 -17758
rect 1093 -18542 1190 -18526
rect 1560 -17232 1657 -17216
rect 1560 -17400 1576 -17232
rect 1610 -17400 1657 -17232
rect 1560 -17416 1657 -17400
rect 2057 -17232 2154 -17216
rect 2057 -17400 2104 -17232
rect 2138 -17400 2154 -17232
rect 2057 -17416 2154 -17400
rect 2196 -17232 2293 -17216
rect 2196 -17400 2212 -17232
rect 2246 -17400 2293 -17232
rect 2196 -17416 2293 -17400
rect 2693 -17232 2790 -17216
rect 2693 -17400 2740 -17232
rect 2774 -17400 2790 -17232
rect 2693 -17416 2790 -17400
rect 1560 -17758 1657 -17742
rect 1560 -18526 1576 -17758
rect 1610 -18526 1657 -17758
rect 1560 -18542 1657 -18526
rect 2057 -17758 2154 -17742
rect 2057 -18526 2104 -17758
rect 2138 -18526 2154 -17758
rect 2057 -18542 2154 -18526
rect 2196 -17758 2293 -17742
rect 2196 -18526 2212 -17758
rect 2246 -18526 2293 -17758
rect 2196 -18542 2293 -18526
rect 2693 -17758 2790 -17742
rect 2693 -18526 2740 -17758
rect 2774 -18526 2790 -17758
rect 2693 -18542 2790 -18526
rect 3160 -17232 3257 -17216
rect 3160 -17400 3176 -17232
rect 3210 -17400 3257 -17232
rect 3160 -17416 3257 -17400
rect 3657 -17232 3754 -17216
rect 3657 -17400 3704 -17232
rect 3738 -17400 3754 -17232
rect 3657 -17416 3754 -17400
rect 3796 -17232 3893 -17216
rect 3796 -17400 3812 -17232
rect 3846 -17400 3893 -17232
rect 3796 -17416 3893 -17400
rect 4293 -17232 4390 -17216
rect 4293 -17400 4340 -17232
rect 4374 -17400 4390 -17232
rect 4293 -17416 4390 -17400
rect 3160 -17758 3257 -17742
rect 3160 -18526 3176 -17758
rect 3210 -18526 3257 -17758
rect 3160 -18542 3257 -18526
rect 3657 -17758 3754 -17742
rect 3657 -18526 3704 -17758
rect 3738 -18526 3754 -17758
rect 3657 -18542 3754 -18526
rect 3796 -17758 3893 -17742
rect 3796 -18526 3812 -17758
rect 3846 -18526 3893 -17758
rect 3796 -18542 3893 -18526
rect 4293 -17758 4390 -17742
rect 4293 -18526 4340 -17758
rect 4374 -18526 4390 -17758
rect 4293 -18542 4390 -18526
rect 4760 -17232 4857 -17216
rect 4760 -17400 4776 -17232
rect 4810 -17400 4857 -17232
rect 4760 -17416 4857 -17400
rect 5257 -17232 5354 -17216
rect 5257 -17400 5304 -17232
rect 5338 -17400 5354 -17232
rect 5257 -17416 5354 -17400
rect 5396 -17232 5493 -17216
rect 5396 -17400 5412 -17232
rect 5446 -17400 5493 -17232
rect 5396 -17416 5493 -17400
rect 5893 -17232 5990 -17216
rect 5893 -17400 5940 -17232
rect 5974 -17400 5990 -17232
rect 5893 -17416 5990 -17400
rect 4760 -17758 4857 -17742
rect 4760 -18526 4776 -17758
rect 4810 -18526 4857 -17758
rect 4760 -18542 4857 -18526
rect 5257 -17758 5354 -17742
rect 5257 -18526 5304 -17758
rect 5338 -18526 5354 -17758
rect 5257 -18542 5354 -18526
rect 5396 -17758 5493 -17742
rect 5396 -18526 5412 -17758
rect 5446 -18526 5493 -17758
rect 5396 -18542 5493 -18526
rect 5893 -17758 5990 -17742
rect 5893 -18526 5940 -17758
rect 5974 -18526 5990 -17758
rect 5893 -18542 5990 -18526
rect 6360 -17232 6457 -17216
rect 6360 -17400 6376 -17232
rect 6410 -17400 6457 -17232
rect 6360 -17416 6457 -17400
rect 6857 -17232 6954 -17216
rect 6857 -17400 6904 -17232
rect 6938 -17400 6954 -17232
rect 6857 -17416 6954 -17400
rect 6996 -17232 7093 -17216
rect 6996 -17400 7012 -17232
rect 7046 -17400 7093 -17232
rect 6996 -17416 7093 -17400
rect 7493 -17232 7590 -17216
rect 7493 -17400 7540 -17232
rect 7574 -17400 7590 -17232
rect 7493 -17416 7590 -17400
rect 6360 -17758 6457 -17742
rect 6360 -18526 6376 -17758
rect 6410 -18526 6457 -17758
rect 6360 -18542 6457 -18526
rect 6857 -17758 6954 -17742
rect 6857 -18526 6904 -17758
rect 6938 -18526 6954 -17758
rect 6857 -18542 6954 -18526
rect 6996 -17758 7093 -17742
rect 6996 -18526 7012 -17758
rect 7046 -18526 7093 -17758
rect 6996 -18542 7093 -18526
rect 7493 -17758 7590 -17742
rect 7493 -18526 7540 -17758
rect 7574 -18526 7590 -17758
rect 7493 -18542 7590 -18526
rect 7960 -17232 8057 -17216
rect 7960 -17400 7976 -17232
rect 8010 -17400 8057 -17232
rect 7960 -17416 8057 -17400
rect 8457 -17232 8554 -17216
rect 8457 -17400 8504 -17232
rect 8538 -17400 8554 -17232
rect 8457 -17416 8554 -17400
rect 8596 -17232 8693 -17216
rect 8596 -17400 8612 -17232
rect 8646 -17400 8693 -17232
rect 8596 -17416 8693 -17400
rect 9093 -17232 9190 -17216
rect 9093 -17400 9140 -17232
rect 9174 -17400 9190 -17232
rect 9093 -17416 9190 -17400
rect 7960 -17758 8057 -17742
rect 7960 -18526 7976 -17758
rect 8010 -18526 8057 -17758
rect 7960 -18542 8057 -18526
rect 8457 -17758 8554 -17742
rect 8457 -18526 8504 -17758
rect 8538 -18526 8554 -17758
rect 8457 -18542 8554 -18526
rect 8596 -17758 8693 -17742
rect 8596 -18526 8612 -17758
rect 8646 -18526 8693 -17758
rect 8596 -18542 8693 -18526
rect 9093 -17758 9190 -17742
rect 9093 -18526 9140 -17758
rect 9174 -18526 9190 -17758
rect 9093 -18542 9190 -18526
rect 9560 -17232 9657 -17216
rect 9560 -17400 9576 -17232
rect 9610 -17400 9657 -17232
rect 9560 -17416 9657 -17400
rect 10057 -17232 10154 -17216
rect 10057 -17400 10104 -17232
rect 10138 -17400 10154 -17232
rect 10057 -17416 10154 -17400
rect 10196 -17232 10293 -17216
rect 10196 -17400 10212 -17232
rect 10246 -17400 10293 -17232
rect 10196 -17416 10293 -17400
rect 10693 -17232 10790 -17216
rect 10693 -17400 10740 -17232
rect 10774 -17400 10790 -17232
rect 10693 -17416 10790 -17400
rect 9560 -17758 9657 -17742
rect 9560 -18526 9576 -17758
rect 9610 -18526 9657 -17758
rect 9560 -18542 9657 -18526
rect 10057 -17758 10154 -17742
rect 10057 -18526 10104 -17758
rect 10138 -18526 10154 -17758
rect 10057 -18542 10154 -18526
rect 10196 -17758 10293 -17742
rect 10196 -18526 10212 -17758
rect 10246 -18526 10293 -17758
rect 10196 -18542 10293 -18526
rect 10693 -17758 10790 -17742
rect 10693 -18526 10740 -17758
rect 10774 -18526 10790 -17758
rect 10693 -18542 10790 -18526
rect 11160 -17232 11257 -17216
rect 11160 -17400 11176 -17232
rect 11210 -17400 11257 -17232
rect 11160 -17416 11257 -17400
rect 11657 -17232 11754 -17216
rect 11657 -17400 11704 -17232
rect 11738 -17400 11754 -17232
rect 11657 -17416 11754 -17400
rect 11796 -17232 11893 -17216
rect 11796 -17400 11812 -17232
rect 11846 -17400 11893 -17232
rect 11796 -17416 11893 -17400
rect 12293 -17232 12390 -17216
rect 12293 -17400 12340 -17232
rect 12374 -17400 12390 -17232
rect 12293 -17416 12390 -17400
rect 11160 -17758 11257 -17742
rect 11160 -18526 11176 -17758
rect 11210 -18526 11257 -17758
rect 11160 -18542 11257 -18526
rect 11657 -17758 11754 -17742
rect 11657 -18526 11704 -17758
rect 11738 -18526 11754 -17758
rect 11657 -18542 11754 -18526
rect 11796 -17758 11893 -17742
rect 11796 -18526 11812 -17758
rect 11846 -18526 11893 -17758
rect 11796 -18542 11893 -18526
rect 12293 -17758 12390 -17742
rect 12293 -18526 12340 -17758
rect 12374 -18526 12390 -17758
rect 12293 -18542 12390 -18526
rect 12760 -17232 12857 -17216
rect 12760 -17400 12776 -17232
rect 12810 -17400 12857 -17232
rect 12760 -17416 12857 -17400
rect 13257 -17232 13354 -17216
rect 13257 -17400 13304 -17232
rect 13338 -17400 13354 -17232
rect 13257 -17416 13354 -17400
rect 13396 -17232 13493 -17216
rect 13396 -17400 13412 -17232
rect 13446 -17400 13493 -17232
rect 13396 -17416 13493 -17400
rect 13893 -17232 13990 -17216
rect 13893 -17400 13940 -17232
rect 13974 -17400 13990 -17232
rect 13893 -17416 13990 -17400
rect 12760 -17758 12857 -17742
rect 12760 -18526 12776 -17758
rect 12810 -18526 12857 -17758
rect 12760 -18542 12857 -18526
rect 13257 -17758 13354 -17742
rect 13257 -18526 13304 -17758
rect 13338 -18526 13354 -17758
rect 13257 -18542 13354 -18526
rect 13396 -17758 13493 -17742
rect 13396 -18526 13412 -17758
rect 13446 -18526 13493 -17758
rect 13396 -18542 13493 -18526
rect 13893 -17758 13990 -17742
rect 13893 -18526 13940 -17758
rect 13974 -18526 13990 -17758
rect 13893 -18542 13990 -18526
rect 14360 -17232 14457 -17216
rect 14360 -17400 14376 -17232
rect 14410 -17400 14457 -17232
rect 14360 -17416 14457 -17400
rect 14857 -17232 14954 -17216
rect 14857 -17400 14904 -17232
rect 14938 -17400 14954 -17232
rect 14857 -17416 14954 -17400
rect 14996 -17232 15093 -17216
rect 14996 -17400 15012 -17232
rect 15046 -17400 15093 -17232
rect 14996 -17416 15093 -17400
rect 15493 -17232 15590 -17216
rect 15493 -17400 15540 -17232
rect 15574 -17400 15590 -17232
rect 15493 -17416 15590 -17400
rect 14360 -17758 14457 -17742
rect 14360 -18526 14376 -17758
rect 14410 -18526 14457 -17758
rect 14360 -18542 14457 -18526
rect 14857 -17758 14954 -17742
rect 14857 -18526 14904 -17758
rect 14938 -18526 14954 -17758
rect 14857 -18542 14954 -18526
rect 14996 -17758 15093 -17742
rect 14996 -18526 15012 -17758
rect 15046 -18526 15093 -17758
rect 14996 -18542 15093 -18526
rect 15493 -17758 15590 -17742
rect 15493 -18526 15540 -17758
rect 15574 -18526 15590 -17758
rect 15493 -18542 15590 -18526
rect 15960 -17232 16057 -17216
rect 15960 -17400 15976 -17232
rect 16010 -17400 16057 -17232
rect 15960 -17416 16057 -17400
rect 16457 -17232 16554 -17216
rect 16457 -17400 16504 -17232
rect 16538 -17400 16554 -17232
rect 16457 -17416 16554 -17400
rect 16596 -17232 16693 -17216
rect 16596 -17400 16612 -17232
rect 16646 -17400 16693 -17232
rect 16596 -17416 16693 -17400
rect 17093 -17232 17190 -17216
rect 17093 -17400 17140 -17232
rect 17174 -17400 17190 -17232
rect 17093 -17416 17190 -17400
rect 15960 -17758 16057 -17742
rect 15960 -18526 15976 -17758
rect 16010 -18526 16057 -17758
rect 15960 -18542 16057 -18526
rect 16457 -17758 16554 -17742
rect 16457 -18526 16504 -17758
rect 16538 -18526 16554 -17758
rect 16457 -18542 16554 -18526
rect 16596 -17758 16693 -17742
rect 16596 -18526 16612 -17758
rect 16646 -18526 16693 -17758
rect 16596 -18542 16693 -18526
rect 17093 -17758 17190 -17742
rect 17093 -18526 17140 -17758
rect 17174 -18526 17190 -17758
rect 17093 -18542 17190 -18526
rect 17560 -17232 17657 -17216
rect 17560 -17400 17576 -17232
rect 17610 -17400 17657 -17232
rect 17560 -17416 17657 -17400
rect 18057 -17232 18154 -17216
rect 18057 -17400 18104 -17232
rect 18138 -17400 18154 -17232
rect 18057 -17416 18154 -17400
rect 18196 -17232 18293 -17216
rect 18196 -17400 18212 -17232
rect 18246 -17400 18293 -17232
rect 18196 -17416 18293 -17400
rect 18693 -17232 18790 -17216
rect 18693 -17400 18740 -17232
rect 18774 -17400 18790 -17232
rect 18693 -17416 18790 -17400
rect 17560 -17758 17657 -17742
rect 17560 -18526 17576 -17758
rect 17610 -18526 17657 -17758
rect 17560 -18542 17657 -18526
rect 18057 -17758 18154 -17742
rect 18057 -18526 18104 -17758
rect 18138 -18526 18154 -17758
rect 18057 -18542 18154 -18526
rect 18196 -17758 18293 -17742
rect 18196 -18526 18212 -17758
rect 18246 -18526 18293 -17758
rect 18196 -18542 18293 -18526
rect 18693 -17758 18790 -17742
rect 18693 -18526 18740 -17758
rect 18774 -18526 18790 -17758
rect 18693 -18542 18790 -18526
rect 19160 -17232 19257 -17216
rect 19160 -17400 19176 -17232
rect 19210 -17400 19257 -17232
rect 19160 -17416 19257 -17400
rect 19657 -17232 19754 -17216
rect 19657 -17400 19704 -17232
rect 19738 -17400 19754 -17232
rect 19657 -17416 19754 -17400
rect 19796 -17232 19893 -17216
rect 19796 -17400 19812 -17232
rect 19846 -17400 19893 -17232
rect 19796 -17416 19893 -17400
rect 20293 -17232 20390 -17216
rect 20293 -17400 20340 -17232
rect 20374 -17400 20390 -17232
rect 20293 -17416 20390 -17400
rect 19160 -17758 19257 -17742
rect 19160 -18526 19176 -17758
rect 19210 -18526 19257 -17758
rect 19160 -18542 19257 -18526
rect 19657 -17758 19754 -17742
rect 19657 -18526 19704 -17758
rect 19738 -18526 19754 -17758
rect 19657 -18542 19754 -18526
rect 19796 -17758 19893 -17742
rect 19796 -18526 19812 -17758
rect 19846 -18526 19893 -17758
rect 19796 -18542 19893 -18526
rect 20293 -17758 20390 -17742
rect 20293 -18526 20340 -17758
rect 20374 -18526 20390 -17758
rect 20293 -18542 20390 -18526
rect 20760 -17232 20857 -17216
rect 20760 -17400 20776 -17232
rect 20810 -17400 20857 -17232
rect 20760 -17416 20857 -17400
rect 21257 -17232 21354 -17216
rect 21257 -17400 21304 -17232
rect 21338 -17400 21354 -17232
rect 21257 -17416 21354 -17400
rect 21396 -17232 21493 -17216
rect 21396 -17400 21412 -17232
rect 21446 -17400 21493 -17232
rect 21396 -17416 21493 -17400
rect 21893 -17232 21990 -17216
rect 21893 -17400 21940 -17232
rect 21974 -17400 21990 -17232
rect 21893 -17416 21990 -17400
rect 20760 -17758 20857 -17742
rect 20760 -18526 20776 -17758
rect 20810 -18526 20857 -17758
rect 20760 -18542 20857 -18526
rect 21257 -17758 21354 -17742
rect 21257 -18526 21304 -17758
rect 21338 -18526 21354 -17758
rect 21257 -18542 21354 -18526
rect 21396 -17758 21493 -17742
rect 21396 -18526 21412 -17758
rect 21446 -18526 21493 -17758
rect 21396 -18542 21493 -18526
rect 21893 -17758 21990 -17742
rect 21893 -18526 21940 -17758
rect 21974 -18526 21990 -17758
rect 21893 -18542 21990 -18526
rect 22360 -17232 22457 -17216
rect 22360 -17400 22376 -17232
rect 22410 -17400 22457 -17232
rect 22360 -17416 22457 -17400
rect 22857 -17232 22954 -17216
rect 22857 -17400 22904 -17232
rect 22938 -17400 22954 -17232
rect 22857 -17416 22954 -17400
rect 22996 -17232 23093 -17216
rect 22996 -17400 23012 -17232
rect 23046 -17400 23093 -17232
rect 22996 -17416 23093 -17400
rect 23493 -17232 23590 -17216
rect 23493 -17400 23540 -17232
rect 23574 -17400 23590 -17232
rect 23493 -17416 23590 -17400
rect 22360 -17758 22457 -17742
rect 22360 -18526 22376 -17758
rect 22410 -18526 22457 -17758
rect 22360 -18542 22457 -18526
rect 22857 -17758 22954 -17742
rect 22857 -18526 22904 -17758
rect 22938 -18526 22954 -17758
rect 22857 -18542 22954 -18526
rect 22996 -17758 23093 -17742
rect 22996 -18526 23012 -17758
rect 23046 -18526 23093 -17758
rect 22996 -18542 23093 -18526
rect 23493 -17758 23590 -17742
rect 23493 -18526 23540 -17758
rect 23574 -18526 23590 -17758
rect 23493 -18542 23590 -18526
rect 23960 -17232 24057 -17216
rect 23960 -17400 23976 -17232
rect 24010 -17400 24057 -17232
rect 23960 -17416 24057 -17400
rect 24457 -17232 24554 -17216
rect 24457 -17400 24504 -17232
rect 24538 -17400 24554 -17232
rect 24457 -17416 24554 -17400
rect 24596 -17232 24693 -17216
rect 24596 -17400 24612 -17232
rect 24646 -17400 24693 -17232
rect 24596 -17416 24693 -17400
rect 25093 -17232 25190 -17216
rect 25093 -17400 25140 -17232
rect 25174 -17400 25190 -17232
rect 25093 -17416 25190 -17400
rect 23960 -17758 24057 -17742
rect 23960 -18526 23976 -17758
rect 24010 -18526 24057 -17758
rect 23960 -18542 24057 -18526
rect 24457 -17758 24554 -17742
rect 24457 -18526 24504 -17758
rect 24538 -18526 24554 -17758
rect 24457 -18542 24554 -18526
rect 24596 -17758 24693 -17742
rect 24596 -18526 24612 -17758
rect 24646 -18526 24693 -17758
rect 24596 -18542 24693 -18526
rect 25093 -17758 25190 -17742
rect 25093 -18526 25140 -17758
rect 25174 -18526 25190 -17758
rect 25093 -18542 25190 -18526
rect 25560 -17232 25657 -17216
rect 25560 -17400 25576 -17232
rect 25610 -17400 25657 -17232
rect 25560 -17416 25657 -17400
rect 26057 -17232 26154 -17216
rect 26057 -17400 26104 -17232
rect 26138 -17400 26154 -17232
rect 26057 -17416 26154 -17400
rect 26196 -17232 26293 -17216
rect 26196 -17400 26212 -17232
rect 26246 -17400 26293 -17232
rect 26196 -17416 26293 -17400
rect 26693 -17232 26790 -17216
rect 26693 -17400 26740 -17232
rect 26774 -17400 26790 -17232
rect 26693 -17416 26790 -17400
rect 25560 -17758 25657 -17742
rect 25560 -18526 25576 -17758
rect 25610 -18526 25657 -17758
rect 25560 -18542 25657 -18526
rect 26057 -17758 26154 -17742
rect 26057 -18526 26104 -17758
rect 26138 -18526 26154 -17758
rect 26057 -18542 26154 -18526
rect 26196 -17758 26293 -17742
rect 26196 -18526 26212 -17758
rect 26246 -18526 26293 -17758
rect 26196 -18542 26293 -18526
rect 26693 -17758 26790 -17742
rect 26693 -18526 26740 -17758
rect 26774 -18526 26790 -17758
rect 26693 -18542 26790 -18526
rect 27160 -17232 27257 -17216
rect 27160 -17400 27176 -17232
rect 27210 -17400 27257 -17232
rect 27160 -17416 27257 -17400
rect 27657 -17232 27754 -17216
rect 27657 -17400 27704 -17232
rect 27738 -17400 27754 -17232
rect 27657 -17416 27754 -17400
rect 27796 -17232 27893 -17216
rect 27796 -17400 27812 -17232
rect 27846 -17400 27893 -17232
rect 27796 -17416 27893 -17400
rect 28293 -17232 28390 -17216
rect 28293 -17400 28340 -17232
rect 28374 -17400 28390 -17232
rect 28293 -17416 28390 -17400
rect 27160 -17758 27257 -17742
rect 27160 -18526 27176 -17758
rect 27210 -18526 27257 -17758
rect 27160 -18542 27257 -18526
rect 27657 -17758 27754 -17742
rect 27657 -18526 27704 -17758
rect 27738 -18526 27754 -17758
rect 27657 -18542 27754 -18526
rect 27796 -17758 27893 -17742
rect 27796 -18526 27812 -17758
rect 27846 -18526 27893 -17758
rect 27796 -18542 27893 -18526
rect 28293 -17758 28390 -17742
rect 28293 -18526 28340 -17758
rect 28374 -18526 28390 -17758
rect 28293 -18542 28390 -18526
rect 28760 -17232 28857 -17216
rect 28760 -17400 28776 -17232
rect 28810 -17400 28857 -17232
rect 28760 -17416 28857 -17400
rect 29257 -17232 29354 -17216
rect 29257 -17400 29304 -17232
rect 29338 -17400 29354 -17232
rect 29257 -17416 29354 -17400
rect 29396 -17232 29493 -17216
rect 29396 -17400 29412 -17232
rect 29446 -17400 29493 -17232
rect 29396 -17416 29493 -17400
rect 29893 -17232 29990 -17216
rect 29893 -17400 29940 -17232
rect 29974 -17400 29990 -17232
rect 29893 -17416 29990 -17400
rect 28760 -17758 28857 -17742
rect 28760 -18526 28776 -17758
rect 28810 -18526 28857 -17758
rect 28760 -18542 28857 -18526
rect 29257 -17758 29354 -17742
rect 29257 -18526 29304 -17758
rect 29338 -18526 29354 -17758
rect 29257 -18542 29354 -18526
rect 29396 -17758 29493 -17742
rect 29396 -18526 29412 -17758
rect 29446 -18526 29493 -17758
rect 29396 -18542 29493 -18526
rect 29893 -17758 29990 -17742
rect 29893 -18526 29940 -17758
rect 29974 -18526 29990 -17758
rect 29893 -18542 29990 -18526
rect 30360 -17232 30457 -17216
rect 30360 -17400 30376 -17232
rect 30410 -17400 30457 -17232
rect 30360 -17416 30457 -17400
rect 30857 -17232 30954 -17216
rect 30857 -17400 30904 -17232
rect 30938 -17400 30954 -17232
rect 30857 -17416 30954 -17400
rect 30996 -17232 31093 -17216
rect 30996 -17400 31012 -17232
rect 31046 -17400 31093 -17232
rect 30996 -17416 31093 -17400
rect 31493 -17232 31590 -17216
rect 31493 -17400 31540 -17232
rect 31574 -17400 31590 -17232
rect 31493 -17416 31590 -17400
rect 30360 -17758 30457 -17742
rect 30360 -18526 30376 -17758
rect 30410 -18526 30457 -17758
rect 30360 -18542 30457 -18526
rect 30857 -17758 30954 -17742
rect 30857 -18526 30904 -17758
rect 30938 -18526 30954 -17758
rect 30857 -18542 30954 -18526
rect 30996 -17758 31093 -17742
rect 30996 -18526 31012 -17758
rect 31046 -18526 31093 -17758
rect 30996 -18542 31093 -18526
rect 31493 -17758 31590 -17742
rect 31493 -18526 31540 -17758
rect 31574 -18526 31590 -17758
rect 31493 -18542 31590 -18526
rect 31960 -17232 32057 -17216
rect 31960 -17400 31976 -17232
rect 32010 -17400 32057 -17232
rect 31960 -17416 32057 -17400
rect 32457 -17232 32554 -17216
rect 32457 -17400 32504 -17232
rect 32538 -17400 32554 -17232
rect 32457 -17416 32554 -17400
rect 32596 -17232 32693 -17216
rect 32596 -17400 32612 -17232
rect 32646 -17400 32693 -17232
rect 32596 -17416 32693 -17400
rect 33093 -17232 33190 -17216
rect 33093 -17400 33140 -17232
rect 33174 -17400 33190 -17232
rect 33093 -17416 33190 -17400
rect 31960 -17758 32057 -17742
rect 31960 -18526 31976 -17758
rect 32010 -18526 32057 -17758
rect 31960 -18542 32057 -18526
rect 32457 -17758 32554 -17742
rect 32457 -18526 32504 -17758
rect 32538 -18526 32554 -17758
rect 32457 -18542 32554 -18526
rect 32596 -17758 32693 -17742
rect 32596 -18526 32612 -17758
rect 32646 -18526 32693 -17758
rect 32596 -18542 32693 -18526
rect 33093 -17758 33190 -17742
rect 33093 -18526 33140 -17758
rect 33174 -18526 33190 -17758
rect 33093 -18542 33190 -18526
rect 33560 -17232 33657 -17216
rect 33560 -17400 33576 -17232
rect 33610 -17400 33657 -17232
rect 33560 -17416 33657 -17400
rect 34057 -17232 34154 -17216
rect 34057 -17400 34104 -17232
rect 34138 -17400 34154 -17232
rect 34057 -17416 34154 -17400
rect 34196 -17232 34293 -17216
rect 34196 -17400 34212 -17232
rect 34246 -17400 34293 -17232
rect 34196 -17416 34293 -17400
rect 34693 -17232 34790 -17216
rect 34693 -17400 34740 -17232
rect 34774 -17400 34790 -17232
rect 34693 -17416 34790 -17400
rect 33560 -17758 33657 -17742
rect 33560 -18526 33576 -17758
rect 33610 -18526 33657 -17758
rect 33560 -18542 33657 -18526
rect 34057 -17758 34154 -17742
rect 34057 -18526 34104 -17758
rect 34138 -18526 34154 -17758
rect 34057 -18542 34154 -18526
rect 34196 -17758 34293 -17742
rect 34196 -18526 34212 -17758
rect 34246 -18526 34293 -17758
rect 34196 -18542 34293 -18526
rect 34693 -17758 34790 -17742
rect 34693 -18526 34740 -17758
rect 34774 -18526 34790 -17758
rect 34693 -18542 34790 -18526
rect 35160 -17232 35257 -17216
rect 35160 -17400 35176 -17232
rect 35210 -17400 35257 -17232
rect 35160 -17416 35257 -17400
rect 35657 -17232 35754 -17216
rect 35657 -17400 35704 -17232
rect 35738 -17400 35754 -17232
rect 35657 -17416 35754 -17400
rect 35796 -17232 35893 -17216
rect 35796 -17400 35812 -17232
rect 35846 -17400 35893 -17232
rect 35796 -17416 35893 -17400
rect 36293 -17232 36390 -17216
rect 36293 -17400 36340 -17232
rect 36374 -17400 36390 -17232
rect 36293 -17416 36390 -17400
rect 35160 -17758 35257 -17742
rect 35160 -18526 35176 -17758
rect 35210 -18526 35257 -17758
rect 35160 -18542 35257 -18526
rect 35657 -17758 35754 -17742
rect 35657 -18526 35704 -17758
rect 35738 -18526 35754 -17758
rect 35657 -18542 35754 -18526
rect 35796 -17758 35893 -17742
rect 35796 -18526 35812 -17758
rect 35846 -18526 35893 -17758
rect 35796 -18542 35893 -18526
rect 36293 -17758 36390 -17742
rect 36293 -18526 36340 -17758
rect 36374 -18526 36390 -17758
rect 36293 -18542 36390 -18526
rect 36760 -17232 36857 -17216
rect 36760 -17400 36776 -17232
rect 36810 -17400 36857 -17232
rect 36760 -17416 36857 -17400
rect 37257 -17232 37354 -17216
rect 37257 -17400 37304 -17232
rect 37338 -17400 37354 -17232
rect 37257 -17416 37354 -17400
rect 37396 -17232 37493 -17216
rect 37396 -17400 37412 -17232
rect 37446 -17400 37493 -17232
rect 37396 -17416 37493 -17400
rect 37893 -17232 37990 -17216
rect 37893 -17400 37940 -17232
rect 37974 -17400 37990 -17232
rect 37893 -17416 37990 -17400
rect 36760 -17758 36857 -17742
rect 36760 -18526 36776 -17758
rect 36810 -18526 36857 -17758
rect 36760 -18542 36857 -18526
rect 37257 -17758 37354 -17742
rect 37257 -18526 37304 -17758
rect 37338 -18526 37354 -17758
rect 37257 -18542 37354 -18526
rect 37396 -17758 37493 -17742
rect 37396 -18526 37412 -17758
rect 37446 -18526 37493 -17758
rect 37396 -18542 37493 -18526
rect 37893 -17758 37990 -17742
rect 37893 -18526 37940 -17758
rect 37974 -18526 37990 -17758
rect 37893 -18542 37990 -18526
rect -40 -19032 57 -19016
rect -40 -19200 -24 -19032
rect 10 -19200 57 -19032
rect -40 -19216 57 -19200
rect 457 -19032 554 -19016
rect 457 -19200 504 -19032
rect 538 -19200 554 -19032
rect 457 -19216 554 -19200
rect 596 -19032 693 -19016
rect 596 -19200 612 -19032
rect 646 -19200 693 -19032
rect 596 -19216 693 -19200
rect 1093 -19032 1190 -19016
rect 1093 -19200 1140 -19032
rect 1174 -19200 1190 -19032
rect 1093 -19216 1190 -19200
rect -40 -19558 57 -19542
rect -40 -20326 -24 -19558
rect 10 -20326 57 -19558
rect -40 -20342 57 -20326
rect 457 -19558 554 -19542
rect 457 -20326 504 -19558
rect 538 -20326 554 -19558
rect 457 -20342 554 -20326
rect 596 -19558 693 -19542
rect 596 -20326 612 -19558
rect 646 -20326 693 -19558
rect 596 -20342 693 -20326
rect 1093 -19558 1190 -19542
rect 1093 -20326 1140 -19558
rect 1174 -20326 1190 -19558
rect 1093 -20342 1190 -20326
rect 1560 -19032 1657 -19016
rect 1560 -19200 1576 -19032
rect 1610 -19200 1657 -19032
rect 1560 -19216 1657 -19200
rect 2057 -19032 2154 -19016
rect 2057 -19200 2104 -19032
rect 2138 -19200 2154 -19032
rect 2057 -19216 2154 -19200
rect 2196 -19032 2293 -19016
rect 2196 -19200 2212 -19032
rect 2246 -19200 2293 -19032
rect 2196 -19216 2293 -19200
rect 2693 -19032 2790 -19016
rect 2693 -19200 2740 -19032
rect 2774 -19200 2790 -19032
rect 2693 -19216 2790 -19200
rect 1560 -19558 1657 -19542
rect 1560 -20326 1576 -19558
rect 1610 -20326 1657 -19558
rect 1560 -20342 1657 -20326
rect 2057 -19558 2154 -19542
rect 2057 -20326 2104 -19558
rect 2138 -20326 2154 -19558
rect 2057 -20342 2154 -20326
rect 2196 -19558 2293 -19542
rect 2196 -20326 2212 -19558
rect 2246 -20326 2293 -19558
rect 2196 -20342 2293 -20326
rect 2693 -19558 2790 -19542
rect 2693 -20326 2740 -19558
rect 2774 -20326 2790 -19558
rect 2693 -20342 2790 -20326
rect 3160 -19032 3257 -19016
rect 3160 -19200 3176 -19032
rect 3210 -19200 3257 -19032
rect 3160 -19216 3257 -19200
rect 3657 -19032 3754 -19016
rect 3657 -19200 3704 -19032
rect 3738 -19200 3754 -19032
rect 3657 -19216 3754 -19200
rect 3796 -19032 3893 -19016
rect 3796 -19200 3812 -19032
rect 3846 -19200 3893 -19032
rect 3796 -19216 3893 -19200
rect 4293 -19032 4390 -19016
rect 4293 -19200 4340 -19032
rect 4374 -19200 4390 -19032
rect 4293 -19216 4390 -19200
rect 3160 -19558 3257 -19542
rect 3160 -20326 3176 -19558
rect 3210 -20326 3257 -19558
rect 3160 -20342 3257 -20326
rect 3657 -19558 3754 -19542
rect 3657 -20326 3704 -19558
rect 3738 -20326 3754 -19558
rect 3657 -20342 3754 -20326
rect 3796 -19558 3893 -19542
rect 3796 -20326 3812 -19558
rect 3846 -20326 3893 -19558
rect 3796 -20342 3893 -20326
rect 4293 -19558 4390 -19542
rect 4293 -20326 4340 -19558
rect 4374 -20326 4390 -19558
rect 4293 -20342 4390 -20326
rect 4760 -19032 4857 -19016
rect 4760 -19200 4776 -19032
rect 4810 -19200 4857 -19032
rect 4760 -19216 4857 -19200
rect 5257 -19032 5354 -19016
rect 5257 -19200 5304 -19032
rect 5338 -19200 5354 -19032
rect 5257 -19216 5354 -19200
rect 5396 -19032 5493 -19016
rect 5396 -19200 5412 -19032
rect 5446 -19200 5493 -19032
rect 5396 -19216 5493 -19200
rect 5893 -19032 5990 -19016
rect 5893 -19200 5940 -19032
rect 5974 -19200 5990 -19032
rect 5893 -19216 5990 -19200
rect 4760 -19558 4857 -19542
rect 4760 -20326 4776 -19558
rect 4810 -20326 4857 -19558
rect 4760 -20342 4857 -20326
rect 5257 -19558 5354 -19542
rect 5257 -20326 5304 -19558
rect 5338 -20326 5354 -19558
rect 5257 -20342 5354 -20326
rect 5396 -19558 5493 -19542
rect 5396 -20326 5412 -19558
rect 5446 -20326 5493 -19558
rect 5396 -20342 5493 -20326
rect 5893 -19558 5990 -19542
rect 5893 -20326 5940 -19558
rect 5974 -20326 5990 -19558
rect 5893 -20342 5990 -20326
rect 6360 -19032 6457 -19016
rect 6360 -19200 6376 -19032
rect 6410 -19200 6457 -19032
rect 6360 -19216 6457 -19200
rect 6857 -19032 6954 -19016
rect 6857 -19200 6904 -19032
rect 6938 -19200 6954 -19032
rect 6857 -19216 6954 -19200
rect 6996 -19032 7093 -19016
rect 6996 -19200 7012 -19032
rect 7046 -19200 7093 -19032
rect 6996 -19216 7093 -19200
rect 7493 -19032 7590 -19016
rect 7493 -19200 7540 -19032
rect 7574 -19200 7590 -19032
rect 7493 -19216 7590 -19200
rect 6360 -19558 6457 -19542
rect 6360 -20326 6376 -19558
rect 6410 -20326 6457 -19558
rect 6360 -20342 6457 -20326
rect 6857 -19558 6954 -19542
rect 6857 -20326 6904 -19558
rect 6938 -20326 6954 -19558
rect 6857 -20342 6954 -20326
rect 6996 -19558 7093 -19542
rect 6996 -20326 7012 -19558
rect 7046 -20326 7093 -19558
rect 6996 -20342 7093 -20326
rect 7493 -19558 7590 -19542
rect 7493 -20326 7540 -19558
rect 7574 -20326 7590 -19558
rect 7493 -20342 7590 -20326
rect 7960 -19032 8057 -19016
rect 7960 -19200 7976 -19032
rect 8010 -19200 8057 -19032
rect 7960 -19216 8057 -19200
rect 8457 -19032 8554 -19016
rect 8457 -19200 8504 -19032
rect 8538 -19200 8554 -19032
rect 8457 -19216 8554 -19200
rect 8596 -19032 8693 -19016
rect 8596 -19200 8612 -19032
rect 8646 -19200 8693 -19032
rect 8596 -19216 8693 -19200
rect 9093 -19032 9190 -19016
rect 9093 -19200 9140 -19032
rect 9174 -19200 9190 -19032
rect 9093 -19216 9190 -19200
rect 7960 -19558 8057 -19542
rect 7960 -20326 7976 -19558
rect 8010 -20326 8057 -19558
rect 7960 -20342 8057 -20326
rect 8457 -19558 8554 -19542
rect 8457 -20326 8504 -19558
rect 8538 -20326 8554 -19558
rect 8457 -20342 8554 -20326
rect 8596 -19558 8693 -19542
rect 8596 -20326 8612 -19558
rect 8646 -20326 8693 -19558
rect 8596 -20342 8693 -20326
rect 9093 -19558 9190 -19542
rect 9093 -20326 9140 -19558
rect 9174 -20326 9190 -19558
rect 9093 -20342 9190 -20326
rect 9560 -19032 9657 -19016
rect 9560 -19200 9576 -19032
rect 9610 -19200 9657 -19032
rect 9560 -19216 9657 -19200
rect 10057 -19032 10154 -19016
rect 10057 -19200 10104 -19032
rect 10138 -19200 10154 -19032
rect 10057 -19216 10154 -19200
rect 10196 -19032 10293 -19016
rect 10196 -19200 10212 -19032
rect 10246 -19200 10293 -19032
rect 10196 -19216 10293 -19200
rect 10693 -19032 10790 -19016
rect 10693 -19200 10740 -19032
rect 10774 -19200 10790 -19032
rect 10693 -19216 10790 -19200
rect 9560 -19558 9657 -19542
rect 9560 -20326 9576 -19558
rect 9610 -20326 9657 -19558
rect 9560 -20342 9657 -20326
rect 10057 -19558 10154 -19542
rect 10057 -20326 10104 -19558
rect 10138 -20326 10154 -19558
rect 10057 -20342 10154 -20326
rect 10196 -19558 10293 -19542
rect 10196 -20326 10212 -19558
rect 10246 -20326 10293 -19558
rect 10196 -20342 10293 -20326
rect 10693 -19558 10790 -19542
rect 10693 -20326 10740 -19558
rect 10774 -20326 10790 -19558
rect 10693 -20342 10790 -20326
rect 11160 -19032 11257 -19016
rect 11160 -19200 11176 -19032
rect 11210 -19200 11257 -19032
rect 11160 -19216 11257 -19200
rect 11657 -19032 11754 -19016
rect 11657 -19200 11704 -19032
rect 11738 -19200 11754 -19032
rect 11657 -19216 11754 -19200
rect 11796 -19032 11893 -19016
rect 11796 -19200 11812 -19032
rect 11846 -19200 11893 -19032
rect 11796 -19216 11893 -19200
rect 12293 -19032 12390 -19016
rect 12293 -19200 12340 -19032
rect 12374 -19200 12390 -19032
rect 12293 -19216 12390 -19200
rect 11160 -19558 11257 -19542
rect 11160 -20326 11176 -19558
rect 11210 -20326 11257 -19558
rect 11160 -20342 11257 -20326
rect 11657 -19558 11754 -19542
rect 11657 -20326 11704 -19558
rect 11738 -20326 11754 -19558
rect 11657 -20342 11754 -20326
rect 11796 -19558 11893 -19542
rect 11796 -20326 11812 -19558
rect 11846 -20326 11893 -19558
rect 11796 -20342 11893 -20326
rect 12293 -19558 12390 -19542
rect 12293 -20326 12340 -19558
rect 12374 -20326 12390 -19558
rect 12293 -20342 12390 -20326
rect 12760 -19032 12857 -19016
rect 12760 -19200 12776 -19032
rect 12810 -19200 12857 -19032
rect 12760 -19216 12857 -19200
rect 13257 -19032 13354 -19016
rect 13257 -19200 13304 -19032
rect 13338 -19200 13354 -19032
rect 13257 -19216 13354 -19200
rect 13396 -19032 13493 -19016
rect 13396 -19200 13412 -19032
rect 13446 -19200 13493 -19032
rect 13396 -19216 13493 -19200
rect 13893 -19032 13990 -19016
rect 13893 -19200 13940 -19032
rect 13974 -19200 13990 -19032
rect 13893 -19216 13990 -19200
rect 12760 -19558 12857 -19542
rect 12760 -20326 12776 -19558
rect 12810 -20326 12857 -19558
rect 12760 -20342 12857 -20326
rect 13257 -19558 13354 -19542
rect 13257 -20326 13304 -19558
rect 13338 -20326 13354 -19558
rect 13257 -20342 13354 -20326
rect 13396 -19558 13493 -19542
rect 13396 -20326 13412 -19558
rect 13446 -20326 13493 -19558
rect 13396 -20342 13493 -20326
rect 13893 -19558 13990 -19542
rect 13893 -20326 13940 -19558
rect 13974 -20326 13990 -19558
rect 13893 -20342 13990 -20326
rect 14360 -19032 14457 -19016
rect 14360 -19200 14376 -19032
rect 14410 -19200 14457 -19032
rect 14360 -19216 14457 -19200
rect 14857 -19032 14954 -19016
rect 14857 -19200 14904 -19032
rect 14938 -19200 14954 -19032
rect 14857 -19216 14954 -19200
rect 14996 -19032 15093 -19016
rect 14996 -19200 15012 -19032
rect 15046 -19200 15093 -19032
rect 14996 -19216 15093 -19200
rect 15493 -19032 15590 -19016
rect 15493 -19200 15540 -19032
rect 15574 -19200 15590 -19032
rect 15493 -19216 15590 -19200
rect 14360 -19558 14457 -19542
rect 14360 -20326 14376 -19558
rect 14410 -20326 14457 -19558
rect 14360 -20342 14457 -20326
rect 14857 -19558 14954 -19542
rect 14857 -20326 14904 -19558
rect 14938 -20326 14954 -19558
rect 14857 -20342 14954 -20326
rect 14996 -19558 15093 -19542
rect 14996 -20326 15012 -19558
rect 15046 -20326 15093 -19558
rect 14996 -20342 15093 -20326
rect 15493 -19558 15590 -19542
rect 15493 -20326 15540 -19558
rect 15574 -20326 15590 -19558
rect 15493 -20342 15590 -20326
rect 15960 -19032 16057 -19016
rect 15960 -19200 15976 -19032
rect 16010 -19200 16057 -19032
rect 15960 -19216 16057 -19200
rect 16457 -19032 16554 -19016
rect 16457 -19200 16504 -19032
rect 16538 -19200 16554 -19032
rect 16457 -19216 16554 -19200
rect 16596 -19032 16693 -19016
rect 16596 -19200 16612 -19032
rect 16646 -19200 16693 -19032
rect 16596 -19216 16693 -19200
rect 17093 -19032 17190 -19016
rect 17093 -19200 17140 -19032
rect 17174 -19200 17190 -19032
rect 17093 -19216 17190 -19200
rect 15960 -19558 16057 -19542
rect 15960 -20326 15976 -19558
rect 16010 -20326 16057 -19558
rect 15960 -20342 16057 -20326
rect 16457 -19558 16554 -19542
rect 16457 -20326 16504 -19558
rect 16538 -20326 16554 -19558
rect 16457 -20342 16554 -20326
rect 16596 -19558 16693 -19542
rect 16596 -20326 16612 -19558
rect 16646 -20326 16693 -19558
rect 16596 -20342 16693 -20326
rect 17093 -19558 17190 -19542
rect 17093 -20326 17140 -19558
rect 17174 -20326 17190 -19558
rect 17093 -20342 17190 -20326
rect 17560 -19032 17657 -19016
rect 17560 -19200 17576 -19032
rect 17610 -19200 17657 -19032
rect 17560 -19216 17657 -19200
rect 18057 -19032 18154 -19016
rect 18057 -19200 18104 -19032
rect 18138 -19200 18154 -19032
rect 18057 -19216 18154 -19200
rect 18196 -19032 18293 -19016
rect 18196 -19200 18212 -19032
rect 18246 -19200 18293 -19032
rect 18196 -19216 18293 -19200
rect 18693 -19032 18790 -19016
rect 18693 -19200 18740 -19032
rect 18774 -19200 18790 -19032
rect 18693 -19216 18790 -19200
rect 17560 -19558 17657 -19542
rect 17560 -20326 17576 -19558
rect 17610 -20326 17657 -19558
rect 17560 -20342 17657 -20326
rect 18057 -19558 18154 -19542
rect 18057 -20326 18104 -19558
rect 18138 -20326 18154 -19558
rect 18057 -20342 18154 -20326
rect 18196 -19558 18293 -19542
rect 18196 -20326 18212 -19558
rect 18246 -20326 18293 -19558
rect 18196 -20342 18293 -20326
rect 18693 -19558 18790 -19542
rect 18693 -20326 18740 -19558
rect 18774 -20326 18790 -19558
rect 18693 -20342 18790 -20326
rect 19160 -19032 19257 -19016
rect 19160 -19200 19176 -19032
rect 19210 -19200 19257 -19032
rect 19160 -19216 19257 -19200
rect 19657 -19032 19754 -19016
rect 19657 -19200 19704 -19032
rect 19738 -19200 19754 -19032
rect 19657 -19216 19754 -19200
rect 19796 -19032 19893 -19016
rect 19796 -19200 19812 -19032
rect 19846 -19200 19893 -19032
rect 19796 -19216 19893 -19200
rect 20293 -19032 20390 -19016
rect 20293 -19200 20340 -19032
rect 20374 -19200 20390 -19032
rect 20293 -19216 20390 -19200
rect 19160 -19558 19257 -19542
rect 19160 -20326 19176 -19558
rect 19210 -20326 19257 -19558
rect 19160 -20342 19257 -20326
rect 19657 -19558 19754 -19542
rect 19657 -20326 19704 -19558
rect 19738 -20326 19754 -19558
rect 19657 -20342 19754 -20326
rect 19796 -19558 19893 -19542
rect 19796 -20326 19812 -19558
rect 19846 -20326 19893 -19558
rect 19796 -20342 19893 -20326
rect 20293 -19558 20390 -19542
rect 20293 -20326 20340 -19558
rect 20374 -20326 20390 -19558
rect 20293 -20342 20390 -20326
rect 20760 -19032 20857 -19016
rect 20760 -19200 20776 -19032
rect 20810 -19200 20857 -19032
rect 20760 -19216 20857 -19200
rect 21257 -19032 21354 -19016
rect 21257 -19200 21304 -19032
rect 21338 -19200 21354 -19032
rect 21257 -19216 21354 -19200
rect 21396 -19032 21493 -19016
rect 21396 -19200 21412 -19032
rect 21446 -19200 21493 -19032
rect 21396 -19216 21493 -19200
rect 21893 -19032 21990 -19016
rect 21893 -19200 21940 -19032
rect 21974 -19200 21990 -19032
rect 21893 -19216 21990 -19200
rect 20760 -19558 20857 -19542
rect 20760 -20326 20776 -19558
rect 20810 -20326 20857 -19558
rect 20760 -20342 20857 -20326
rect 21257 -19558 21354 -19542
rect 21257 -20326 21304 -19558
rect 21338 -20326 21354 -19558
rect 21257 -20342 21354 -20326
rect 21396 -19558 21493 -19542
rect 21396 -20326 21412 -19558
rect 21446 -20326 21493 -19558
rect 21396 -20342 21493 -20326
rect 21893 -19558 21990 -19542
rect 21893 -20326 21940 -19558
rect 21974 -20326 21990 -19558
rect 21893 -20342 21990 -20326
rect 22360 -19032 22457 -19016
rect 22360 -19200 22376 -19032
rect 22410 -19200 22457 -19032
rect 22360 -19216 22457 -19200
rect 22857 -19032 22954 -19016
rect 22857 -19200 22904 -19032
rect 22938 -19200 22954 -19032
rect 22857 -19216 22954 -19200
rect 22996 -19032 23093 -19016
rect 22996 -19200 23012 -19032
rect 23046 -19200 23093 -19032
rect 22996 -19216 23093 -19200
rect 23493 -19032 23590 -19016
rect 23493 -19200 23540 -19032
rect 23574 -19200 23590 -19032
rect 23493 -19216 23590 -19200
rect 22360 -19558 22457 -19542
rect 22360 -20326 22376 -19558
rect 22410 -20326 22457 -19558
rect 22360 -20342 22457 -20326
rect 22857 -19558 22954 -19542
rect 22857 -20326 22904 -19558
rect 22938 -20326 22954 -19558
rect 22857 -20342 22954 -20326
rect 22996 -19558 23093 -19542
rect 22996 -20326 23012 -19558
rect 23046 -20326 23093 -19558
rect 22996 -20342 23093 -20326
rect 23493 -19558 23590 -19542
rect 23493 -20326 23540 -19558
rect 23574 -20326 23590 -19558
rect 23493 -20342 23590 -20326
rect 23960 -19032 24057 -19016
rect 23960 -19200 23976 -19032
rect 24010 -19200 24057 -19032
rect 23960 -19216 24057 -19200
rect 24457 -19032 24554 -19016
rect 24457 -19200 24504 -19032
rect 24538 -19200 24554 -19032
rect 24457 -19216 24554 -19200
rect 24596 -19032 24693 -19016
rect 24596 -19200 24612 -19032
rect 24646 -19200 24693 -19032
rect 24596 -19216 24693 -19200
rect 25093 -19032 25190 -19016
rect 25093 -19200 25140 -19032
rect 25174 -19200 25190 -19032
rect 25093 -19216 25190 -19200
rect 23960 -19558 24057 -19542
rect 23960 -20326 23976 -19558
rect 24010 -20326 24057 -19558
rect 23960 -20342 24057 -20326
rect 24457 -19558 24554 -19542
rect 24457 -20326 24504 -19558
rect 24538 -20326 24554 -19558
rect 24457 -20342 24554 -20326
rect 24596 -19558 24693 -19542
rect 24596 -20326 24612 -19558
rect 24646 -20326 24693 -19558
rect 24596 -20342 24693 -20326
rect 25093 -19558 25190 -19542
rect 25093 -20326 25140 -19558
rect 25174 -20326 25190 -19558
rect 25093 -20342 25190 -20326
rect 25560 -19032 25657 -19016
rect 25560 -19200 25576 -19032
rect 25610 -19200 25657 -19032
rect 25560 -19216 25657 -19200
rect 26057 -19032 26154 -19016
rect 26057 -19200 26104 -19032
rect 26138 -19200 26154 -19032
rect 26057 -19216 26154 -19200
rect 26196 -19032 26293 -19016
rect 26196 -19200 26212 -19032
rect 26246 -19200 26293 -19032
rect 26196 -19216 26293 -19200
rect 26693 -19032 26790 -19016
rect 26693 -19200 26740 -19032
rect 26774 -19200 26790 -19032
rect 26693 -19216 26790 -19200
rect 25560 -19558 25657 -19542
rect 25560 -20326 25576 -19558
rect 25610 -20326 25657 -19558
rect 25560 -20342 25657 -20326
rect 26057 -19558 26154 -19542
rect 26057 -20326 26104 -19558
rect 26138 -20326 26154 -19558
rect 26057 -20342 26154 -20326
rect 26196 -19558 26293 -19542
rect 26196 -20326 26212 -19558
rect 26246 -20326 26293 -19558
rect 26196 -20342 26293 -20326
rect 26693 -19558 26790 -19542
rect 26693 -20326 26740 -19558
rect 26774 -20326 26790 -19558
rect 26693 -20342 26790 -20326
rect 27160 -19032 27257 -19016
rect 27160 -19200 27176 -19032
rect 27210 -19200 27257 -19032
rect 27160 -19216 27257 -19200
rect 27657 -19032 27754 -19016
rect 27657 -19200 27704 -19032
rect 27738 -19200 27754 -19032
rect 27657 -19216 27754 -19200
rect 27796 -19032 27893 -19016
rect 27796 -19200 27812 -19032
rect 27846 -19200 27893 -19032
rect 27796 -19216 27893 -19200
rect 28293 -19032 28390 -19016
rect 28293 -19200 28340 -19032
rect 28374 -19200 28390 -19032
rect 28293 -19216 28390 -19200
rect 27160 -19558 27257 -19542
rect 27160 -20326 27176 -19558
rect 27210 -20326 27257 -19558
rect 27160 -20342 27257 -20326
rect 27657 -19558 27754 -19542
rect 27657 -20326 27704 -19558
rect 27738 -20326 27754 -19558
rect 27657 -20342 27754 -20326
rect 27796 -19558 27893 -19542
rect 27796 -20326 27812 -19558
rect 27846 -20326 27893 -19558
rect 27796 -20342 27893 -20326
rect 28293 -19558 28390 -19542
rect 28293 -20326 28340 -19558
rect 28374 -20326 28390 -19558
rect 28293 -20342 28390 -20326
rect 28760 -19032 28857 -19016
rect 28760 -19200 28776 -19032
rect 28810 -19200 28857 -19032
rect 28760 -19216 28857 -19200
rect 29257 -19032 29354 -19016
rect 29257 -19200 29304 -19032
rect 29338 -19200 29354 -19032
rect 29257 -19216 29354 -19200
rect 29396 -19032 29493 -19016
rect 29396 -19200 29412 -19032
rect 29446 -19200 29493 -19032
rect 29396 -19216 29493 -19200
rect 29893 -19032 29990 -19016
rect 29893 -19200 29940 -19032
rect 29974 -19200 29990 -19032
rect 29893 -19216 29990 -19200
rect 28760 -19558 28857 -19542
rect 28760 -20326 28776 -19558
rect 28810 -20326 28857 -19558
rect 28760 -20342 28857 -20326
rect 29257 -19558 29354 -19542
rect 29257 -20326 29304 -19558
rect 29338 -20326 29354 -19558
rect 29257 -20342 29354 -20326
rect 29396 -19558 29493 -19542
rect 29396 -20326 29412 -19558
rect 29446 -20326 29493 -19558
rect 29396 -20342 29493 -20326
rect 29893 -19558 29990 -19542
rect 29893 -20326 29940 -19558
rect 29974 -20326 29990 -19558
rect 29893 -20342 29990 -20326
rect 30360 -19032 30457 -19016
rect 30360 -19200 30376 -19032
rect 30410 -19200 30457 -19032
rect 30360 -19216 30457 -19200
rect 30857 -19032 30954 -19016
rect 30857 -19200 30904 -19032
rect 30938 -19200 30954 -19032
rect 30857 -19216 30954 -19200
rect 30996 -19032 31093 -19016
rect 30996 -19200 31012 -19032
rect 31046 -19200 31093 -19032
rect 30996 -19216 31093 -19200
rect 31493 -19032 31590 -19016
rect 31493 -19200 31540 -19032
rect 31574 -19200 31590 -19032
rect 31493 -19216 31590 -19200
rect 30360 -19558 30457 -19542
rect 30360 -20326 30376 -19558
rect 30410 -20326 30457 -19558
rect 30360 -20342 30457 -20326
rect 30857 -19558 30954 -19542
rect 30857 -20326 30904 -19558
rect 30938 -20326 30954 -19558
rect 30857 -20342 30954 -20326
rect 30996 -19558 31093 -19542
rect 30996 -20326 31012 -19558
rect 31046 -20326 31093 -19558
rect 30996 -20342 31093 -20326
rect 31493 -19558 31590 -19542
rect 31493 -20326 31540 -19558
rect 31574 -20326 31590 -19558
rect 31493 -20342 31590 -20326
rect 31960 -19032 32057 -19016
rect 31960 -19200 31976 -19032
rect 32010 -19200 32057 -19032
rect 31960 -19216 32057 -19200
rect 32457 -19032 32554 -19016
rect 32457 -19200 32504 -19032
rect 32538 -19200 32554 -19032
rect 32457 -19216 32554 -19200
rect 32596 -19032 32693 -19016
rect 32596 -19200 32612 -19032
rect 32646 -19200 32693 -19032
rect 32596 -19216 32693 -19200
rect 33093 -19032 33190 -19016
rect 33093 -19200 33140 -19032
rect 33174 -19200 33190 -19032
rect 33093 -19216 33190 -19200
rect 31960 -19558 32057 -19542
rect 31960 -20326 31976 -19558
rect 32010 -20326 32057 -19558
rect 31960 -20342 32057 -20326
rect 32457 -19558 32554 -19542
rect 32457 -20326 32504 -19558
rect 32538 -20326 32554 -19558
rect 32457 -20342 32554 -20326
rect 32596 -19558 32693 -19542
rect 32596 -20326 32612 -19558
rect 32646 -20326 32693 -19558
rect 32596 -20342 32693 -20326
rect 33093 -19558 33190 -19542
rect 33093 -20326 33140 -19558
rect 33174 -20326 33190 -19558
rect 33093 -20342 33190 -20326
rect 33560 -19032 33657 -19016
rect 33560 -19200 33576 -19032
rect 33610 -19200 33657 -19032
rect 33560 -19216 33657 -19200
rect 34057 -19032 34154 -19016
rect 34057 -19200 34104 -19032
rect 34138 -19200 34154 -19032
rect 34057 -19216 34154 -19200
rect 34196 -19032 34293 -19016
rect 34196 -19200 34212 -19032
rect 34246 -19200 34293 -19032
rect 34196 -19216 34293 -19200
rect 34693 -19032 34790 -19016
rect 34693 -19200 34740 -19032
rect 34774 -19200 34790 -19032
rect 34693 -19216 34790 -19200
rect 33560 -19558 33657 -19542
rect 33560 -20326 33576 -19558
rect 33610 -20326 33657 -19558
rect 33560 -20342 33657 -20326
rect 34057 -19558 34154 -19542
rect 34057 -20326 34104 -19558
rect 34138 -20326 34154 -19558
rect 34057 -20342 34154 -20326
rect 34196 -19558 34293 -19542
rect 34196 -20326 34212 -19558
rect 34246 -20326 34293 -19558
rect 34196 -20342 34293 -20326
rect 34693 -19558 34790 -19542
rect 34693 -20326 34740 -19558
rect 34774 -20326 34790 -19558
rect 34693 -20342 34790 -20326
rect 35160 -19032 35257 -19016
rect 35160 -19200 35176 -19032
rect 35210 -19200 35257 -19032
rect 35160 -19216 35257 -19200
rect 35657 -19032 35754 -19016
rect 35657 -19200 35704 -19032
rect 35738 -19200 35754 -19032
rect 35657 -19216 35754 -19200
rect 35796 -19032 35893 -19016
rect 35796 -19200 35812 -19032
rect 35846 -19200 35893 -19032
rect 35796 -19216 35893 -19200
rect 36293 -19032 36390 -19016
rect 36293 -19200 36340 -19032
rect 36374 -19200 36390 -19032
rect 36293 -19216 36390 -19200
rect 35160 -19558 35257 -19542
rect 35160 -20326 35176 -19558
rect 35210 -20326 35257 -19558
rect 35160 -20342 35257 -20326
rect 35657 -19558 35754 -19542
rect 35657 -20326 35704 -19558
rect 35738 -20326 35754 -19558
rect 35657 -20342 35754 -20326
rect 35796 -19558 35893 -19542
rect 35796 -20326 35812 -19558
rect 35846 -20326 35893 -19558
rect 35796 -20342 35893 -20326
rect 36293 -19558 36390 -19542
rect 36293 -20326 36340 -19558
rect 36374 -20326 36390 -19558
rect 36293 -20342 36390 -20326
rect 36760 -19032 36857 -19016
rect 36760 -19200 36776 -19032
rect 36810 -19200 36857 -19032
rect 36760 -19216 36857 -19200
rect 37257 -19032 37354 -19016
rect 37257 -19200 37304 -19032
rect 37338 -19200 37354 -19032
rect 37257 -19216 37354 -19200
rect 37396 -19032 37493 -19016
rect 37396 -19200 37412 -19032
rect 37446 -19200 37493 -19032
rect 37396 -19216 37493 -19200
rect 37893 -19032 37990 -19016
rect 37893 -19200 37940 -19032
rect 37974 -19200 37990 -19032
rect 37893 -19216 37990 -19200
rect 36760 -19558 36857 -19542
rect 36760 -20326 36776 -19558
rect 36810 -20326 36857 -19558
rect 36760 -20342 36857 -20326
rect 37257 -19558 37354 -19542
rect 37257 -20326 37304 -19558
rect 37338 -20326 37354 -19558
rect 37257 -20342 37354 -20326
rect 37396 -19558 37493 -19542
rect 37396 -20326 37412 -19558
rect 37446 -20326 37493 -19558
rect 37396 -20342 37493 -20326
rect 37893 -19558 37990 -19542
rect 37893 -20326 37940 -19558
rect 37974 -20326 37990 -19558
rect 37893 -20342 37990 -20326
rect -40 -20832 57 -20816
rect -40 -21000 -24 -20832
rect 10 -21000 57 -20832
rect -40 -21016 57 -21000
rect 457 -20832 554 -20816
rect 457 -21000 504 -20832
rect 538 -21000 554 -20832
rect 457 -21016 554 -21000
rect 596 -20832 693 -20816
rect 596 -21000 612 -20832
rect 646 -21000 693 -20832
rect 596 -21016 693 -21000
rect 1093 -20832 1190 -20816
rect 1093 -21000 1140 -20832
rect 1174 -21000 1190 -20832
rect 1093 -21016 1190 -21000
rect -40 -21358 57 -21342
rect -40 -22126 -24 -21358
rect 10 -22126 57 -21358
rect -40 -22142 57 -22126
rect 457 -21358 554 -21342
rect 457 -22126 504 -21358
rect 538 -22126 554 -21358
rect 457 -22142 554 -22126
rect 596 -21358 693 -21342
rect 596 -22126 612 -21358
rect 646 -22126 693 -21358
rect 596 -22142 693 -22126
rect 1093 -21358 1190 -21342
rect 1093 -22126 1140 -21358
rect 1174 -22126 1190 -21358
rect 1093 -22142 1190 -22126
rect 1560 -20832 1657 -20816
rect 1560 -21000 1576 -20832
rect 1610 -21000 1657 -20832
rect 1560 -21016 1657 -21000
rect 2057 -20832 2154 -20816
rect 2057 -21000 2104 -20832
rect 2138 -21000 2154 -20832
rect 2057 -21016 2154 -21000
rect 2196 -20832 2293 -20816
rect 2196 -21000 2212 -20832
rect 2246 -21000 2293 -20832
rect 2196 -21016 2293 -21000
rect 2693 -20832 2790 -20816
rect 2693 -21000 2740 -20832
rect 2774 -21000 2790 -20832
rect 2693 -21016 2790 -21000
rect 1560 -21358 1657 -21342
rect 1560 -22126 1576 -21358
rect 1610 -22126 1657 -21358
rect 1560 -22142 1657 -22126
rect 2057 -21358 2154 -21342
rect 2057 -22126 2104 -21358
rect 2138 -22126 2154 -21358
rect 2057 -22142 2154 -22126
rect 2196 -21358 2293 -21342
rect 2196 -22126 2212 -21358
rect 2246 -22126 2293 -21358
rect 2196 -22142 2293 -22126
rect 2693 -21358 2790 -21342
rect 2693 -22126 2740 -21358
rect 2774 -22126 2790 -21358
rect 2693 -22142 2790 -22126
rect 3160 -20832 3257 -20816
rect 3160 -21000 3176 -20832
rect 3210 -21000 3257 -20832
rect 3160 -21016 3257 -21000
rect 3657 -20832 3754 -20816
rect 3657 -21000 3704 -20832
rect 3738 -21000 3754 -20832
rect 3657 -21016 3754 -21000
rect 3796 -20832 3893 -20816
rect 3796 -21000 3812 -20832
rect 3846 -21000 3893 -20832
rect 3796 -21016 3893 -21000
rect 4293 -20832 4390 -20816
rect 4293 -21000 4340 -20832
rect 4374 -21000 4390 -20832
rect 4293 -21016 4390 -21000
rect 3160 -21358 3257 -21342
rect 3160 -22126 3176 -21358
rect 3210 -22126 3257 -21358
rect 3160 -22142 3257 -22126
rect 3657 -21358 3754 -21342
rect 3657 -22126 3704 -21358
rect 3738 -22126 3754 -21358
rect 3657 -22142 3754 -22126
rect 3796 -21358 3893 -21342
rect 3796 -22126 3812 -21358
rect 3846 -22126 3893 -21358
rect 3796 -22142 3893 -22126
rect 4293 -21358 4390 -21342
rect 4293 -22126 4340 -21358
rect 4374 -22126 4390 -21358
rect 4293 -22142 4390 -22126
rect 4760 -20832 4857 -20816
rect 4760 -21000 4776 -20832
rect 4810 -21000 4857 -20832
rect 4760 -21016 4857 -21000
rect 5257 -20832 5354 -20816
rect 5257 -21000 5304 -20832
rect 5338 -21000 5354 -20832
rect 5257 -21016 5354 -21000
rect 5396 -20832 5493 -20816
rect 5396 -21000 5412 -20832
rect 5446 -21000 5493 -20832
rect 5396 -21016 5493 -21000
rect 5893 -20832 5990 -20816
rect 5893 -21000 5940 -20832
rect 5974 -21000 5990 -20832
rect 5893 -21016 5990 -21000
rect 4760 -21358 4857 -21342
rect 4760 -22126 4776 -21358
rect 4810 -22126 4857 -21358
rect 4760 -22142 4857 -22126
rect 5257 -21358 5354 -21342
rect 5257 -22126 5304 -21358
rect 5338 -22126 5354 -21358
rect 5257 -22142 5354 -22126
rect 5396 -21358 5493 -21342
rect 5396 -22126 5412 -21358
rect 5446 -22126 5493 -21358
rect 5396 -22142 5493 -22126
rect 5893 -21358 5990 -21342
rect 5893 -22126 5940 -21358
rect 5974 -22126 5990 -21358
rect 5893 -22142 5990 -22126
rect 6360 -20832 6457 -20816
rect 6360 -21000 6376 -20832
rect 6410 -21000 6457 -20832
rect 6360 -21016 6457 -21000
rect 6857 -20832 6954 -20816
rect 6857 -21000 6904 -20832
rect 6938 -21000 6954 -20832
rect 6857 -21016 6954 -21000
rect 6996 -20832 7093 -20816
rect 6996 -21000 7012 -20832
rect 7046 -21000 7093 -20832
rect 6996 -21016 7093 -21000
rect 7493 -20832 7590 -20816
rect 7493 -21000 7540 -20832
rect 7574 -21000 7590 -20832
rect 7493 -21016 7590 -21000
rect 6360 -21358 6457 -21342
rect 6360 -22126 6376 -21358
rect 6410 -22126 6457 -21358
rect 6360 -22142 6457 -22126
rect 6857 -21358 6954 -21342
rect 6857 -22126 6904 -21358
rect 6938 -22126 6954 -21358
rect 6857 -22142 6954 -22126
rect 6996 -21358 7093 -21342
rect 6996 -22126 7012 -21358
rect 7046 -22126 7093 -21358
rect 6996 -22142 7093 -22126
rect 7493 -21358 7590 -21342
rect 7493 -22126 7540 -21358
rect 7574 -22126 7590 -21358
rect 7493 -22142 7590 -22126
rect 7960 -20832 8057 -20816
rect 7960 -21000 7976 -20832
rect 8010 -21000 8057 -20832
rect 7960 -21016 8057 -21000
rect 8457 -20832 8554 -20816
rect 8457 -21000 8504 -20832
rect 8538 -21000 8554 -20832
rect 8457 -21016 8554 -21000
rect 8596 -20832 8693 -20816
rect 8596 -21000 8612 -20832
rect 8646 -21000 8693 -20832
rect 8596 -21016 8693 -21000
rect 9093 -20832 9190 -20816
rect 9093 -21000 9140 -20832
rect 9174 -21000 9190 -20832
rect 9093 -21016 9190 -21000
rect 7960 -21358 8057 -21342
rect 7960 -22126 7976 -21358
rect 8010 -22126 8057 -21358
rect 7960 -22142 8057 -22126
rect 8457 -21358 8554 -21342
rect 8457 -22126 8504 -21358
rect 8538 -22126 8554 -21358
rect 8457 -22142 8554 -22126
rect 8596 -21358 8693 -21342
rect 8596 -22126 8612 -21358
rect 8646 -22126 8693 -21358
rect 8596 -22142 8693 -22126
rect 9093 -21358 9190 -21342
rect 9093 -22126 9140 -21358
rect 9174 -22126 9190 -21358
rect 9093 -22142 9190 -22126
rect 9560 -20832 9657 -20816
rect 9560 -21000 9576 -20832
rect 9610 -21000 9657 -20832
rect 9560 -21016 9657 -21000
rect 10057 -20832 10154 -20816
rect 10057 -21000 10104 -20832
rect 10138 -21000 10154 -20832
rect 10057 -21016 10154 -21000
rect 10196 -20832 10293 -20816
rect 10196 -21000 10212 -20832
rect 10246 -21000 10293 -20832
rect 10196 -21016 10293 -21000
rect 10693 -20832 10790 -20816
rect 10693 -21000 10740 -20832
rect 10774 -21000 10790 -20832
rect 10693 -21016 10790 -21000
rect 9560 -21358 9657 -21342
rect 9560 -22126 9576 -21358
rect 9610 -22126 9657 -21358
rect 9560 -22142 9657 -22126
rect 10057 -21358 10154 -21342
rect 10057 -22126 10104 -21358
rect 10138 -22126 10154 -21358
rect 10057 -22142 10154 -22126
rect 10196 -21358 10293 -21342
rect 10196 -22126 10212 -21358
rect 10246 -22126 10293 -21358
rect 10196 -22142 10293 -22126
rect 10693 -21358 10790 -21342
rect 10693 -22126 10740 -21358
rect 10774 -22126 10790 -21358
rect 10693 -22142 10790 -22126
rect 11160 -20832 11257 -20816
rect 11160 -21000 11176 -20832
rect 11210 -21000 11257 -20832
rect 11160 -21016 11257 -21000
rect 11657 -20832 11754 -20816
rect 11657 -21000 11704 -20832
rect 11738 -21000 11754 -20832
rect 11657 -21016 11754 -21000
rect 11796 -20832 11893 -20816
rect 11796 -21000 11812 -20832
rect 11846 -21000 11893 -20832
rect 11796 -21016 11893 -21000
rect 12293 -20832 12390 -20816
rect 12293 -21000 12340 -20832
rect 12374 -21000 12390 -20832
rect 12293 -21016 12390 -21000
rect 11160 -21358 11257 -21342
rect 11160 -22126 11176 -21358
rect 11210 -22126 11257 -21358
rect 11160 -22142 11257 -22126
rect 11657 -21358 11754 -21342
rect 11657 -22126 11704 -21358
rect 11738 -22126 11754 -21358
rect 11657 -22142 11754 -22126
rect 11796 -21358 11893 -21342
rect 11796 -22126 11812 -21358
rect 11846 -22126 11893 -21358
rect 11796 -22142 11893 -22126
rect 12293 -21358 12390 -21342
rect 12293 -22126 12340 -21358
rect 12374 -22126 12390 -21358
rect 12293 -22142 12390 -22126
rect 12760 -20832 12857 -20816
rect 12760 -21000 12776 -20832
rect 12810 -21000 12857 -20832
rect 12760 -21016 12857 -21000
rect 13257 -20832 13354 -20816
rect 13257 -21000 13304 -20832
rect 13338 -21000 13354 -20832
rect 13257 -21016 13354 -21000
rect 13396 -20832 13493 -20816
rect 13396 -21000 13412 -20832
rect 13446 -21000 13493 -20832
rect 13396 -21016 13493 -21000
rect 13893 -20832 13990 -20816
rect 13893 -21000 13940 -20832
rect 13974 -21000 13990 -20832
rect 13893 -21016 13990 -21000
rect 12760 -21358 12857 -21342
rect 12760 -22126 12776 -21358
rect 12810 -22126 12857 -21358
rect 12760 -22142 12857 -22126
rect 13257 -21358 13354 -21342
rect 13257 -22126 13304 -21358
rect 13338 -22126 13354 -21358
rect 13257 -22142 13354 -22126
rect 13396 -21358 13493 -21342
rect 13396 -22126 13412 -21358
rect 13446 -22126 13493 -21358
rect 13396 -22142 13493 -22126
rect 13893 -21358 13990 -21342
rect 13893 -22126 13940 -21358
rect 13974 -22126 13990 -21358
rect 13893 -22142 13990 -22126
rect 14360 -20832 14457 -20816
rect 14360 -21000 14376 -20832
rect 14410 -21000 14457 -20832
rect 14360 -21016 14457 -21000
rect 14857 -20832 14954 -20816
rect 14857 -21000 14904 -20832
rect 14938 -21000 14954 -20832
rect 14857 -21016 14954 -21000
rect 14996 -20832 15093 -20816
rect 14996 -21000 15012 -20832
rect 15046 -21000 15093 -20832
rect 14996 -21016 15093 -21000
rect 15493 -20832 15590 -20816
rect 15493 -21000 15540 -20832
rect 15574 -21000 15590 -20832
rect 15493 -21016 15590 -21000
rect 14360 -21358 14457 -21342
rect 14360 -22126 14376 -21358
rect 14410 -22126 14457 -21358
rect 14360 -22142 14457 -22126
rect 14857 -21358 14954 -21342
rect 14857 -22126 14904 -21358
rect 14938 -22126 14954 -21358
rect 14857 -22142 14954 -22126
rect 14996 -21358 15093 -21342
rect 14996 -22126 15012 -21358
rect 15046 -22126 15093 -21358
rect 14996 -22142 15093 -22126
rect 15493 -21358 15590 -21342
rect 15493 -22126 15540 -21358
rect 15574 -22126 15590 -21358
rect 15493 -22142 15590 -22126
rect 15960 -20832 16057 -20816
rect 15960 -21000 15976 -20832
rect 16010 -21000 16057 -20832
rect 15960 -21016 16057 -21000
rect 16457 -20832 16554 -20816
rect 16457 -21000 16504 -20832
rect 16538 -21000 16554 -20832
rect 16457 -21016 16554 -21000
rect 16596 -20832 16693 -20816
rect 16596 -21000 16612 -20832
rect 16646 -21000 16693 -20832
rect 16596 -21016 16693 -21000
rect 17093 -20832 17190 -20816
rect 17093 -21000 17140 -20832
rect 17174 -21000 17190 -20832
rect 17093 -21016 17190 -21000
rect 15960 -21358 16057 -21342
rect 15960 -22126 15976 -21358
rect 16010 -22126 16057 -21358
rect 15960 -22142 16057 -22126
rect 16457 -21358 16554 -21342
rect 16457 -22126 16504 -21358
rect 16538 -22126 16554 -21358
rect 16457 -22142 16554 -22126
rect 16596 -21358 16693 -21342
rect 16596 -22126 16612 -21358
rect 16646 -22126 16693 -21358
rect 16596 -22142 16693 -22126
rect 17093 -21358 17190 -21342
rect 17093 -22126 17140 -21358
rect 17174 -22126 17190 -21358
rect 17093 -22142 17190 -22126
rect 17560 -20832 17657 -20816
rect 17560 -21000 17576 -20832
rect 17610 -21000 17657 -20832
rect 17560 -21016 17657 -21000
rect 18057 -20832 18154 -20816
rect 18057 -21000 18104 -20832
rect 18138 -21000 18154 -20832
rect 18057 -21016 18154 -21000
rect 18196 -20832 18293 -20816
rect 18196 -21000 18212 -20832
rect 18246 -21000 18293 -20832
rect 18196 -21016 18293 -21000
rect 18693 -20832 18790 -20816
rect 18693 -21000 18740 -20832
rect 18774 -21000 18790 -20832
rect 18693 -21016 18790 -21000
rect 17560 -21358 17657 -21342
rect 17560 -22126 17576 -21358
rect 17610 -22126 17657 -21358
rect 17560 -22142 17657 -22126
rect 18057 -21358 18154 -21342
rect 18057 -22126 18104 -21358
rect 18138 -22126 18154 -21358
rect 18057 -22142 18154 -22126
rect 18196 -21358 18293 -21342
rect 18196 -22126 18212 -21358
rect 18246 -22126 18293 -21358
rect 18196 -22142 18293 -22126
rect 18693 -21358 18790 -21342
rect 18693 -22126 18740 -21358
rect 18774 -22126 18790 -21358
rect 18693 -22142 18790 -22126
rect 19160 -20832 19257 -20816
rect 19160 -21000 19176 -20832
rect 19210 -21000 19257 -20832
rect 19160 -21016 19257 -21000
rect 19657 -20832 19754 -20816
rect 19657 -21000 19704 -20832
rect 19738 -21000 19754 -20832
rect 19657 -21016 19754 -21000
rect 19796 -20832 19893 -20816
rect 19796 -21000 19812 -20832
rect 19846 -21000 19893 -20832
rect 19796 -21016 19893 -21000
rect 20293 -20832 20390 -20816
rect 20293 -21000 20340 -20832
rect 20374 -21000 20390 -20832
rect 20293 -21016 20390 -21000
rect 19160 -21358 19257 -21342
rect 19160 -22126 19176 -21358
rect 19210 -22126 19257 -21358
rect 19160 -22142 19257 -22126
rect 19657 -21358 19754 -21342
rect 19657 -22126 19704 -21358
rect 19738 -22126 19754 -21358
rect 19657 -22142 19754 -22126
rect 19796 -21358 19893 -21342
rect 19796 -22126 19812 -21358
rect 19846 -22126 19893 -21358
rect 19796 -22142 19893 -22126
rect 20293 -21358 20390 -21342
rect 20293 -22126 20340 -21358
rect 20374 -22126 20390 -21358
rect 20293 -22142 20390 -22126
rect 20760 -20832 20857 -20816
rect 20760 -21000 20776 -20832
rect 20810 -21000 20857 -20832
rect 20760 -21016 20857 -21000
rect 21257 -20832 21354 -20816
rect 21257 -21000 21304 -20832
rect 21338 -21000 21354 -20832
rect 21257 -21016 21354 -21000
rect 21396 -20832 21493 -20816
rect 21396 -21000 21412 -20832
rect 21446 -21000 21493 -20832
rect 21396 -21016 21493 -21000
rect 21893 -20832 21990 -20816
rect 21893 -21000 21940 -20832
rect 21974 -21000 21990 -20832
rect 21893 -21016 21990 -21000
rect 20760 -21358 20857 -21342
rect 20760 -22126 20776 -21358
rect 20810 -22126 20857 -21358
rect 20760 -22142 20857 -22126
rect 21257 -21358 21354 -21342
rect 21257 -22126 21304 -21358
rect 21338 -22126 21354 -21358
rect 21257 -22142 21354 -22126
rect 21396 -21358 21493 -21342
rect 21396 -22126 21412 -21358
rect 21446 -22126 21493 -21358
rect 21396 -22142 21493 -22126
rect 21893 -21358 21990 -21342
rect 21893 -22126 21940 -21358
rect 21974 -22126 21990 -21358
rect 21893 -22142 21990 -22126
rect 22360 -20832 22457 -20816
rect 22360 -21000 22376 -20832
rect 22410 -21000 22457 -20832
rect 22360 -21016 22457 -21000
rect 22857 -20832 22954 -20816
rect 22857 -21000 22904 -20832
rect 22938 -21000 22954 -20832
rect 22857 -21016 22954 -21000
rect 22996 -20832 23093 -20816
rect 22996 -21000 23012 -20832
rect 23046 -21000 23093 -20832
rect 22996 -21016 23093 -21000
rect 23493 -20832 23590 -20816
rect 23493 -21000 23540 -20832
rect 23574 -21000 23590 -20832
rect 23493 -21016 23590 -21000
rect 22360 -21358 22457 -21342
rect 22360 -22126 22376 -21358
rect 22410 -22126 22457 -21358
rect 22360 -22142 22457 -22126
rect 22857 -21358 22954 -21342
rect 22857 -22126 22904 -21358
rect 22938 -22126 22954 -21358
rect 22857 -22142 22954 -22126
rect 22996 -21358 23093 -21342
rect 22996 -22126 23012 -21358
rect 23046 -22126 23093 -21358
rect 22996 -22142 23093 -22126
rect 23493 -21358 23590 -21342
rect 23493 -22126 23540 -21358
rect 23574 -22126 23590 -21358
rect 23493 -22142 23590 -22126
rect 23960 -20832 24057 -20816
rect 23960 -21000 23976 -20832
rect 24010 -21000 24057 -20832
rect 23960 -21016 24057 -21000
rect 24457 -20832 24554 -20816
rect 24457 -21000 24504 -20832
rect 24538 -21000 24554 -20832
rect 24457 -21016 24554 -21000
rect 24596 -20832 24693 -20816
rect 24596 -21000 24612 -20832
rect 24646 -21000 24693 -20832
rect 24596 -21016 24693 -21000
rect 25093 -20832 25190 -20816
rect 25093 -21000 25140 -20832
rect 25174 -21000 25190 -20832
rect 25093 -21016 25190 -21000
rect 23960 -21358 24057 -21342
rect 23960 -22126 23976 -21358
rect 24010 -22126 24057 -21358
rect 23960 -22142 24057 -22126
rect 24457 -21358 24554 -21342
rect 24457 -22126 24504 -21358
rect 24538 -22126 24554 -21358
rect 24457 -22142 24554 -22126
rect 24596 -21358 24693 -21342
rect 24596 -22126 24612 -21358
rect 24646 -22126 24693 -21358
rect 24596 -22142 24693 -22126
rect 25093 -21358 25190 -21342
rect 25093 -22126 25140 -21358
rect 25174 -22126 25190 -21358
rect 25093 -22142 25190 -22126
rect 25560 -20832 25657 -20816
rect 25560 -21000 25576 -20832
rect 25610 -21000 25657 -20832
rect 25560 -21016 25657 -21000
rect 26057 -20832 26154 -20816
rect 26057 -21000 26104 -20832
rect 26138 -21000 26154 -20832
rect 26057 -21016 26154 -21000
rect 26196 -20832 26293 -20816
rect 26196 -21000 26212 -20832
rect 26246 -21000 26293 -20832
rect 26196 -21016 26293 -21000
rect 26693 -20832 26790 -20816
rect 26693 -21000 26740 -20832
rect 26774 -21000 26790 -20832
rect 26693 -21016 26790 -21000
rect 25560 -21358 25657 -21342
rect 25560 -22126 25576 -21358
rect 25610 -22126 25657 -21358
rect 25560 -22142 25657 -22126
rect 26057 -21358 26154 -21342
rect 26057 -22126 26104 -21358
rect 26138 -22126 26154 -21358
rect 26057 -22142 26154 -22126
rect 26196 -21358 26293 -21342
rect 26196 -22126 26212 -21358
rect 26246 -22126 26293 -21358
rect 26196 -22142 26293 -22126
rect 26693 -21358 26790 -21342
rect 26693 -22126 26740 -21358
rect 26774 -22126 26790 -21358
rect 26693 -22142 26790 -22126
rect 27160 -20832 27257 -20816
rect 27160 -21000 27176 -20832
rect 27210 -21000 27257 -20832
rect 27160 -21016 27257 -21000
rect 27657 -20832 27754 -20816
rect 27657 -21000 27704 -20832
rect 27738 -21000 27754 -20832
rect 27657 -21016 27754 -21000
rect 27796 -20832 27893 -20816
rect 27796 -21000 27812 -20832
rect 27846 -21000 27893 -20832
rect 27796 -21016 27893 -21000
rect 28293 -20832 28390 -20816
rect 28293 -21000 28340 -20832
rect 28374 -21000 28390 -20832
rect 28293 -21016 28390 -21000
rect 27160 -21358 27257 -21342
rect 27160 -22126 27176 -21358
rect 27210 -22126 27257 -21358
rect 27160 -22142 27257 -22126
rect 27657 -21358 27754 -21342
rect 27657 -22126 27704 -21358
rect 27738 -22126 27754 -21358
rect 27657 -22142 27754 -22126
rect 27796 -21358 27893 -21342
rect 27796 -22126 27812 -21358
rect 27846 -22126 27893 -21358
rect 27796 -22142 27893 -22126
rect 28293 -21358 28390 -21342
rect 28293 -22126 28340 -21358
rect 28374 -22126 28390 -21358
rect 28293 -22142 28390 -22126
rect 28760 -20832 28857 -20816
rect 28760 -21000 28776 -20832
rect 28810 -21000 28857 -20832
rect 28760 -21016 28857 -21000
rect 29257 -20832 29354 -20816
rect 29257 -21000 29304 -20832
rect 29338 -21000 29354 -20832
rect 29257 -21016 29354 -21000
rect 29396 -20832 29493 -20816
rect 29396 -21000 29412 -20832
rect 29446 -21000 29493 -20832
rect 29396 -21016 29493 -21000
rect 29893 -20832 29990 -20816
rect 29893 -21000 29940 -20832
rect 29974 -21000 29990 -20832
rect 29893 -21016 29990 -21000
rect 28760 -21358 28857 -21342
rect 28760 -22126 28776 -21358
rect 28810 -22126 28857 -21358
rect 28760 -22142 28857 -22126
rect 29257 -21358 29354 -21342
rect 29257 -22126 29304 -21358
rect 29338 -22126 29354 -21358
rect 29257 -22142 29354 -22126
rect 29396 -21358 29493 -21342
rect 29396 -22126 29412 -21358
rect 29446 -22126 29493 -21358
rect 29396 -22142 29493 -22126
rect 29893 -21358 29990 -21342
rect 29893 -22126 29940 -21358
rect 29974 -22126 29990 -21358
rect 29893 -22142 29990 -22126
rect 30360 -20832 30457 -20816
rect 30360 -21000 30376 -20832
rect 30410 -21000 30457 -20832
rect 30360 -21016 30457 -21000
rect 30857 -20832 30954 -20816
rect 30857 -21000 30904 -20832
rect 30938 -21000 30954 -20832
rect 30857 -21016 30954 -21000
rect 30996 -20832 31093 -20816
rect 30996 -21000 31012 -20832
rect 31046 -21000 31093 -20832
rect 30996 -21016 31093 -21000
rect 31493 -20832 31590 -20816
rect 31493 -21000 31540 -20832
rect 31574 -21000 31590 -20832
rect 31493 -21016 31590 -21000
rect 30360 -21358 30457 -21342
rect 30360 -22126 30376 -21358
rect 30410 -22126 30457 -21358
rect 30360 -22142 30457 -22126
rect 30857 -21358 30954 -21342
rect 30857 -22126 30904 -21358
rect 30938 -22126 30954 -21358
rect 30857 -22142 30954 -22126
rect 30996 -21358 31093 -21342
rect 30996 -22126 31012 -21358
rect 31046 -22126 31093 -21358
rect 30996 -22142 31093 -22126
rect 31493 -21358 31590 -21342
rect 31493 -22126 31540 -21358
rect 31574 -22126 31590 -21358
rect 31493 -22142 31590 -22126
rect 31960 -20832 32057 -20816
rect 31960 -21000 31976 -20832
rect 32010 -21000 32057 -20832
rect 31960 -21016 32057 -21000
rect 32457 -20832 32554 -20816
rect 32457 -21000 32504 -20832
rect 32538 -21000 32554 -20832
rect 32457 -21016 32554 -21000
rect 32596 -20832 32693 -20816
rect 32596 -21000 32612 -20832
rect 32646 -21000 32693 -20832
rect 32596 -21016 32693 -21000
rect 33093 -20832 33190 -20816
rect 33093 -21000 33140 -20832
rect 33174 -21000 33190 -20832
rect 33093 -21016 33190 -21000
rect 31960 -21358 32057 -21342
rect 31960 -22126 31976 -21358
rect 32010 -22126 32057 -21358
rect 31960 -22142 32057 -22126
rect 32457 -21358 32554 -21342
rect 32457 -22126 32504 -21358
rect 32538 -22126 32554 -21358
rect 32457 -22142 32554 -22126
rect 32596 -21358 32693 -21342
rect 32596 -22126 32612 -21358
rect 32646 -22126 32693 -21358
rect 32596 -22142 32693 -22126
rect 33093 -21358 33190 -21342
rect 33093 -22126 33140 -21358
rect 33174 -22126 33190 -21358
rect 33093 -22142 33190 -22126
rect 33560 -20832 33657 -20816
rect 33560 -21000 33576 -20832
rect 33610 -21000 33657 -20832
rect 33560 -21016 33657 -21000
rect 34057 -20832 34154 -20816
rect 34057 -21000 34104 -20832
rect 34138 -21000 34154 -20832
rect 34057 -21016 34154 -21000
rect 34196 -20832 34293 -20816
rect 34196 -21000 34212 -20832
rect 34246 -21000 34293 -20832
rect 34196 -21016 34293 -21000
rect 34693 -20832 34790 -20816
rect 34693 -21000 34740 -20832
rect 34774 -21000 34790 -20832
rect 34693 -21016 34790 -21000
rect 33560 -21358 33657 -21342
rect 33560 -22126 33576 -21358
rect 33610 -22126 33657 -21358
rect 33560 -22142 33657 -22126
rect 34057 -21358 34154 -21342
rect 34057 -22126 34104 -21358
rect 34138 -22126 34154 -21358
rect 34057 -22142 34154 -22126
rect 34196 -21358 34293 -21342
rect 34196 -22126 34212 -21358
rect 34246 -22126 34293 -21358
rect 34196 -22142 34293 -22126
rect 34693 -21358 34790 -21342
rect 34693 -22126 34740 -21358
rect 34774 -22126 34790 -21358
rect 34693 -22142 34790 -22126
rect 35160 -20832 35257 -20816
rect 35160 -21000 35176 -20832
rect 35210 -21000 35257 -20832
rect 35160 -21016 35257 -21000
rect 35657 -20832 35754 -20816
rect 35657 -21000 35704 -20832
rect 35738 -21000 35754 -20832
rect 35657 -21016 35754 -21000
rect 35796 -20832 35893 -20816
rect 35796 -21000 35812 -20832
rect 35846 -21000 35893 -20832
rect 35796 -21016 35893 -21000
rect 36293 -20832 36390 -20816
rect 36293 -21000 36340 -20832
rect 36374 -21000 36390 -20832
rect 36293 -21016 36390 -21000
rect 35160 -21358 35257 -21342
rect 35160 -22126 35176 -21358
rect 35210 -22126 35257 -21358
rect 35160 -22142 35257 -22126
rect 35657 -21358 35754 -21342
rect 35657 -22126 35704 -21358
rect 35738 -22126 35754 -21358
rect 35657 -22142 35754 -22126
rect 35796 -21358 35893 -21342
rect 35796 -22126 35812 -21358
rect 35846 -22126 35893 -21358
rect 35796 -22142 35893 -22126
rect 36293 -21358 36390 -21342
rect 36293 -22126 36340 -21358
rect 36374 -22126 36390 -21358
rect 36293 -22142 36390 -22126
rect 36760 -20832 36857 -20816
rect 36760 -21000 36776 -20832
rect 36810 -21000 36857 -20832
rect 36760 -21016 36857 -21000
rect 37257 -20832 37354 -20816
rect 37257 -21000 37304 -20832
rect 37338 -21000 37354 -20832
rect 37257 -21016 37354 -21000
rect 37396 -20832 37493 -20816
rect 37396 -21000 37412 -20832
rect 37446 -21000 37493 -20832
rect 37396 -21016 37493 -21000
rect 37893 -20832 37990 -20816
rect 37893 -21000 37940 -20832
rect 37974 -21000 37990 -20832
rect 37893 -21016 37990 -21000
rect 36760 -21358 36857 -21342
rect 36760 -22126 36776 -21358
rect 36810 -22126 36857 -21358
rect 36760 -22142 36857 -22126
rect 37257 -21358 37354 -21342
rect 37257 -22126 37304 -21358
rect 37338 -22126 37354 -21358
rect 37257 -22142 37354 -22126
rect 37396 -21358 37493 -21342
rect 37396 -22126 37412 -21358
rect 37446 -22126 37493 -21358
rect 37396 -22142 37493 -22126
rect 37893 -21358 37990 -21342
rect 37893 -22126 37940 -21358
rect 37974 -22126 37990 -21358
rect 37893 -22142 37990 -22126
rect 28398 -22672 28498 -22646
rect 28556 -22672 28656 -22646
rect 28714 -22672 28814 -22646
rect 28872 -22672 28972 -22646
rect 28398 -23519 28498 -23472
rect 28398 -23553 28414 -23519
rect 28482 -23553 28498 -23519
rect 28398 -23569 28498 -23553
rect 28556 -23519 28656 -23472
rect 28556 -23553 28572 -23519
rect 28640 -23553 28656 -23519
rect 28556 -23569 28656 -23553
rect 28714 -23519 28814 -23472
rect 28714 -23553 28730 -23519
rect 28798 -23553 28814 -23519
rect 28714 -23569 28814 -23553
rect 28872 -23519 28972 -23472
rect 28872 -23553 28888 -23519
rect 28956 -23553 28972 -23519
rect 28872 -23569 28972 -23553
rect 32678 -22542 32778 -22526
rect 32678 -22576 32694 -22542
rect 32762 -22576 32778 -22542
rect 32678 -22623 32778 -22576
rect 32836 -22542 32936 -22526
rect 32836 -22576 32852 -22542
rect 32920 -22576 32936 -22542
rect 32836 -22623 32936 -22576
rect 32994 -22542 33094 -22526
rect 32994 -22576 33010 -22542
rect 33078 -22576 33094 -22542
rect 32994 -22623 33094 -22576
rect 33152 -22542 33252 -22526
rect 33152 -22576 33168 -22542
rect 33236 -22576 33252 -22542
rect 33152 -22623 33252 -22576
rect 32678 -23070 32778 -23023
rect 32678 -23104 32694 -23070
rect 32762 -23104 32778 -23070
rect 32678 -23120 32778 -23104
rect 32836 -23070 32936 -23023
rect 32836 -23104 32852 -23070
rect 32920 -23104 32936 -23070
rect 32836 -23120 32936 -23104
rect 32994 -23070 33094 -23023
rect 32994 -23104 33010 -23070
rect 33078 -23104 33094 -23070
rect 32994 -23120 33094 -23104
rect 33152 -23070 33252 -23023
rect 33152 -23104 33168 -23070
rect 33236 -23104 33252 -23070
rect 33152 -23120 33252 -23104
rect 34048 -22562 34148 -22546
rect 34048 -22596 34064 -22562
rect 34132 -22596 34148 -22562
rect 34048 -22643 34148 -22596
rect 34206 -22562 34306 -22546
rect 34206 -22596 34222 -22562
rect 34290 -22596 34306 -22562
rect 34206 -22643 34306 -22596
rect 34048 -23090 34148 -23043
rect 34048 -23124 34064 -23090
rect 34132 -23124 34148 -23090
rect 34048 -23140 34148 -23124
rect 34206 -23090 34306 -23043
rect 34206 -23124 34222 -23090
rect 34290 -23124 34306 -23090
rect 34206 -23140 34306 -23124
rect 170 -24368 267 -24352
rect 170 -24636 186 -24368
rect 220 -24636 267 -24368
rect 170 -24652 267 -24636
rect 1867 -24368 1964 -24352
rect 1867 -24636 1914 -24368
rect 1948 -24636 1964 -24368
rect 1867 -24652 1964 -24636
rect 2370 -24368 2467 -24352
rect 2370 -24636 2386 -24368
rect 2420 -24636 2467 -24368
rect 2370 -24652 2467 -24636
rect 4067 -24368 4164 -24352
rect 4067 -24636 4114 -24368
rect 4148 -24636 4164 -24368
rect 4067 -24652 4164 -24636
rect 4570 -24368 4667 -24352
rect 4570 -24636 4586 -24368
rect 4620 -24636 4667 -24368
rect 4570 -24652 4667 -24636
rect 6267 -24368 6364 -24352
rect 6267 -24636 6314 -24368
rect 6348 -24636 6364 -24368
rect 6267 -24652 6364 -24636
rect 6770 -24368 6867 -24352
rect 6770 -24636 6786 -24368
rect 6820 -24636 6867 -24368
rect 6770 -24652 6867 -24636
rect 8467 -24368 8564 -24352
rect 8467 -24636 8514 -24368
rect 8548 -24636 8564 -24368
rect 8467 -24652 8564 -24636
rect 8970 -24368 9067 -24352
rect 8970 -24636 8986 -24368
rect 9020 -24636 9067 -24368
rect 8970 -24652 9067 -24636
rect 10667 -24368 10764 -24352
rect 10667 -24636 10714 -24368
rect 10748 -24636 10764 -24368
rect 10667 -24652 10764 -24636
rect 11170 -24368 11267 -24352
rect 11170 -24636 11186 -24368
rect 11220 -24636 11267 -24368
rect 11170 -24652 11267 -24636
rect 12867 -24368 12964 -24352
rect 12867 -24636 12914 -24368
rect 12948 -24636 12964 -24368
rect 12867 -24652 12964 -24636
rect 13370 -24368 13467 -24352
rect 13370 -24636 13386 -24368
rect 13420 -24636 13467 -24368
rect 13370 -24652 13467 -24636
rect 15067 -24368 15164 -24352
rect 15067 -24636 15114 -24368
rect 15148 -24636 15164 -24368
rect 15067 -24652 15164 -24636
rect 15570 -24368 15667 -24352
rect 15570 -24636 15586 -24368
rect 15620 -24636 15667 -24368
rect 15570 -24652 15667 -24636
rect 17267 -24368 17364 -24352
rect 17267 -24636 17314 -24368
rect 17348 -24636 17364 -24368
rect 17267 -24652 17364 -24636
rect 17770 -24368 17867 -24352
rect 17770 -24636 17786 -24368
rect 17820 -24636 17867 -24368
rect 17770 -24652 17867 -24636
rect 19467 -24368 19564 -24352
rect 19467 -24636 19514 -24368
rect 19548 -24636 19564 -24368
rect 19467 -24652 19564 -24636
rect 19970 -24368 20067 -24352
rect 19970 -24636 19986 -24368
rect 20020 -24636 20067 -24368
rect 19970 -24652 20067 -24636
rect 21667 -24368 21764 -24352
rect 21667 -24636 21714 -24368
rect 21748 -24636 21764 -24368
rect 21667 -24652 21764 -24636
rect 33216 -23684 33316 -23668
rect 33216 -23718 33232 -23684
rect 33300 -23718 33316 -23684
rect 33216 -23765 33316 -23718
rect 33374 -23684 33474 -23668
rect 33374 -23718 33390 -23684
rect 33458 -23718 33474 -23684
rect 33374 -23765 33474 -23718
rect 33532 -23684 33632 -23668
rect 33532 -23718 33548 -23684
rect 33616 -23718 33632 -23684
rect 33532 -23765 33632 -23718
rect 33690 -23684 33790 -23668
rect 33690 -23718 33706 -23684
rect 33774 -23718 33790 -23684
rect 33690 -23765 33790 -23718
rect 33848 -23684 33948 -23668
rect 33848 -23718 33864 -23684
rect 33932 -23718 33948 -23684
rect 33848 -23765 33948 -23718
rect 34006 -23684 34106 -23668
rect 34006 -23718 34022 -23684
rect 34090 -23718 34106 -23684
rect 34006 -23765 34106 -23718
rect 33216 -24212 33316 -24165
rect 33216 -24246 33232 -24212
rect 33300 -24246 33316 -24212
rect 33216 -24262 33316 -24246
rect 33374 -24212 33474 -24165
rect 33374 -24246 33390 -24212
rect 33458 -24246 33474 -24212
rect 33374 -24262 33474 -24246
rect 33532 -24212 33632 -24165
rect 33532 -24246 33548 -24212
rect 33616 -24246 33632 -24212
rect 33532 -24262 33632 -24246
rect 33690 -24212 33790 -24165
rect 33690 -24246 33706 -24212
rect 33774 -24246 33790 -24212
rect 33690 -24262 33790 -24246
rect 33848 -24212 33948 -24165
rect 33848 -24246 33864 -24212
rect 33932 -24246 33948 -24212
rect 33848 -24262 33948 -24246
rect 34006 -24212 34106 -24165
rect 34006 -24246 34022 -24212
rect 34090 -24246 34106 -24212
rect 34006 -24262 34106 -24246
rect 34588 -23682 34688 -23666
rect 34588 -23716 34604 -23682
rect 34672 -23716 34688 -23682
rect 34588 -23763 34688 -23716
rect 34746 -23682 34846 -23666
rect 34746 -23716 34762 -23682
rect 34830 -23716 34846 -23682
rect 34746 -23763 34846 -23716
rect 34904 -23682 35004 -23666
rect 34904 -23716 34920 -23682
rect 34988 -23716 35004 -23682
rect 34904 -23763 35004 -23716
rect 35062 -23682 35162 -23666
rect 35062 -23716 35078 -23682
rect 35146 -23716 35162 -23682
rect 35062 -23763 35162 -23716
rect 35220 -23682 35320 -23666
rect 35220 -23716 35236 -23682
rect 35304 -23716 35320 -23682
rect 35220 -23763 35320 -23716
rect 35378 -23682 35478 -23666
rect 35378 -23716 35394 -23682
rect 35462 -23716 35478 -23682
rect 35378 -23763 35478 -23716
rect 35536 -23682 35636 -23666
rect 35536 -23716 35552 -23682
rect 35620 -23716 35636 -23682
rect 35536 -23763 35636 -23716
rect 35694 -23682 35794 -23666
rect 35694 -23716 35710 -23682
rect 35778 -23716 35794 -23682
rect 35694 -23763 35794 -23716
rect 35852 -23682 35952 -23666
rect 35852 -23716 35868 -23682
rect 35936 -23716 35952 -23682
rect 35852 -23763 35952 -23716
rect 36010 -23682 36110 -23666
rect 36010 -23716 36026 -23682
rect 36094 -23716 36110 -23682
rect 36010 -23763 36110 -23716
rect 36168 -23682 36268 -23666
rect 36168 -23716 36184 -23682
rect 36252 -23716 36268 -23682
rect 36168 -23763 36268 -23716
rect 36326 -23682 36426 -23666
rect 36326 -23716 36342 -23682
rect 36410 -23716 36426 -23682
rect 36326 -23763 36426 -23716
rect 36484 -23682 36584 -23666
rect 36484 -23716 36500 -23682
rect 36568 -23716 36584 -23682
rect 36484 -23763 36584 -23716
rect 36642 -23682 36742 -23666
rect 36642 -23716 36658 -23682
rect 36726 -23716 36742 -23682
rect 36642 -23763 36742 -23716
rect 36800 -23682 36900 -23666
rect 36800 -23716 36816 -23682
rect 36884 -23716 36900 -23682
rect 36800 -23763 36900 -23716
rect 36958 -23682 37058 -23666
rect 36958 -23716 36974 -23682
rect 37042 -23716 37058 -23682
rect 36958 -23763 37058 -23716
rect 34588 -24210 34688 -24163
rect 34588 -24244 34604 -24210
rect 34672 -24244 34688 -24210
rect 34588 -24260 34688 -24244
rect 34746 -24210 34846 -24163
rect 34746 -24244 34762 -24210
rect 34830 -24244 34846 -24210
rect 34746 -24260 34846 -24244
rect 34904 -24210 35004 -24163
rect 34904 -24244 34920 -24210
rect 34988 -24244 35004 -24210
rect 34904 -24260 35004 -24244
rect 35062 -24210 35162 -24163
rect 35062 -24244 35078 -24210
rect 35146 -24244 35162 -24210
rect 35062 -24260 35162 -24244
rect 35220 -24210 35320 -24163
rect 35220 -24244 35236 -24210
rect 35304 -24244 35320 -24210
rect 35220 -24260 35320 -24244
rect 35378 -24210 35478 -24163
rect 35378 -24244 35394 -24210
rect 35462 -24244 35478 -24210
rect 35378 -24260 35478 -24244
rect 35536 -24210 35636 -24163
rect 35536 -24244 35552 -24210
rect 35620 -24244 35636 -24210
rect 35536 -24260 35636 -24244
rect 35694 -24210 35794 -24163
rect 35694 -24244 35710 -24210
rect 35778 -24244 35794 -24210
rect 35694 -24260 35794 -24244
rect 35852 -24210 35952 -24163
rect 35852 -24244 35868 -24210
rect 35936 -24244 35952 -24210
rect 35852 -24260 35952 -24244
rect 36010 -24210 36110 -24163
rect 36010 -24244 36026 -24210
rect 36094 -24244 36110 -24210
rect 36010 -24260 36110 -24244
rect 36168 -24210 36268 -24163
rect 36168 -24244 36184 -24210
rect 36252 -24244 36268 -24210
rect 36168 -24260 36268 -24244
rect 36326 -24210 36426 -24163
rect 36326 -24244 36342 -24210
rect 36410 -24244 36426 -24210
rect 36326 -24260 36426 -24244
rect 36484 -24210 36584 -24163
rect 36484 -24244 36500 -24210
rect 36568 -24244 36584 -24210
rect 36484 -24260 36584 -24244
rect 36642 -24210 36742 -24163
rect 36642 -24244 36658 -24210
rect 36726 -24244 36742 -24210
rect 36642 -24260 36742 -24244
rect 36800 -24210 36900 -24163
rect 36800 -24244 36816 -24210
rect 36884 -24244 36900 -24210
rect 36800 -24260 36900 -24244
rect 36958 -24210 37058 -24163
rect 36958 -24244 36974 -24210
rect 37042 -24244 37058 -24210
rect 36958 -24260 37058 -24244
rect 170 -25168 267 -25152
rect 170 -25436 186 -25168
rect 220 -25436 267 -25168
rect 170 -25452 267 -25436
rect 1867 -25168 1964 -25152
rect 1867 -25436 1914 -25168
rect 1948 -25436 1964 -25168
rect 1867 -25452 1964 -25436
rect 2370 -25168 2467 -25152
rect 2370 -25436 2386 -25168
rect 2420 -25436 2467 -25168
rect 2370 -25452 2467 -25436
rect 4067 -25168 4164 -25152
rect 4067 -25436 4114 -25168
rect 4148 -25436 4164 -25168
rect 4067 -25452 4164 -25436
rect 4570 -25168 4667 -25152
rect 4570 -25436 4586 -25168
rect 4620 -25436 4667 -25168
rect 4570 -25452 4667 -25436
rect 6267 -25168 6364 -25152
rect 6267 -25436 6314 -25168
rect 6348 -25436 6364 -25168
rect 6267 -25452 6364 -25436
rect 6770 -25168 6867 -25152
rect 6770 -25436 6786 -25168
rect 6820 -25436 6867 -25168
rect 6770 -25452 6867 -25436
rect 8467 -25168 8564 -25152
rect 8467 -25436 8514 -25168
rect 8548 -25436 8564 -25168
rect 8467 -25452 8564 -25436
rect 8970 -25168 9067 -25152
rect 8970 -25436 8986 -25168
rect 9020 -25436 9067 -25168
rect 8970 -25452 9067 -25436
rect 10667 -25168 10764 -25152
rect 10667 -25436 10714 -25168
rect 10748 -25436 10764 -25168
rect 10667 -25452 10764 -25436
rect 11170 -25168 11267 -25152
rect 11170 -25436 11186 -25168
rect 11220 -25436 11267 -25168
rect 11170 -25452 11267 -25436
rect 12867 -25168 12964 -25152
rect 12867 -25436 12914 -25168
rect 12948 -25436 12964 -25168
rect 12867 -25452 12964 -25436
rect 13370 -25168 13467 -25152
rect 13370 -25436 13386 -25168
rect 13420 -25436 13467 -25168
rect 13370 -25452 13467 -25436
rect 15067 -25168 15164 -25152
rect 15067 -25436 15114 -25168
rect 15148 -25436 15164 -25168
rect 15067 -25452 15164 -25436
rect 15570 -25168 15667 -25152
rect 15570 -25436 15586 -25168
rect 15620 -25436 15667 -25168
rect 15570 -25452 15667 -25436
rect 17267 -25168 17364 -25152
rect 17267 -25436 17314 -25168
rect 17348 -25436 17364 -25168
rect 17267 -25452 17364 -25436
rect 17770 -25168 17867 -25152
rect 17770 -25436 17786 -25168
rect 17820 -25436 17867 -25168
rect 17770 -25452 17867 -25436
rect 19467 -25168 19564 -25152
rect 19467 -25436 19514 -25168
rect 19548 -25436 19564 -25168
rect 19467 -25452 19564 -25436
rect 19970 -25168 20067 -25152
rect 19970 -25436 19986 -25168
rect 20020 -25436 20067 -25168
rect 19970 -25452 20067 -25436
rect 21667 -25168 21764 -25152
rect 21667 -25436 21714 -25168
rect 21748 -25436 21764 -25168
rect 21667 -25452 21764 -25436
rect 170 -25968 267 -25952
rect 170 -26236 186 -25968
rect 220 -26236 267 -25968
rect 170 -26252 267 -26236
rect 1867 -25968 1964 -25952
rect 1867 -26236 1914 -25968
rect 1948 -26236 1964 -25968
rect 1867 -26252 1964 -26236
rect 2370 -25968 2467 -25952
rect 2370 -26236 2386 -25968
rect 2420 -26236 2467 -25968
rect 2370 -26252 2467 -26236
rect 4067 -25968 4164 -25952
rect 4067 -26236 4114 -25968
rect 4148 -26236 4164 -25968
rect 4067 -26252 4164 -26236
rect 4570 -25968 4667 -25952
rect 4570 -26236 4586 -25968
rect 4620 -26236 4667 -25968
rect 4570 -26252 4667 -26236
rect 6267 -25968 6364 -25952
rect 6267 -26236 6314 -25968
rect 6348 -26236 6364 -25968
rect 6267 -26252 6364 -26236
rect 6770 -25968 6867 -25952
rect 6770 -26236 6786 -25968
rect 6820 -26236 6867 -25968
rect 6770 -26252 6867 -26236
rect 8467 -25968 8564 -25952
rect 8467 -26236 8514 -25968
rect 8548 -26236 8564 -25968
rect 8467 -26252 8564 -26236
rect 8970 -25968 9067 -25952
rect 8970 -26236 8986 -25968
rect 9020 -26236 9067 -25968
rect 8970 -26252 9067 -26236
rect 10667 -25968 10764 -25952
rect 10667 -26236 10714 -25968
rect 10748 -26236 10764 -25968
rect 10667 -26252 10764 -26236
rect 11170 -25968 11267 -25952
rect 11170 -26236 11186 -25968
rect 11220 -26236 11267 -25968
rect 11170 -26252 11267 -26236
rect 12867 -25968 12964 -25952
rect 12867 -26236 12914 -25968
rect 12948 -26236 12964 -25968
rect 12867 -26252 12964 -26236
rect 13370 -25968 13467 -25952
rect 13370 -26236 13386 -25968
rect 13420 -26236 13467 -25968
rect 13370 -26252 13467 -26236
rect 15067 -25968 15164 -25952
rect 15067 -26236 15114 -25968
rect 15148 -26236 15164 -25968
rect 15067 -26252 15164 -26236
rect 15570 -25968 15667 -25952
rect 15570 -26236 15586 -25968
rect 15620 -26236 15667 -25968
rect 15570 -26252 15667 -26236
rect 17267 -25968 17364 -25952
rect 17267 -26236 17314 -25968
rect 17348 -26236 17364 -25968
rect 17267 -26252 17364 -26236
rect 17770 -25968 17867 -25952
rect 17770 -26236 17786 -25968
rect 17820 -26236 17867 -25968
rect 17770 -26252 17867 -26236
rect 19467 -25968 19564 -25952
rect 19467 -26236 19514 -25968
rect 19548 -26236 19564 -25968
rect 19467 -26252 19564 -26236
rect 19970 -25968 20067 -25952
rect 19970 -26236 19986 -25968
rect 20020 -26236 20067 -25968
rect 19970 -26252 20067 -26236
rect 21667 -25968 21764 -25952
rect 21667 -26236 21714 -25968
rect 21748 -26236 21764 -25968
rect 21667 -26252 21764 -26236
rect 170 -26768 267 -26752
rect 170 -27036 186 -26768
rect 220 -27036 267 -26768
rect 170 -27052 267 -27036
rect 1867 -26768 1964 -26752
rect 1867 -27036 1914 -26768
rect 1948 -27036 1964 -26768
rect 1867 -27052 1964 -27036
rect 2370 -26768 2467 -26752
rect 2370 -27036 2386 -26768
rect 2420 -27036 2467 -26768
rect 2370 -27052 2467 -27036
rect 4067 -26768 4164 -26752
rect 4067 -27036 4114 -26768
rect 4148 -27036 4164 -26768
rect 4067 -27052 4164 -27036
rect 4570 -26768 4667 -26752
rect 4570 -27036 4586 -26768
rect 4620 -27036 4667 -26768
rect 4570 -27052 4667 -27036
rect 6267 -26768 6364 -26752
rect 6267 -27036 6314 -26768
rect 6348 -27036 6364 -26768
rect 6267 -27052 6364 -27036
rect 6770 -26768 6867 -26752
rect 6770 -27036 6786 -26768
rect 6820 -27036 6867 -26768
rect 6770 -27052 6867 -27036
rect 8467 -26768 8564 -26752
rect 8467 -27036 8514 -26768
rect 8548 -27036 8564 -26768
rect 8467 -27052 8564 -27036
rect 8970 -26768 9067 -26752
rect 8970 -27036 8986 -26768
rect 9020 -27036 9067 -26768
rect 8970 -27052 9067 -27036
rect 10667 -26768 10764 -26752
rect 10667 -27036 10714 -26768
rect 10748 -27036 10764 -26768
rect 10667 -27052 10764 -27036
rect 11170 -26768 11267 -26752
rect 11170 -27036 11186 -26768
rect 11220 -27036 11267 -26768
rect 11170 -27052 11267 -27036
rect 12867 -26768 12964 -26752
rect 12867 -27036 12914 -26768
rect 12948 -27036 12964 -26768
rect 12867 -27052 12964 -27036
rect 13370 -26768 13467 -26752
rect 13370 -27036 13386 -26768
rect 13420 -27036 13467 -26768
rect 13370 -27052 13467 -27036
rect 15067 -26768 15164 -26752
rect 15067 -27036 15114 -26768
rect 15148 -27036 15164 -26768
rect 15067 -27052 15164 -27036
rect 15570 -26768 15667 -26752
rect 15570 -27036 15586 -26768
rect 15620 -27036 15667 -26768
rect 15570 -27052 15667 -27036
rect 17267 -26768 17364 -26752
rect 17267 -27036 17314 -26768
rect 17348 -27036 17364 -26768
rect 17267 -27052 17364 -27036
rect 17770 -26768 17867 -26752
rect 17770 -27036 17786 -26768
rect 17820 -27036 17867 -26768
rect 17770 -27052 17867 -27036
rect 19467 -26768 19564 -26752
rect 19467 -27036 19514 -26768
rect 19548 -27036 19564 -26768
rect 19467 -27052 19564 -27036
rect 19970 -26768 20067 -26752
rect 19970 -27036 19986 -26768
rect 20020 -27036 20067 -26768
rect 19970 -27052 20067 -27036
rect 21667 -26768 21764 -26752
rect 21667 -27036 21714 -26768
rect 21748 -27036 21764 -26768
rect 21667 -27052 21764 -27036
rect 170 -27568 267 -27552
rect 170 -27836 186 -27568
rect 220 -27836 267 -27568
rect 170 -27852 267 -27836
rect 1867 -27568 1964 -27552
rect 1867 -27836 1914 -27568
rect 1948 -27836 1964 -27568
rect 1867 -27852 1964 -27836
rect 2370 -27568 2467 -27552
rect 2370 -27836 2386 -27568
rect 2420 -27836 2467 -27568
rect 2370 -27852 2467 -27836
rect 4067 -27568 4164 -27552
rect 4067 -27836 4114 -27568
rect 4148 -27836 4164 -27568
rect 4067 -27852 4164 -27836
rect 4570 -27568 4667 -27552
rect 4570 -27836 4586 -27568
rect 4620 -27836 4667 -27568
rect 4570 -27852 4667 -27836
rect 6267 -27568 6364 -27552
rect 6267 -27836 6314 -27568
rect 6348 -27836 6364 -27568
rect 6267 -27852 6364 -27836
rect 6770 -27568 6867 -27552
rect 6770 -27836 6786 -27568
rect 6820 -27836 6867 -27568
rect 6770 -27852 6867 -27836
rect 8467 -27568 8564 -27552
rect 8467 -27836 8514 -27568
rect 8548 -27836 8564 -27568
rect 8467 -27852 8564 -27836
rect 8970 -27568 9067 -27552
rect 8970 -27836 8986 -27568
rect 9020 -27836 9067 -27568
rect 8970 -27852 9067 -27836
rect 10667 -27568 10764 -27552
rect 10667 -27836 10714 -27568
rect 10748 -27836 10764 -27568
rect 10667 -27852 10764 -27836
rect 11170 -27568 11267 -27552
rect 11170 -27836 11186 -27568
rect 11220 -27836 11267 -27568
rect 11170 -27852 11267 -27836
rect 12867 -27568 12964 -27552
rect 12867 -27836 12914 -27568
rect 12948 -27836 12964 -27568
rect 12867 -27852 12964 -27836
rect 13370 -27568 13467 -27552
rect 13370 -27836 13386 -27568
rect 13420 -27836 13467 -27568
rect 13370 -27852 13467 -27836
rect 15067 -27568 15164 -27552
rect 15067 -27836 15114 -27568
rect 15148 -27836 15164 -27568
rect 15067 -27852 15164 -27836
rect 15570 -27568 15667 -27552
rect 15570 -27836 15586 -27568
rect 15620 -27836 15667 -27568
rect 15570 -27852 15667 -27836
rect 17267 -27568 17364 -27552
rect 17267 -27836 17314 -27568
rect 17348 -27836 17364 -27568
rect 17267 -27852 17364 -27836
rect 17770 -27568 17867 -27552
rect 17770 -27836 17786 -27568
rect 17820 -27836 17867 -27568
rect 17770 -27852 17867 -27836
rect 19467 -27568 19564 -27552
rect 19467 -27836 19514 -27568
rect 19548 -27836 19564 -27568
rect 19467 -27852 19564 -27836
rect 19970 -27568 20067 -27552
rect 19970 -27836 19986 -27568
rect 20020 -27836 20067 -27568
rect 19970 -27852 20067 -27836
rect 21667 -27568 21764 -27552
rect 21667 -27836 21714 -27568
rect 21748 -27836 21764 -27568
rect 21667 -27852 21764 -27836
rect 170 -28368 267 -28352
rect 170 -28636 186 -28368
rect 220 -28636 267 -28368
rect 170 -28652 267 -28636
rect 1867 -28368 1964 -28352
rect 1867 -28636 1914 -28368
rect 1948 -28636 1964 -28368
rect 1867 -28652 1964 -28636
rect 2370 -28368 2467 -28352
rect 2370 -28636 2386 -28368
rect 2420 -28636 2467 -28368
rect 2370 -28652 2467 -28636
rect 4067 -28368 4164 -28352
rect 4067 -28636 4114 -28368
rect 4148 -28636 4164 -28368
rect 4067 -28652 4164 -28636
rect 4570 -28368 4667 -28352
rect 4570 -28636 4586 -28368
rect 4620 -28636 4667 -28368
rect 4570 -28652 4667 -28636
rect 6267 -28368 6364 -28352
rect 6267 -28636 6314 -28368
rect 6348 -28636 6364 -28368
rect 6267 -28652 6364 -28636
rect 6770 -28368 6867 -28352
rect 6770 -28636 6786 -28368
rect 6820 -28636 6867 -28368
rect 6770 -28652 6867 -28636
rect 8467 -28368 8564 -28352
rect 8467 -28636 8514 -28368
rect 8548 -28636 8564 -28368
rect 8467 -28652 8564 -28636
rect 8970 -28368 9067 -28352
rect 8970 -28636 8986 -28368
rect 9020 -28636 9067 -28368
rect 8970 -28652 9067 -28636
rect 10667 -28368 10764 -28352
rect 10667 -28636 10714 -28368
rect 10748 -28636 10764 -28368
rect 10667 -28652 10764 -28636
rect 11170 -28368 11267 -28352
rect 11170 -28636 11186 -28368
rect 11220 -28636 11267 -28368
rect 11170 -28652 11267 -28636
rect 12867 -28368 12964 -28352
rect 12867 -28636 12914 -28368
rect 12948 -28636 12964 -28368
rect 12867 -28652 12964 -28636
rect 13370 -28368 13467 -28352
rect 13370 -28636 13386 -28368
rect 13420 -28636 13467 -28368
rect 13370 -28652 13467 -28636
rect 15067 -28368 15164 -28352
rect 15067 -28636 15114 -28368
rect 15148 -28636 15164 -28368
rect 15067 -28652 15164 -28636
rect 15570 -28368 15667 -28352
rect 15570 -28636 15586 -28368
rect 15620 -28636 15667 -28368
rect 15570 -28652 15667 -28636
rect 17267 -28368 17364 -28352
rect 17267 -28636 17314 -28368
rect 17348 -28636 17364 -28368
rect 17267 -28652 17364 -28636
rect 17770 -28368 17867 -28352
rect 17770 -28636 17786 -28368
rect 17820 -28636 17867 -28368
rect 17770 -28652 17867 -28636
rect 19467 -28368 19564 -28352
rect 19467 -28636 19514 -28368
rect 19548 -28636 19564 -28368
rect 19467 -28652 19564 -28636
rect 19970 -28368 20067 -28352
rect 19970 -28636 19986 -28368
rect 20020 -28636 20067 -28368
rect 19970 -28652 20067 -28636
rect 21667 -28368 21764 -28352
rect 21667 -28636 21714 -28368
rect 21748 -28636 21764 -28368
rect 21667 -28652 21764 -28636
rect 170 -29168 267 -29152
rect 170 -29436 186 -29168
rect 220 -29436 267 -29168
rect 170 -29452 267 -29436
rect 1867 -29168 1964 -29152
rect 1867 -29436 1914 -29168
rect 1948 -29436 1964 -29168
rect 1867 -29452 1964 -29436
rect 2370 -29168 2467 -29152
rect 2370 -29436 2386 -29168
rect 2420 -29436 2467 -29168
rect 2370 -29452 2467 -29436
rect 4067 -29168 4164 -29152
rect 4067 -29436 4114 -29168
rect 4148 -29436 4164 -29168
rect 4067 -29452 4164 -29436
rect 4570 -29168 4667 -29152
rect 4570 -29436 4586 -29168
rect 4620 -29436 4667 -29168
rect 4570 -29452 4667 -29436
rect 6267 -29168 6364 -29152
rect 6267 -29436 6314 -29168
rect 6348 -29436 6364 -29168
rect 6267 -29452 6364 -29436
rect 6770 -29168 6867 -29152
rect 6770 -29436 6786 -29168
rect 6820 -29436 6867 -29168
rect 6770 -29452 6867 -29436
rect 8467 -29168 8564 -29152
rect 8467 -29436 8514 -29168
rect 8548 -29436 8564 -29168
rect 8467 -29452 8564 -29436
rect 8970 -29168 9067 -29152
rect 8970 -29436 8986 -29168
rect 9020 -29436 9067 -29168
rect 8970 -29452 9067 -29436
rect 10667 -29168 10764 -29152
rect 10667 -29436 10714 -29168
rect 10748 -29436 10764 -29168
rect 10667 -29452 10764 -29436
rect 11170 -29168 11267 -29152
rect 11170 -29436 11186 -29168
rect 11220 -29436 11267 -29168
rect 11170 -29452 11267 -29436
rect 12867 -29168 12964 -29152
rect 12867 -29436 12914 -29168
rect 12948 -29436 12964 -29168
rect 12867 -29452 12964 -29436
rect 13370 -29168 13467 -29152
rect 13370 -29436 13386 -29168
rect 13420 -29436 13467 -29168
rect 13370 -29452 13467 -29436
rect 15067 -29168 15164 -29152
rect 15067 -29436 15114 -29168
rect 15148 -29436 15164 -29168
rect 15067 -29452 15164 -29436
rect 15570 -29168 15667 -29152
rect 15570 -29436 15586 -29168
rect 15620 -29436 15667 -29168
rect 15570 -29452 15667 -29436
rect 17267 -29168 17364 -29152
rect 17267 -29436 17314 -29168
rect 17348 -29436 17364 -29168
rect 17267 -29452 17364 -29436
rect 17770 -29168 17867 -29152
rect 17770 -29436 17786 -29168
rect 17820 -29436 17867 -29168
rect 17770 -29452 17867 -29436
rect 19467 -29168 19564 -29152
rect 19467 -29436 19514 -29168
rect 19548 -29436 19564 -29168
rect 19467 -29452 19564 -29436
rect 19970 -29168 20067 -29152
rect 19970 -29436 19986 -29168
rect 20020 -29436 20067 -29168
rect 19970 -29452 20067 -29436
rect 21667 -29168 21764 -29152
rect 21667 -29436 21714 -29168
rect 21748 -29436 21764 -29168
rect 21667 -29452 21764 -29436
rect 170 -29968 267 -29952
rect 170 -30236 186 -29968
rect 220 -30236 267 -29968
rect 170 -30252 267 -30236
rect 1867 -29968 1964 -29952
rect 1867 -30236 1914 -29968
rect 1948 -30236 1964 -29968
rect 1867 -30252 1964 -30236
rect 2370 -29968 2467 -29952
rect 2370 -30236 2386 -29968
rect 2420 -30236 2467 -29968
rect 2370 -30252 2467 -30236
rect 4067 -29968 4164 -29952
rect 4067 -30236 4114 -29968
rect 4148 -30236 4164 -29968
rect 4067 -30252 4164 -30236
rect 4570 -29968 4667 -29952
rect 4570 -30236 4586 -29968
rect 4620 -30236 4667 -29968
rect 4570 -30252 4667 -30236
rect 6267 -29968 6364 -29952
rect 6267 -30236 6314 -29968
rect 6348 -30236 6364 -29968
rect 6267 -30252 6364 -30236
rect 6770 -29968 6867 -29952
rect 6770 -30236 6786 -29968
rect 6820 -30236 6867 -29968
rect 6770 -30252 6867 -30236
rect 8467 -29968 8564 -29952
rect 8467 -30236 8514 -29968
rect 8548 -30236 8564 -29968
rect 8467 -30252 8564 -30236
rect 8970 -29968 9067 -29952
rect 8970 -30236 8986 -29968
rect 9020 -30236 9067 -29968
rect 8970 -30252 9067 -30236
rect 10667 -29968 10764 -29952
rect 10667 -30236 10714 -29968
rect 10748 -30236 10764 -29968
rect 10667 -30252 10764 -30236
rect 11170 -29968 11267 -29952
rect 11170 -30236 11186 -29968
rect 11220 -30236 11267 -29968
rect 11170 -30252 11267 -30236
rect 12867 -29968 12964 -29952
rect 12867 -30236 12914 -29968
rect 12948 -30236 12964 -29968
rect 12867 -30252 12964 -30236
rect 13370 -29968 13467 -29952
rect 13370 -30236 13386 -29968
rect 13420 -30236 13467 -29968
rect 13370 -30252 13467 -30236
rect 15067 -29968 15164 -29952
rect 15067 -30236 15114 -29968
rect 15148 -30236 15164 -29968
rect 15067 -30252 15164 -30236
rect 15570 -29968 15667 -29952
rect 15570 -30236 15586 -29968
rect 15620 -30236 15667 -29968
rect 15570 -30252 15667 -30236
rect 17267 -29968 17364 -29952
rect 17267 -30236 17314 -29968
rect 17348 -30236 17364 -29968
rect 17267 -30252 17364 -30236
rect 17770 -29968 17867 -29952
rect 17770 -30236 17786 -29968
rect 17820 -30236 17867 -29968
rect 17770 -30252 17867 -30236
rect 19467 -29968 19564 -29952
rect 19467 -30236 19514 -29968
rect 19548 -30236 19564 -29968
rect 19467 -30252 19564 -30236
rect 19970 -29968 20067 -29952
rect 19970 -30236 19986 -29968
rect 20020 -30236 20067 -29968
rect 19970 -30252 20067 -30236
rect 21667 -29968 21764 -29952
rect 21667 -30236 21714 -29968
rect 21748 -30236 21764 -29968
rect 21667 -30252 21764 -30236
rect 170 -30768 267 -30752
rect 170 -31036 186 -30768
rect 220 -31036 267 -30768
rect 170 -31052 267 -31036
rect 1867 -30768 1964 -30752
rect 1867 -31036 1914 -30768
rect 1948 -31036 1964 -30768
rect 1867 -31052 1964 -31036
rect 2370 -30768 2467 -30752
rect 2370 -31036 2386 -30768
rect 2420 -31036 2467 -30768
rect 2370 -31052 2467 -31036
rect 4067 -30768 4164 -30752
rect 4067 -31036 4114 -30768
rect 4148 -31036 4164 -30768
rect 4067 -31052 4164 -31036
rect 4570 -30768 4667 -30752
rect 4570 -31036 4586 -30768
rect 4620 -31036 4667 -30768
rect 4570 -31052 4667 -31036
rect 6267 -30768 6364 -30752
rect 6267 -31036 6314 -30768
rect 6348 -31036 6364 -30768
rect 6267 -31052 6364 -31036
rect 6770 -30768 6867 -30752
rect 6770 -31036 6786 -30768
rect 6820 -31036 6867 -30768
rect 6770 -31052 6867 -31036
rect 8467 -30768 8564 -30752
rect 8467 -31036 8514 -30768
rect 8548 -31036 8564 -30768
rect 8467 -31052 8564 -31036
rect 8970 -30768 9067 -30752
rect 8970 -31036 8986 -30768
rect 9020 -31036 9067 -30768
rect 8970 -31052 9067 -31036
rect 10667 -30768 10764 -30752
rect 10667 -31036 10714 -30768
rect 10748 -31036 10764 -30768
rect 10667 -31052 10764 -31036
rect 11170 -30768 11267 -30752
rect 11170 -31036 11186 -30768
rect 11220 -31036 11267 -30768
rect 11170 -31052 11267 -31036
rect 12867 -30768 12964 -30752
rect 12867 -31036 12914 -30768
rect 12948 -31036 12964 -30768
rect 12867 -31052 12964 -31036
rect 13370 -30768 13467 -30752
rect 13370 -31036 13386 -30768
rect 13420 -31036 13467 -30768
rect 13370 -31052 13467 -31036
rect 15067 -30768 15164 -30752
rect 15067 -31036 15114 -30768
rect 15148 -31036 15164 -30768
rect 15067 -31052 15164 -31036
rect 15570 -30768 15667 -30752
rect 15570 -31036 15586 -30768
rect 15620 -31036 15667 -30768
rect 15570 -31052 15667 -31036
rect 17267 -30768 17364 -30752
rect 17267 -31036 17314 -30768
rect 17348 -31036 17364 -30768
rect 17267 -31052 17364 -31036
rect 17770 -30768 17867 -30752
rect 17770 -31036 17786 -30768
rect 17820 -31036 17867 -30768
rect 17770 -31052 17867 -31036
rect 19467 -30768 19564 -30752
rect 19467 -31036 19514 -30768
rect 19548 -31036 19564 -30768
rect 19467 -31052 19564 -31036
rect 19970 -30768 20067 -30752
rect 19970 -31036 19986 -30768
rect 20020 -31036 20067 -30768
rect 19970 -31052 20067 -31036
rect 21667 -30768 21764 -30752
rect 21667 -31036 21714 -30768
rect 21748 -31036 21764 -30768
rect 21667 -31052 21764 -31036
rect 170 -31568 267 -31552
rect 170 -31836 186 -31568
rect 220 -31836 267 -31568
rect 170 -31852 267 -31836
rect 1867 -31568 1964 -31552
rect 1867 -31836 1914 -31568
rect 1948 -31836 1964 -31568
rect 1867 -31852 1964 -31836
rect 2370 -31568 2467 -31552
rect 2370 -31836 2386 -31568
rect 2420 -31836 2467 -31568
rect 2370 -31852 2467 -31836
rect 4067 -31568 4164 -31552
rect 4067 -31836 4114 -31568
rect 4148 -31836 4164 -31568
rect 4067 -31852 4164 -31836
rect 4570 -31568 4667 -31552
rect 4570 -31836 4586 -31568
rect 4620 -31836 4667 -31568
rect 4570 -31852 4667 -31836
rect 6267 -31568 6364 -31552
rect 6267 -31836 6314 -31568
rect 6348 -31836 6364 -31568
rect 6267 -31852 6364 -31836
rect 6770 -31568 6867 -31552
rect 6770 -31836 6786 -31568
rect 6820 -31836 6867 -31568
rect 6770 -31852 6867 -31836
rect 8467 -31568 8564 -31552
rect 8467 -31836 8514 -31568
rect 8548 -31836 8564 -31568
rect 8467 -31852 8564 -31836
rect 8970 -31568 9067 -31552
rect 8970 -31836 8986 -31568
rect 9020 -31836 9067 -31568
rect 8970 -31852 9067 -31836
rect 10667 -31568 10764 -31552
rect 10667 -31836 10714 -31568
rect 10748 -31836 10764 -31568
rect 10667 -31852 10764 -31836
rect 11170 -31568 11267 -31552
rect 11170 -31836 11186 -31568
rect 11220 -31836 11267 -31568
rect 11170 -31852 11267 -31836
rect 12867 -31568 12964 -31552
rect 12867 -31836 12914 -31568
rect 12948 -31836 12964 -31568
rect 12867 -31852 12964 -31836
rect 13370 -31568 13467 -31552
rect 13370 -31836 13386 -31568
rect 13420 -31836 13467 -31568
rect 13370 -31852 13467 -31836
rect 15067 -31568 15164 -31552
rect 15067 -31836 15114 -31568
rect 15148 -31836 15164 -31568
rect 15067 -31852 15164 -31836
rect 15570 -31568 15667 -31552
rect 15570 -31836 15586 -31568
rect 15620 -31836 15667 -31568
rect 15570 -31852 15667 -31836
rect 17267 -31568 17364 -31552
rect 17267 -31836 17314 -31568
rect 17348 -31836 17364 -31568
rect 17267 -31852 17364 -31836
rect 17770 -31568 17867 -31552
rect 17770 -31836 17786 -31568
rect 17820 -31836 17867 -31568
rect 17770 -31852 17867 -31836
rect 19467 -31568 19564 -31552
rect 19467 -31836 19514 -31568
rect 19548 -31836 19564 -31568
rect 19467 -31852 19564 -31836
rect 19970 -31568 20067 -31552
rect 19970 -31836 19986 -31568
rect 20020 -31836 20067 -31568
rect 19970 -31852 20067 -31836
rect 21667 -31568 21764 -31552
rect 21667 -31836 21714 -31568
rect 21748 -31836 21764 -31568
rect 21667 -31852 21764 -31836
rect 27968 -24640 28768 -24624
rect 27968 -24674 27984 -24640
rect 28752 -24674 28768 -24640
rect 27968 -24712 28768 -24674
rect 27968 -25150 28768 -25112
rect 27968 -25184 27984 -25150
rect 28752 -25184 28768 -25150
rect 27968 -25200 28768 -25184
rect 27910 -25688 27936 -25588
rect 28736 -25604 28824 -25588
rect 28736 -25672 28774 -25604
rect 28808 -25672 28824 -25604
rect 28736 -25688 28824 -25672
rect 27910 -25846 27936 -25746
rect 28736 -25762 28824 -25746
rect 28736 -25830 28774 -25762
rect 28808 -25830 28824 -25762
rect 28736 -25846 28824 -25830
rect 27910 -26004 27936 -25904
rect 28736 -25920 28824 -25904
rect 28736 -25988 28774 -25920
rect 28808 -25988 28824 -25920
rect 28736 -26004 28824 -25988
rect 27910 -26162 27936 -26062
rect 28736 -26078 28824 -26062
rect 28736 -26146 28774 -26078
rect 28808 -26146 28824 -26078
rect 28736 -26162 28824 -26146
rect 27910 -26728 27936 -26628
rect 28736 -26644 28824 -26628
rect 28736 -26712 28774 -26644
rect 28808 -26712 28824 -26644
rect 28736 -26728 28824 -26712
rect 27910 -26886 27936 -26786
rect 28736 -26802 28824 -26786
rect 28736 -26870 28774 -26802
rect 28808 -26870 28824 -26802
rect 28736 -26886 28824 -26870
rect 27910 -27044 27936 -26944
rect 28736 -26960 28824 -26944
rect 28736 -27028 28774 -26960
rect 28808 -27028 28824 -26960
rect 28736 -27044 28824 -27028
rect 27910 -27202 27936 -27102
rect 28736 -27118 28824 -27102
rect 28736 -27186 28774 -27118
rect 28808 -27186 28824 -27118
rect 28736 -27202 28824 -27186
rect 34880 -24892 34977 -24876
rect 34880 -25060 34896 -24892
rect 34930 -25060 34977 -24892
rect 34880 -25076 34977 -25060
rect 35777 -24892 35874 -24876
rect 35777 -25060 35824 -24892
rect 35858 -25060 35874 -24892
rect 35777 -25076 35874 -25060
rect 34880 -25150 34977 -25134
rect 34880 -25318 34896 -25150
rect 34930 -25318 34977 -25150
rect 34880 -25334 34977 -25318
rect 35777 -25150 35874 -25134
rect 35777 -25318 35824 -25150
rect 35858 -25318 35874 -25150
rect 35777 -25334 35874 -25318
rect 34880 -25408 34977 -25392
rect 34880 -25576 34896 -25408
rect 34930 -25576 34977 -25408
rect 34880 -25592 34977 -25576
rect 35777 -25408 35874 -25392
rect 35777 -25576 35824 -25408
rect 35858 -25576 35874 -25408
rect 35777 -25592 35874 -25576
rect 34880 -25666 34977 -25650
rect 34880 -25834 34896 -25666
rect 34930 -25834 34977 -25666
rect 34880 -25850 34977 -25834
rect 35777 -25666 35874 -25650
rect 35777 -25834 35824 -25666
rect 35858 -25834 35874 -25666
rect 35777 -25850 35874 -25834
rect 34880 -25924 34977 -25908
rect 34880 -26092 34896 -25924
rect 34930 -26092 34977 -25924
rect 34880 -26108 34977 -26092
rect 35777 -25924 35874 -25908
rect 35777 -26092 35824 -25924
rect 35858 -26092 35874 -25924
rect 35777 -26108 35874 -26092
rect 34880 -26182 34977 -26166
rect 34880 -26350 34896 -26182
rect 34930 -26350 34977 -26182
rect 34880 -26366 34977 -26350
rect 35777 -26182 35874 -26166
rect 35777 -26350 35824 -26182
rect 35858 -26350 35874 -26182
rect 35777 -26366 35874 -26350
rect 34880 -26440 34977 -26424
rect 34880 -26608 34896 -26440
rect 34930 -26608 34977 -26440
rect 34880 -26624 34977 -26608
rect 35777 -26440 35874 -26424
rect 35777 -26608 35824 -26440
rect 35858 -26608 35874 -26440
rect 35777 -26624 35874 -26608
rect 34880 -26698 34977 -26682
rect 34880 -26866 34896 -26698
rect 34930 -26866 34977 -26698
rect 34880 -26882 34977 -26866
rect 35777 -26698 35874 -26682
rect 35777 -26866 35824 -26698
rect 35858 -26866 35874 -26698
rect 35777 -26882 35874 -26866
rect 36220 -24892 36317 -24876
rect 36220 -25060 36236 -24892
rect 36270 -25060 36317 -24892
rect 36220 -25076 36317 -25060
rect 37117 -24892 37214 -24876
rect 37117 -25060 37164 -24892
rect 37198 -25060 37214 -24892
rect 37117 -25076 37214 -25060
rect 36220 -25150 36317 -25134
rect 36220 -25318 36236 -25150
rect 36270 -25318 36317 -25150
rect 36220 -25334 36317 -25318
rect 37117 -25150 37214 -25134
rect 37117 -25318 37164 -25150
rect 37198 -25318 37214 -25150
rect 37117 -25334 37214 -25318
rect 36220 -25408 36317 -25392
rect 36220 -25576 36236 -25408
rect 36270 -25576 36317 -25408
rect 36220 -25592 36317 -25576
rect 37117 -25408 37214 -25392
rect 37117 -25576 37164 -25408
rect 37198 -25576 37214 -25408
rect 37117 -25592 37214 -25576
rect 36220 -25666 36317 -25650
rect 36220 -25834 36236 -25666
rect 36270 -25834 36317 -25666
rect 36220 -25850 36317 -25834
rect 37117 -25666 37214 -25650
rect 37117 -25834 37164 -25666
rect 37198 -25834 37214 -25666
rect 37117 -25850 37214 -25834
rect 36220 -25924 36317 -25908
rect 36220 -26092 36236 -25924
rect 36270 -26092 36317 -25924
rect 36220 -26108 36317 -26092
rect 37117 -25924 37214 -25908
rect 37117 -26092 37164 -25924
rect 37198 -26092 37214 -25924
rect 37117 -26108 37214 -26092
rect 36220 -26182 36317 -26166
rect 36220 -26350 36236 -26182
rect 36270 -26350 36317 -26182
rect 36220 -26366 36317 -26350
rect 37117 -26182 37214 -26166
rect 37117 -26350 37164 -26182
rect 37198 -26350 37214 -26182
rect 37117 -26366 37214 -26350
rect 36220 -26440 36317 -26424
rect 36220 -26608 36236 -26440
rect 36270 -26608 36317 -26440
rect 36220 -26624 36317 -26608
rect 37117 -26440 37214 -26424
rect 37117 -26608 37164 -26440
rect 37198 -26608 37214 -26440
rect 37117 -26624 37214 -26608
rect 36220 -26698 36317 -26682
rect 36220 -26866 36236 -26698
rect 36270 -26866 36317 -26698
rect 36220 -26882 36317 -26866
rect 37117 -26698 37214 -26682
rect 37117 -26866 37164 -26698
rect 37198 -26866 37214 -26698
rect 37117 -26882 37214 -26866
rect 27910 -27768 27936 -27668
rect 28736 -27684 28824 -27668
rect 28736 -27752 28774 -27684
rect 28808 -27752 28824 -27684
rect 28736 -27768 28824 -27752
rect 27910 -27926 27936 -27826
rect 28736 -27842 28824 -27826
rect 28736 -27910 28774 -27842
rect 28808 -27910 28824 -27842
rect 28736 -27926 28824 -27910
rect 27910 -28084 27936 -27984
rect 28736 -28000 28824 -27984
rect 28736 -28068 28774 -28000
rect 28808 -28068 28824 -28000
rect 28736 -28084 28824 -28068
rect 27910 -28242 27936 -28142
rect 28736 -28158 28824 -28142
rect 28736 -28226 28774 -28158
rect 28808 -28226 28824 -28158
rect 28736 -28242 28824 -28226
rect 27910 -28808 27936 -28708
rect 28736 -28724 28824 -28708
rect 28736 -28792 28774 -28724
rect 28808 -28792 28824 -28724
rect 28736 -28808 28824 -28792
rect 27910 -28966 27936 -28866
rect 28736 -28882 28824 -28866
rect 28736 -28950 28774 -28882
rect 28808 -28950 28824 -28882
rect 28736 -28966 28824 -28950
rect 27910 -29124 27936 -29024
rect 28736 -29040 28824 -29024
rect 28736 -29108 28774 -29040
rect 28808 -29108 28824 -29040
rect 28736 -29124 28824 -29108
rect 27910 -29282 27936 -29182
rect 28736 -29198 28824 -29182
rect 28736 -29266 28774 -29198
rect 28808 -29266 28824 -29198
rect 28736 -29282 28824 -29266
rect 31858 -28440 31958 -28424
rect 31858 -28474 31874 -28440
rect 31942 -28474 31958 -28440
rect 31858 -28521 31958 -28474
rect 31858 -28968 31958 -28921
rect 31858 -29002 31874 -28968
rect 31942 -29002 31958 -28968
rect 31858 -29018 31958 -29002
rect 32298 -28440 32398 -28424
rect 32298 -28474 32314 -28440
rect 32382 -28474 32398 -28440
rect 32298 -28521 32398 -28474
rect 32298 -28968 32398 -28921
rect 32298 -29002 32314 -28968
rect 32382 -29002 32398 -28968
rect 32298 -29018 32398 -29002
rect 32738 -28440 32838 -28424
rect 32738 -28474 32754 -28440
rect 32822 -28474 32838 -28440
rect 32738 -28521 32838 -28474
rect 32738 -28968 32838 -28921
rect 32738 -29002 32754 -28968
rect 32822 -29002 32838 -28968
rect 32738 -29018 32838 -29002
rect 33152 -28740 33552 -28724
rect 33152 -28774 33168 -28740
rect 33536 -28774 33552 -28740
rect 33152 -28821 33552 -28774
rect 33152 -28968 33552 -28921
rect 33152 -29002 33168 -28968
rect 33536 -29002 33552 -28968
rect 33152 -29018 33552 -29002
rect 34058 -28440 34158 -28424
rect 34058 -28474 34074 -28440
rect 34142 -28474 34158 -28440
rect 34058 -28521 34158 -28474
rect 34058 -28968 34158 -28921
rect 34058 -29002 34074 -28968
rect 34142 -29002 34158 -28968
rect 34058 -29018 34158 -29002
rect 34498 -28440 34598 -28424
rect 34498 -28474 34514 -28440
rect 34582 -28474 34598 -28440
rect 34498 -28521 34598 -28474
rect 34498 -28968 34598 -28921
rect 34498 -29002 34514 -28968
rect 34582 -29002 34598 -28968
rect 34498 -29018 34598 -29002
rect 34938 -28440 35038 -28424
rect 34938 -28474 34954 -28440
rect 35022 -28474 35038 -28440
rect 34938 -28521 35038 -28474
rect 34938 -28968 35038 -28921
rect 34938 -29002 34954 -28968
rect 35022 -29002 35038 -28968
rect 34938 -29018 35038 -29002
rect 35352 -28740 35752 -28724
rect 35352 -28774 35368 -28740
rect 35736 -28774 35752 -28740
rect 35352 -28821 35752 -28774
rect 35352 -28968 35752 -28921
rect 35352 -29002 35368 -28968
rect 35736 -29002 35752 -28968
rect 35352 -29018 35752 -29002
rect 36258 -28440 36358 -28424
rect 36258 -28474 36274 -28440
rect 36342 -28474 36358 -28440
rect 36258 -28521 36358 -28474
rect 36258 -28968 36358 -28921
rect 36258 -29002 36274 -28968
rect 36342 -29002 36358 -28968
rect 36258 -29018 36358 -29002
rect 36698 -28440 36798 -28424
rect 36698 -28474 36714 -28440
rect 36782 -28474 36798 -28440
rect 36698 -28521 36798 -28474
rect 36698 -28968 36798 -28921
rect 36698 -29002 36714 -28968
rect 36782 -29002 36798 -28968
rect 36698 -29018 36798 -29002
rect 37138 -28440 37238 -28424
rect 37138 -28474 37154 -28440
rect 37222 -28474 37238 -28440
rect 37138 -28521 37238 -28474
rect 37138 -28968 37238 -28921
rect 37138 -29002 37154 -28968
rect 37222 -29002 37238 -28968
rect 37138 -29018 37238 -29002
rect 37552 -28740 37952 -28724
rect 37552 -28774 37568 -28740
rect 37936 -28774 37952 -28740
rect 37552 -28821 37952 -28774
rect 37552 -28968 37952 -28921
rect 37552 -29002 37568 -28968
rect 37936 -29002 37952 -28968
rect 37552 -29018 37952 -29002
rect 27910 -29848 27936 -29748
rect 28736 -29764 28824 -29748
rect 28736 -29832 28774 -29764
rect 28808 -29832 28824 -29764
rect 28736 -29848 28824 -29832
rect 27910 -30006 27936 -29906
rect 28736 -29922 28824 -29906
rect 28736 -29990 28774 -29922
rect 28808 -29990 28824 -29922
rect 28736 -30006 28824 -29990
rect 27910 -30164 27936 -30064
rect 28736 -30080 28824 -30064
rect 28736 -30148 28774 -30080
rect 28808 -30148 28824 -30080
rect 28736 -30164 28824 -30148
rect 27910 -30322 27936 -30222
rect 28736 -30238 28824 -30222
rect 28736 -30306 28774 -30238
rect 28808 -30306 28824 -30238
rect 28736 -30322 28824 -30306
rect 31859 -29469 31959 -29453
rect 31859 -29503 31875 -29469
rect 31943 -29503 31959 -29469
rect 31859 -29541 31959 -29503
rect 31859 -29779 31959 -29741
rect 31859 -29813 31875 -29779
rect 31943 -29813 31959 -29779
rect 31859 -29829 31959 -29813
rect 32299 -29469 32399 -29453
rect 32299 -29503 32315 -29469
rect 32383 -29503 32399 -29469
rect 32299 -29541 32399 -29503
rect 32299 -29779 32399 -29741
rect 32299 -29813 32315 -29779
rect 32383 -29813 32399 -29779
rect 32299 -29829 32399 -29813
rect 32739 -29469 32839 -29453
rect 32739 -29503 32755 -29469
rect 32823 -29503 32839 -29469
rect 32739 -29541 32839 -29503
rect 32739 -29779 32839 -29741
rect 32739 -29813 32755 -29779
rect 32823 -29813 32839 -29779
rect 32739 -29829 32839 -29813
rect 33178 -29469 33278 -29453
rect 33178 -29503 33194 -29469
rect 33262 -29503 33278 -29469
rect 33178 -29541 33278 -29503
rect 33336 -29469 33436 -29453
rect 33336 -29503 33352 -29469
rect 33420 -29503 33436 -29469
rect 33336 -29541 33436 -29503
rect 33494 -29469 33594 -29453
rect 33494 -29503 33510 -29469
rect 33578 -29503 33594 -29469
rect 33494 -29541 33594 -29503
rect 33178 -29779 33278 -29741
rect 33178 -29813 33194 -29779
rect 33262 -29813 33278 -29779
rect 33178 -29829 33278 -29813
rect 33336 -29779 33436 -29741
rect 33336 -29813 33352 -29779
rect 33420 -29813 33436 -29779
rect 33336 -29829 33436 -29813
rect 33494 -29779 33594 -29741
rect 33494 -29813 33510 -29779
rect 33578 -29813 33594 -29779
rect 33494 -29829 33594 -29813
rect 34059 -29469 34159 -29453
rect 34059 -29503 34075 -29469
rect 34143 -29503 34159 -29469
rect 34059 -29541 34159 -29503
rect 34059 -29779 34159 -29741
rect 34059 -29813 34075 -29779
rect 34143 -29813 34159 -29779
rect 34059 -29829 34159 -29813
rect 34499 -29469 34599 -29453
rect 34499 -29503 34515 -29469
rect 34583 -29503 34599 -29469
rect 34499 -29541 34599 -29503
rect 34499 -29779 34599 -29741
rect 34499 -29813 34515 -29779
rect 34583 -29813 34599 -29779
rect 34499 -29829 34599 -29813
rect 34939 -29469 35039 -29453
rect 34939 -29503 34955 -29469
rect 35023 -29503 35039 -29469
rect 34939 -29541 35039 -29503
rect 34939 -29779 35039 -29741
rect 34939 -29813 34955 -29779
rect 35023 -29813 35039 -29779
rect 34939 -29829 35039 -29813
rect 35378 -29469 35478 -29453
rect 35378 -29503 35394 -29469
rect 35462 -29503 35478 -29469
rect 35378 -29541 35478 -29503
rect 35536 -29469 35636 -29453
rect 35536 -29503 35552 -29469
rect 35620 -29503 35636 -29469
rect 35536 -29541 35636 -29503
rect 35694 -29469 35794 -29453
rect 35694 -29503 35710 -29469
rect 35778 -29503 35794 -29469
rect 35694 -29541 35794 -29503
rect 35378 -29779 35478 -29741
rect 35378 -29813 35394 -29779
rect 35462 -29813 35478 -29779
rect 35378 -29829 35478 -29813
rect 35536 -29779 35636 -29741
rect 35536 -29813 35552 -29779
rect 35620 -29813 35636 -29779
rect 35536 -29829 35636 -29813
rect 35694 -29779 35794 -29741
rect 35694 -29813 35710 -29779
rect 35778 -29813 35794 -29779
rect 35694 -29829 35794 -29813
rect 36259 -29469 36359 -29453
rect 36259 -29503 36275 -29469
rect 36343 -29503 36359 -29469
rect 36259 -29541 36359 -29503
rect 36259 -29779 36359 -29741
rect 36259 -29813 36275 -29779
rect 36343 -29813 36359 -29779
rect 36259 -29829 36359 -29813
rect 36699 -29469 36799 -29453
rect 36699 -29503 36715 -29469
rect 36783 -29503 36799 -29469
rect 36699 -29541 36799 -29503
rect 36699 -29779 36799 -29741
rect 36699 -29813 36715 -29779
rect 36783 -29813 36799 -29779
rect 36699 -29829 36799 -29813
rect 37139 -29469 37239 -29453
rect 37139 -29503 37155 -29469
rect 37223 -29503 37239 -29469
rect 37139 -29541 37239 -29503
rect 37139 -29779 37239 -29741
rect 37139 -29813 37155 -29779
rect 37223 -29813 37239 -29779
rect 37139 -29829 37239 -29813
rect 37578 -29469 37678 -29453
rect 37578 -29503 37594 -29469
rect 37662 -29503 37678 -29469
rect 37578 -29541 37678 -29503
rect 37736 -29469 37836 -29453
rect 37736 -29503 37752 -29469
rect 37820 -29503 37836 -29469
rect 37736 -29541 37836 -29503
rect 37894 -29469 37994 -29453
rect 37894 -29503 37910 -29469
rect 37978 -29503 37994 -29469
rect 37894 -29541 37994 -29503
rect 37578 -29779 37678 -29741
rect 37578 -29813 37594 -29779
rect 37662 -29813 37678 -29779
rect 37578 -29829 37678 -29813
rect 37736 -29779 37836 -29741
rect 37736 -29813 37752 -29779
rect 37820 -29813 37836 -29779
rect 37736 -29829 37836 -29813
rect 37894 -29779 37994 -29741
rect 37894 -29813 37910 -29779
rect 37978 -29813 37994 -29779
rect 37894 -29829 37994 -29813
rect 27910 -30888 27936 -30788
rect 28736 -30804 28824 -30788
rect 28736 -30872 28774 -30804
rect 28808 -30872 28824 -30804
rect 28736 -30888 28824 -30872
rect 27910 -31046 27936 -30946
rect 28736 -30962 28824 -30946
rect 28736 -31030 28774 -30962
rect 28808 -31030 28824 -30962
rect 28736 -31046 28824 -31030
rect 27910 -31204 27936 -31104
rect 28736 -31120 28824 -31104
rect 28736 -31188 28774 -31120
rect 28808 -31188 28824 -31120
rect 28736 -31204 28824 -31188
rect 27910 -31362 27936 -31262
rect 28736 -31278 28824 -31262
rect 28736 -31346 28774 -31278
rect 28808 -31346 28824 -31278
rect 28736 -31362 28824 -31346
rect 31828 -30211 31928 -30195
rect 31828 -30245 31844 -30211
rect 31912 -30245 31928 -30211
rect 31828 -30283 31928 -30245
rect 31986 -30211 32086 -30195
rect 31986 -30245 32002 -30211
rect 32070 -30245 32086 -30211
rect 31986 -30283 32086 -30245
rect 32144 -30211 32244 -30195
rect 32144 -30245 32160 -30211
rect 32228 -30245 32244 -30211
rect 32144 -30283 32244 -30245
rect 31828 -30521 31928 -30483
rect 31828 -30555 31844 -30521
rect 31912 -30555 31928 -30521
rect 31828 -30571 31928 -30555
rect 31986 -30521 32086 -30483
rect 31986 -30555 32002 -30521
rect 32070 -30555 32086 -30521
rect 31986 -30571 32086 -30555
rect 32144 -30521 32244 -30483
rect 32144 -30555 32160 -30521
rect 32228 -30555 32244 -30521
rect 32144 -30571 32244 -30555
rect 32583 -30211 32683 -30195
rect 32583 -30245 32599 -30211
rect 32667 -30245 32683 -30211
rect 32583 -30283 32683 -30245
rect 32583 -30521 32683 -30483
rect 32583 -30555 32599 -30521
rect 32667 -30555 32683 -30521
rect 32583 -30571 32683 -30555
rect 33023 -30211 33123 -30195
rect 33023 -30245 33039 -30211
rect 33107 -30245 33123 -30211
rect 33023 -30283 33123 -30245
rect 33023 -30521 33123 -30483
rect 33023 -30555 33039 -30521
rect 33107 -30555 33123 -30521
rect 33023 -30571 33123 -30555
rect 33463 -30211 33563 -30195
rect 33463 -30245 33479 -30211
rect 33547 -30245 33563 -30211
rect 33463 -30283 33563 -30245
rect 33463 -30521 33563 -30483
rect 33463 -30555 33479 -30521
rect 33547 -30555 33563 -30521
rect 33463 -30571 33563 -30555
rect 34028 -30211 34128 -30195
rect 34028 -30245 34044 -30211
rect 34112 -30245 34128 -30211
rect 34028 -30283 34128 -30245
rect 34186 -30211 34286 -30195
rect 34186 -30245 34202 -30211
rect 34270 -30245 34286 -30211
rect 34186 -30283 34286 -30245
rect 34344 -30211 34444 -30195
rect 34344 -30245 34360 -30211
rect 34428 -30245 34444 -30211
rect 34344 -30283 34444 -30245
rect 34028 -30521 34128 -30483
rect 34028 -30555 34044 -30521
rect 34112 -30555 34128 -30521
rect 34028 -30571 34128 -30555
rect 34186 -30521 34286 -30483
rect 34186 -30555 34202 -30521
rect 34270 -30555 34286 -30521
rect 34186 -30571 34286 -30555
rect 34344 -30521 34444 -30483
rect 34344 -30555 34360 -30521
rect 34428 -30555 34444 -30521
rect 34344 -30571 34444 -30555
rect 34783 -30211 34883 -30195
rect 34783 -30245 34799 -30211
rect 34867 -30245 34883 -30211
rect 34783 -30283 34883 -30245
rect 34783 -30521 34883 -30483
rect 34783 -30555 34799 -30521
rect 34867 -30555 34883 -30521
rect 34783 -30571 34883 -30555
rect 35223 -30211 35323 -30195
rect 35223 -30245 35239 -30211
rect 35307 -30245 35323 -30211
rect 35223 -30283 35323 -30245
rect 35223 -30521 35323 -30483
rect 35223 -30555 35239 -30521
rect 35307 -30555 35323 -30521
rect 35223 -30571 35323 -30555
rect 35663 -30211 35763 -30195
rect 35663 -30245 35679 -30211
rect 35747 -30245 35763 -30211
rect 35663 -30283 35763 -30245
rect 35663 -30521 35763 -30483
rect 35663 -30555 35679 -30521
rect 35747 -30555 35763 -30521
rect 35663 -30571 35763 -30555
rect 36228 -30211 36328 -30195
rect 36228 -30245 36244 -30211
rect 36312 -30245 36328 -30211
rect 36228 -30283 36328 -30245
rect 36386 -30211 36486 -30195
rect 36386 -30245 36402 -30211
rect 36470 -30245 36486 -30211
rect 36386 -30283 36486 -30245
rect 36544 -30211 36644 -30195
rect 36544 -30245 36560 -30211
rect 36628 -30245 36644 -30211
rect 36544 -30283 36644 -30245
rect 36228 -30521 36328 -30483
rect 36228 -30555 36244 -30521
rect 36312 -30555 36328 -30521
rect 36228 -30571 36328 -30555
rect 36386 -30521 36486 -30483
rect 36386 -30555 36402 -30521
rect 36470 -30555 36486 -30521
rect 36386 -30571 36486 -30555
rect 36544 -30521 36644 -30483
rect 36544 -30555 36560 -30521
rect 36628 -30555 36644 -30521
rect 36544 -30571 36644 -30555
rect 36983 -30211 37083 -30195
rect 36983 -30245 36999 -30211
rect 37067 -30245 37083 -30211
rect 36983 -30283 37083 -30245
rect 36983 -30521 37083 -30483
rect 36983 -30555 36999 -30521
rect 37067 -30555 37083 -30521
rect 36983 -30571 37083 -30555
rect 37423 -30211 37523 -30195
rect 37423 -30245 37439 -30211
rect 37507 -30245 37523 -30211
rect 37423 -30283 37523 -30245
rect 37423 -30521 37523 -30483
rect 37423 -30555 37439 -30521
rect 37507 -30555 37523 -30521
rect 37423 -30571 37523 -30555
rect 37863 -30211 37963 -30195
rect 37863 -30245 37879 -30211
rect 37947 -30245 37963 -30211
rect 37863 -30283 37963 -30245
rect 37863 -30521 37963 -30483
rect 37863 -30555 37879 -30521
rect 37947 -30555 37963 -30521
rect 37863 -30571 37963 -30555
rect 31870 -31022 32270 -31006
rect 31870 -31056 31886 -31022
rect 32254 -31056 32270 -31022
rect 31870 -31103 32270 -31056
rect 31870 -31250 32270 -31203
rect 31870 -31284 31886 -31250
rect 32254 -31284 32270 -31250
rect 31870 -31300 32270 -31284
rect 32584 -31022 32684 -31006
rect 32584 -31056 32600 -31022
rect 32668 -31056 32684 -31022
rect 32584 -31103 32684 -31056
rect 32584 -31550 32684 -31503
rect 32584 -31584 32600 -31550
rect 32668 -31584 32684 -31550
rect 32584 -31600 32684 -31584
rect 33024 -31022 33124 -31006
rect 33024 -31056 33040 -31022
rect 33108 -31056 33124 -31022
rect 33024 -31103 33124 -31056
rect 33024 -31550 33124 -31503
rect 33024 -31584 33040 -31550
rect 33108 -31584 33124 -31550
rect 33024 -31600 33124 -31584
rect 33464 -31022 33564 -31006
rect 33464 -31056 33480 -31022
rect 33548 -31056 33564 -31022
rect 33464 -31103 33564 -31056
rect 33464 -31550 33564 -31503
rect 33464 -31584 33480 -31550
rect 33548 -31584 33564 -31550
rect 33464 -31600 33564 -31584
rect 34070 -31022 34470 -31006
rect 34070 -31056 34086 -31022
rect 34454 -31056 34470 -31022
rect 34070 -31103 34470 -31056
rect 34070 -31250 34470 -31203
rect 34070 -31284 34086 -31250
rect 34454 -31284 34470 -31250
rect 34070 -31300 34470 -31284
rect 34784 -31022 34884 -31006
rect 34784 -31056 34800 -31022
rect 34868 -31056 34884 -31022
rect 34784 -31103 34884 -31056
rect 34784 -31550 34884 -31503
rect 34784 -31584 34800 -31550
rect 34868 -31584 34884 -31550
rect 34784 -31600 34884 -31584
rect 35224 -31022 35324 -31006
rect 35224 -31056 35240 -31022
rect 35308 -31056 35324 -31022
rect 35224 -31103 35324 -31056
rect 35224 -31550 35324 -31503
rect 35224 -31584 35240 -31550
rect 35308 -31584 35324 -31550
rect 35224 -31600 35324 -31584
rect 35664 -31022 35764 -31006
rect 35664 -31056 35680 -31022
rect 35748 -31056 35764 -31022
rect 35664 -31103 35764 -31056
rect 35664 -31550 35764 -31503
rect 35664 -31584 35680 -31550
rect 35748 -31584 35764 -31550
rect 35664 -31600 35764 -31584
rect 36270 -31022 36670 -31006
rect 36270 -31056 36286 -31022
rect 36654 -31056 36670 -31022
rect 36270 -31103 36670 -31056
rect 36270 -31250 36670 -31203
rect 36270 -31284 36286 -31250
rect 36654 -31284 36670 -31250
rect 36270 -31300 36670 -31284
rect 36984 -31022 37084 -31006
rect 36984 -31056 37000 -31022
rect 37068 -31056 37084 -31022
rect 36984 -31103 37084 -31056
rect 36984 -31550 37084 -31503
rect 36984 -31584 37000 -31550
rect 37068 -31584 37084 -31550
rect 36984 -31600 37084 -31584
rect 37424 -31022 37524 -31006
rect 37424 -31056 37440 -31022
rect 37508 -31056 37524 -31022
rect 37424 -31103 37524 -31056
rect 37424 -31550 37524 -31503
rect 37424 -31584 37440 -31550
rect 37508 -31584 37524 -31550
rect 37424 -31600 37524 -31584
rect 37864 -31022 37964 -31006
rect 37864 -31056 37880 -31022
rect 37948 -31056 37964 -31022
rect 37864 -31103 37964 -31056
rect 37864 -31550 37964 -31503
rect 37864 -31584 37880 -31550
rect 37948 -31584 37964 -31550
rect 37864 -31600 37964 -31584
<< polycont >>
rect 187 11445 221 11713
rect 1897 11445 1931 11713
rect 2387 11445 2421 11713
rect 4097 11445 4131 11713
rect 4587 11445 4621 11713
rect 6297 11445 6331 11713
rect 6787 11445 6821 11713
rect 8497 11445 8531 11713
rect 8987 11445 9021 11713
rect 10697 11445 10731 11713
rect 11187 11445 11221 11713
rect 12897 11445 12931 11713
rect 13387 11445 13421 11713
rect 15097 11445 15131 11713
rect 15587 11445 15621 11713
rect 17297 11445 17331 11713
rect 17787 11445 17821 11713
rect 19497 11445 19531 11713
rect 19987 11445 20021 11713
rect 21697 11445 21731 11713
rect 187 10645 221 10913
rect 1897 10645 1931 10913
rect 2386 10644 2420 10912
rect 4096 10644 4130 10912
rect 4586 10644 4620 10912
rect 6296 10644 6330 10912
rect 6786 10644 6820 10912
rect 8496 10644 8530 10912
rect 8986 10644 9020 10912
rect 10696 10644 10730 10912
rect 11186 10644 11220 10912
rect 12896 10644 12930 10912
rect 13386 10644 13420 10912
rect 15096 10644 15130 10912
rect 15586 10644 15620 10912
rect 17296 10644 17330 10912
rect 17786 10644 17820 10912
rect 19496 10644 19530 10912
rect 19987 10645 20021 10913
rect 21697 10645 21731 10913
rect 187 9845 221 10113
rect 1897 9845 1931 10113
rect 2386 9844 2420 10112
rect 4096 9844 4130 10112
rect 4586 9844 4620 10112
rect 6296 9844 6330 10112
rect 6786 9844 6820 10112
rect 8496 9844 8530 10112
rect 8986 9844 9020 10112
rect 10696 9844 10730 10112
rect 11186 9844 11220 10112
rect 12896 9844 12930 10112
rect 13386 9844 13420 10112
rect 15096 9844 15130 10112
rect 15586 9844 15620 10112
rect 17296 9844 17330 10112
rect 17786 9844 17820 10112
rect 19496 9844 19530 10112
rect 19987 9845 20021 10113
rect 21697 9845 21731 10113
rect 187 9045 221 9313
rect 1897 9045 1931 9313
rect 2386 9044 2420 9312
rect 4096 9044 4130 9312
rect 4586 9044 4620 9312
rect 6296 9044 6330 9312
rect 6786 9044 6820 9312
rect 8496 9044 8530 9312
rect 8986 9044 9020 9312
rect 10696 9044 10730 9312
rect 11186 9044 11220 9312
rect 12896 9044 12930 9312
rect 13386 9044 13420 9312
rect 15096 9044 15130 9312
rect 15586 9044 15620 9312
rect 17296 9044 17330 9312
rect 17786 9044 17820 9312
rect 19496 9044 19530 9312
rect 19987 9045 20021 9313
rect 21697 9045 21731 9313
rect 187 8245 221 8513
rect 1897 8245 1931 8513
rect 2386 8244 2420 8512
rect 4096 8244 4130 8512
rect 4586 8244 4620 8512
rect 6296 8244 6330 8512
rect 6786 8244 6820 8512
rect 8496 8244 8530 8512
rect 8986 8244 9020 8512
rect 10696 8244 10730 8512
rect 11186 8244 11220 8512
rect 12896 8244 12930 8512
rect 13386 8244 13420 8512
rect 15096 8244 15130 8512
rect 15586 8244 15620 8512
rect 17296 8244 17330 8512
rect 17786 8244 17820 8512
rect 19496 8244 19530 8512
rect 19987 8245 20021 8513
rect 21697 8245 21731 8513
rect 187 7445 221 7713
rect 1897 7445 1931 7713
rect 2386 7444 2420 7712
rect 4096 7444 4130 7712
rect 4586 7444 4620 7712
rect 6296 7444 6330 7712
rect 6786 7444 6820 7712
rect 8496 7444 8530 7712
rect 8986 7444 9020 7712
rect 10696 7444 10730 7712
rect 11186 7444 11220 7712
rect 12896 7444 12930 7712
rect 13386 7444 13420 7712
rect 15096 7444 15130 7712
rect 15586 7444 15620 7712
rect 17296 7444 17330 7712
rect 17786 7444 17820 7712
rect 19496 7444 19530 7712
rect 19987 7445 20021 7713
rect 21697 7445 21731 7713
rect 187 6645 221 6913
rect 1897 6645 1931 6913
rect 2386 6644 2420 6912
rect 4096 6644 4130 6912
rect 4586 6644 4620 6912
rect 6296 6644 6330 6912
rect 6786 6644 6820 6912
rect 8496 6644 8530 6912
rect 8986 6644 9020 6912
rect 10696 6644 10730 6912
rect 11186 6644 11220 6912
rect 12896 6644 12930 6912
rect 13386 6644 13420 6912
rect 15096 6644 15130 6912
rect 15586 6644 15620 6912
rect 17296 6644 17330 6912
rect 17786 6644 17820 6912
rect 19496 6644 19530 6912
rect 19987 6645 20021 6913
rect 21697 6645 21731 6913
rect 187 5845 221 6113
rect 1897 5845 1931 6113
rect 2386 5844 2420 6112
rect 4096 5844 4130 6112
rect 4586 5844 4620 6112
rect 6296 5844 6330 6112
rect 6786 5844 6820 6112
rect 8496 5844 8530 6112
rect 8986 5844 9020 6112
rect 10696 5844 10730 6112
rect 11186 5844 11220 6112
rect 12896 5844 12930 6112
rect 13386 5844 13420 6112
rect 15096 5844 15130 6112
rect 15586 5844 15620 6112
rect 17296 5844 17330 6112
rect 17786 5844 17820 6112
rect 19496 5844 19530 6112
rect 19987 5845 20021 6113
rect 21697 5845 21731 6113
rect 187 5045 221 5313
rect 1897 5045 1931 5313
rect 2386 5044 2420 5312
rect 4096 5044 4130 5312
rect 4586 5044 4620 5312
rect 6296 5044 6330 5312
rect 6786 5044 6820 5312
rect 8496 5044 8530 5312
rect 8986 5044 9020 5312
rect 10696 5044 10730 5312
rect 11186 5044 11220 5312
rect 12896 5044 12930 5312
rect 13386 5044 13420 5312
rect 15096 5044 15130 5312
rect 15586 5044 15620 5312
rect 17296 5044 17330 5312
rect 17786 5044 17820 5312
rect 19496 5044 19530 5312
rect 19987 5045 20021 5313
rect 21697 5045 21731 5313
rect 187 4245 221 4513
rect 1897 4245 1931 4513
rect 2387 4245 2421 4513
rect 4097 4245 4131 4513
rect 4587 4245 4621 4513
rect 6297 4245 6331 4513
rect 6787 4245 6821 4513
rect 8497 4245 8531 4513
rect 8988 4246 9022 4514
rect 10698 4246 10732 4514
rect 11188 4246 11222 4514
rect 12898 4246 12932 4514
rect 13387 4245 13421 4513
rect 15097 4245 15131 4513
rect 15587 4245 15621 4513
rect 17297 4245 17331 4513
rect 17787 4245 17821 4513
rect 19497 4245 19531 4513
rect 19987 4245 20021 4513
rect 21697 4245 21731 4513
rect 28773 11328 28807 11396
rect 28773 11170 28807 11238
rect 28773 11012 28807 11080
rect 28773 10854 28807 10922
rect 30164 11765 30232 11799
rect 30322 11765 30390 11799
rect 30480 11765 30548 11799
rect 30164 11455 30232 11489
rect 30322 11455 30390 11489
rect 30480 11455 30548 11489
rect 30919 11765 30987 11799
rect 30919 11455 30987 11489
rect 31359 11765 31427 11799
rect 31359 11455 31427 11489
rect 31799 11765 31867 11799
rect 31799 11455 31867 11489
rect 32364 11765 32432 11799
rect 32522 11765 32590 11799
rect 32680 11765 32748 11799
rect 32364 11455 32432 11489
rect 32522 11455 32590 11489
rect 32680 11455 32748 11489
rect 33119 11765 33187 11799
rect 33119 11455 33187 11489
rect 33559 11765 33627 11799
rect 33559 11455 33627 11489
rect 33999 11765 34067 11799
rect 33999 11455 34067 11489
rect 34564 11765 34632 11799
rect 34722 11765 34790 11799
rect 34880 11765 34948 11799
rect 34564 11455 34632 11489
rect 34722 11455 34790 11489
rect 34880 11455 34948 11489
rect 35319 11765 35387 11799
rect 35319 11455 35387 11489
rect 35759 11765 35827 11799
rect 35759 11455 35827 11489
rect 36199 11765 36267 11799
rect 36199 11455 36267 11489
rect 30206 10954 30574 10988
rect 30206 10726 30574 10760
rect 30920 10954 30988 10988
rect 28773 10288 28807 10356
rect 28773 10130 28807 10198
rect 28773 9972 28807 10040
rect 28773 9814 28807 9882
rect 30920 10426 30988 10460
rect 31360 10954 31428 10988
rect 31360 10426 31428 10460
rect 31800 10954 31868 10988
rect 31800 10426 31868 10460
rect 32406 10954 32774 10988
rect 32406 10726 32774 10760
rect 33120 10954 33188 10988
rect 33120 10426 33188 10460
rect 33560 10954 33628 10988
rect 33560 10426 33628 10460
rect 34000 10954 34068 10988
rect 34000 10426 34068 10460
rect 34606 10954 34974 10988
rect 34606 10726 34974 10760
rect 35320 10954 35388 10988
rect 35320 10426 35388 10460
rect 35760 10954 35828 10988
rect 35760 10426 35828 10460
rect 36200 10954 36268 10988
rect 36200 10426 36268 10460
rect 28773 9248 28807 9316
rect 28773 9090 28807 9158
rect 28773 8932 28807 9000
rect 28773 8774 28807 8842
rect 29794 9644 30562 9678
rect 30652 9644 31420 9678
rect 29794 9116 30562 9150
rect 30652 9116 31420 9150
rect 28773 8208 28807 8276
rect 28773 8050 28807 8118
rect 28773 7892 28807 7960
rect 28773 7734 28807 7802
rect 28773 7168 28807 7236
rect 28773 7010 28807 7078
rect 28773 6852 28807 6920
rect 28773 6694 28807 6762
rect 29794 8640 30562 8674
rect 30652 8640 31420 8674
rect 29794 8112 30562 8146
rect 30652 8112 31420 8146
rect 29794 8004 30562 8038
rect 30652 8004 31420 8038
rect 29794 7476 30562 7510
rect 30652 7476 31420 7510
rect 32972 8906 33140 8940
rect 33230 8906 33398 8940
rect 32972 7978 33140 8012
rect 33230 7978 33398 8012
rect 33812 8906 33980 8940
rect 34070 8906 34238 8940
rect 33812 7978 33980 8012
rect 34070 7978 34238 8012
rect 34634 8686 34668 8720
rect 34634 8158 34668 8192
rect 35054 8686 35088 8720
rect 35054 8158 35088 8192
rect 35474 8686 35508 8720
rect 35474 8158 35508 8192
rect 29676 6834 29710 7002
rect 30604 6834 30638 7002
rect 31016 6834 31050 7002
rect 31944 6834 31978 7002
rect 33534 7476 33602 7510
rect 33692 7476 33760 7510
rect 33850 7476 33918 7510
rect 34008 7476 34076 7510
rect 33534 6966 33602 7000
rect 33692 6966 33760 7000
rect 33850 6966 33918 7000
rect 34008 6966 34076 7000
rect 34634 7368 34668 7402
rect 34634 7058 34668 7092
rect 35054 7368 35088 7402
rect 35054 7058 35088 7092
rect 35474 7368 35508 7402
rect 35474 7058 35508 7092
rect 28773 6128 28807 6196
rect 28773 5970 28807 6038
rect 28773 5812 28807 5880
rect 28773 5654 28807 5722
rect 29686 6004 29720 6172
rect 30596 6004 30630 6172
rect 31026 6004 31060 6172
rect 31936 6004 31970 6172
rect 27974 5204 28742 5238
rect 27974 4276 28742 4310
rect 29984 5546 30352 5580
rect 29984 5336 30352 5370
rect 31294 5546 31662 5580
rect 31294 5336 31662 5370
rect 29686 4744 29720 4912
rect 30596 4744 30630 4912
rect 31026 4744 31060 4912
rect 31936 4744 31970 4912
rect 17164 3354 17232 3388
rect 17322 3354 17390 3388
rect 17480 3354 17548 3388
rect 17638 3354 17706 3388
rect 32784 3996 32852 4030
rect 32942 3996 33010 4030
rect 33100 3996 33168 4030
rect 33258 3996 33326 4030
rect 33416 3996 33484 4030
rect 33574 3996 33642 4030
rect 33732 3996 33800 4030
rect 33890 3996 33958 4030
rect 32784 3486 32852 3520
rect 32942 3486 33010 3520
rect 33100 3486 33168 3520
rect 33258 3486 33326 3520
rect 33416 3486 33484 3520
rect 33574 3486 33642 3520
rect 33732 3486 33800 3520
rect 33890 3486 33958 3520
rect 34974 3996 35042 4030
rect 35132 3996 35200 4030
rect 35290 3996 35358 4030
rect 34974 3486 35042 3520
rect 35132 3486 35200 3520
rect 35290 3486 35358 3520
rect 36376 5770 36410 5938
rect 36886 5770 36920 5938
rect 36376 5512 36410 5680
rect 36886 5512 36920 5680
rect 36376 5254 36410 5422
rect 36886 5254 36920 5422
rect 36376 4996 36410 5164
rect 36886 4996 36920 5164
rect 36376 4738 36410 4906
rect 36886 4738 36920 4906
rect 36376 4480 36410 4648
rect 36886 4480 36920 4648
rect 36376 4222 36410 4390
rect 36886 4222 36920 4390
rect 36376 3964 36410 4132
rect 36886 3964 36920 4132
rect 37162 5770 37196 5938
rect 37672 5770 37706 5938
rect 37162 5512 37196 5680
rect 37672 5512 37706 5680
rect 37162 5254 37196 5422
rect 37672 5254 37706 5422
rect 37162 4996 37196 5164
rect 37672 4996 37706 5164
rect 37162 4738 37196 4906
rect 37672 4738 37706 4906
rect 37162 4480 37196 4648
rect 37672 4480 37706 4648
rect 37162 4222 37196 4390
rect 37672 4222 37706 4390
rect 37162 3964 37196 4132
rect 37672 3964 37706 4132
rect 32454 3066 32522 3100
rect 32612 3066 32680 3100
rect 32454 2556 32522 2590
rect 32612 2556 32680 2590
rect 34054 3066 34122 3100
rect 34212 3066 34280 3100
rect 34054 2556 34122 2590
rect 34212 2556 34280 2590
rect 35654 3066 35722 3100
rect 35812 3066 35880 3100
rect 35654 2556 35722 2590
rect 35812 2556 35880 2590
rect -13 1265 21 2033
rect 497 1265 531 2033
rect 605 1265 639 2033
rect 1115 1265 1149 2033
rect -13 719 21 887
rect 497 719 531 887
rect 605 719 639 887
rect 1115 719 1149 887
rect 1587 1265 1621 2033
rect 2097 1265 2131 2033
rect 2205 1265 2239 2033
rect 2715 1265 2749 2033
rect 1587 719 1621 887
rect 2097 719 2131 887
rect 2205 719 2239 887
rect 2715 719 2749 887
rect 3187 1265 3221 2033
rect 3697 1265 3731 2033
rect 3805 1265 3839 2033
rect 4315 1265 4349 2033
rect 3187 719 3221 887
rect 3697 719 3731 887
rect 3805 719 3839 887
rect 4315 719 4349 887
rect 4787 1265 4821 2033
rect 5297 1265 5331 2033
rect 5405 1265 5439 2033
rect 5915 1265 5949 2033
rect 4787 719 4821 887
rect 5297 719 5331 887
rect 5405 719 5439 887
rect 5915 719 5949 887
rect 6387 1265 6421 2033
rect 6897 1265 6931 2033
rect 7005 1265 7039 2033
rect 7515 1265 7549 2033
rect 6387 719 6421 887
rect 6897 719 6931 887
rect 7005 719 7039 887
rect 7515 719 7549 887
rect 7987 1265 8021 2033
rect 8497 1265 8531 2033
rect 8605 1265 8639 2033
rect 9115 1265 9149 2033
rect 7987 719 8021 887
rect 8497 719 8531 887
rect 8605 719 8639 887
rect 9115 719 9149 887
rect 9587 1265 9621 2033
rect 10097 1265 10131 2033
rect 10205 1265 10239 2033
rect 10715 1265 10749 2033
rect 9587 719 9621 887
rect 10097 719 10131 887
rect 10205 719 10239 887
rect 10715 719 10749 887
rect 11187 1265 11221 2033
rect 11697 1265 11731 2033
rect 11805 1265 11839 2033
rect 12315 1265 12349 2033
rect 11187 719 11221 887
rect 11697 719 11731 887
rect 11805 719 11839 887
rect 12315 719 12349 887
rect 12787 1265 12821 2033
rect 13297 1265 13331 2033
rect 13405 1265 13439 2033
rect 13915 1265 13949 2033
rect 12787 719 12821 887
rect 13297 719 13331 887
rect 13405 719 13439 887
rect 13915 719 13949 887
rect 14387 1265 14421 2033
rect 14897 1265 14931 2033
rect 15005 1265 15039 2033
rect 15515 1265 15549 2033
rect 14387 719 14421 887
rect 14897 719 14931 887
rect 15005 719 15039 887
rect 15515 719 15549 887
rect 15987 1265 16021 2033
rect 16497 1265 16531 2033
rect 16605 1265 16639 2033
rect 17115 1265 17149 2033
rect 15987 719 16021 887
rect 16497 719 16531 887
rect 16605 719 16639 887
rect 17115 719 17149 887
rect 17587 1265 17621 2033
rect 18097 1265 18131 2033
rect 18205 1265 18239 2033
rect 18715 1265 18749 2033
rect 17587 719 17621 887
rect 18097 719 18131 887
rect 18205 719 18239 887
rect 18715 719 18749 887
rect 19187 1265 19221 2033
rect 19697 1265 19731 2033
rect 19805 1265 19839 2033
rect 20315 1265 20349 2033
rect 19187 719 19221 887
rect 19697 719 19731 887
rect 19805 719 19839 887
rect 20315 719 20349 887
rect 20787 1265 20821 2033
rect 21297 1265 21331 2033
rect 21405 1265 21439 2033
rect 21915 1265 21949 2033
rect 20787 719 20821 887
rect 21297 719 21331 887
rect 21405 719 21439 887
rect 21915 719 21949 887
rect 22387 1265 22421 2033
rect 22897 1265 22931 2033
rect 23005 1265 23039 2033
rect 23515 1265 23549 2033
rect 22387 719 22421 887
rect 22897 719 22931 887
rect 23005 719 23039 887
rect 23515 719 23549 887
rect 23987 1265 24021 2033
rect 24497 1265 24531 2033
rect 24605 1265 24639 2033
rect 25115 1265 25149 2033
rect 23987 719 24021 887
rect 24497 719 24531 887
rect 24605 719 24639 887
rect 25115 719 25149 887
rect 25587 1265 25621 2033
rect 26097 1265 26131 2033
rect 26205 1265 26239 2033
rect 26715 1265 26749 2033
rect 25587 719 25621 887
rect 26097 719 26131 887
rect 26205 719 26239 887
rect 26715 719 26749 887
rect 27187 1265 27221 2033
rect 27697 1265 27731 2033
rect 27805 1265 27839 2033
rect 28315 1265 28349 2033
rect 27187 719 27221 887
rect 27697 719 27731 887
rect 27805 719 27839 887
rect 28315 719 28349 887
rect 28787 1265 28821 2033
rect 29297 1265 29331 2033
rect 29405 1265 29439 2033
rect 29915 1265 29949 2033
rect 28787 719 28821 887
rect 29297 719 29331 887
rect 29405 719 29439 887
rect 29915 719 29949 887
rect 30387 1265 30421 2033
rect 30897 1265 30931 2033
rect 31005 1265 31039 2033
rect 31515 1265 31549 2033
rect 30387 719 30421 887
rect 30897 719 30931 887
rect 31005 719 31039 887
rect 31515 719 31549 887
rect 31987 1265 32021 2033
rect 32497 1265 32531 2033
rect 32605 1265 32639 2033
rect 33115 1265 33149 2033
rect 31987 719 32021 887
rect 32497 719 32531 887
rect 32605 719 32639 887
rect 33115 719 33149 887
rect 33587 1265 33621 2033
rect 34097 1265 34131 2033
rect 34205 1265 34239 2033
rect 34715 1265 34749 2033
rect 33587 719 33621 887
rect 34097 719 34131 887
rect 34205 719 34239 887
rect 34715 719 34749 887
rect 35187 1265 35221 2033
rect 35697 1265 35731 2033
rect 35805 1265 35839 2033
rect 36315 1265 36349 2033
rect 35187 719 35221 887
rect 35697 719 35731 887
rect 35805 719 35839 887
rect 36315 719 36349 887
rect 36787 1265 36821 2033
rect 37297 1265 37331 2033
rect 37405 1265 37439 2033
rect 37915 1265 37949 2033
rect 36787 719 36821 887
rect 37297 719 37331 887
rect 37405 719 37439 887
rect 37915 719 37949 887
rect -13 -535 21 233
rect 497 -535 531 233
rect 605 -535 639 233
rect 1115 -535 1149 233
rect -13 -1081 21 -913
rect 497 -1081 531 -913
rect 605 -1081 639 -913
rect 1115 -1081 1149 -913
rect 1587 -535 1621 233
rect 2097 -535 2131 233
rect 2205 -535 2239 233
rect 2715 -535 2749 233
rect 1587 -1081 1621 -913
rect 2097 -1081 2131 -913
rect 2205 -1081 2239 -913
rect 2715 -1081 2749 -913
rect 3187 -535 3221 233
rect 3697 -535 3731 233
rect 3805 -535 3839 233
rect 4315 -535 4349 233
rect 3187 -1081 3221 -913
rect 3697 -1081 3731 -913
rect 3805 -1081 3839 -913
rect 4315 -1081 4349 -913
rect 4787 -535 4821 233
rect 5297 -535 5331 233
rect 5405 -535 5439 233
rect 5915 -535 5949 233
rect 4787 -1081 4821 -913
rect 5297 -1081 5331 -913
rect 5405 -1081 5439 -913
rect 5915 -1081 5949 -913
rect 6387 -535 6421 233
rect 6897 -535 6931 233
rect 7005 -535 7039 233
rect 7515 -535 7549 233
rect 6387 -1081 6421 -913
rect 6897 -1081 6931 -913
rect 7005 -1081 7039 -913
rect 7515 -1081 7549 -913
rect 7987 -535 8021 233
rect 8497 -535 8531 233
rect 8605 -535 8639 233
rect 9115 -535 9149 233
rect 7987 -1081 8021 -913
rect 8497 -1081 8531 -913
rect 8605 -1081 8639 -913
rect 9115 -1081 9149 -913
rect 9587 -535 9621 233
rect 10097 -535 10131 233
rect 10205 -535 10239 233
rect 10715 -535 10749 233
rect 9587 -1081 9621 -913
rect 10097 -1081 10131 -913
rect 10205 -1081 10239 -913
rect 10715 -1081 10749 -913
rect 11187 -535 11221 233
rect 11697 -535 11731 233
rect 11805 -535 11839 233
rect 12315 -535 12349 233
rect 11187 -1081 11221 -913
rect 11697 -1081 11731 -913
rect 11805 -1081 11839 -913
rect 12315 -1081 12349 -913
rect 12787 -535 12821 233
rect 13297 -535 13331 233
rect 13405 -535 13439 233
rect 13915 -535 13949 233
rect 12787 -1081 12821 -913
rect 13297 -1081 13331 -913
rect 13405 -1081 13439 -913
rect 13915 -1081 13949 -913
rect 14387 -535 14421 233
rect 14897 -535 14931 233
rect 15005 -535 15039 233
rect 15515 -535 15549 233
rect 14387 -1081 14421 -913
rect 14897 -1081 14931 -913
rect 15005 -1081 15039 -913
rect 15515 -1081 15549 -913
rect 15987 -535 16021 233
rect 16497 -535 16531 233
rect 16605 -535 16639 233
rect 17115 -535 17149 233
rect 15987 -1081 16021 -913
rect 16497 -1081 16531 -913
rect 16605 -1081 16639 -913
rect 17115 -1081 17149 -913
rect 17587 -535 17621 233
rect 18097 -535 18131 233
rect 18205 -535 18239 233
rect 18715 -535 18749 233
rect 17587 -1081 17621 -913
rect 18097 -1081 18131 -913
rect 18205 -1081 18239 -913
rect 18715 -1081 18749 -913
rect 19187 -535 19221 233
rect 19697 -535 19731 233
rect 19805 -535 19839 233
rect 20315 -535 20349 233
rect 19187 -1081 19221 -913
rect 19697 -1081 19731 -913
rect 19805 -1081 19839 -913
rect 20315 -1081 20349 -913
rect 20787 -535 20821 233
rect 21297 -535 21331 233
rect 21405 -535 21439 233
rect 21915 -535 21949 233
rect 20787 -1081 20821 -913
rect 21297 -1081 21331 -913
rect 21405 -1081 21439 -913
rect 21915 -1081 21949 -913
rect 22387 -535 22421 233
rect 22897 -535 22931 233
rect 23005 -535 23039 233
rect 23515 -535 23549 233
rect 22387 -1081 22421 -913
rect 22897 -1081 22931 -913
rect 23005 -1081 23039 -913
rect 23515 -1081 23549 -913
rect 23987 -535 24021 233
rect 24497 -535 24531 233
rect 24605 -535 24639 233
rect 25115 -535 25149 233
rect 23987 -1081 24021 -913
rect 24497 -1081 24531 -913
rect 24605 -1081 24639 -913
rect 25115 -1081 25149 -913
rect 25587 -535 25621 233
rect 26097 -535 26131 233
rect 26205 -535 26239 233
rect 26715 -535 26749 233
rect 25587 -1081 25621 -913
rect 26097 -1081 26131 -913
rect 26205 -1081 26239 -913
rect 26715 -1081 26749 -913
rect 27187 -535 27221 233
rect 27697 -535 27731 233
rect 27805 -535 27839 233
rect 28315 -535 28349 233
rect 27187 -1081 27221 -913
rect 27697 -1081 27731 -913
rect 27805 -1081 27839 -913
rect 28315 -1081 28349 -913
rect 28787 -535 28821 233
rect 29297 -535 29331 233
rect 29405 -535 29439 233
rect 29915 -535 29949 233
rect 28787 -1081 28821 -913
rect 29297 -1081 29331 -913
rect 29405 -1081 29439 -913
rect 29915 -1081 29949 -913
rect 30387 -535 30421 233
rect 30897 -535 30931 233
rect 31005 -535 31039 233
rect 31515 -535 31549 233
rect 30387 -1081 30421 -913
rect 30897 -1081 30931 -913
rect 31005 -1081 31039 -913
rect 31515 -1081 31549 -913
rect 31987 -535 32021 233
rect 32497 -535 32531 233
rect 32605 -535 32639 233
rect 33115 -535 33149 233
rect 31987 -1081 32021 -913
rect 32497 -1081 32531 -913
rect 32605 -1081 32639 -913
rect 33115 -1081 33149 -913
rect 33587 -535 33621 233
rect 34097 -535 34131 233
rect 34205 -535 34239 233
rect 34715 -535 34749 233
rect 33587 -1081 33621 -913
rect 34097 -1081 34131 -913
rect 34205 -1081 34239 -913
rect 34715 -1081 34749 -913
rect 35187 -535 35221 233
rect 35697 -535 35731 233
rect 35805 -535 35839 233
rect 36315 -535 36349 233
rect 35187 -1081 35221 -913
rect 35697 -1081 35731 -913
rect 35805 -1081 35839 -913
rect 36315 -1081 36349 -913
rect 36787 -535 36821 233
rect 37297 -535 37331 233
rect 37405 -535 37439 233
rect 37915 -535 37949 233
rect 36787 -1081 36821 -913
rect 37297 -1081 37331 -913
rect 37405 -1081 37439 -913
rect 37915 -1081 37949 -913
rect -13 -2335 21 -1567
rect 497 -2335 531 -1567
rect 605 -2335 639 -1567
rect 1115 -2335 1149 -1567
rect -13 -2881 21 -2713
rect 497 -2881 531 -2713
rect 605 -2881 639 -2713
rect 1115 -2881 1149 -2713
rect 1587 -2335 1621 -1567
rect 2097 -2335 2131 -1567
rect 2205 -2335 2239 -1567
rect 2715 -2335 2749 -1567
rect 1587 -2881 1621 -2713
rect 2097 -2881 2131 -2713
rect 2205 -2881 2239 -2713
rect 2715 -2881 2749 -2713
rect 3187 -2335 3221 -1567
rect 3697 -2335 3731 -1567
rect 3805 -2335 3839 -1567
rect 4315 -2335 4349 -1567
rect 3187 -2881 3221 -2713
rect 3697 -2881 3731 -2713
rect 3805 -2881 3839 -2713
rect 4315 -2881 4349 -2713
rect 4787 -2335 4821 -1567
rect 5297 -2335 5331 -1567
rect 5405 -2335 5439 -1567
rect 5915 -2335 5949 -1567
rect 4787 -2881 4821 -2713
rect 5297 -2881 5331 -2713
rect 5405 -2881 5439 -2713
rect 5915 -2881 5949 -2713
rect 6387 -2335 6421 -1567
rect 6897 -2335 6931 -1567
rect 7005 -2335 7039 -1567
rect 7515 -2335 7549 -1567
rect 6387 -2881 6421 -2713
rect 6897 -2881 6931 -2713
rect 7005 -2881 7039 -2713
rect 7515 -2881 7549 -2713
rect 7987 -2335 8021 -1567
rect 8497 -2335 8531 -1567
rect 8605 -2335 8639 -1567
rect 9115 -2335 9149 -1567
rect 7987 -2881 8021 -2713
rect 8497 -2881 8531 -2713
rect 8605 -2881 8639 -2713
rect 9115 -2881 9149 -2713
rect 9587 -2335 9621 -1567
rect 10097 -2335 10131 -1567
rect 10205 -2335 10239 -1567
rect 10715 -2335 10749 -1567
rect 9587 -2881 9621 -2713
rect 10097 -2881 10131 -2713
rect 10205 -2881 10239 -2713
rect 10715 -2881 10749 -2713
rect 11187 -2335 11221 -1567
rect 11697 -2335 11731 -1567
rect 11805 -2335 11839 -1567
rect 12315 -2335 12349 -1567
rect 11187 -2881 11221 -2713
rect 11697 -2881 11731 -2713
rect 11805 -2881 11839 -2713
rect 12315 -2881 12349 -2713
rect 12787 -2335 12821 -1567
rect 13297 -2335 13331 -1567
rect 13405 -2335 13439 -1567
rect 13915 -2335 13949 -1567
rect 12787 -2881 12821 -2713
rect 13297 -2881 13331 -2713
rect 13405 -2881 13439 -2713
rect 13915 -2881 13949 -2713
rect 14387 -2335 14421 -1567
rect 14897 -2335 14931 -1567
rect 15005 -2335 15039 -1567
rect 15515 -2335 15549 -1567
rect 14387 -2881 14421 -2713
rect 14897 -2881 14931 -2713
rect 15005 -2881 15039 -2713
rect 15515 -2881 15549 -2713
rect 15987 -2335 16021 -1567
rect 16497 -2335 16531 -1567
rect 16605 -2335 16639 -1567
rect 17115 -2335 17149 -1567
rect 15987 -2881 16021 -2713
rect 16497 -2881 16531 -2713
rect 16605 -2881 16639 -2713
rect 17115 -2881 17149 -2713
rect 17587 -2335 17621 -1567
rect 18097 -2335 18131 -1567
rect 18205 -2335 18239 -1567
rect 18715 -2335 18749 -1567
rect 17587 -2881 17621 -2713
rect 18097 -2881 18131 -2713
rect 18205 -2881 18239 -2713
rect 18715 -2881 18749 -2713
rect 19187 -2335 19221 -1567
rect 19697 -2335 19731 -1567
rect 19805 -2335 19839 -1567
rect 20315 -2335 20349 -1567
rect 19187 -2881 19221 -2713
rect 19697 -2881 19731 -2713
rect 19805 -2881 19839 -2713
rect 20315 -2881 20349 -2713
rect 20787 -2335 20821 -1567
rect 21297 -2335 21331 -1567
rect 21405 -2335 21439 -1567
rect 21915 -2335 21949 -1567
rect 20787 -2881 20821 -2713
rect 21297 -2881 21331 -2713
rect 21405 -2881 21439 -2713
rect 21915 -2881 21949 -2713
rect 22387 -2335 22421 -1567
rect 22897 -2335 22931 -1567
rect 23005 -2335 23039 -1567
rect 23515 -2335 23549 -1567
rect 22387 -2881 22421 -2713
rect 22897 -2881 22931 -2713
rect 23005 -2881 23039 -2713
rect 23515 -2881 23549 -2713
rect 23987 -2335 24021 -1567
rect 24497 -2335 24531 -1567
rect 24605 -2335 24639 -1567
rect 25115 -2335 25149 -1567
rect 23987 -2881 24021 -2713
rect 24497 -2881 24531 -2713
rect 24605 -2881 24639 -2713
rect 25115 -2881 25149 -2713
rect 25587 -2335 25621 -1567
rect 26097 -2335 26131 -1567
rect 26205 -2335 26239 -1567
rect 26715 -2335 26749 -1567
rect 25587 -2881 25621 -2713
rect 26097 -2881 26131 -2713
rect 26205 -2881 26239 -2713
rect 26715 -2881 26749 -2713
rect 27187 -2335 27221 -1567
rect 27697 -2335 27731 -1567
rect 27805 -2335 27839 -1567
rect 28315 -2335 28349 -1567
rect 27187 -2881 27221 -2713
rect 27697 -2881 27731 -2713
rect 27805 -2881 27839 -2713
rect 28315 -2881 28349 -2713
rect 28787 -2335 28821 -1567
rect 29297 -2335 29331 -1567
rect 29405 -2335 29439 -1567
rect 29915 -2335 29949 -1567
rect 28787 -2881 28821 -2713
rect 29297 -2881 29331 -2713
rect 29405 -2881 29439 -2713
rect 29915 -2881 29949 -2713
rect 30387 -2335 30421 -1567
rect 30897 -2335 30931 -1567
rect 31005 -2335 31039 -1567
rect 31515 -2335 31549 -1567
rect 30387 -2881 30421 -2713
rect 30897 -2881 30931 -2713
rect 31005 -2881 31039 -2713
rect 31515 -2881 31549 -2713
rect 31987 -2335 32021 -1567
rect 32497 -2335 32531 -1567
rect 32605 -2335 32639 -1567
rect 33115 -2335 33149 -1567
rect 31987 -2881 32021 -2713
rect 32497 -2881 32531 -2713
rect 32605 -2881 32639 -2713
rect 33115 -2881 33149 -2713
rect 33587 -2335 33621 -1567
rect 34097 -2335 34131 -1567
rect 34205 -2335 34239 -1567
rect 34715 -2335 34749 -1567
rect 33587 -2881 33621 -2713
rect 34097 -2881 34131 -2713
rect 34205 -2881 34239 -2713
rect 34715 -2881 34749 -2713
rect 35187 -2335 35221 -1567
rect 35697 -2335 35731 -1567
rect 35805 -2335 35839 -1567
rect 36315 -2335 36349 -1567
rect 35187 -2881 35221 -2713
rect 35697 -2881 35731 -2713
rect 35805 -2881 35839 -2713
rect 36315 -2881 36349 -2713
rect 36787 -2335 36821 -1567
rect 37297 -2335 37331 -1567
rect 37405 -2335 37439 -1567
rect 37915 -2335 37949 -1567
rect 36787 -2881 36821 -2713
rect 37297 -2881 37331 -2713
rect 37405 -2881 37439 -2713
rect 37915 -2881 37949 -2713
rect -13 -4135 21 -3367
rect 497 -4135 531 -3367
rect 605 -4135 639 -3367
rect 1115 -4135 1149 -3367
rect -13 -4681 21 -4513
rect 497 -4681 531 -4513
rect 605 -4681 639 -4513
rect 1115 -4681 1149 -4513
rect 1587 -4135 1621 -3367
rect 2097 -4135 2131 -3367
rect 2205 -4135 2239 -3367
rect 2715 -4135 2749 -3367
rect 1587 -4681 1621 -4513
rect 2097 -4681 2131 -4513
rect 2205 -4681 2239 -4513
rect 2715 -4681 2749 -4513
rect 3187 -4135 3221 -3367
rect 3697 -4135 3731 -3367
rect 3805 -4135 3839 -3367
rect 4315 -4135 4349 -3367
rect 3187 -4681 3221 -4513
rect 3697 -4681 3731 -4513
rect 3805 -4681 3839 -4513
rect 4315 -4681 4349 -4513
rect 4787 -4135 4821 -3367
rect 5297 -4135 5331 -3367
rect 5405 -4135 5439 -3367
rect 5915 -4135 5949 -3367
rect 4787 -4681 4821 -4513
rect 5297 -4681 5331 -4513
rect 5405 -4681 5439 -4513
rect 5915 -4681 5949 -4513
rect 6387 -4135 6421 -3367
rect 6897 -4135 6931 -3367
rect 7005 -4135 7039 -3367
rect 7515 -4135 7549 -3367
rect 6387 -4681 6421 -4513
rect 6897 -4681 6931 -4513
rect 7005 -4681 7039 -4513
rect 7515 -4681 7549 -4513
rect 7987 -4135 8021 -3367
rect 8497 -4135 8531 -3367
rect 8605 -4135 8639 -3367
rect 9115 -4135 9149 -3367
rect 7987 -4681 8021 -4513
rect 8497 -4681 8531 -4513
rect 8605 -4681 8639 -4513
rect 9115 -4681 9149 -4513
rect 9587 -4135 9621 -3367
rect 10097 -4135 10131 -3367
rect 10205 -4135 10239 -3367
rect 10715 -4135 10749 -3367
rect 9587 -4681 9621 -4513
rect 10097 -4681 10131 -4513
rect 10205 -4681 10239 -4513
rect 10715 -4681 10749 -4513
rect 11187 -4135 11221 -3367
rect 11697 -4135 11731 -3367
rect 11805 -4135 11839 -3367
rect 12315 -4135 12349 -3367
rect 11187 -4681 11221 -4513
rect 11697 -4681 11731 -4513
rect 11805 -4681 11839 -4513
rect 12315 -4681 12349 -4513
rect 12787 -4135 12821 -3367
rect 13297 -4135 13331 -3367
rect 13405 -4135 13439 -3367
rect 13915 -4135 13949 -3367
rect 12787 -4681 12821 -4513
rect 13297 -4681 13331 -4513
rect 13405 -4681 13439 -4513
rect 13915 -4681 13949 -4513
rect 14387 -4135 14421 -3367
rect 14897 -4135 14931 -3367
rect 15005 -4135 15039 -3367
rect 15515 -4135 15549 -3367
rect 14387 -4681 14421 -4513
rect 14897 -4681 14931 -4513
rect 15005 -4681 15039 -4513
rect 15515 -4681 15549 -4513
rect 15987 -4135 16021 -3367
rect 16497 -4135 16531 -3367
rect 16605 -4135 16639 -3367
rect 17115 -4135 17149 -3367
rect 15987 -4681 16021 -4513
rect 16497 -4681 16531 -4513
rect 16605 -4681 16639 -4513
rect 17115 -4681 17149 -4513
rect 17587 -4135 17621 -3367
rect 18097 -4135 18131 -3367
rect 18205 -4135 18239 -3367
rect 18715 -4135 18749 -3367
rect 17587 -4681 17621 -4513
rect 18097 -4681 18131 -4513
rect 18205 -4681 18239 -4513
rect 18715 -4681 18749 -4513
rect 19187 -4135 19221 -3367
rect 19697 -4135 19731 -3367
rect 19805 -4135 19839 -3367
rect 20315 -4135 20349 -3367
rect 19187 -4681 19221 -4513
rect 19697 -4681 19731 -4513
rect 19805 -4681 19839 -4513
rect 20315 -4681 20349 -4513
rect 20787 -4135 20821 -3367
rect 21297 -4135 21331 -3367
rect 21405 -4135 21439 -3367
rect 21915 -4135 21949 -3367
rect 20787 -4681 20821 -4513
rect 21297 -4681 21331 -4513
rect 21405 -4681 21439 -4513
rect 21915 -4681 21949 -4513
rect 22387 -4135 22421 -3367
rect 22897 -4135 22931 -3367
rect 23005 -4135 23039 -3367
rect 23515 -4135 23549 -3367
rect 22387 -4681 22421 -4513
rect 22897 -4681 22931 -4513
rect 23005 -4681 23039 -4513
rect 23515 -4681 23549 -4513
rect 23987 -4135 24021 -3367
rect 24497 -4135 24531 -3367
rect 24605 -4135 24639 -3367
rect 25115 -4135 25149 -3367
rect 23987 -4681 24021 -4513
rect 24497 -4681 24531 -4513
rect 24605 -4681 24639 -4513
rect 25115 -4681 25149 -4513
rect 25587 -4135 25621 -3367
rect 26097 -4135 26131 -3367
rect 26205 -4135 26239 -3367
rect 26715 -4135 26749 -3367
rect 25587 -4681 25621 -4513
rect 26097 -4681 26131 -4513
rect 26205 -4681 26239 -4513
rect 26715 -4681 26749 -4513
rect 27187 -4135 27221 -3367
rect 27697 -4135 27731 -3367
rect 27805 -4135 27839 -3367
rect 28315 -4135 28349 -3367
rect 27187 -4681 27221 -4513
rect 27697 -4681 27731 -4513
rect 27805 -4681 27839 -4513
rect 28315 -4681 28349 -4513
rect 28787 -4135 28821 -3367
rect 29297 -4135 29331 -3367
rect 29405 -4135 29439 -3367
rect 29915 -4135 29949 -3367
rect 28787 -4681 28821 -4513
rect 29297 -4681 29331 -4513
rect 29405 -4681 29439 -4513
rect 29915 -4681 29949 -4513
rect 30387 -4135 30421 -3367
rect 30897 -4135 30931 -3367
rect 31005 -4135 31039 -3367
rect 31515 -4135 31549 -3367
rect 30387 -4681 30421 -4513
rect 30897 -4681 30931 -4513
rect 31005 -4681 31039 -4513
rect 31515 -4681 31549 -4513
rect 31987 -4135 32021 -3367
rect 32497 -4135 32531 -3367
rect 32605 -4135 32639 -3367
rect 33115 -4135 33149 -3367
rect 31987 -4681 32021 -4513
rect 32497 -4681 32531 -4513
rect 32605 -4681 32639 -4513
rect 33115 -4681 33149 -4513
rect 33587 -4135 33621 -3367
rect 34097 -4135 34131 -3367
rect 34205 -4135 34239 -3367
rect 34715 -4135 34749 -3367
rect 33587 -4681 33621 -4513
rect 34097 -4681 34131 -4513
rect 34205 -4681 34239 -4513
rect 34715 -4681 34749 -4513
rect 35187 -4135 35221 -3367
rect 35697 -4135 35731 -3367
rect 35805 -4135 35839 -3367
rect 36315 -4135 36349 -3367
rect 35187 -4681 35221 -4513
rect 35697 -4681 35731 -4513
rect 35805 -4681 35839 -4513
rect 36315 -4681 36349 -4513
rect 36787 -4135 36821 -3367
rect 37297 -4135 37331 -3367
rect 37405 -4135 37439 -3367
rect 37915 -4135 37949 -3367
rect 36787 -4681 36821 -4513
rect 37297 -4681 37331 -4513
rect 37405 -4681 37439 -4513
rect 37915 -4681 37949 -4513
rect -24 -8400 10 -8232
rect 504 -8400 538 -8232
rect 612 -8400 646 -8232
rect 1140 -8400 1174 -8232
rect -24 -9526 10 -8758
rect 504 -9526 538 -8758
rect 612 -9526 646 -8758
rect 1140 -9526 1174 -8758
rect 1576 -8400 1610 -8232
rect 2104 -8400 2138 -8232
rect 2212 -8400 2246 -8232
rect 2740 -8400 2774 -8232
rect 1576 -9526 1610 -8758
rect 2104 -9526 2138 -8758
rect 2212 -9526 2246 -8758
rect 2740 -9526 2774 -8758
rect 3176 -8400 3210 -8232
rect 3704 -8400 3738 -8232
rect 3812 -8400 3846 -8232
rect 4340 -8400 4374 -8232
rect 3176 -9526 3210 -8758
rect 3704 -9526 3738 -8758
rect 3812 -9526 3846 -8758
rect 4340 -9526 4374 -8758
rect 4776 -8400 4810 -8232
rect 5304 -8400 5338 -8232
rect 5412 -8400 5446 -8232
rect 5940 -8400 5974 -8232
rect 4776 -9526 4810 -8758
rect 5304 -9526 5338 -8758
rect 5412 -9526 5446 -8758
rect 5940 -9526 5974 -8758
rect 6376 -8400 6410 -8232
rect 6904 -8400 6938 -8232
rect 7012 -8400 7046 -8232
rect 7540 -8400 7574 -8232
rect 6376 -9526 6410 -8758
rect 6904 -9526 6938 -8758
rect 7012 -9526 7046 -8758
rect 7540 -9526 7574 -8758
rect 7976 -8400 8010 -8232
rect 8504 -8400 8538 -8232
rect 8612 -8400 8646 -8232
rect 9140 -8400 9174 -8232
rect 7976 -9526 8010 -8758
rect 8504 -9526 8538 -8758
rect 8612 -9526 8646 -8758
rect 9140 -9526 9174 -8758
rect 9576 -8400 9610 -8232
rect 10104 -8400 10138 -8232
rect 10212 -8400 10246 -8232
rect 10740 -8400 10774 -8232
rect 9576 -9526 9610 -8758
rect 10104 -9526 10138 -8758
rect 10212 -9526 10246 -8758
rect 10740 -9526 10774 -8758
rect 11176 -8400 11210 -8232
rect 11704 -8400 11738 -8232
rect 11812 -8400 11846 -8232
rect 12340 -8400 12374 -8232
rect 11176 -9526 11210 -8758
rect 11704 -9526 11738 -8758
rect 11812 -9526 11846 -8758
rect 12340 -9526 12374 -8758
rect 12776 -8400 12810 -8232
rect 13304 -8400 13338 -8232
rect 13412 -8400 13446 -8232
rect 13940 -8400 13974 -8232
rect 12776 -9526 12810 -8758
rect 13304 -9526 13338 -8758
rect 13412 -9526 13446 -8758
rect 13940 -9526 13974 -8758
rect 14376 -8400 14410 -8232
rect 14904 -8400 14938 -8232
rect 15012 -8400 15046 -8232
rect 15540 -8400 15574 -8232
rect 14376 -9526 14410 -8758
rect 14904 -9526 14938 -8758
rect 15012 -9526 15046 -8758
rect 15540 -9526 15574 -8758
rect 15976 -8400 16010 -8232
rect 16504 -8400 16538 -8232
rect 16612 -8400 16646 -8232
rect 17140 -8400 17174 -8232
rect 15976 -9526 16010 -8758
rect 16504 -9526 16538 -8758
rect 16612 -9526 16646 -8758
rect 17140 -9526 17174 -8758
rect 17576 -8400 17610 -8232
rect 18104 -8400 18138 -8232
rect 18212 -8400 18246 -8232
rect 18740 -8400 18774 -8232
rect 17576 -9526 17610 -8758
rect 18104 -9526 18138 -8758
rect 18212 -9526 18246 -8758
rect 18740 -9526 18774 -8758
rect 19176 -8400 19210 -8232
rect 19704 -8400 19738 -8232
rect 19812 -8400 19846 -8232
rect 20340 -8400 20374 -8232
rect 19176 -9526 19210 -8758
rect 19704 -9526 19738 -8758
rect 19812 -9526 19846 -8758
rect 20340 -9526 20374 -8758
rect 20776 -8400 20810 -8232
rect 21304 -8400 21338 -8232
rect 21412 -8400 21446 -8232
rect 21940 -8400 21974 -8232
rect 20776 -9526 20810 -8758
rect 21304 -9526 21338 -8758
rect 21412 -9526 21446 -8758
rect 21940 -9526 21974 -8758
rect 22376 -8400 22410 -8232
rect 22904 -8400 22938 -8232
rect 23012 -8400 23046 -8232
rect 23540 -8400 23574 -8232
rect 22376 -9526 22410 -8758
rect 22904 -9526 22938 -8758
rect 23012 -9526 23046 -8758
rect 23540 -9526 23574 -8758
rect 23976 -8400 24010 -8232
rect 24504 -8400 24538 -8232
rect 24612 -8400 24646 -8232
rect 25140 -8400 25174 -8232
rect 23976 -9526 24010 -8758
rect 24504 -9526 24538 -8758
rect 24612 -9526 24646 -8758
rect 25140 -9526 25174 -8758
rect 25576 -8400 25610 -8232
rect 26104 -8400 26138 -8232
rect 26212 -8400 26246 -8232
rect 26740 -8400 26774 -8232
rect 25576 -9526 25610 -8758
rect 26104 -9526 26138 -8758
rect 26212 -9526 26246 -8758
rect 26740 -9526 26774 -8758
rect 27176 -8400 27210 -8232
rect 27704 -8400 27738 -8232
rect 27812 -8400 27846 -8232
rect 28340 -8400 28374 -8232
rect 27176 -9526 27210 -8758
rect 27704 -9526 27738 -8758
rect 27812 -9526 27846 -8758
rect 28340 -9526 28374 -8758
rect 28776 -8400 28810 -8232
rect 29304 -8400 29338 -8232
rect 29412 -8400 29446 -8232
rect 29940 -8400 29974 -8232
rect 28776 -9526 28810 -8758
rect 29304 -9526 29338 -8758
rect 29412 -9526 29446 -8758
rect 29940 -9526 29974 -8758
rect 30376 -8400 30410 -8232
rect 30904 -8400 30938 -8232
rect 31012 -8400 31046 -8232
rect 31540 -8400 31574 -8232
rect 30376 -9526 30410 -8758
rect 30904 -9526 30938 -8758
rect 31012 -9526 31046 -8758
rect 31540 -9526 31574 -8758
rect 31976 -8400 32010 -8232
rect 32504 -8400 32538 -8232
rect 32612 -8400 32646 -8232
rect 33140 -8400 33174 -8232
rect 31976 -9526 32010 -8758
rect 32504 -9526 32538 -8758
rect 32612 -9526 32646 -8758
rect 33140 -9526 33174 -8758
rect 33576 -8400 33610 -8232
rect 34104 -8400 34138 -8232
rect 34212 -8400 34246 -8232
rect 34740 -8400 34774 -8232
rect 33576 -9526 33610 -8758
rect 34104 -9526 34138 -8758
rect 34212 -9526 34246 -8758
rect 34740 -9526 34774 -8758
rect 35176 -8400 35210 -8232
rect 35704 -8400 35738 -8232
rect 35812 -8400 35846 -8232
rect 36340 -8400 36374 -8232
rect 35176 -9526 35210 -8758
rect 35704 -9526 35738 -8758
rect 35812 -9526 35846 -8758
rect 36340 -9526 36374 -8758
rect 36776 -8400 36810 -8232
rect 37304 -8400 37338 -8232
rect 37412 -8400 37446 -8232
rect 37940 -8400 37974 -8232
rect 36776 -9526 36810 -8758
rect 37304 -9526 37338 -8758
rect 37412 -9526 37446 -8758
rect 37940 -9526 37974 -8758
rect -24 -10200 10 -10032
rect 504 -10200 538 -10032
rect 612 -10200 646 -10032
rect 1140 -10200 1174 -10032
rect -24 -11326 10 -10558
rect 504 -11326 538 -10558
rect 612 -11326 646 -10558
rect 1140 -11326 1174 -10558
rect 1576 -10200 1610 -10032
rect 2104 -10200 2138 -10032
rect 2212 -10200 2246 -10032
rect 2740 -10200 2774 -10032
rect 1576 -11326 1610 -10558
rect 2104 -11326 2138 -10558
rect 2212 -11326 2246 -10558
rect 2740 -11326 2774 -10558
rect 3176 -10200 3210 -10032
rect 3704 -10200 3738 -10032
rect 3812 -10200 3846 -10032
rect 4340 -10200 4374 -10032
rect 3176 -11326 3210 -10558
rect 3704 -11326 3738 -10558
rect 3812 -11326 3846 -10558
rect 4340 -11326 4374 -10558
rect 4776 -10200 4810 -10032
rect 5304 -10200 5338 -10032
rect 5412 -10200 5446 -10032
rect 5940 -10200 5974 -10032
rect 4776 -11326 4810 -10558
rect 5304 -11326 5338 -10558
rect 5412 -11326 5446 -10558
rect 5940 -11326 5974 -10558
rect 6376 -10200 6410 -10032
rect 6904 -10200 6938 -10032
rect 7012 -10200 7046 -10032
rect 7540 -10200 7574 -10032
rect 6376 -11326 6410 -10558
rect 6904 -11326 6938 -10558
rect 7012 -11326 7046 -10558
rect 7540 -11326 7574 -10558
rect 7976 -10200 8010 -10032
rect 8504 -10200 8538 -10032
rect 8612 -10200 8646 -10032
rect 9140 -10200 9174 -10032
rect 7976 -11326 8010 -10558
rect 8504 -11326 8538 -10558
rect 8612 -11326 8646 -10558
rect 9140 -11326 9174 -10558
rect 9576 -10200 9610 -10032
rect 10104 -10200 10138 -10032
rect 10212 -10200 10246 -10032
rect 10740 -10200 10774 -10032
rect 9576 -11326 9610 -10558
rect 10104 -11326 10138 -10558
rect 10212 -11326 10246 -10558
rect 10740 -11326 10774 -10558
rect 11176 -10200 11210 -10032
rect 11704 -10200 11738 -10032
rect 11812 -10200 11846 -10032
rect 12340 -10200 12374 -10032
rect 11176 -11326 11210 -10558
rect 11704 -11326 11738 -10558
rect 11812 -11326 11846 -10558
rect 12340 -11326 12374 -10558
rect 12776 -10200 12810 -10032
rect 13304 -10200 13338 -10032
rect 13412 -10200 13446 -10032
rect 13940 -10200 13974 -10032
rect 12776 -11326 12810 -10558
rect 13304 -11326 13338 -10558
rect 13412 -11326 13446 -10558
rect 13940 -11326 13974 -10558
rect 14376 -10200 14410 -10032
rect 14904 -10200 14938 -10032
rect 15012 -10200 15046 -10032
rect 15540 -10200 15574 -10032
rect 14376 -11326 14410 -10558
rect 14904 -11326 14938 -10558
rect 15012 -11326 15046 -10558
rect 15540 -11326 15574 -10558
rect 15976 -10200 16010 -10032
rect 16504 -10200 16538 -10032
rect 16612 -10200 16646 -10032
rect 17140 -10200 17174 -10032
rect 15976 -11326 16010 -10558
rect 16504 -11326 16538 -10558
rect 16612 -11326 16646 -10558
rect 17140 -11326 17174 -10558
rect 17576 -10200 17610 -10032
rect 18104 -10200 18138 -10032
rect 18212 -10200 18246 -10032
rect 18740 -10200 18774 -10032
rect 17576 -11326 17610 -10558
rect 18104 -11326 18138 -10558
rect 18212 -11326 18246 -10558
rect 18740 -11326 18774 -10558
rect 19176 -10200 19210 -10032
rect 19704 -10200 19738 -10032
rect 19812 -10200 19846 -10032
rect 20340 -10200 20374 -10032
rect 19176 -11326 19210 -10558
rect 19704 -11326 19738 -10558
rect 19812 -11326 19846 -10558
rect 20340 -11326 20374 -10558
rect 20776 -10200 20810 -10032
rect 21304 -10200 21338 -10032
rect 21412 -10200 21446 -10032
rect 21940 -10200 21974 -10032
rect 20776 -11326 20810 -10558
rect 21304 -11326 21338 -10558
rect 21412 -11326 21446 -10558
rect 21940 -11326 21974 -10558
rect 22376 -10200 22410 -10032
rect 22904 -10200 22938 -10032
rect 23012 -10200 23046 -10032
rect 23540 -10200 23574 -10032
rect 22376 -11326 22410 -10558
rect 22904 -11326 22938 -10558
rect 23012 -11326 23046 -10558
rect 23540 -11326 23574 -10558
rect 23976 -10200 24010 -10032
rect 24504 -10200 24538 -10032
rect 24612 -10200 24646 -10032
rect 25140 -10200 25174 -10032
rect 23976 -11326 24010 -10558
rect 24504 -11326 24538 -10558
rect 24612 -11326 24646 -10558
rect 25140 -11326 25174 -10558
rect 25576 -10200 25610 -10032
rect 26104 -10200 26138 -10032
rect 26212 -10200 26246 -10032
rect 26740 -10200 26774 -10032
rect 25576 -11326 25610 -10558
rect 26104 -11326 26138 -10558
rect 26212 -11326 26246 -10558
rect 26740 -11326 26774 -10558
rect 27176 -10200 27210 -10032
rect 27704 -10200 27738 -10032
rect 27812 -10200 27846 -10032
rect 28340 -10200 28374 -10032
rect 27176 -11326 27210 -10558
rect 27704 -11326 27738 -10558
rect 27812 -11326 27846 -10558
rect 28340 -11326 28374 -10558
rect 28776 -10200 28810 -10032
rect 29304 -10200 29338 -10032
rect 29412 -10200 29446 -10032
rect 29940 -10200 29974 -10032
rect 28776 -11326 28810 -10558
rect 29304 -11326 29338 -10558
rect 29412 -11326 29446 -10558
rect 29940 -11326 29974 -10558
rect 30376 -10200 30410 -10032
rect 30904 -10200 30938 -10032
rect 31012 -10200 31046 -10032
rect 31540 -10200 31574 -10032
rect 30376 -11326 30410 -10558
rect 30904 -11326 30938 -10558
rect 31012 -11326 31046 -10558
rect 31540 -11326 31574 -10558
rect 31976 -10200 32010 -10032
rect 32504 -10200 32538 -10032
rect 32612 -10200 32646 -10032
rect 33140 -10200 33174 -10032
rect 31976 -11326 32010 -10558
rect 32504 -11326 32538 -10558
rect 32612 -11326 32646 -10558
rect 33140 -11326 33174 -10558
rect 33576 -10200 33610 -10032
rect 34104 -10200 34138 -10032
rect 34212 -10200 34246 -10032
rect 34740 -10200 34774 -10032
rect 33576 -11326 33610 -10558
rect 34104 -11326 34138 -10558
rect 34212 -11326 34246 -10558
rect 34740 -11326 34774 -10558
rect 35176 -10200 35210 -10032
rect 35704 -10200 35738 -10032
rect 35812 -10200 35846 -10032
rect 36340 -10200 36374 -10032
rect 35176 -11326 35210 -10558
rect 35704 -11326 35738 -10558
rect 35812 -11326 35846 -10558
rect 36340 -11326 36374 -10558
rect 36776 -10200 36810 -10032
rect 37304 -10200 37338 -10032
rect 37412 -10200 37446 -10032
rect 37940 -10200 37974 -10032
rect 36776 -11326 36810 -10558
rect 37304 -11326 37338 -10558
rect 37412 -11326 37446 -10558
rect 37940 -11326 37974 -10558
rect -24 -12000 10 -11832
rect 504 -12000 538 -11832
rect 612 -12000 646 -11832
rect 1140 -12000 1174 -11832
rect -24 -13126 10 -12358
rect 504 -13126 538 -12358
rect 612 -13126 646 -12358
rect 1140 -13126 1174 -12358
rect 1576 -12000 1610 -11832
rect 2104 -12000 2138 -11832
rect 2212 -12000 2246 -11832
rect 2740 -12000 2774 -11832
rect 1576 -13126 1610 -12358
rect 2104 -13126 2138 -12358
rect 2212 -13126 2246 -12358
rect 2740 -13126 2774 -12358
rect 3176 -12000 3210 -11832
rect 3704 -12000 3738 -11832
rect 3812 -12000 3846 -11832
rect 4340 -12000 4374 -11832
rect 3176 -13126 3210 -12358
rect 3704 -13126 3738 -12358
rect 3812 -13126 3846 -12358
rect 4340 -13126 4374 -12358
rect 4776 -12000 4810 -11832
rect 5304 -12000 5338 -11832
rect 5412 -12000 5446 -11832
rect 5940 -12000 5974 -11832
rect 4776 -13126 4810 -12358
rect 5304 -13126 5338 -12358
rect 5412 -13126 5446 -12358
rect 5940 -13126 5974 -12358
rect 6376 -12000 6410 -11832
rect 6904 -12000 6938 -11832
rect 7012 -12000 7046 -11832
rect 7540 -12000 7574 -11832
rect 6376 -13126 6410 -12358
rect 6904 -13126 6938 -12358
rect 7012 -13126 7046 -12358
rect 7540 -13126 7574 -12358
rect 7976 -12000 8010 -11832
rect 8504 -12000 8538 -11832
rect 8612 -12000 8646 -11832
rect 9140 -12000 9174 -11832
rect 7976 -13126 8010 -12358
rect 8504 -13126 8538 -12358
rect 8612 -13126 8646 -12358
rect 9140 -13126 9174 -12358
rect 9576 -12000 9610 -11832
rect 10104 -12000 10138 -11832
rect 10212 -12000 10246 -11832
rect 10740 -12000 10774 -11832
rect 9576 -13126 9610 -12358
rect 10104 -13126 10138 -12358
rect 10212 -13126 10246 -12358
rect 10740 -13126 10774 -12358
rect 11176 -12000 11210 -11832
rect 11704 -12000 11738 -11832
rect 11812 -12000 11846 -11832
rect 12340 -12000 12374 -11832
rect 11176 -13126 11210 -12358
rect 11704 -13126 11738 -12358
rect 11812 -13126 11846 -12358
rect 12340 -13126 12374 -12358
rect 12776 -12000 12810 -11832
rect 13304 -12000 13338 -11832
rect 13412 -12000 13446 -11832
rect 13940 -12000 13974 -11832
rect 12776 -13126 12810 -12358
rect 13304 -13126 13338 -12358
rect 13412 -13126 13446 -12358
rect 13940 -13126 13974 -12358
rect 14376 -12000 14410 -11832
rect 14904 -12000 14938 -11832
rect 15012 -12000 15046 -11832
rect 15540 -12000 15574 -11832
rect 14376 -13126 14410 -12358
rect 14904 -13126 14938 -12358
rect 15012 -13126 15046 -12358
rect 15540 -13126 15574 -12358
rect 15976 -12000 16010 -11832
rect 16504 -12000 16538 -11832
rect 16612 -12000 16646 -11832
rect 17140 -12000 17174 -11832
rect 15976 -13126 16010 -12358
rect 16504 -13126 16538 -12358
rect 16612 -13126 16646 -12358
rect 17140 -13126 17174 -12358
rect 17576 -12000 17610 -11832
rect 18104 -12000 18138 -11832
rect 18212 -12000 18246 -11832
rect 18740 -12000 18774 -11832
rect 17576 -13126 17610 -12358
rect 18104 -13126 18138 -12358
rect 18212 -13126 18246 -12358
rect 18740 -13126 18774 -12358
rect 19176 -12000 19210 -11832
rect 19704 -12000 19738 -11832
rect 19812 -12000 19846 -11832
rect 20340 -12000 20374 -11832
rect 19176 -13126 19210 -12358
rect 19704 -13126 19738 -12358
rect 19812 -13126 19846 -12358
rect 20340 -13126 20374 -12358
rect 20776 -12000 20810 -11832
rect 21304 -12000 21338 -11832
rect 21412 -12000 21446 -11832
rect 21940 -12000 21974 -11832
rect 20776 -13126 20810 -12358
rect 21304 -13126 21338 -12358
rect 21412 -13126 21446 -12358
rect 21940 -13126 21974 -12358
rect 22376 -12000 22410 -11832
rect 22904 -12000 22938 -11832
rect 23012 -12000 23046 -11832
rect 23540 -12000 23574 -11832
rect 22376 -13126 22410 -12358
rect 22904 -13126 22938 -12358
rect 23012 -13126 23046 -12358
rect 23540 -13126 23574 -12358
rect 23976 -12000 24010 -11832
rect 24504 -12000 24538 -11832
rect 24612 -12000 24646 -11832
rect 25140 -12000 25174 -11832
rect 23976 -13126 24010 -12358
rect 24504 -13126 24538 -12358
rect 24612 -13126 24646 -12358
rect 25140 -13126 25174 -12358
rect 25576 -12000 25610 -11832
rect 26104 -12000 26138 -11832
rect 26212 -12000 26246 -11832
rect 26740 -12000 26774 -11832
rect 25576 -13126 25610 -12358
rect 26104 -13126 26138 -12358
rect 26212 -13126 26246 -12358
rect 26740 -13126 26774 -12358
rect 27176 -12000 27210 -11832
rect 27704 -12000 27738 -11832
rect 27812 -12000 27846 -11832
rect 28340 -12000 28374 -11832
rect 27176 -13126 27210 -12358
rect 27704 -13126 27738 -12358
rect 27812 -13126 27846 -12358
rect 28340 -13126 28374 -12358
rect 28776 -12000 28810 -11832
rect 29304 -12000 29338 -11832
rect 29412 -12000 29446 -11832
rect 29940 -12000 29974 -11832
rect 28776 -13126 28810 -12358
rect 29304 -13126 29338 -12358
rect 29412 -13126 29446 -12358
rect 29940 -13126 29974 -12358
rect 30376 -12000 30410 -11832
rect 30904 -12000 30938 -11832
rect 31012 -12000 31046 -11832
rect 31540 -12000 31574 -11832
rect 30376 -13126 30410 -12358
rect 30904 -13126 30938 -12358
rect 31012 -13126 31046 -12358
rect 31540 -13126 31574 -12358
rect 31976 -12000 32010 -11832
rect 32504 -12000 32538 -11832
rect 32612 -12000 32646 -11832
rect 33140 -12000 33174 -11832
rect 31976 -13126 32010 -12358
rect 32504 -13126 32538 -12358
rect 32612 -13126 32646 -12358
rect 33140 -13126 33174 -12358
rect 33576 -12000 33610 -11832
rect 34104 -12000 34138 -11832
rect 34212 -12000 34246 -11832
rect 34740 -12000 34774 -11832
rect 33576 -13126 33610 -12358
rect 34104 -13126 34138 -12358
rect 34212 -13126 34246 -12358
rect 34740 -13126 34774 -12358
rect 35176 -12000 35210 -11832
rect 35704 -12000 35738 -11832
rect 35812 -12000 35846 -11832
rect 36340 -12000 36374 -11832
rect 35176 -13126 35210 -12358
rect 35704 -13126 35738 -12358
rect 35812 -13126 35846 -12358
rect 36340 -13126 36374 -12358
rect 36776 -12000 36810 -11832
rect 37304 -12000 37338 -11832
rect 37412 -12000 37446 -11832
rect 37940 -12000 37974 -11832
rect 36776 -13126 36810 -12358
rect 37304 -13126 37338 -12358
rect 37412 -13126 37446 -12358
rect 37940 -13126 37974 -12358
rect -24 -13800 10 -13632
rect 504 -13800 538 -13632
rect 612 -13800 646 -13632
rect 1140 -13800 1174 -13632
rect -24 -14926 10 -14158
rect 504 -14926 538 -14158
rect 612 -14926 646 -14158
rect 1140 -14926 1174 -14158
rect 1576 -13800 1610 -13632
rect 2104 -13800 2138 -13632
rect 2212 -13800 2246 -13632
rect 2740 -13800 2774 -13632
rect 1576 -14926 1610 -14158
rect 2104 -14926 2138 -14158
rect 2212 -14926 2246 -14158
rect 2740 -14926 2774 -14158
rect 3176 -13800 3210 -13632
rect 3704 -13800 3738 -13632
rect 3812 -13800 3846 -13632
rect 4340 -13800 4374 -13632
rect 3176 -14926 3210 -14158
rect 3704 -14926 3738 -14158
rect 3812 -14926 3846 -14158
rect 4340 -14926 4374 -14158
rect 4776 -13800 4810 -13632
rect 5304 -13800 5338 -13632
rect 5412 -13800 5446 -13632
rect 5940 -13800 5974 -13632
rect 4776 -14926 4810 -14158
rect 5304 -14926 5338 -14158
rect 5412 -14926 5446 -14158
rect 5940 -14926 5974 -14158
rect 6376 -13800 6410 -13632
rect 6904 -13800 6938 -13632
rect 7012 -13800 7046 -13632
rect 7540 -13800 7574 -13632
rect 6376 -14926 6410 -14158
rect 6904 -14926 6938 -14158
rect 7012 -14926 7046 -14158
rect 7540 -14926 7574 -14158
rect 7976 -13800 8010 -13632
rect 8504 -13800 8538 -13632
rect 8612 -13800 8646 -13632
rect 9140 -13800 9174 -13632
rect 7976 -14926 8010 -14158
rect 8504 -14926 8538 -14158
rect 8612 -14926 8646 -14158
rect 9140 -14926 9174 -14158
rect 9576 -13800 9610 -13632
rect 10104 -13800 10138 -13632
rect 10212 -13800 10246 -13632
rect 10740 -13800 10774 -13632
rect 9576 -14926 9610 -14158
rect 10104 -14926 10138 -14158
rect 10212 -14926 10246 -14158
rect 10740 -14926 10774 -14158
rect 11176 -13800 11210 -13632
rect 11704 -13800 11738 -13632
rect 11812 -13800 11846 -13632
rect 12340 -13800 12374 -13632
rect 11176 -14926 11210 -14158
rect 11704 -14926 11738 -14158
rect 11812 -14926 11846 -14158
rect 12340 -14926 12374 -14158
rect 12776 -13800 12810 -13632
rect 13304 -13800 13338 -13632
rect 13412 -13800 13446 -13632
rect 13940 -13800 13974 -13632
rect 12776 -14926 12810 -14158
rect 13304 -14926 13338 -14158
rect 13412 -14926 13446 -14158
rect 13940 -14926 13974 -14158
rect 14376 -13800 14410 -13632
rect 14904 -13800 14938 -13632
rect 15012 -13800 15046 -13632
rect 15540 -13800 15574 -13632
rect 14376 -14926 14410 -14158
rect 14904 -14926 14938 -14158
rect 15012 -14926 15046 -14158
rect 15540 -14926 15574 -14158
rect 15976 -13800 16010 -13632
rect 16504 -13800 16538 -13632
rect 16612 -13800 16646 -13632
rect 17140 -13800 17174 -13632
rect 15976 -14926 16010 -14158
rect 16504 -14926 16538 -14158
rect 16612 -14926 16646 -14158
rect 17140 -14926 17174 -14158
rect 17576 -13800 17610 -13632
rect 18104 -13800 18138 -13632
rect 18212 -13800 18246 -13632
rect 18740 -13800 18774 -13632
rect 17576 -14926 17610 -14158
rect 18104 -14926 18138 -14158
rect 18212 -14926 18246 -14158
rect 18740 -14926 18774 -14158
rect 19176 -13800 19210 -13632
rect 19704 -13800 19738 -13632
rect 19812 -13800 19846 -13632
rect 20340 -13800 20374 -13632
rect 19176 -14926 19210 -14158
rect 19704 -14926 19738 -14158
rect 19812 -14926 19846 -14158
rect 20340 -14926 20374 -14158
rect 20776 -13800 20810 -13632
rect 21304 -13800 21338 -13632
rect 21412 -13800 21446 -13632
rect 21940 -13800 21974 -13632
rect 20776 -14926 20810 -14158
rect 21304 -14926 21338 -14158
rect 21412 -14926 21446 -14158
rect 21940 -14926 21974 -14158
rect 22376 -13800 22410 -13632
rect 22904 -13800 22938 -13632
rect 23012 -13800 23046 -13632
rect 23540 -13800 23574 -13632
rect 22376 -14926 22410 -14158
rect 22904 -14926 22938 -14158
rect 23012 -14926 23046 -14158
rect 23540 -14926 23574 -14158
rect 23976 -13800 24010 -13632
rect 24504 -13800 24538 -13632
rect 24612 -13800 24646 -13632
rect 25140 -13800 25174 -13632
rect 23976 -14926 24010 -14158
rect 24504 -14926 24538 -14158
rect 24612 -14926 24646 -14158
rect 25140 -14926 25174 -14158
rect 25576 -13800 25610 -13632
rect 26104 -13800 26138 -13632
rect 26212 -13800 26246 -13632
rect 26740 -13800 26774 -13632
rect 25576 -14926 25610 -14158
rect 26104 -14926 26138 -14158
rect 26212 -14926 26246 -14158
rect 26740 -14926 26774 -14158
rect 27176 -13800 27210 -13632
rect 27704 -13800 27738 -13632
rect 27812 -13800 27846 -13632
rect 28340 -13800 28374 -13632
rect 27176 -14926 27210 -14158
rect 27704 -14926 27738 -14158
rect 27812 -14926 27846 -14158
rect 28340 -14926 28374 -14158
rect 28776 -13800 28810 -13632
rect 29304 -13800 29338 -13632
rect 29412 -13800 29446 -13632
rect 29940 -13800 29974 -13632
rect 28776 -14926 28810 -14158
rect 29304 -14926 29338 -14158
rect 29412 -14926 29446 -14158
rect 29940 -14926 29974 -14158
rect 30376 -13800 30410 -13632
rect 30904 -13800 30938 -13632
rect 31012 -13800 31046 -13632
rect 31540 -13800 31574 -13632
rect 30376 -14926 30410 -14158
rect 30904 -14926 30938 -14158
rect 31012 -14926 31046 -14158
rect 31540 -14926 31574 -14158
rect 31976 -13800 32010 -13632
rect 32504 -13800 32538 -13632
rect 32612 -13800 32646 -13632
rect 33140 -13800 33174 -13632
rect 31976 -14926 32010 -14158
rect 32504 -14926 32538 -14158
rect 32612 -14926 32646 -14158
rect 33140 -14926 33174 -14158
rect 33576 -13800 33610 -13632
rect 34104 -13800 34138 -13632
rect 34212 -13800 34246 -13632
rect 34740 -13800 34774 -13632
rect 33576 -14926 33610 -14158
rect 34104 -14926 34138 -14158
rect 34212 -14926 34246 -14158
rect 34740 -14926 34774 -14158
rect 35176 -13800 35210 -13632
rect 35704 -13800 35738 -13632
rect 35812 -13800 35846 -13632
rect 36340 -13800 36374 -13632
rect 35176 -14926 35210 -14158
rect 35704 -14926 35738 -14158
rect 35812 -14926 35846 -14158
rect 36340 -14926 36374 -14158
rect 36776 -13800 36810 -13632
rect 37304 -13800 37338 -13632
rect 37412 -13800 37446 -13632
rect 37940 -13800 37974 -13632
rect 36776 -14926 36810 -14158
rect 37304 -14926 37338 -14158
rect 37412 -14926 37446 -14158
rect 37940 -14926 37974 -14158
rect -24 -15600 10 -15432
rect 504 -15600 538 -15432
rect 612 -15600 646 -15432
rect 1140 -15600 1174 -15432
rect -24 -16726 10 -15958
rect 504 -16726 538 -15958
rect 612 -16726 646 -15958
rect 1140 -16726 1174 -15958
rect 1576 -15600 1610 -15432
rect 2104 -15600 2138 -15432
rect 2212 -15600 2246 -15432
rect 2740 -15600 2774 -15432
rect 1576 -16726 1610 -15958
rect 2104 -16726 2138 -15958
rect 2212 -16726 2246 -15958
rect 2740 -16726 2774 -15958
rect 3176 -15600 3210 -15432
rect 3704 -15600 3738 -15432
rect 3812 -15600 3846 -15432
rect 4340 -15600 4374 -15432
rect 3176 -16726 3210 -15958
rect 3704 -16726 3738 -15958
rect 3812 -16726 3846 -15958
rect 4340 -16726 4374 -15958
rect 4776 -15600 4810 -15432
rect 5304 -15600 5338 -15432
rect 5412 -15600 5446 -15432
rect 5940 -15600 5974 -15432
rect 4776 -16726 4810 -15958
rect 5304 -16726 5338 -15958
rect 5412 -16726 5446 -15958
rect 5940 -16726 5974 -15958
rect 6376 -15600 6410 -15432
rect 6904 -15600 6938 -15432
rect 7012 -15600 7046 -15432
rect 7540 -15600 7574 -15432
rect 6376 -16726 6410 -15958
rect 6904 -16726 6938 -15958
rect 7012 -16726 7046 -15958
rect 7540 -16726 7574 -15958
rect 7976 -15600 8010 -15432
rect 8504 -15600 8538 -15432
rect 8612 -15600 8646 -15432
rect 9140 -15600 9174 -15432
rect 7976 -16726 8010 -15958
rect 8504 -16726 8538 -15958
rect 8612 -16726 8646 -15958
rect 9140 -16726 9174 -15958
rect 9576 -15600 9610 -15432
rect 10104 -15600 10138 -15432
rect 10212 -15600 10246 -15432
rect 10740 -15600 10774 -15432
rect 9576 -16726 9610 -15958
rect 10104 -16726 10138 -15958
rect 10212 -16726 10246 -15958
rect 10740 -16726 10774 -15958
rect 11176 -15600 11210 -15432
rect 11704 -15600 11738 -15432
rect 11812 -15600 11846 -15432
rect 12340 -15600 12374 -15432
rect 11176 -16726 11210 -15958
rect 11704 -16726 11738 -15958
rect 11812 -16726 11846 -15958
rect 12340 -16726 12374 -15958
rect 12776 -15600 12810 -15432
rect 13304 -15600 13338 -15432
rect 13412 -15600 13446 -15432
rect 13940 -15600 13974 -15432
rect 12776 -16726 12810 -15958
rect 13304 -16726 13338 -15958
rect 13412 -16726 13446 -15958
rect 13940 -16726 13974 -15958
rect 14376 -15600 14410 -15432
rect 14904 -15600 14938 -15432
rect 15012 -15600 15046 -15432
rect 15540 -15600 15574 -15432
rect 14376 -16726 14410 -15958
rect 14904 -16726 14938 -15958
rect 15012 -16726 15046 -15958
rect 15540 -16726 15574 -15958
rect 15976 -15600 16010 -15432
rect 16504 -15600 16538 -15432
rect 16612 -15600 16646 -15432
rect 17140 -15600 17174 -15432
rect 15976 -16726 16010 -15958
rect 16504 -16726 16538 -15958
rect 16612 -16726 16646 -15958
rect 17140 -16726 17174 -15958
rect 17576 -15600 17610 -15432
rect 18104 -15600 18138 -15432
rect 18212 -15600 18246 -15432
rect 18740 -15600 18774 -15432
rect 17576 -16726 17610 -15958
rect 18104 -16726 18138 -15958
rect 18212 -16726 18246 -15958
rect 18740 -16726 18774 -15958
rect 19176 -15600 19210 -15432
rect 19704 -15600 19738 -15432
rect 19812 -15600 19846 -15432
rect 20340 -15600 20374 -15432
rect 19176 -16726 19210 -15958
rect 19704 -16726 19738 -15958
rect 19812 -16726 19846 -15958
rect 20340 -16726 20374 -15958
rect 20776 -15600 20810 -15432
rect 21304 -15600 21338 -15432
rect 21412 -15600 21446 -15432
rect 21940 -15600 21974 -15432
rect 20776 -16726 20810 -15958
rect 21304 -16726 21338 -15958
rect 21412 -16726 21446 -15958
rect 21940 -16726 21974 -15958
rect 22376 -15600 22410 -15432
rect 22904 -15600 22938 -15432
rect 23012 -15600 23046 -15432
rect 23540 -15600 23574 -15432
rect 22376 -16726 22410 -15958
rect 22904 -16726 22938 -15958
rect 23012 -16726 23046 -15958
rect 23540 -16726 23574 -15958
rect 23976 -15600 24010 -15432
rect 24504 -15600 24538 -15432
rect 24612 -15600 24646 -15432
rect 25140 -15600 25174 -15432
rect 23976 -16726 24010 -15958
rect 24504 -16726 24538 -15958
rect 24612 -16726 24646 -15958
rect 25140 -16726 25174 -15958
rect 25576 -15600 25610 -15432
rect 26104 -15600 26138 -15432
rect 26212 -15600 26246 -15432
rect 26740 -15600 26774 -15432
rect 25576 -16726 25610 -15958
rect 26104 -16726 26138 -15958
rect 26212 -16726 26246 -15958
rect 26740 -16726 26774 -15958
rect 27176 -15600 27210 -15432
rect 27704 -15600 27738 -15432
rect 27812 -15600 27846 -15432
rect 28340 -15600 28374 -15432
rect 27176 -16726 27210 -15958
rect 27704 -16726 27738 -15958
rect 27812 -16726 27846 -15958
rect 28340 -16726 28374 -15958
rect 28776 -15600 28810 -15432
rect 29304 -15600 29338 -15432
rect 29412 -15600 29446 -15432
rect 29940 -15600 29974 -15432
rect 28776 -16726 28810 -15958
rect 29304 -16726 29338 -15958
rect 29412 -16726 29446 -15958
rect 29940 -16726 29974 -15958
rect 30376 -15600 30410 -15432
rect 30904 -15600 30938 -15432
rect 31012 -15600 31046 -15432
rect 31540 -15600 31574 -15432
rect 30376 -16726 30410 -15958
rect 30904 -16726 30938 -15958
rect 31012 -16726 31046 -15958
rect 31540 -16726 31574 -15958
rect 31976 -15600 32010 -15432
rect 32504 -15600 32538 -15432
rect 32612 -15600 32646 -15432
rect 33140 -15600 33174 -15432
rect 31976 -16726 32010 -15958
rect 32504 -16726 32538 -15958
rect 32612 -16726 32646 -15958
rect 33140 -16726 33174 -15958
rect 33576 -15600 33610 -15432
rect 34104 -15600 34138 -15432
rect 34212 -15600 34246 -15432
rect 34740 -15600 34774 -15432
rect 33576 -16726 33610 -15958
rect 34104 -16726 34138 -15958
rect 34212 -16726 34246 -15958
rect 34740 -16726 34774 -15958
rect 35176 -15600 35210 -15432
rect 35704 -15600 35738 -15432
rect 35812 -15600 35846 -15432
rect 36340 -15600 36374 -15432
rect 35176 -16726 35210 -15958
rect 35704 -16726 35738 -15958
rect 35812 -16726 35846 -15958
rect 36340 -16726 36374 -15958
rect 36776 -15600 36810 -15432
rect 37304 -15600 37338 -15432
rect 37412 -15600 37446 -15432
rect 37940 -15600 37974 -15432
rect 36776 -16726 36810 -15958
rect 37304 -16726 37338 -15958
rect 37412 -16726 37446 -15958
rect 37940 -16726 37974 -15958
rect -24 -17400 10 -17232
rect 504 -17400 538 -17232
rect 612 -17400 646 -17232
rect 1140 -17400 1174 -17232
rect -24 -18526 10 -17758
rect 504 -18526 538 -17758
rect 612 -18526 646 -17758
rect 1140 -18526 1174 -17758
rect 1576 -17400 1610 -17232
rect 2104 -17400 2138 -17232
rect 2212 -17400 2246 -17232
rect 2740 -17400 2774 -17232
rect 1576 -18526 1610 -17758
rect 2104 -18526 2138 -17758
rect 2212 -18526 2246 -17758
rect 2740 -18526 2774 -17758
rect 3176 -17400 3210 -17232
rect 3704 -17400 3738 -17232
rect 3812 -17400 3846 -17232
rect 4340 -17400 4374 -17232
rect 3176 -18526 3210 -17758
rect 3704 -18526 3738 -17758
rect 3812 -18526 3846 -17758
rect 4340 -18526 4374 -17758
rect 4776 -17400 4810 -17232
rect 5304 -17400 5338 -17232
rect 5412 -17400 5446 -17232
rect 5940 -17400 5974 -17232
rect 4776 -18526 4810 -17758
rect 5304 -18526 5338 -17758
rect 5412 -18526 5446 -17758
rect 5940 -18526 5974 -17758
rect 6376 -17400 6410 -17232
rect 6904 -17400 6938 -17232
rect 7012 -17400 7046 -17232
rect 7540 -17400 7574 -17232
rect 6376 -18526 6410 -17758
rect 6904 -18526 6938 -17758
rect 7012 -18526 7046 -17758
rect 7540 -18526 7574 -17758
rect 7976 -17400 8010 -17232
rect 8504 -17400 8538 -17232
rect 8612 -17400 8646 -17232
rect 9140 -17400 9174 -17232
rect 7976 -18526 8010 -17758
rect 8504 -18526 8538 -17758
rect 8612 -18526 8646 -17758
rect 9140 -18526 9174 -17758
rect 9576 -17400 9610 -17232
rect 10104 -17400 10138 -17232
rect 10212 -17400 10246 -17232
rect 10740 -17400 10774 -17232
rect 9576 -18526 9610 -17758
rect 10104 -18526 10138 -17758
rect 10212 -18526 10246 -17758
rect 10740 -18526 10774 -17758
rect 11176 -17400 11210 -17232
rect 11704 -17400 11738 -17232
rect 11812 -17400 11846 -17232
rect 12340 -17400 12374 -17232
rect 11176 -18526 11210 -17758
rect 11704 -18526 11738 -17758
rect 11812 -18526 11846 -17758
rect 12340 -18526 12374 -17758
rect 12776 -17400 12810 -17232
rect 13304 -17400 13338 -17232
rect 13412 -17400 13446 -17232
rect 13940 -17400 13974 -17232
rect 12776 -18526 12810 -17758
rect 13304 -18526 13338 -17758
rect 13412 -18526 13446 -17758
rect 13940 -18526 13974 -17758
rect 14376 -17400 14410 -17232
rect 14904 -17400 14938 -17232
rect 15012 -17400 15046 -17232
rect 15540 -17400 15574 -17232
rect 14376 -18526 14410 -17758
rect 14904 -18526 14938 -17758
rect 15012 -18526 15046 -17758
rect 15540 -18526 15574 -17758
rect 15976 -17400 16010 -17232
rect 16504 -17400 16538 -17232
rect 16612 -17400 16646 -17232
rect 17140 -17400 17174 -17232
rect 15976 -18526 16010 -17758
rect 16504 -18526 16538 -17758
rect 16612 -18526 16646 -17758
rect 17140 -18526 17174 -17758
rect 17576 -17400 17610 -17232
rect 18104 -17400 18138 -17232
rect 18212 -17400 18246 -17232
rect 18740 -17400 18774 -17232
rect 17576 -18526 17610 -17758
rect 18104 -18526 18138 -17758
rect 18212 -18526 18246 -17758
rect 18740 -18526 18774 -17758
rect 19176 -17400 19210 -17232
rect 19704 -17400 19738 -17232
rect 19812 -17400 19846 -17232
rect 20340 -17400 20374 -17232
rect 19176 -18526 19210 -17758
rect 19704 -18526 19738 -17758
rect 19812 -18526 19846 -17758
rect 20340 -18526 20374 -17758
rect 20776 -17400 20810 -17232
rect 21304 -17400 21338 -17232
rect 21412 -17400 21446 -17232
rect 21940 -17400 21974 -17232
rect 20776 -18526 20810 -17758
rect 21304 -18526 21338 -17758
rect 21412 -18526 21446 -17758
rect 21940 -18526 21974 -17758
rect 22376 -17400 22410 -17232
rect 22904 -17400 22938 -17232
rect 23012 -17400 23046 -17232
rect 23540 -17400 23574 -17232
rect 22376 -18526 22410 -17758
rect 22904 -18526 22938 -17758
rect 23012 -18526 23046 -17758
rect 23540 -18526 23574 -17758
rect 23976 -17400 24010 -17232
rect 24504 -17400 24538 -17232
rect 24612 -17400 24646 -17232
rect 25140 -17400 25174 -17232
rect 23976 -18526 24010 -17758
rect 24504 -18526 24538 -17758
rect 24612 -18526 24646 -17758
rect 25140 -18526 25174 -17758
rect 25576 -17400 25610 -17232
rect 26104 -17400 26138 -17232
rect 26212 -17400 26246 -17232
rect 26740 -17400 26774 -17232
rect 25576 -18526 25610 -17758
rect 26104 -18526 26138 -17758
rect 26212 -18526 26246 -17758
rect 26740 -18526 26774 -17758
rect 27176 -17400 27210 -17232
rect 27704 -17400 27738 -17232
rect 27812 -17400 27846 -17232
rect 28340 -17400 28374 -17232
rect 27176 -18526 27210 -17758
rect 27704 -18526 27738 -17758
rect 27812 -18526 27846 -17758
rect 28340 -18526 28374 -17758
rect 28776 -17400 28810 -17232
rect 29304 -17400 29338 -17232
rect 29412 -17400 29446 -17232
rect 29940 -17400 29974 -17232
rect 28776 -18526 28810 -17758
rect 29304 -18526 29338 -17758
rect 29412 -18526 29446 -17758
rect 29940 -18526 29974 -17758
rect 30376 -17400 30410 -17232
rect 30904 -17400 30938 -17232
rect 31012 -17400 31046 -17232
rect 31540 -17400 31574 -17232
rect 30376 -18526 30410 -17758
rect 30904 -18526 30938 -17758
rect 31012 -18526 31046 -17758
rect 31540 -18526 31574 -17758
rect 31976 -17400 32010 -17232
rect 32504 -17400 32538 -17232
rect 32612 -17400 32646 -17232
rect 33140 -17400 33174 -17232
rect 31976 -18526 32010 -17758
rect 32504 -18526 32538 -17758
rect 32612 -18526 32646 -17758
rect 33140 -18526 33174 -17758
rect 33576 -17400 33610 -17232
rect 34104 -17400 34138 -17232
rect 34212 -17400 34246 -17232
rect 34740 -17400 34774 -17232
rect 33576 -18526 33610 -17758
rect 34104 -18526 34138 -17758
rect 34212 -18526 34246 -17758
rect 34740 -18526 34774 -17758
rect 35176 -17400 35210 -17232
rect 35704 -17400 35738 -17232
rect 35812 -17400 35846 -17232
rect 36340 -17400 36374 -17232
rect 35176 -18526 35210 -17758
rect 35704 -18526 35738 -17758
rect 35812 -18526 35846 -17758
rect 36340 -18526 36374 -17758
rect 36776 -17400 36810 -17232
rect 37304 -17400 37338 -17232
rect 37412 -17400 37446 -17232
rect 37940 -17400 37974 -17232
rect 36776 -18526 36810 -17758
rect 37304 -18526 37338 -17758
rect 37412 -18526 37446 -17758
rect 37940 -18526 37974 -17758
rect -24 -19200 10 -19032
rect 504 -19200 538 -19032
rect 612 -19200 646 -19032
rect 1140 -19200 1174 -19032
rect -24 -20326 10 -19558
rect 504 -20326 538 -19558
rect 612 -20326 646 -19558
rect 1140 -20326 1174 -19558
rect 1576 -19200 1610 -19032
rect 2104 -19200 2138 -19032
rect 2212 -19200 2246 -19032
rect 2740 -19200 2774 -19032
rect 1576 -20326 1610 -19558
rect 2104 -20326 2138 -19558
rect 2212 -20326 2246 -19558
rect 2740 -20326 2774 -19558
rect 3176 -19200 3210 -19032
rect 3704 -19200 3738 -19032
rect 3812 -19200 3846 -19032
rect 4340 -19200 4374 -19032
rect 3176 -20326 3210 -19558
rect 3704 -20326 3738 -19558
rect 3812 -20326 3846 -19558
rect 4340 -20326 4374 -19558
rect 4776 -19200 4810 -19032
rect 5304 -19200 5338 -19032
rect 5412 -19200 5446 -19032
rect 5940 -19200 5974 -19032
rect 4776 -20326 4810 -19558
rect 5304 -20326 5338 -19558
rect 5412 -20326 5446 -19558
rect 5940 -20326 5974 -19558
rect 6376 -19200 6410 -19032
rect 6904 -19200 6938 -19032
rect 7012 -19200 7046 -19032
rect 7540 -19200 7574 -19032
rect 6376 -20326 6410 -19558
rect 6904 -20326 6938 -19558
rect 7012 -20326 7046 -19558
rect 7540 -20326 7574 -19558
rect 7976 -19200 8010 -19032
rect 8504 -19200 8538 -19032
rect 8612 -19200 8646 -19032
rect 9140 -19200 9174 -19032
rect 7976 -20326 8010 -19558
rect 8504 -20326 8538 -19558
rect 8612 -20326 8646 -19558
rect 9140 -20326 9174 -19558
rect 9576 -19200 9610 -19032
rect 10104 -19200 10138 -19032
rect 10212 -19200 10246 -19032
rect 10740 -19200 10774 -19032
rect 9576 -20326 9610 -19558
rect 10104 -20326 10138 -19558
rect 10212 -20326 10246 -19558
rect 10740 -20326 10774 -19558
rect 11176 -19200 11210 -19032
rect 11704 -19200 11738 -19032
rect 11812 -19200 11846 -19032
rect 12340 -19200 12374 -19032
rect 11176 -20326 11210 -19558
rect 11704 -20326 11738 -19558
rect 11812 -20326 11846 -19558
rect 12340 -20326 12374 -19558
rect 12776 -19200 12810 -19032
rect 13304 -19200 13338 -19032
rect 13412 -19200 13446 -19032
rect 13940 -19200 13974 -19032
rect 12776 -20326 12810 -19558
rect 13304 -20326 13338 -19558
rect 13412 -20326 13446 -19558
rect 13940 -20326 13974 -19558
rect 14376 -19200 14410 -19032
rect 14904 -19200 14938 -19032
rect 15012 -19200 15046 -19032
rect 15540 -19200 15574 -19032
rect 14376 -20326 14410 -19558
rect 14904 -20326 14938 -19558
rect 15012 -20326 15046 -19558
rect 15540 -20326 15574 -19558
rect 15976 -19200 16010 -19032
rect 16504 -19200 16538 -19032
rect 16612 -19200 16646 -19032
rect 17140 -19200 17174 -19032
rect 15976 -20326 16010 -19558
rect 16504 -20326 16538 -19558
rect 16612 -20326 16646 -19558
rect 17140 -20326 17174 -19558
rect 17576 -19200 17610 -19032
rect 18104 -19200 18138 -19032
rect 18212 -19200 18246 -19032
rect 18740 -19200 18774 -19032
rect 17576 -20326 17610 -19558
rect 18104 -20326 18138 -19558
rect 18212 -20326 18246 -19558
rect 18740 -20326 18774 -19558
rect 19176 -19200 19210 -19032
rect 19704 -19200 19738 -19032
rect 19812 -19200 19846 -19032
rect 20340 -19200 20374 -19032
rect 19176 -20326 19210 -19558
rect 19704 -20326 19738 -19558
rect 19812 -20326 19846 -19558
rect 20340 -20326 20374 -19558
rect 20776 -19200 20810 -19032
rect 21304 -19200 21338 -19032
rect 21412 -19200 21446 -19032
rect 21940 -19200 21974 -19032
rect 20776 -20326 20810 -19558
rect 21304 -20326 21338 -19558
rect 21412 -20326 21446 -19558
rect 21940 -20326 21974 -19558
rect 22376 -19200 22410 -19032
rect 22904 -19200 22938 -19032
rect 23012 -19200 23046 -19032
rect 23540 -19200 23574 -19032
rect 22376 -20326 22410 -19558
rect 22904 -20326 22938 -19558
rect 23012 -20326 23046 -19558
rect 23540 -20326 23574 -19558
rect 23976 -19200 24010 -19032
rect 24504 -19200 24538 -19032
rect 24612 -19200 24646 -19032
rect 25140 -19200 25174 -19032
rect 23976 -20326 24010 -19558
rect 24504 -20326 24538 -19558
rect 24612 -20326 24646 -19558
rect 25140 -20326 25174 -19558
rect 25576 -19200 25610 -19032
rect 26104 -19200 26138 -19032
rect 26212 -19200 26246 -19032
rect 26740 -19200 26774 -19032
rect 25576 -20326 25610 -19558
rect 26104 -20326 26138 -19558
rect 26212 -20326 26246 -19558
rect 26740 -20326 26774 -19558
rect 27176 -19200 27210 -19032
rect 27704 -19200 27738 -19032
rect 27812 -19200 27846 -19032
rect 28340 -19200 28374 -19032
rect 27176 -20326 27210 -19558
rect 27704 -20326 27738 -19558
rect 27812 -20326 27846 -19558
rect 28340 -20326 28374 -19558
rect 28776 -19200 28810 -19032
rect 29304 -19200 29338 -19032
rect 29412 -19200 29446 -19032
rect 29940 -19200 29974 -19032
rect 28776 -20326 28810 -19558
rect 29304 -20326 29338 -19558
rect 29412 -20326 29446 -19558
rect 29940 -20326 29974 -19558
rect 30376 -19200 30410 -19032
rect 30904 -19200 30938 -19032
rect 31012 -19200 31046 -19032
rect 31540 -19200 31574 -19032
rect 30376 -20326 30410 -19558
rect 30904 -20326 30938 -19558
rect 31012 -20326 31046 -19558
rect 31540 -20326 31574 -19558
rect 31976 -19200 32010 -19032
rect 32504 -19200 32538 -19032
rect 32612 -19200 32646 -19032
rect 33140 -19200 33174 -19032
rect 31976 -20326 32010 -19558
rect 32504 -20326 32538 -19558
rect 32612 -20326 32646 -19558
rect 33140 -20326 33174 -19558
rect 33576 -19200 33610 -19032
rect 34104 -19200 34138 -19032
rect 34212 -19200 34246 -19032
rect 34740 -19200 34774 -19032
rect 33576 -20326 33610 -19558
rect 34104 -20326 34138 -19558
rect 34212 -20326 34246 -19558
rect 34740 -20326 34774 -19558
rect 35176 -19200 35210 -19032
rect 35704 -19200 35738 -19032
rect 35812 -19200 35846 -19032
rect 36340 -19200 36374 -19032
rect 35176 -20326 35210 -19558
rect 35704 -20326 35738 -19558
rect 35812 -20326 35846 -19558
rect 36340 -20326 36374 -19558
rect 36776 -19200 36810 -19032
rect 37304 -19200 37338 -19032
rect 37412 -19200 37446 -19032
rect 37940 -19200 37974 -19032
rect 36776 -20326 36810 -19558
rect 37304 -20326 37338 -19558
rect 37412 -20326 37446 -19558
rect 37940 -20326 37974 -19558
rect -24 -21000 10 -20832
rect 504 -21000 538 -20832
rect 612 -21000 646 -20832
rect 1140 -21000 1174 -20832
rect -24 -22126 10 -21358
rect 504 -22126 538 -21358
rect 612 -22126 646 -21358
rect 1140 -22126 1174 -21358
rect 1576 -21000 1610 -20832
rect 2104 -21000 2138 -20832
rect 2212 -21000 2246 -20832
rect 2740 -21000 2774 -20832
rect 1576 -22126 1610 -21358
rect 2104 -22126 2138 -21358
rect 2212 -22126 2246 -21358
rect 2740 -22126 2774 -21358
rect 3176 -21000 3210 -20832
rect 3704 -21000 3738 -20832
rect 3812 -21000 3846 -20832
rect 4340 -21000 4374 -20832
rect 3176 -22126 3210 -21358
rect 3704 -22126 3738 -21358
rect 3812 -22126 3846 -21358
rect 4340 -22126 4374 -21358
rect 4776 -21000 4810 -20832
rect 5304 -21000 5338 -20832
rect 5412 -21000 5446 -20832
rect 5940 -21000 5974 -20832
rect 4776 -22126 4810 -21358
rect 5304 -22126 5338 -21358
rect 5412 -22126 5446 -21358
rect 5940 -22126 5974 -21358
rect 6376 -21000 6410 -20832
rect 6904 -21000 6938 -20832
rect 7012 -21000 7046 -20832
rect 7540 -21000 7574 -20832
rect 6376 -22126 6410 -21358
rect 6904 -22126 6938 -21358
rect 7012 -22126 7046 -21358
rect 7540 -22126 7574 -21358
rect 7976 -21000 8010 -20832
rect 8504 -21000 8538 -20832
rect 8612 -21000 8646 -20832
rect 9140 -21000 9174 -20832
rect 7976 -22126 8010 -21358
rect 8504 -22126 8538 -21358
rect 8612 -22126 8646 -21358
rect 9140 -22126 9174 -21358
rect 9576 -21000 9610 -20832
rect 10104 -21000 10138 -20832
rect 10212 -21000 10246 -20832
rect 10740 -21000 10774 -20832
rect 9576 -22126 9610 -21358
rect 10104 -22126 10138 -21358
rect 10212 -22126 10246 -21358
rect 10740 -22126 10774 -21358
rect 11176 -21000 11210 -20832
rect 11704 -21000 11738 -20832
rect 11812 -21000 11846 -20832
rect 12340 -21000 12374 -20832
rect 11176 -22126 11210 -21358
rect 11704 -22126 11738 -21358
rect 11812 -22126 11846 -21358
rect 12340 -22126 12374 -21358
rect 12776 -21000 12810 -20832
rect 13304 -21000 13338 -20832
rect 13412 -21000 13446 -20832
rect 13940 -21000 13974 -20832
rect 12776 -22126 12810 -21358
rect 13304 -22126 13338 -21358
rect 13412 -22126 13446 -21358
rect 13940 -22126 13974 -21358
rect 14376 -21000 14410 -20832
rect 14904 -21000 14938 -20832
rect 15012 -21000 15046 -20832
rect 15540 -21000 15574 -20832
rect 14376 -22126 14410 -21358
rect 14904 -22126 14938 -21358
rect 15012 -22126 15046 -21358
rect 15540 -22126 15574 -21358
rect 15976 -21000 16010 -20832
rect 16504 -21000 16538 -20832
rect 16612 -21000 16646 -20832
rect 17140 -21000 17174 -20832
rect 15976 -22126 16010 -21358
rect 16504 -22126 16538 -21358
rect 16612 -22126 16646 -21358
rect 17140 -22126 17174 -21358
rect 17576 -21000 17610 -20832
rect 18104 -21000 18138 -20832
rect 18212 -21000 18246 -20832
rect 18740 -21000 18774 -20832
rect 17576 -22126 17610 -21358
rect 18104 -22126 18138 -21358
rect 18212 -22126 18246 -21358
rect 18740 -22126 18774 -21358
rect 19176 -21000 19210 -20832
rect 19704 -21000 19738 -20832
rect 19812 -21000 19846 -20832
rect 20340 -21000 20374 -20832
rect 19176 -22126 19210 -21358
rect 19704 -22126 19738 -21358
rect 19812 -22126 19846 -21358
rect 20340 -22126 20374 -21358
rect 20776 -21000 20810 -20832
rect 21304 -21000 21338 -20832
rect 21412 -21000 21446 -20832
rect 21940 -21000 21974 -20832
rect 20776 -22126 20810 -21358
rect 21304 -22126 21338 -21358
rect 21412 -22126 21446 -21358
rect 21940 -22126 21974 -21358
rect 22376 -21000 22410 -20832
rect 22904 -21000 22938 -20832
rect 23012 -21000 23046 -20832
rect 23540 -21000 23574 -20832
rect 22376 -22126 22410 -21358
rect 22904 -22126 22938 -21358
rect 23012 -22126 23046 -21358
rect 23540 -22126 23574 -21358
rect 23976 -21000 24010 -20832
rect 24504 -21000 24538 -20832
rect 24612 -21000 24646 -20832
rect 25140 -21000 25174 -20832
rect 23976 -22126 24010 -21358
rect 24504 -22126 24538 -21358
rect 24612 -22126 24646 -21358
rect 25140 -22126 25174 -21358
rect 25576 -21000 25610 -20832
rect 26104 -21000 26138 -20832
rect 26212 -21000 26246 -20832
rect 26740 -21000 26774 -20832
rect 25576 -22126 25610 -21358
rect 26104 -22126 26138 -21358
rect 26212 -22126 26246 -21358
rect 26740 -22126 26774 -21358
rect 27176 -21000 27210 -20832
rect 27704 -21000 27738 -20832
rect 27812 -21000 27846 -20832
rect 28340 -21000 28374 -20832
rect 27176 -22126 27210 -21358
rect 27704 -22126 27738 -21358
rect 27812 -22126 27846 -21358
rect 28340 -22126 28374 -21358
rect 28776 -21000 28810 -20832
rect 29304 -21000 29338 -20832
rect 29412 -21000 29446 -20832
rect 29940 -21000 29974 -20832
rect 28776 -22126 28810 -21358
rect 29304 -22126 29338 -21358
rect 29412 -22126 29446 -21358
rect 29940 -22126 29974 -21358
rect 30376 -21000 30410 -20832
rect 30904 -21000 30938 -20832
rect 31012 -21000 31046 -20832
rect 31540 -21000 31574 -20832
rect 30376 -22126 30410 -21358
rect 30904 -22126 30938 -21358
rect 31012 -22126 31046 -21358
rect 31540 -22126 31574 -21358
rect 31976 -21000 32010 -20832
rect 32504 -21000 32538 -20832
rect 32612 -21000 32646 -20832
rect 33140 -21000 33174 -20832
rect 31976 -22126 32010 -21358
rect 32504 -22126 32538 -21358
rect 32612 -22126 32646 -21358
rect 33140 -22126 33174 -21358
rect 33576 -21000 33610 -20832
rect 34104 -21000 34138 -20832
rect 34212 -21000 34246 -20832
rect 34740 -21000 34774 -20832
rect 33576 -22126 33610 -21358
rect 34104 -22126 34138 -21358
rect 34212 -22126 34246 -21358
rect 34740 -22126 34774 -21358
rect 35176 -21000 35210 -20832
rect 35704 -21000 35738 -20832
rect 35812 -21000 35846 -20832
rect 36340 -21000 36374 -20832
rect 35176 -22126 35210 -21358
rect 35704 -22126 35738 -21358
rect 35812 -22126 35846 -21358
rect 36340 -22126 36374 -21358
rect 36776 -21000 36810 -20832
rect 37304 -21000 37338 -20832
rect 37412 -21000 37446 -20832
rect 37940 -21000 37974 -20832
rect 36776 -22126 36810 -21358
rect 37304 -22126 37338 -21358
rect 37412 -22126 37446 -21358
rect 37940 -22126 37974 -21358
rect 28414 -23553 28482 -23519
rect 28572 -23553 28640 -23519
rect 28730 -23553 28798 -23519
rect 28888 -23553 28956 -23519
rect 32694 -22576 32762 -22542
rect 32852 -22576 32920 -22542
rect 33010 -22576 33078 -22542
rect 33168 -22576 33236 -22542
rect 32694 -23104 32762 -23070
rect 32852 -23104 32920 -23070
rect 33010 -23104 33078 -23070
rect 33168 -23104 33236 -23070
rect 34064 -22596 34132 -22562
rect 34222 -22596 34290 -22562
rect 34064 -23124 34132 -23090
rect 34222 -23124 34290 -23090
rect 186 -24636 220 -24368
rect 1914 -24636 1948 -24368
rect 2386 -24636 2420 -24368
rect 4114 -24636 4148 -24368
rect 4586 -24636 4620 -24368
rect 6314 -24636 6348 -24368
rect 6786 -24636 6820 -24368
rect 8514 -24636 8548 -24368
rect 8986 -24636 9020 -24368
rect 10714 -24636 10748 -24368
rect 11186 -24636 11220 -24368
rect 12914 -24636 12948 -24368
rect 13386 -24636 13420 -24368
rect 15114 -24636 15148 -24368
rect 15586 -24636 15620 -24368
rect 17314 -24636 17348 -24368
rect 17786 -24636 17820 -24368
rect 19514 -24636 19548 -24368
rect 19986 -24636 20020 -24368
rect 21714 -24636 21748 -24368
rect 33232 -23718 33300 -23684
rect 33390 -23718 33458 -23684
rect 33548 -23718 33616 -23684
rect 33706 -23718 33774 -23684
rect 33864 -23718 33932 -23684
rect 34022 -23718 34090 -23684
rect 33232 -24246 33300 -24212
rect 33390 -24246 33458 -24212
rect 33548 -24246 33616 -24212
rect 33706 -24246 33774 -24212
rect 33864 -24246 33932 -24212
rect 34022 -24246 34090 -24212
rect 34604 -23716 34672 -23682
rect 34762 -23716 34830 -23682
rect 34920 -23716 34988 -23682
rect 35078 -23716 35146 -23682
rect 35236 -23716 35304 -23682
rect 35394 -23716 35462 -23682
rect 35552 -23716 35620 -23682
rect 35710 -23716 35778 -23682
rect 35868 -23716 35936 -23682
rect 36026 -23716 36094 -23682
rect 36184 -23716 36252 -23682
rect 36342 -23716 36410 -23682
rect 36500 -23716 36568 -23682
rect 36658 -23716 36726 -23682
rect 36816 -23716 36884 -23682
rect 36974 -23716 37042 -23682
rect 34604 -24244 34672 -24210
rect 34762 -24244 34830 -24210
rect 34920 -24244 34988 -24210
rect 35078 -24244 35146 -24210
rect 35236 -24244 35304 -24210
rect 35394 -24244 35462 -24210
rect 35552 -24244 35620 -24210
rect 35710 -24244 35778 -24210
rect 35868 -24244 35936 -24210
rect 36026 -24244 36094 -24210
rect 36184 -24244 36252 -24210
rect 36342 -24244 36410 -24210
rect 36500 -24244 36568 -24210
rect 36658 -24244 36726 -24210
rect 36816 -24244 36884 -24210
rect 36974 -24244 37042 -24210
rect 186 -25436 220 -25168
rect 1914 -25436 1948 -25168
rect 2386 -25436 2420 -25168
rect 4114 -25436 4148 -25168
rect 4586 -25436 4620 -25168
rect 6314 -25436 6348 -25168
rect 6786 -25436 6820 -25168
rect 8514 -25436 8548 -25168
rect 8986 -25436 9020 -25168
rect 10714 -25436 10748 -25168
rect 11186 -25436 11220 -25168
rect 12914 -25436 12948 -25168
rect 13386 -25436 13420 -25168
rect 15114 -25436 15148 -25168
rect 15586 -25436 15620 -25168
rect 17314 -25436 17348 -25168
rect 17786 -25436 17820 -25168
rect 19514 -25436 19548 -25168
rect 19986 -25436 20020 -25168
rect 21714 -25436 21748 -25168
rect 186 -26236 220 -25968
rect 1914 -26236 1948 -25968
rect 2386 -26236 2420 -25968
rect 4114 -26236 4148 -25968
rect 4586 -26236 4620 -25968
rect 6314 -26236 6348 -25968
rect 6786 -26236 6820 -25968
rect 8514 -26236 8548 -25968
rect 8986 -26236 9020 -25968
rect 10714 -26236 10748 -25968
rect 11186 -26236 11220 -25968
rect 12914 -26236 12948 -25968
rect 13386 -26236 13420 -25968
rect 15114 -26236 15148 -25968
rect 15586 -26236 15620 -25968
rect 17314 -26236 17348 -25968
rect 17786 -26236 17820 -25968
rect 19514 -26236 19548 -25968
rect 19986 -26236 20020 -25968
rect 21714 -26236 21748 -25968
rect 186 -27036 220 -26768
rect 1914 -27036 1948 -26768
rect 2386 -27036 2420 -26768
rect 4114 -27036 4148 -26768
rect 4586 -27036 4620 -26768
rect 6314 -27036 6348 -26768
rect 6786 -27036 6820 -26768
rect 8514 -27036 8548 -26768
rect 8986 -27036 9020 -26768
rect 10714 -27036 10748 -26768
rect 11186 -27036 11220 -26768
rect 12914 -27036 12948 -26768
rect 13386 -27036 13420 -26768
rect 15114 -27036 15148 -26768
rect 15586 -27036 15620 -26768
rect 17314 -27036 17348 -26768
rect 17786 -27036 17820 -26768
rect 19514 -27036 19548 -26768
rect 19986 -27036 20020 -26768
rect 21714 -27036 21748 -26768
rect 186 -27836 220 -27568
rect 1914 -27836 1948 -27568
rect 2386 -27836 2420 -27568
rect 4114 -27836 4148 -27568
rect 4586 -27836 4620 -27568
rect 6314 -27836 6348 -27568
rect 6786 -27836 6820 -27568
rect 8514 -27836 8548 -27568
rect 8986 -27836 9020 -27568
rect 10714 -27836 10748 -27568
rect 11186 -27836 11220 -27568
rect 12914 -27836 12948 -27568
rect 13386 -27836 13420 -27568
rect 15114 -27836 15148 -27568
rect 15586 -27836 15620 -27568
rect 17314 -27836 17348 -27568
rect 17786 -27836 17820 -27568
rect 19514 -27836 19548 -27568
rect 19986 -27836 20020 -27568
rect 21714 -27836 21748 -27568
rect 186 -28636 220 -28368
rect 1914 -28636 1948 -28368
rect 2386 -28636 2420 -28368
rect 4114 -28636 4148 -28368
rect 4586 -28636 4620 -28368
rect 6314 -28636 6348 -28368
rect 6786 -28636 6820 -28368
rect 8514 -28636 8548 -28368
rect 8986 -28636 9020 -28368
rect 10714 -28636 10748 -28368
rect 11186 -28636 11220 -28368
rect 12914 -28636 12948 -28368
rect 13386 -28636 13420 -28368
rect 15114 -28636 15148 -28368
rect 15586 -28636 15620 -28368
rect 17314 -28636 17348 -28368
rect 17786 -28636 17820 -28368
rect 19514 -28636 19548 -28368
rect 19986 -28636 20020 -28368
rect 21714 -28636 21748 -28368
rect 186 -29436 220 -29168
rect 1914 -29436 1948 -29168
rect 2386 -29436 2420 -29168
rect 4114 -29436 4148 -29168
rect 4586 -29436 4620 -29168
rect 6314 -29436 6348 -29168
rect 6786 -29436 6820 -29168
rect 8514 -29436 8548 -29168
rect 8986 -29436 9020 -29168
rect 10714 -29436 10748 -29168
rect 11186 -29436 11220 -29168
rect 12914 -29436 12948 -29168
rect 13386 -29436 13420 -29168
rect 15114 -29436 15148 -29168
rect 15586 -29436 15620 -29168
rect 17314 -29436 17348 -29168
rect 17786 -29436 17820 -29168
rect 19514 -29436 19548 -29168
rect 19986 -29436 20020 -29168
rect 21714 -29436 21748 -29168
rect 186 -30236 220 -29968
rect 1914 -30236 1948 -29968
rect 2386 -30236 2420 -29968
rect 4114 -30236 4148 -29968
rect 4586 -30236 4620 -29968
rect 6314 -30236 6348 -29968
rect 6786 -30236 6820 -29968
rect 8514 -30236 8548 -29968
rect 8986 -30236 9020 -29968
rect 10714 -30236 10748 -29968
rect 11186 -30236 11220 -29968
rect 12914 -30236 12948 -29968
rect 13386 -30236 13420 -29968
rect 15114 -30236 15148 -29968
rect 15586 -30236 15620 -29968
rect 17314 -30236 17348 -29968
rect 17786 -30236 17820 -29968
rect 19514 -30236 19548 -29968
rect 19986 -30236 20020 -29968
rect 21714 -30236 21748 -29968
rect 186 -31036 220 -30768
rect 1914 -31036 1948 -30768
rect 2386 -31036 2420 -30768
rect 4114 -31036 4148 -30768
rect 4586 -31036 4620 -30768
rect 6314 -31036 6348 -30768
rect 6786 -31036 6820 -30768
rect 8514 -31036 8548 -30768
rect 8986 -31036 9020 -30768
rect 10714 -31036 10748 -30768
rect 11186 -31036 11220 -30768
rect 12914 -31036 12948 -30768
rect 13386 -31036 13420 -30768
rect 15114 -31036 15148 -30768
rect 15586 -31036 15620 -30768
rect 17314 -31036 17348 -30768
rect 17786 -31036 17820 -30768
rect 19514 -31036 19548 -30768
rect 19986 -31036 20020 -30768
rect 21714 -31036 21748 -30768
rect 186 -31836 220 -31568
rect 1914 -31836 1948 -31568
rect 2386 -31836 2420 -31568
rect 4114 -31836 4148 -31568
rect 4586 -31836 4620 -31568
rect 6314 -31836 6348 -31568
rect 6786 -31836 6820 -31568
rect 8514 -31836 8548 -31568
rect 8986 -31836 9020 -31568
rect 10714 -31836 10748 -31568
rect 11186 -31836 11220 -31568
rect 12914 -31836 12948 -31568
rect 13386 -31836 13420 -31568
rect 15114 -31836 15148 -31568
rect 15586 -31836 15620 -31568
rect 17314 -31836 17348 -31568
rect 17786 -31836 17820 -31568
rect 19514 -31836 19548 -31568
rect 19986 -31836 20020 -31568
rect 21714 -31836 21748 -31568
rect 27984 -24674 28752 -24640
rect 27984 -25184 28752 -25150
rect 28774 -25672 28808 -25604
rect 28774 -25830 28808 -25762
rect 28774 -25988 28808 -25920
rect 28774 -26146 28808 -26078
rect 28774 -26712 28808 -26644
rect 28774 -26870 28808 -26802
rect 28774 -27028 28808 -26960
rect 28774 -27186 28808 -27118
rect 34896 -25060 34930 -24892
rect 35824 -25060 35858 -24892
rect 34896 -25318 34930 -25150
rect 35824 -25318 35858 -25150
rect 34896 -25576 34930 -25408
rect 35824 -25576 35858 -25408
rect 34896 -25834 34930 -25666
rect 35824 -25834 35858 -25666
rect 34896 -26092 34930 -25924
rect 35824 -26092 35858 -25924
rect 34896 -26350 34930 -26182
rect 35824 -26350 35858 -26182
rect 34896 -26608 34930 -26440
rect 35824 -26608 35858 -26440
rect 34896 -26866 34930 -26698
rect 35824 -26866 35858 -26698
rect 36236 -25060 36270 -24892
rect 37164 -25060 37198 -24892
rect 36236 -25318 36270 -25150
rect 37164 -25318 37198 -25150
rect 36236 -25576 36270 -25408
rect 37164 -25576 37198 -25408
rect 36236 -25834 36270 -25666
rect 37164 -25834 37198 -25666
rect 36236 -26092 36270 -25924
rect 37164 -26092 37198 -25924
rect 36236 -26350 36270 -26182
rect 37164 -26350 37198 -26182
rect 36236 -26608 36270 -26440
rect 37164 -26608 37198 -26440
rect 36236 -26866 36270 -26698
rect 37164 -26866 37198 -26698
rect 28774 -27752 28808 -27684
rect 28774 -27910 28808 -27842
rect 28774 -28068 28808 -28000
rect 28774 -28226 28808 -28158
rect 28774 -28792 28808 -28724
rect 28774 -28950 28808 -28882
rect 28774 -29108 28808 -29040
rect 28774 -29266 28808 -29198
rect 31874 -28474 31942 -28440
rect 31874 -29002 31942 -28968
rect 32314 -28474 32382 -28440
rect 32314 -29002 32382 -28968
rect 32754 -28474 32822 -28440
rect 32754 -29002 32822 -28968
rect 33168 -28774 33536 -28740
rect 33168 -29002 33536 -28968
rect 34074 -28474 34142 -28440
rect 34074 -29002 34142 -28968
rect 34514 -28474 34582 -28440
rect 34514 -29002 34582 -28968
rect 34954 -28474 35022 -28440
rect 34954 -29002 35022 -28968
rect 35368 -28774 35736 -28740
rect 35368 -29002 35736 -28968
rect 36274 -28474 36342 -28440
rect 36274 -29002 36342 -28968
rect 36714 -28474 36782 -28440
rect 36714 -29002 36782 -28968
rect 37154 -28474 37222 -28440
rect 37154 -29002 37222 -28968
rect 37568 -28774 37936 -28740
rect 37568 -29002 37936 -28968
rect 28774 -29832 28808 -29764
rect 28774 -29990 28808 -29922
rect 28774 -30148 28808 -30080
rect 28774 -30306 28808 -30238
rect 31875 -29503 31943 -29469
rect 31875 -29813 31943 -29779
rect 32315 -29503 32383 -29469
rect 32315 -29813 32383 -29779
rect 32755 -29503 32823 -29469
rect 32755 -29813 32823 -29779
rect 33194 -29503 33262 -29469
rect 33352 -29503 33420 -29469
rect 33510 -29503 33578 -29469
rect 33194 -29813 33262 -29779
rect 33352 -29813 33420 -29779
rect 33510 -29813 33578 -29779
rect 34075 -29503 34143 -29469
rect 34075 -29813 34143 -29779
rect 34515 -29503 34583 -29469
rect 34515 -29813 34583 -29779
rect 34955 -29503 35023 -29469
rect 34955 -29813 35023 -29779
rect 35394 -29503 35462 -29469
rect 35552 -29503 35620 -29469
rect 35710 -29503 35778 -29469
rect 35394 -29813 35462 -29779
rect 35552 -29813 35620 -29779
rect 35710 -29813 35778 -29779
rect 36275 -29503 36343 -29469
rect 36275 -29813 36343 -29779
rect 36715 -29503 36783 -29469
rect 36715 -29813 36783 -29779
rect 37155 -29503 37223 -29469
rect 37155 -29813 37223 -29779
rect 37594 -29503 37662 -29469
rect 37752 -29503 37820 -29469
rect 37910 -29503 37978 -29469
rect 37594 -29813 37662 -29779
rect 37752 -29813 37820 -29779
rect 37910 -29813 37978 -29779
rect 28774 -30872 28808 -30804
rect 28774 -31030 28808 -30962
rect 28774 -31188 28808 -31120
rect 28774 -31346 28808 -31278
rect 31844 -30245 31912 -30211
rect 32002 -30245 32070 -30211
rect 32160 -30245 32228 -30211
rect 31844 -30555 31912 -30521
rect 32002 -30555 32070 -30521
rect 32160 -30555 32228 -30521
rect 32599 -30245 32667 -30211
rect 32599 -30555 32667 -30521
rect 33039 -30245 33107 -30211
rect 33039 -30555 33107 -30521
rect 33479 -30245 33547 -30211
rect 33479 -30555 33547 -30521
rect 34044 -30245 34112 -30211
rect 34202 -30245 34270 -30211
rect 34360 -30245 34428 -30211
rect 34044 -30555 34112 -30521
rect 34202 -30555 34270 -30521
rect 34360 -30555 34428 -30521
rect 34799 -30245 34867 -30211
rect 34799 -30555 34867 -30521
rect 35239 -30245 35307 -30211
rect 35239 -30555 35307 -30521
rect 35679 -30245 35747 -30211
rect 35679 -30555 35747 -30521
rect 36244 -30245 36312 -30211
rect 36402 -30245 36470 -30211
rect 36560 -30245 36628 -30211
rect 36244 -30555 36312 -30521
rect 36402 -30555 36470 -30521
rect 36560 -30555 36628 -30521
rect 36999 -30245 37067 -30211
rect 36999 -30555 37067 -30521
rect 37439 -30245 37507 -30211
rect 37439 -30555 37507 -30521
rect 37879 -30245 37947 -30211
rect 37879 -30555 37947 -30521
rect 31886 -31056 32254 -31022
rect 31886 -31284 32254 -31250
rect 32600 -31056 32668 -31022
rect 32600 -31584 32668 -31550
rect 33040 -31056 33108 -31022
rect 33040 -31584 33108 -31550
rect 33480 -31056 33548 -31022
rect 33480 -31584 33548 -31550
rect 34086 -31056 34454 -31022
rect 34086 -31284 34454 -31250
rect 34800 -31056 34868 -31022
rect 34800 -31584 34868 -31550
rect 35240 -31056 35308 -31022
rect 35240 -31584 35308 -31550
rect 35680 -31056 35748 -31022
rect 35680 -31584 35748 -31550
rect 36286 -31056 36654 -31022
rect 36286 -31284 36654 -31250
rect 37000 -31056 37068 -31022
rect 37000 -31584 37068 -31550
rect 37440 -31056 37508 -31022
rect 37440 -31584 37508 -31550
rect 37880 -31056 37948 -31022
rect 37880 -31584 37948 -31550
<< xpolycontact >>
rect 22366 11382 22936 11814
rect 22366 4566 22936 4998
rect 23032 11382 23602 11814
rect 23032 4566 23602 4998
rect 23698 11382 24268 11814
rect 23698 4566 24268 4998
rect 24364 11382 24934 11814
rect 24364 4566 24934 4998
rect 25030 11382 25600 11814
rect 25030 4566 25600 4998
rect 25696 11382 26266 11814
rect 25696 4566 26266 4998
rect 26362 11382 26932 11814
rect 26362 4566 26932 4998
rect 22347 -25097 22917 -24665
rect 22347 -31913 22917 -31481
rect 23013 -25097 23583 -24665
rect 23013 -31913 23583 -31481
rect 23679 -25097 24249 -24665
rect 23679 -31913 24249 -31481
rect 24345 -25097 24915 -24665
rect 24345 -31913 24915 -31481
rect 25011 -25097 25581 -24665
rect 25011 -31913 25581 -31481
rect 25677 -25097 26247 -24665
rect 25677 -31913 26247 -31481
rect 26343 -25097 26913 -24665
rect 26343 -31913 26913 -31481
<< ppolyres >>
rect 22366 4998 22936 11382
rect 23032 4998 23602 11382
rect 23698 4998 24268 11382
rect 24364 4998 24934 11382
rect 25030 4998 25600 11382
rect 25696 4998 26266 11382
rect 26362 4998 26932 11382
rect 22347 -31481 22917 -25097
rect 23013 -31481 23583 -25097
rect 23679 -31481 24249 -25097
rect 24345 -31481 24915 -25097
rect 25011 -31481 25581 -25097
rect 25677 -31481 26247 -25097
rect 26343 -31481 26913 -25097
<< locali >>
rect -300 11944 27280 12100
rect -300 11910 22332 11944
rect 26966 11910 27280 11944
rect 29960 11937 36840 12040
rect 29960 11920 30064 11937
rect -300 11909 22920 11910
rect -300 11875 145 11909
rect 1973 11875 2345 11909
rect 4173 11875 4545 11909
rect 6373 11875 6745 11909
rect 8573 11875 8945 11909
rect 10773 11875 11145 11909
rect 12973 11875 13345 11909
rect 15173 11875 15545 11909
rect 17373 11875 17745 11909
rect 19573 11875 19945 11909
rect 21773 11875 22920 11909
rect -300 11813 83 11875
rect -300 11345 49 11813
rect 300 11775 500 11875
rect 960 11775 1160 11875
rect 1620 11775 1820 11875
rect 2035 11813 2283 11875
rect 255 11741 271 11775
rect 1847 11741 1863 11775
rect 187 11713 221 11729
rect 83 11520 187 11620
rect 187 11429 221 11445
rect 1897 11713 1931 11729
rect 1931 11520 2035 11620
rect 1897 11429 1931 11445
rect 255 11383 271 11417
rect 1847 11383 1863 11417
rect -300 11283 83 11345
rect 280 11283 480 11383
rect 960 11283 1160 11383
rect 1620 11283 1820 11383
rect 2069 11345 2249 11813
rect 2500 11775 2700 11875
rect 3160 11775 3360 11875
rect 3820 11775 4020 11875
rect 4235 11813 4483 11875
rect 2455 11741 2471 11775
rect 4047 11741 4063 11775
rect 2387 11713 2421 11729
rect 2283 11520 2387 11620
rect 2387 11429 2421 11445
rect 4097 11713 4131 11729
rect 4131 11520 4235 11620
rect 4097 11429 4131 11445
rect 2455 11383 2471 11417
rect 4047 11383 4063 11417
rect 2035 11283 2283 11345
rect 2480 11283 2680 11383
rect 3160 11283 3360 11383
rect 3820 11283 4020 11383
rect 4269 11345 4449 11813
rect 4700 11775 4900 11875
rect 5360 11775 5560 11875
rect 6020 11775 6220 11875
rect 6435 11813 6683 11875
rect 4655 11741 4671 11775
rect 6247 11741 6263 11775
rect 4587 11713 4621 11729
rect 4483 11520 4587 11620
rect 4587 11429 4621 11445
rect 6297 11713 6331 11729
rect 6331 11520 6435 11620
rect 6297 11429 6331 11445
rect 4655 11383 4671 11417
rect 6247 11383 6263 11417
rect 4235 11283 4483 11345
rect 4680 11283 4880 11383
rect 5360 11283 5560 11383
rect 6020 11283 6220 11383
rect 6469 11345 6649 11813
rect 6900 11775 7100 11875
rect 7560 11775 7760 11875
rect 8220 11775 8420 11875
rect 8635 11813 8883 11875
rect 6855 11741 6871 11775
rect 8447 11741 8463 11775
rect 6787 11713 6821 11729
rect 6683 11520 6787 11620
rect 6787 11429 6821 11445
rect 8497 11713 8531 11729
rect 8531 11520 8635 11620
rect 8497 11429 8531 11445
rect 6855 11383 6871 11417
rect 8447 11383 8463 11417
rect 6435 11283 6683 11345
rect 6880 11283 7080 11383
rect 7560 11283 7760 11383
rect 8220 11283 8420 11383
rect 8669 11345 8849 11813
rect 9100 11775 9300 11875
rect 9760 11775 9960 11875
rect 10420 11775 10620 11875
rect 10835 11813 11083 11875
rect 9055 11741 9071 11775
rect 10647 11741 10663 11775
rect 8987 11713 9021 11729
rect 8883 11520 8987 11620
rect 8987 11429 9021 11445
rect 10697 11713 10731 11729
rect 10731 11520 10835 11620
rect 10697 11429 10731 11445
rect 9055 11383 9071 11417
rect 10647 11383 10663 11417
rect 8635 11283 8883 11345
rect 9080 11283 9280 11383
rect 9760 11283 9960 11383
rect 10420 11283 10620 11383
rect 10869 11345 11049 11813
rect 11300 11775 11500 11875
rect 11960 11775 12160 11875
rect 12620 11775 12820 11875
rect 13035 11813 13283 11875
rect 11255 11741 11271 11775
rect 12847 11741 12863 11775
rect 11187 11713 11221 11729
rect 11083 11520 11187 11620
rect 11187 11429 11221 11445
rect 12897 11713 12931 11729
rect 12931 11520 13035 11620
rect 12897 11429 12931 11445
rect 11255 11383 11271 11417
rect 12847 11383 12863 11417
rect 10835 11283 11083 11345
rect 11280 11283 11480 11383
rect 11960 11283 12160 11383
rect 12620 11283 12820 11383
rect 13069 11345 13249 11813
rect 13500 11775 13700 11875
rect 14160 11775 14360 11875
rect 14820 11775 15020 11875
rect 15235 11813 15483 11875
rect 13455 11741 13471 11775
rect 15047 11741 15063 11775
rect 13387 11713 13421 11729
rect 13283 11520 13387 11620
rect 13387 11429 13421 11445
rect 15097 11713 15131 11729
rect 15131 11520 15235 11620
rect 15097 11429 15131 11445
rect 13455 11383 13471 11417
rect 15047 11383 15063 11417
rect 13035 11283 13283 11345
rect 13480 11283 13680 11383
rect 14160 11283 14360 11383
rect 14820 11283 15020 11383
rect 15269 11345 15449 11813
rect 15700 11775 15900 11875
rect 16360 11775 16560 11875
rect 17020 11775 17220 11875
rect 17435 11813 17683 11875
rect 15655 11741 15671 11775
rect 17247 11741 17263 11775
rect 15587 11713 15621 11729
rect 15483 11520 15587 11620
rect 15587 11429 15621 11445
rect 17297 11713 17331 11729
rect 17331 11520 17435 11620
rect 17297 11429 17331 11445
rect 15655 11383 15671 11417
rect 17247 11383 17263 11417
rect 15235 11283 15483 11345
rect 15680 11283 15880 11383
rect 16360 11283 16560 11383
rect 17020 11283 17220 11383
rect 17469 11345 17649 11813
rect 17900 11775 18100 11875
rect 18560 11775 18760 11875
rect 19220 11775 19420 11875
rect 19635 11813 19883 11875
rect 17855 11741 17871 11775
rect 19447 11741 19463 11775
rect 17787 11713 17821 11729
rect 17683 11520 17787 11620
rect 17787 11429 17821 11445
rect 19497 11713 19531 11729
rect 19531 11520 19635 11620
rect 19497 11429 19531 11445
rect 17855 11383 17871 11417
rect 19447 11383 19463 11417
rect 17435 11283 17683 11345
rect 17880 11283 18080 11383
rect 18560 11283 18760 11383
rect 19220 11283 19420 11383
rect 19669 11345 19849 11813
rect 20100 11775 20300 11875
rect 20760 11775 20960 11875
rect 21420 11775 21620 11875
rect 21835 11848 22920 11875
rect 21835 11813 22236 11848
rect 20055 11741 20071 11775
rect 21647 11741 21663 11775
rect 19987 11713 20021 11729
rect 19883 11520 19987 11620
rect 19987 11429 20021 11445
rect 21697 11713 21731 11729
rect 21731 11520 21835 11620
rect 21697 11429 21731 11445
rect 20055 11383 20071 11417
rect 21647 11383 21663 11417
rect 19635 11283 19883 11345
rect 20080 11283 20280 11383
rect 20760 11283 20960 11383
rect 21420 11283 21620 11383
rect 21869 11345 22236 11813
rect 22270 11814 22920 11848
rect 26380 11848 27280 11910
rect 26380 11814 27028 11848
rect 21835 11283 22236 11345
rect -300 11249 145 11283
rect 1973 11249 2345 11283
rect 4173 11249 4545 11283
rect 6373 11249 6745 11283
rect 8573 11249 8945 11283
rect 10773 11249 11145 11283
rect 12973 11249 13345 11283
rect 15173 11249 15545 11283
rect 17373 11249 17745 11283
rect 19573 11249 19945 11283
rect 21773 11249 22236 11283
rect -300 11109 22236 11249
rect -300 11075 145 11109
rect 1973 11108 19945 11109
rect 1973 11075 2344 11108
rect -300 11013 83 11075
rect -300 10930 49 11013
rect -300 10870 -70 10930
rect -10 10870 49 10930
rect -300 10545 49 10870
rect 300 10975 500 11075
rect 960 10975 1160 11075
rect 1620 10975 1820 11075
rect 2035 11074 2344 11075
rect 4172 11074 4544 11108
rect 6372 11074 6744 11108
rect 8572 11074 8944 11108
rect 10772 11074 11144 11108
rect 12972 11074 13344 11108
rect 15172 11074 15544 11108
rect 17372 11074 17744 11108
rect 19572 11075 19945 11108
rect 21773 11075 22236 11109
rect 19572 11074 19883 11075
rect 2035 11013 2282 11074
rect 255 10941 271 10975
rect 1847 10941 1863 10975
rect 187 10913 221 10929
rect 83 10720 187 10820
rect 187 10629 221 10645
rect 1897 10913 1931 10929
rect 1931 10720 2035 10820
rect 1897 10629 1931 10645
rect 255 10583 271 10617
rect 1847 10583 1863 10617
rect -300 10483 83 10545
rect 280 10483 480 10583
rect 960 10483 1160 10583
rect 1620 10483 1820 10583
rect 2069 11012 2282 11013
rect 2069 10930 2248 11012
rect 2069 10870 2130 10930
rect 2190 10870 2248 10930
rect 2069 10545 2248 10870
rect 2035 10544 2248 10545
rect 4234 11012 4482 11074
rect 2454 10940 2470 10974
rect 4046 10940 4062 10974
rect 2386 10912 2420 10928
rect 2386 10628 2420 10644
rect 4096 10912 4130 10928
rect 4096 10628 4130 10644
rect 2454 10582 2470 10616
rect 4046 10582 4062 10616
rect 2035 10483 2282 10544
rect -300 10449 145 10483
rect 1973 10482 2282 10483
rect 4268 10930 4448 11012
rect 4268 10870 4330 10930
rect 4390 10870 4448 10930
rect 4268 10544 4448 10870
rect 6434 11012 6682 11074
rect 4654 10940 4670 10974
rect 6246 10940 6262 10974
rect 4586 10912 4620 10928
rect 4586 10628 4620 10644
rect 6296 10912 6330 10928
rect 6296 10628 6330 10644
rect 4654 10582 4670 10616
rect 6246 10582 6262 10616
rect 4234 10482 4482 10544
rect 6468 10930 6648 11012
rect 6468 10870 6530 10930
rect 6590 10870 6648 10930
rect 6468 10544 6648 10870
rect 8634 11012 8882 11074
rect 6854 10940 6870 10974
rect 8446 10940 8462 10974
rect 6786 10912 6820 10928
rect 6786 10628 6820 10644
rect 8496 10912 8530 10928
rect 8496 10628 8530 10644
rect 6854 10582 6870 10616
rect 8446 10582 8462 10616
rect 6434 10482 6682 10544
rect 8668 10930 8848 11012
rect 8668 10870 8730 10930
rect 8790 10870 8848 10930
rect 8668 10544 8848 10870
rect 10834 11012 11082 11074
rect 9054 10940 9070 10974
rect 10646 10940 10662 10974
rect 8986 10912 9020 10928
rect 8986 10628 9020 10644
rect 10696 10912 10730 10928
rect 10696 10628 10730 10644
rect 9054 10582 9070 10616
rect 10646 10582 10662 10616
rect 8634 10482 8882 10544
rect 10868 10930 11048 11012
rect 10868 10870 10930 10930
rect 10990 10870 11048 10930
rect 10868 10544 11048 10870
rect 13034 11012 13282 11074
rect 11254 10940 11270 10974
rect 12846 10940 12862 10974
rect 11186 10912 11220 10928
rect 11186 10628 11220 10644
rect 12896 10912 12930 10928
rect 12896 10628 12930 10644
rect 11254 10582 11270 10616
rect 12846 10582 12862 10616
rect 10834 10482 11082 10544
rect 13068 10930 13248 11012
rect 13068 10870 13130 10930
rect 13190 10870 13248 10930
rect 13068 10544 13248 10870
rect 15234 11012 15482 11074
rect 13454 10940 13470 10974
rect 15046 10940 15062 10974
rect 13386 10912 13420 10928
rect 13386 10628 13420 10644
rect 15096 10912 15130 10928
rect 15096 10628 15130 10644
rect 13454 10582 13470 10616
rect 15046 10582 15062 10616
rect 13034 10482 13282 10544
rect 15268 10930 15448 11012
rect 15268 10870 15330 10930
rect 15390 10870 15448 10930
rect 15268 10544 15448 10870
rect 17434 11012 17682 11074
rect 15654 10940 15670 10974
rect 17246 10940 17262 10974
rect 15586 10912 15620 10928
rect 15586 10628 15620 10644
rect 17296 10912 17330 10928
rect 17296 10628 17330 10644
rect 15654 10582 15670 10616
rect 17246 10582 17262 10616
rect 15234 10482 15482 10544
rect 17468 10930 17648 11012
rect 17468 10870 17530 10930
rect 17590 10870 17648 10930
rect 17468 10544 17648 10870
rect 19634 11013 19883 11074
rect 19634 11012 19849 11013
rect 17854 10940 17870 10974
rect 19446 10940 19462 10974
rect 17786 10912 17820 10928
rect 17786 10628 17820 10644
rect 19496 10912 19530 10928
rect 19496 10628 19530 10644
rect 17854 10582 17870 10616
rect 19446 10582 19462 10616
rect 17434 10482 17682 10544
rect 19668 10930 19849 11012
rect 19668 10870 19730 10930
rect 19790 10870 19849 10930
rect 19668 10545 19849 10870
rect 20100 10975 20300 11075
rect 20760 10975 20960 11075
rect 21420 10975 21620 11075
rect 21835 11013 22236 11075
rect 20055 10941 20071 10975
rect 21647 10941 21663 10975
rect 19987 10913 20021 10929
rect 19883 10720 19987 10820
rect 19987 10629 20021 10645
rect 21697 10913 21731 10929
rect 21731 10720 21835 10820
rect 21697 10629 21731 10645
rect 20055 10583 20071 10617
rect 21647 10583 21663 10617
rect 19668 10544 19883 10545
rect 19634 10483 19883 10544
rect 20080 10483 20280 10583
rect 20760 10483 20960 10583
rect 21420 10483 21620 10583
rect 21869 10930 22236 11013
rect 21869 10870 21930 10930
rect 21990 10870 22236 10930
rect 21869 10545 22236 10870
rect 21835 10483 22236 10545
rect 19634 10482 19945 10483
rect 1973 10449 2344 10482
rect -300 10448 2344 10449
rect 4172 10448 4544 10482
rect 6372 10448 6744 10482
rect 8572 10448 8944 10482
rect 10772 10448 11144 10482
rect 12972 10448 13344 10482
rect 15172 10448 15544 10482
rect 17372 10448 17744 10482
rect 19572 10449 19945 10482
rect 21773 10449 22236 10483
rect 19572 10448 22236 10449
rect -300 10309 22236 10448
rect -300 10275 145 10309
rect 1973 10308 19945 10309
rect 1973 10275 2344 10308
rect -300 10213 83 10275
rect -300 10130 49 10213
rect -300 10070 -70 10130
rect -10 10070 49 10130
rect -300 9745 49 10070
rect 300 10175 500 10275
rect 960 10175 1160 10275
rect 1620 10175 1820 10275
rect 2035 10274 2344 10275
rect 4172 10274 4544 10308
rect 6372 10274 6744 10308
rect 8572 10274 8944 10308
rect 10772 10274 11144 10308
rect 12972 10274 13344 10308
rect 15172 10274 15544 10308
rect 17372 10274 17744 10308
rect 19572 10275 19945 10308
rect 21773 10275 22236 10309
rect 19572 10274 19883 10275
rect 2035 10213 2282 10274
rect 255 10141 271 10175
rect 1847 10141 1863 10175
rect 187 10113 221 10129
rect 83 9920 187 10020
rect 187 9829 221 9845
rect 1897 10113 1931 10129
rect 1931 9920 2035 10020
rect 1897 9829 1931 9845
rect 255 9783 271 9817
rect 1847 9783 1863 9817
rect -300 9683 83 9745
rect 280 9683 480 9783
rect 960 9683 1160 9783
rect 1620 9683 1820 9783
rect 2069 10212 2282 10213
rect 2069 10130 2248 10212
rect 2069 10070 2130 10130
rect 2190 10070 2248 10130
rect 2069 9745 2248 10070
rect 2035 9744 2248 9745
rect 4234 10212 4482 10274
rect 2454 10140 2470 10174
rect 4046 10140 4062 10174
rect 2386 10112 2420 10128
rect 2386 9828 2420 9844
rect 4096 10112 4130 10128
rect 4096 9828 4130 9844
rect 2454 9782 2470 9816
rect 4046 9782 4062 9816
rect 2035 9683 2282 9744
rect -300 9649 145 9683
rect 1973 9682 2282 9683
rect 4268 10130 4448 10212
rect 4268 10070 4330 10130
rect 4390 10070 4448 10130
rect 4268 9744 4448 10070
rect 6434 10212 6682 10274
rect 4654 10140 4670 10174
rect 6246 10140 6262 10174
rect 4586 10112 4620 10128
rect 4586 9828 4620 9844
rect 6296 10112 6330 10128
rect 6296 9828 6330 9844
rect 4654 9782 4670 9816
rect 6246 9782 6262 9816
rect 4234 9682 4482 9744
rect 6468 10130 6648 10212
rect 6468 10070 6530 10130
rect 6590 10070 6648 10130
rect 6468 9744 6648 10070
rect 8634 10212 8882 10274
rect 6854 10140 6870 10174
rect 8446 10140 8462 10174
rect 6786 10112 6820 10128
rect 6786 9828 6820 9844
rect 8496 10112 8530 10128
rect 8496 9828 8530 9844
rect 6854 9782 6870 9816
rect 8446 9782 8462 9816
rect 6434 9682 6682 9744
rect 8668 10130 8848 10212
rect 8668 10070 8730 10130
rect 8790 10070 8848 10130
rect 8668 9744 8848 10070
rect 10834 10212 11082 10274
rect 9054 10140 9070 10174
rect 10646 10140 10662 10174
rect 8986 10112 9020 10128
rect 8986 9828 9020 9844
rect 10696 10112 10730 10128
rect 10696 9828 10730 9844
rect 9054 9782 9070 9816
rect 10646 9782 10662 9816
rect 8634 9682 8882 9744
rect 10868 10130 11048 10212
rect 10868 10070 10930 10130
rect 10990 10070 11048 10130
rect 10868 9744 11048 10070
rect 13034 10212 13282 10274
rect 11254 10140 11270 10174
rect 12846 10140 12862 10174
rect 11186 10112 11220 10128
rect 11186 9828 11220 9844
rect 12896 10112 12930 10128
rect 12896 9828 12930 9844
rect 11254 9782 11270 9816
rect 12846 9782 12862 9816
rect 10834 9682 11082 9744
rect 13068 10130 13248 10212
rect 13068 10070 13130 10130
rect 13190 10070 13248 10130
rect 13068 9744 13248 10070
rect 15234 10212 15482 10274
rect 13454 10140 13470 10174
rect 15046 10140 15062 10174
rect 13386 10112 13420 10128
rect 13386 9828 13420 9844
rect 15096 10112 15130 10128
rect 15096 9828 15130 9844
rect 13454 9782 13470 9816
rect 15046 9782 15062 9816
rect 13034 9682 13282 9744
rect 15268 10130 15448 10212
rect 15268 10070 15330 10130
rect 15390 10070 15448 10130
rect 15268 9744 15448 10070
rect 17434 10212 17682 10274
rect 15654 10140 15670 10174
rect 17246 10140 17262 10174
rect 15586 10112 15620 10128
rect 15586 9828 15620 9844
rect 17296 10112 17330 10128
rect 17296 9828 17330 9844
rect 15654 9782 15670 9816
rect 17246 9782 17262 9816
rect 15234 9682 15482 9744
rect 17468 10130 17648 10212
rect 17468 10070 17530 10130
rect 17590 10070 17648 10130
rect 17468 9744 17648 10070
rect 19634 10213 19883 10274
rect 19634 10212 19849 10213
rect 17854 10140 17870 10174
rect 19446 10140 19462 10174
rect 17786 10112 17820 10128
rect 17786 9828 17820 9844
rect 19496 10112 19530 10128
rect 19496 9828 19530 9844
rect 17854 9782 17870 9816
rect 19446 9782 19462 9816
rect 17434 9682 17682 9744
rect 19668 10130 19849 10212
rect 19668 10070 19730 10130
rect 19790 10070 19849 10130
rect 19668 9745 19849 10070
rect 20100 10175 20300 10275
rect 20760 10175 20960 10275
rect 21420 10175 21620 10275
rect 21835 10213 22236 10275
rect 20055 10141 20071 10175
rect 21647 10141 21663 10175
rect 19987 10113 20021 10129
rect 19883 9920 19987 10020
rect 19987 9829 20021 9845
rect 21697 10113 21731 10129
rect 21731 9920 21835 10020
rect 21697 9829 21731 9845
rect 20055 9783 20071 9817
rect 21647 9783 21663 9817
rect 19668 9744 19883 9745
rect 19634 9683 19883 9744
rect 20080 9683 20280 9783
rect 20760 9683 20960 9783
rect 21420 9683 21620 9783
rect 21869 10130 22236 10213
rect 21869 10070 21930 10130
rect 21990 10070 22236 10130
rect 21869 9745 22236 10070
rect 21835 9683 22236 9745
rect 19634 9682 19945 9683
rect 1973 9649 2344 9682
rect -300 9648 2344 9649
rect 4172 9648 4544 9682
rect 6372 9648 6744 9682
rect 8572 9648 8944 9682
rect 10772 9648 11144 9682
rect 12972 9648 13344 9682
rect 15172 9648 15544 9682
rect 17372 9648 17744 9682
rect 19572 9649 19945 9682
rect 21773 9649 22236 9683
rect 19572 9648 22236 9649
rect -300 9509 22236 9648
rect -300 9475 145 9509
rect 1973 9508 19945 9509
rect 1973 9475 2344 9508
rect -300 9413 83 9475
rect -300 9330 49 9413
rect -300 9270 -70 9330
rect -10 9270 49 9330
rect -300 8945 49 9270
rect 300 9375 500 9475
rect 960 9375 1160 9475
rect 1620 9375 1820 9475
rect 2035 9474 2344 9475
rect 4172 9474 4544 9508
rect 6372 9474 6744 9508
rect 8572 9474 8944 9508
rect 10772 9474 11144 9508
rect 12972 9474 13344 9508
rect 15172 9474 15544 9508
rect 17372 9474 17744 9508
rect 19572 9475 19945 9508
rect 21773 9475 22236 9509
rect 19572 9474 19883 9475
rect 2035 9413 2282 9474
rect 255 9341 271 9375
rect 1847 9341 1863 9375
rect 187 9313 221 9329
rect 83 9120 187 9220
rect 187 9029 221 9045
rect 1897 9313 1931 9329
rect 1931 9120 2035 9220
rect 1897 9029 1931 9045
rect 255 8983 271 9017
rect 1847 8983 1863 9017
rect -300 8883 83 8945
rect 280 8883 480 8983
rect 960 8883 1160 8983
rect 1620 8883 1820 8983
rect 2069 9412 2282 9413
rect 2069 9330 2248 9412
rect 2069 9270 2130 9330
rect 2190 9270 2248 9330
rect 2069 8945 2248 9270
rect 2035 8944 2248 8945
rect 4234 9412 4482 9474
rect 2454 9340 2470 9374
rect 4046 9340 4062 9374
rect 2386 9312 2420 9328
rect 2386 9028 2420 9044
rect 4096 9312 4130 9328
rect 4096 9028 4130 9044
rect 2454 8982 2470 9016
rect 4046 8982 4062 9016
rect 2035 8883 2282 8944
rect -300 8849 145 8883
rect 1973 8882 2282 8883
rect 4268 9330 4448 9412
rect 4268 9270 4330 9330
rect 4390 9270 4448 9330
rect 4268 8944 4448 9270
rect 6434 9412 6682 9474
rect 4654 9340 4670 9374
rect 6246 9340 6262 9374
rect 4586 9312 4620 9328
rect 4586 9028 4620 9044
rect 6296 9312 6330 9328
rect 6296 9028 6330 9044
rect 4654 8982 4670 9016
rect 6246 8982 6262 9016
rect 4234 8882 4482 8944
rect 6468 9330 6648 9412
rect 6468 9270 6530 9330
rect 6590 9270 6648 9330
rect 6468 8944 6648 9270
rect 8634 9412 8882 9474
rect 6854 9340 6870 9374
rect 8446 9340 8462 9374
rect 6786 9312 6820 9328
rect 6786 9028 6820 9044
rect 8496 9312 8530 9328
rect 8496 9028 8530 9044
rect 6854 8982 6870 9016
rect 8446 8982 8462 9016
rect 6434 8882 6682 8944
rect 8668 9330 8848 9412
rect 8668 9270 8730 9330
rect 8790 9270 8848 9330
rect 8668 8944 8848 9270
rect 10834 9412 11082 9474
rect 9054 9340 9070 9374
rect 10646 9340 10662 9374
rect 8986 9312 9020 9328
rect 8986 9028 9020 9044
rect 10696 9312 10730 9328
rect 10696 9028 10730 9044
rect 9054 8982 9070 9016
rect 10646 8982 10662 9016
rect 8634 8882 8882 8944
rect 10868 9330 11048 9412
rect 10868 9270 10930 9330
rect 10990 9270 11048 9330
rect 10868 8944 11048 9270
rect 13034 9412 13282 9474
rect 11254 9340 11270 9374
rect 12846 9340 12862 9374
rect 11186 9312 11220 9328
rect 11186 9028 11220 9044
rect 12896 9312 12930 9328
rect 12896 9028 12930 9044
rect 11254 8982 11270 9016
rect 12846 8982 12862 9016
rect 10834 8882 11082 8944
rect 13068 9330 13248 9412
rect 13068 9270 13130 9330
rect 13190 9270 13248 9330
rect 13068 8944 13248 9270
rect 15234 9412 15482 9474
rect 13454 9340 13470 9374
rect 15046 9340 15062 9374
rect 13386 9312 13420 9328
rect 13386 9028 13420 9044
rect 15096 9312 15130 9328
rect 15096 9028 15130 9044
rect 13454 8982 13470 9016
rect 15046 8982 15062 9016
rect 13034 8882 13282 8944
rect 15268 9330 15448 9412
rect 15268 9270 15330 9330
rect 15390 9270 15448 9330
rect 15268 8944 15448 9270
rect 17434 9412 17682 9474
rect 15654 9340 15670 9374
rect 17246 9340 17262 9374
rect 15586 9312 15620 9328
rect 15586 9028 15620 9044
rect 17296 9312 17330 9328
rect 17296 9028 17330 9044
rect 15654 8982 15670 9016
rect 17246 8982 17262 9016
rect 15234 8882 15482 8944
rect 17468 9330 17648 9412
rect 17468 9270 17530 9330
rect 17590 9270 17648 9330
rect 17468 8944 17648 9270
rect 19634 9413 19883 9474
rect 19634 9412 19849 9413
rect 17854 9340 17870 9374
rect 19446 9340 19462 9374
rect 17786 9312 17820 9328
rect 17786 9028 17820 9044
rect 19496 9312 19530 9328
rect 19496 9028 19530 9044
rect 17854 8982 17870 9016
rect 19446 8982 19462 9016
rect 17434 8882 17682 8944
rect 19668 9330 19849 9412
rect 19668 9270 19730 9330
rect 19790 9270 19849 9330
rect 19668 8945 19849 9270
rect 20100 9375 20300 9475
rect 20760 9375 20960 9475
rect 21420 9375 21620 9475
rect 21835 9413 22236 9475
rect 20055 9341 20071 9375
rect 21647 9341 21663 9375
rect 19987 9313 20021 9329
rect 19883 9120 19987 9220
rect 19987 9029 20021 9045
rect 21697 9313 21731 9329
rect 21731 9120 21835 9220
rect 21697 9029 21731 9045
rect 20055 8983 20071 9017
rect 21647 8983 21663 9017
rect 19668 8944 19883 8945
rect 19634 8883 19883 8944
rect 20080 8883 20280 8983
rect 20760 8883 20960 8983
rect 21420 8883 21620 8983
rect 21869 9330 22236 9413
rect 21869 9270 21930 9330
rect 21990 9270 22236 9330
rect 21869 8945 22236 9270
rect 21835 8883 22236 8945
rect 19634 8882 19945 8883
rect 1973 8849 2344 8882
rect -300 8848 2344 8849
rect 4172 8848 4544 8882
rect 6372 8848 6744 8882
rect 8572 8848 8944 8882
rect 10772 8848 11144 8882
rect 12972 8848 13344 8882
rect 15172 8848 15544 8882
rect 17372 8848 17744 8882
rect 19572 8849 19945 8882
rect 21773 8849 22236 8883
rect 19572 8848 22236 8849
rect -300 8709 22236 8848
rect -300 8675 145 8709
rect 1973 8708 19945 8709
rect 1973 8675 2344 8708
rect -300 8613 83 8675
rect -300 8530 49 8613
rect -300 8470 -70 8530
rect -10 8470 49 8530
rect -300 8145 49 8470
rect 300 8575 500 8675
rect 960 8575 1160 8675
rect 1620 8575 1820 8675
rect 2035 8674 2344 8675
rect 4172 8674 4544 8708
rect 6372 8674 6744 8708
rect 8572 8674 8944 8708
rect 10772 8674 11144 8708
rect 12972 8674 13344 8708
rect 15172 8674 15544 8708
rect 17372 8674 17744 8708
rect 19572 8675 19945 8708
rect 21773 8675 22236 8709
rect 19572 8674 19883 8675
rect 2035 8613 2282 8674
rect 255 8541 271 8575
rect 1847 8541 1863 8575
rect 187 8513 221 8529
rect 83 8320 187 8420
rect 187 8229 221 8245
rect 1897 8513 1931 8529
rect 1931 8320 2035 8420
rect 1897 8229 1931 8245
rect 255 8183 271 8217
rect 1847 8183 1863 8217
rect -300 8083 83 8145
rect 280 8083 480 8183
rect 960 8083 1160 8183
rect 1620 8083 1820 8183
rect 2069 8612 2282 8613
rect 2069 8530 2248 8612
rect 2069 8470 2130 8530
rect 2190 8470 2248 8530
rect 2069 8145 2248 8470
rect 2035 8144 2248 8145
rect 4234 8612 4482 8674
rect 2454 8540 2470 8574
rect 4046 8540 4062 8574
rect 2386 8512 2420 8528
rect 2386 8228 2420 8244
rect 4096 8512 4130 8528
rect 4096 8228 4130 8244
rect 2454 8182 2470 8216
rect 4046 8182 4062 8216
rect 2035 8083 2282 8144
rect -300 8049 145 8083
rect 1973 8082 2282 8083
rect 4268 8530 4448 8612
rect 4268 8470 4330 8530
rect 4390 8470 4448 8530
rect 4268 8144 4448 8470
rect 6434 8612 6682 8674
rect 4654 8540 4670 8574
rect 6246 8540 6262 8574
rect 4586 8512 4620 8528
rect 4586 8228 4620 8244
rect 6296 8512 6330 8528
rect 6296 8228 6330 8244
rect 4654 8182 4670 8216
rect 6246 8182 6262 8216
rect 4234 8082 4482 8144
rect 6468 8530 6648 8612
rect 6468 8470 6530 8530
rect 6590 8470 6648 8530
rect 6468 8144 6648 8470
rect 8634 8612 8882 8674
rect 6854 8540 6870 8574
rect 8446 8540 8462 8574
rect 6786 8512 6820 8528
rect 6786 8228 6820 8244
rect 8496 8512 8530 8528
rect 8496 8228 8530 8244
rect 6854 8182 6870 8216
rect 8446 8182 8462 8216
rect 6434 8082 6682 8144
rect 8668 8530 8848 8612
rect 8668 8470 8730 8530
rect 8790 8470 8848 8530
rect 8668 8144 8848 8470
rect 10834 8612 11082 8674
rect 9054 8540 9070 8574
rect 10646 8540 10662 8574
rect 8986 8512 9020 8528
rect 8986 8228 9020 8244
rect 10696 8512 10730 8528
rect 10696 8228 10730 8244
rect 9054 8182 9070 8216
rect 10646 8182 10662 8216
rect 8634 8082 8882 8144
rect 10868 8530 11048 8612
rect 10868 8470 10930 8530
rect 10990 8470 11048 8530
rect 10868 8144 11048 8470
rect 13034 8612 13282 8674
rect 11254 8540 11270 8574
rect 12846 8540 12862 8574
rect 11186 8512 11220 8528
rect 11186 8228 11220 8244
rect 12896 8512 12930 8528
rect 12896 8228 12930 8244
rect 11254 8182 11270 8216
rect 12846 8182 12862 8216
rect 10834 8082 11082 8144
rect 13068 8530 13248 8612
rect 13068 8470 13130 8530
rect 13190 8470 13248 8530
rect 13068 8144 13248 8470
rect 15234 8612 15482 8674
rect 13454 8540 13470 8574
rect 15046 8540 15062 8574
rect 13386 8512 13420 8528
rect 13386 8228 13420 8244
rect 15096 8512 15130 8528
rect 15096 8228 15130 8244
rect 13454 8182 13470 8216
rect 15046 8182 15062 8216
rect 13034 8082 13282 8144
rect 15268 8530 15448 8612
rect 15268 8470 15330 8530
rect 15390 8470 15448 8530
rect 15268 8144 15448 8470
rect 17434 8612 17682 8674
rect 15654 8540 15670 8574
rect 17246 8540 17262 8574
rect 15586 8512 15620 8528
rect 15586 8228 15620 8244
rect 17296 8512 17330 8528
rect 17296 8228 17330 8244
rect 15654 8182 15670 8216
rect 17246 8182 17262 8216
rect 15234 8082 15482 8144
rect 17468 8530 17648 8612
rect 17468 8470 17530 8530
rect 17590 8470 17648 8530
rect 17468 8144 17648 8470
rect 19634 8613 19883 8674
rect 19634 8612 19849 8613
rect 17854 8540 17870 8574
rect 19446 8540 19462 8574
rect 17786 8512 17820 8528
rect 17786 8228 17820 8244
rect 19496 8512 19530 8528
rect 19496 8228 19530 8244
rect 17854 8182 17870 8216
rect 19446 8182 19462 8216
rect 17434 8082 17682 8144
rect 19668 8530 19849 8612
rect 19668 8470 19730 8530
rect 19790 8470 19849 8530
rect 19668 8145 19849 8470
rect 20100 8575 20300 8675
rect 20760 8575 20960 8675
rect 21420 8575 21620 8675
rect 21835 8613 22236 8675
rect 20055 8541 20071 8575
rect 21647 8541 21663 8575
rect 19987 8513 20021 8529
rect 19883 8320 19987 8420
rect 19987 8229 20021 8245
rect 21697 8513 21731 8529
rect 21731 8320 21835 8420
rect 21697 8229 21731 8245
rect 20055 8183 20071 8217
rect 21647 8183 21663 8217
rect 19668 8144 19883 8145
rect 19634 8083 19883 8144
rect 20080 8083 20280 8183
rect 20760 8083 20960 8183
rect 21420 8083 21620 8183
rect 21869 8530 22236 8613
rect 21869 8470 21930 8530
rect 21990 8470 22236 8530
rect 21869 8145 22236 8470
rect 21835 8083 22236 8145
rect 19634 8082 19945 8083
rect 1973 8049 2344 8082
rect -300 8048 2344 8049
rect 4172 8048 4544 8082
rect 6372 8048 6744 8082
rect 8572 8048 8944 8082
rect 10772 8048 11144 8082
rect 12972 8048 13344 8082
rect 15172 8048 15544 8082
rect 17372 8048 17744 8082
rect 19572 8049 19945 8082
rect 21773 8049 22236 8083
rect 19572 8048 22236 8049
rect -300 7909 22236 8048
rect -300 7875 145 7909
rect 1973 7908 19945 7909
rect 1973 7875 2344 7908
rect -300 7813 83 7875
rect -300 7730 49 7813
rect -300 7670 -70 7730
rect -10 7670 49 7730
rect -300 7345 49 7670
rect 300 7775 500 7875
rect 960 7775 1160 7875
rect 1620 7775 1820 7875
rect 2035 7874 2344 7875
rect 4172 7874 4544 7908
rect 6372 7874 6744 7908
rect 8572 7874 8944 7908
rect 10772 7874 11144 7908
rect 12972 7874 13344 7908
rect 15172 7874 15544 7908
rect 17372 7874 17744 7908
rect 19572 7875 19945 7908
rect 21773 7875 22236 7909
rect 19572 7874 19883 7875
rect 2035 7813 2282 7874
rect 255 7741 271 7775
rect 1847 7741 1863 7775
rect 187 7713 221 7729
rect 83 7520 187 7620
rect 187 7429 221 7445
rect 1897 7713 1931 7729
rect 1931 7520 2035 7620
rect 1897 7429 1931 7445
rect 255 7383 271 7417
rect 1847 7383 1863 7417
rect -300 7283 83 7345
rect 280 7283 480 7383
rect 960 7283 1160 7383
rect 1620 7283 1820 7383
rect 2069 7812 2282 7813
rect 2069 7730 2248 7812
rect 2069 7670 2130 7730
rect 2190 7670 2248 7730
rect 2069 7345 2248 7670
rect 2035 7344 2248 7345
rect 4234 7812 4482 7874
rect 2454 7740 2470 7774
rect 4046 7740 4062 7774
rect 2386 7712 2420 7728
rect 2386 7428 2420 7444
rect 4096 7712 4130 7728
rect 4096 7428 4130 7444
rect 2454 7382 2470 7416
rect 4046 7382 4062 7416
rect 2035 7283 2282 7344
rect -300 7249 145 7283
rect 1973 7282 2282 7283
rect 4268 7730 4448 7812
rect 4268 7670 4330 7730
rect 4390 7670 4448 7730
rect 4268 7344 4448 7670
rect 6434 7812 6682 7874
rect 4654 7740 4670 7774
rect 6246 7740 6262 7774
rect 4586 7712 4620 7728
rect 4586 7428 4620 7444
rect 6296 7712 6330 7728
rect 6296 7428 6330 7444
rect 4654 7382 4670 7416
rect 6246 7382 6262 7416
rect 4234 7282 4482 7344
rect 6468 7730 6648 7812
rect 6468 7670 6530 7730
rect 6590 7670 6648 7730
rect 6468 7344 6648 7670
rect 8634 7812 8882 7874
rect 6854 7740 6870 7774
rect 8446 7740 8462 7774
rect 6786 7712 6820 7728
rect 6786 7428 6820 7444
rect 8496 7712 8530 7728
rect 8496 7428 8530 7444
rect 6854 7382 6870 7416
rect 8446 7382 8462 7416
rect 6434 7282 6682 7344
rect 8668 7730 8848 7812
rect 8668 7670 8730 7730
rect 8790 7670 8848 7730
rect 8668 7344 8848 7670
rect 10834 7812 11082 7874
rect 9054 7740 9070 7774
rect 10646 7740 10662 7774
rect 8986 7712 9020 7728
rect 8986 7428 9020 7444
rect 10696 7712 10730 7728
rect 10696 7428 10730 7444
rect 9054 7382 9070 7416
rect 10646 7382 10662 7416
rect 8634 7282 8882 7344
rect 10868 7730 11048 7812
rect 10868 7670 10930 7730
rect 10990 7670 11048 7730
rect 10868 7344 11048 7670
rect 13034 7812 13282 7874
rect 11254 7740 11270 7774
rect 12846 7740 12862 7774
rect 11186 7712 11220 7728
rect 11186 7428 11220 7444
rect 12896 7712 12930 7728
rect 12896 7428 12930 7444
rect 11254 7382 11270 7416
rect 12846 7382 12862 7416
rect 10834 7282 11082 7344
rect 13068 7730 13248 7812
rect 13068 7670 13130 7730
rect 13190 7670 13248 7730
rect 13068 7344 13248 7670
rect 15234 7812 15482 7874
rect 13454 7740 13470 7774
rect 15046 7740 15062 7774
rect 13386 7712 13420 7728
rect 13386 7428 13420 7444
rect 15096 7712 15130 7728
rect 15096 7428 15130 7444
rect 13454 7382 13470 7416
rect 15046 7382 15062 7416
rect 13034 7282 13282 7344
rect 15268 7730 15448 7812
rect 15268 7670 15330 7730
rect 15390 7670 15448 7730
rect 15268 7344 15448 7670
rect 17434 7812 17682 7874
rect 15654 7740 15670 7774
rect 17246 7740 17262 7774
rect 15586 7712 15620 7728
rect 15586 7428 15620 7444
rect 17296 7712 17330 7728
rect 17296 7428 17330 7444
rect 15654 7382 15670 7416
rect 17246 7382 17262 7416
rect 15234 7282 15482 7344
rect 17468 7730 17648 7812
rect 17468 7670 17530 7730
rect 17590 7670 17648 7730
rect 17468 7344 17648 7670
rect 19634 7813 19883 7874
rect 19634 7812 19849 7813
rect 17854 7740 17870 7774
rect 19446 7740 19462 7774
rect 17786 7712 17820 7728
rect 17786 7428 17820 7444
rect 19496 7712 19530 7728
rect 19496 7428 19530 7444
rect 17854 7382 17870 7416
rect 19446 7382 19462 7416
rect 17434 7282 17682 7344
rect 19668 7730 19849 7812
rect 19668 7670 19730 7730
rect 19790 7670 19849 7730
rect 19668 7345 19849 7670
rect 20100 7775 20300 7875
rect 20760 7775 20960 7875
rect 21420 7775 21620 7875
rect 21835 7813 22236 7875
rect 20055 7741 20071 7775
rect 21647 7741 21663 7775
rect 19987 7713 20021 7729
rect 19883 7520 19987 7620
rect 19987 7429 20021 7445
rect 21697 7713 21731 7729
rect 21731 7520 21835 7620
rect 21697 7429 21731 7445
rect 20055 7383 20071 7417
rect 21647 7383 21663 7417
rect 19668 7344 19883 7345
rect 19634 7283 19883 7344
rect 20080 7283 20280 7383
rect 20760 7283 20960 7383
rect 21420 7283 21620 7383
rect 21869 7730 22236 7813
rect 21869 7670 21930 7730
rect 21990 7670 22236 7730
rect 21869 7345 22236 7670
rect 21835 7283 22236 7345
rect 19634 7282 19945 7283
rect 1973 7249 2344 7282
rect -300 7248 2344 7249
rect 4172 7248 4544 7282
rect 6372 7248 6744 7282
rect 8572 7248 8944 7282
rect 10772 7248 11144 7282
rect 12972 7248 13344 7282
rect 15172 7248 15544 7282
rect 17372 7248 17744 7282
rect 19572 7249 19945 7282
rect 21773 7249 22236 7283
rect 19572 7248 22236 7249
rect -300 7109 22236 7248
rect -300 7075 145 7109
rect 1973 7108 19945 7109
rect 1973 7075 2344 7108
rect -300 7013 83 7075
rect -300 6930 49 7013
rect -300 6870 -70 6930
rect -10 6870 49 6930
rect -300 6545 49 6870
rect 300 6975 500 7075
rect 960 6975 1160 7075
rect 1620 6975 1820 7075
rect 2035 7074 2344 7075
rect 4172 7074 4544 7108
rect 6372 7074 6744 7108
rect 8572 7074 8944 7108
rect 10772 7074 11144 7108
rect 12972 7074 13344 7108
rect 15172 7074 15544 7108
rect 17372 7074 17744 7108
rect 19572 7075 19945 7108
rect 21773 7075 22236 7109
rect 19572 7074 19883 7075
rect 2035 7013 2282 7074
rect 255 6941 271 6975
rect 1847 6941 1863 6975
rect 187 6913 221 6929
rect 83 6720 187 6820
rect 187 6629 221 6645
rect 1897 6913 1931 6929
rect 1931 6720 2035 6820
rect 1897 6629 1931 6645
rect 255 6583 271 6617
rect 1847 6583 1863 6617
rect -300 6483 83 6545
rect 280 6483 480 6583
rect 960 6483 1160 6583
rect 1620 6483 1820 6583
rect 2069 7012 2282 7013
rect 2069 6930 2248 7012
rect 2069 6870 2130 6930
rect 2190 6870 2248 6930
rect 2069 6545 2248 6870
rect 2035 6544 2248 6545
rect 4234 7012 4482 7074
rect 2454 6940 2470 6974
rect 4046 6940 4062 6974
rect 2386 6912 2420 6928
rect 2386 6628 2420 6644
rect 4096 6912 4130 6928
rect 4096 6628 4130 6644
rect 2454 6582 2470 6616
rect 4046 6582 4062 6616
rect 2035 6483 2282 6544
rect -300 6449 145 6483
rect 1973 6482 2282 6483
rect 4268 6930 4448 7012
rect 4268 6870 4330 6930
rect 4390 6870 4448 6930
rect 4268 6544 4448 6870
rect 6434 7012 6682 7074
rect 4654 6940 4670 6974
rect 6246 6940 6262 6974
rect 4586 6912 4620 6928
rect 4586 6628 4620 6644
rect 6296 6912 6330 6928
rect 6296 6628 6330 6644
rect 4654 6582 4670 6616
rect 6246 6582 6262 6616
rect 4234 6482 4482 6544
rect 6468 6930 6648 7012
rect 6468 6870 6530 6930
rect 6590 6870 6648 6930
rect 6468 6544 6648 6870
rect 8634 7012 8882 7074
rect 6854 6940 6870 6974
rect 8446 6940 8462 6974
rect 6786 6912 6820 6928
rect 6786 6628 6820 6644
rect 8496 6912 8530 6928
rect 8496 6628 8530 6644
rect 6854 6582 6870 6616
rect 8446 6582 8462 6616
rect 6434 6482 6682 6544
rect 8668 6930 8848 7012
rect 8668 6870 8730 6930
rect 8790 6870 8848 6930
rect 8668 6544 8848 6870
rect 10834 7012 11082 7074
rect 9054 6940 9070 6974
rect 10646 6940 10662 6974
rect 8986 6912 9020 6928
rect 8986 6628 9020 6644
rect 10696 6912 10730 6928
rect 10696 6628 10730 6644
rect 9054 6582 9070 6616
rect 10646 6582 10662 6616
rect 8634 6482 8882 6544
rect 10868 6930 11048 7012
rect 10868 6870 10930 6930
rect 10990 6870 11048 6930
rect 10868 6544 11048 6870
rect 13034 7012 13282 7074
rect 11254 6940 11270 6974
rect 12846 6940 12862 6974
rect 11186 6912 11220 6928
rect 11186 6628 11220 6644
rect 12896 6912 12930 6928
rect 12896 6628 12930 6644
rect 11254 6582 11270 6616
rect 12846 6582 12862 6616
rect 10834 6482 11082 6544
rect 13068 6930 13248 7012
rect 13068 6870 13130 6930
rect 13190 6870 13248 6930
rect 13068 6544 13248 6870
rect 15234 7012 15482 7074
rect 13454 6940 13470 6974
rect 15046 6940 15062 6974
rect 13386 6912 13420 6928
rect 13386 6628 13420 6644
rect 15096 6912 15130 6928
rect 15096 6628 15130 6644
rect 13454 6582 13470 6616
rect 15046 6582 15062 6616
rect 13034 6482 13282 6544
rect 15268 6930 15448 7012
rect 15268 6870 15330 6930
rect 15390 6870 15448 6930
rect 15268 6544 15448 6870
rect 17434 7012 17682 7074
rect 15654 6940 15670 6974
rect 17246 6940 17262 6974
rect 15586 6912 15620 6928
rect 15586 6628 15620 6644
rect 17296 6912 17330 6928
rect 17296 6628 17330 6644
rect 15654 6582 15670 6616
rect 17246 6582 17262 6616
rect 15234 6482 15482 6544
rect 17468 6930 17648 7012
rect 17468 6870 17530 6930
rect 17590 6870 17648 6930
rect 17468 6544 17648 6870
rect 19634 7013 19883 7074
rect 19634 7012 19849 7013
rect 17854 6940 17870 6974
rect 19446 6940 19462 6974
rect 17786 6912 17820 6928
rect 17786 6628 17820 6644
rect 19496 6912 19530 6928
rect 19496 6628 19530 6644
rect 17854 6582 17870 6616
rect 19446 6582 19462 6616
rect 17434 6482 17682 6544
rect 19668 6930 19849 7012
rect 19668 6870 19730 6930
rect 19790 6870 19849 6930
rect 19668 6545 19849 6870
rect 20100 6975 20300 7075
rect 20760 6975 20960 7075
rect 21420 6975 21620 7075
rect 21835 7013 22236 7075
rect 20055 6941 20071 6975
rect 21647 6941 21663 6975
rect 19987 6913 20021 6929
rect 19883 6720 19987 6820
rect 19987 6629 20021 6645
rect 21697 6913 21731 6929
rect 21731 6720 21835 6820
rect 21697 6629 21731 6645
rect 20055 6583 20071 6617
rect 21647 6583 21663 6617
rect 19668 6544 19883 6545
rect 19634 6483 19883 6544
rect 20080 6483 20280 6583
rect 20760 6483 20960 6583
rect 21420 6483 21620 6583
rect 21869 6930 22236 7013
rect 21869 6870 21930 6930
rect 21990 6870 22236 6930
rect 21869 6545 22236 6870
rect 21835 6483 22236 6545
rect 19634 6482 19945 6483
rect 1973 6449 2344 6482
rect -300 6448 2344 6449
rect 4172 6448 4544 6482
rect 6372 6448 6744 6482
rect 8572 6448 8944 6482
rect 10772 6448 11144 6482
rect 12972 6448 13344 6482
rect 15172 6448 15544 6482
rect 17372 6448 17744 6482
rect 19572 6449 19945 6482
rect 21773 6449 22236 6483
rect 19572 6448 22236 6449
rect -300 6309 22236 6448
rect -300 6275 145 6309
rect 1973 6308 19945 6309
rect 1973 6275 2344 6308
rect -300 6213 83 6275
rect -300 6130 49 6213
rect -300 6070 -70 6130
rect -10 6070 49 6130
rect -300 5745 49 6070
rect 300 6175 500 6275
rect 960 6175 1160 6275
rect 1620 6175 1820 6275
rect 2035 6274 2344 6275
rect 4172 6274 4544 6308
rect 6372 6274 6744 6308
rect 8572 6274 8944 6308
rect 10772 6274 11144 6308
rect 12972 6274 13344 6308
rect 15172 6274 15544 6308
rect 17372 6274 17744 6308
rect 19572 6275 19945 6308
rect 21773 6275 22236 6309
rect 19572 6274 19883 6275
rect 2035 6213 2282 6274
rect 255 6141 271 6175
rect 1847 6141 1863 6175
rect 187 6113 221 6129
rect 83 5920 187 6020
rect 187 5829 221 5845
rect 1897 6113 1931 6129
rect 1931 5920 2035 6020
rect 1897 5829 1931 5845
rect 255 5783 271 5817
rect 1847 5783 1863 5817
rect -300 5683 83 5745
rect 280 5683 480 5783
rect 960 5683 1160 5783
rect 1620 5683 1820 5783
rect 2069 6212 2282 6213
rect 2069 6130 2248 6212
rect 2069 6070 2130 6130
rect 2190 6070 2248 6130
rect 2069 5745 2248 6070
rect 2035 5744 2248 5745
rect 4234 6212 4482 6274
rect 2454 6140 2470 6174
rect 4046 6140 4062 6174
rect 2386 6112 2420 6128
rect 2386 5828 2420 5844
rect 4096 6112 4130 6128
rect 4096 5828 4130 5844
rect 2454 5782 2470 5816
rect 4046 5782 4062 5816
rect 2035 5683 2282 5744
rect -300 5649 145 5683
rect 1973 5682 2282 5683
rect 4268 6130 4448 6212
rect 4268 6070 4330 6130
rect 4390 6070 4448 6130
rect 4268 5744 4448 6070
rect 6434 6212 6682 6274
rect 4654 6140 4670 6174
rect 6246 6140 6262 6174
rect 4586 6112 4620 6128
rect 4586 5828 4620 5844
rect 6296 6112 6330 6128
rect 6296 5828 6330 5844
rect 4654 5782 4670 5816
rect 6246 5782 6262 5816
rect 4234 5682 4482 5744
rect 6468 6130 6648 6212
rect 6468 6070 6530 6130
rect 6590 6070 6648 6130
rect 6468 5744 6648 6070
rect 8634 6212 8882 6274
rect 6854 6140 6870 6174
rect 8446 6140 8462 6174
rect 6786 6112 6820 6128
rect 6786 5828 6820 5844
rect 8496 6112 8530 6128
rect 8496 5828 8530 5844
rect 6854 5782 6870 5816
rect 8446 5782 8462 5816
rect 6434 5682 6682 5744
rect 8668 6130 8848 6212
rect 8668 6070 8730 6130
rect 8790 6070 8848 6130
rect 8668 5744 8848 6070
rect 10834 6212 11082 6274
rect 9054 6140 9070 6174
rect 10646 6140 10662 6174
rect 8986 6112 9020 6128
rect 8986 5828 9020 5844
rect 10696 6112 10730 6128
rect 10696 5828 10730 5844
rect 9054 5782 9070 5816
rect 10646 5782 10662 5816
rect 8634 5682 8882 5744
rect 10868 6130 11048 6212
rect 10868 6070 10930 6130
rect 10990 6070 11048 6130
rect 10868 5744 11048 6070
rect 13034 6212 13282 6274
rect 11254 6140 11270 6174
rect 12846 6140 12862 6174
rect 11186 6112 11220 6128
rect 11186 5828 11220 5844
rect 12896 6112 12930 6128
rect 12896 5828 12930 5844
rect 11254 5782 11270 5816
rect 12846 5782 12862 5816
rect 10834 5682 11082 5744
rect 13068 6130 13248 6212
rect 13068 6070 13130 6130
rect 13190 6070 13248 6130
rect 13068 5744 13248 6070
rect 15234 6212 15482 6274
rect 13454 6140 13470 6174
rect 15046 6140 15062 6174
rect 13386 6112 13420 6128
rect 13386 5828 13420 5844
rect 15096 6112 15130 6128
rect 15096 5828 15130 5844
rect 13454 5782 13470 5816
rect 15046 5782 15062 5816
rect 13034 5682 13282 5744
rect 15268 6130 15448 6212
rect 15268 6070 15330 6130
rect 15390 6070 15448 6130
rect 15268 5744 15448 6070
rect 17434 6212 17682 6274
rect 15654 6140 15670 6174
rect 17246 6140 17262 6174
rect 15586 6112 15620 6128
rect 15586 5828 15620 5844
rect 17296 6112 17330 6128
rect 17296 5828 17330 5844
rect 15654 5782 15670 5816
rect 17246 5782 17262 5816
rect 15234 5682 15482 5744
rect 17468 6130 17648 6212
rect 17468 6070 17530 6130
rect 17590 6070 17648 6130
rect 17468 5744 17648 6070
rect 19634 6213 19883 6274
rect 19634 6212 19849 6213
rect 17854 6140 17870 6174
rect 19446 6140 19462 6174
rect 17786 6112 17820 6128
rect 17786 5828 17820 5844
rect 19496 6112 19530 6128
rect 19496 5828 19530 5844
rect 17854 5782 17870 5816
rect 19446 5782 19462 5816
rect 17434 5682 17682 5744
rect 19668 6130 19849 6212
rect 19668 6070 19730 6130
rect 19790 6070 19849 6130
rect 19668 5745 19849 6070
rect 20100 6175 20300 6275
rect 20760 6175 20960 6275
rect 21420 6175 21620 6275
rect 21835 6213 22236 6275
rect 20055 6141 20071 6175
rect 21647 6141 21663 6175
rect 19987 6113 20021 6129
rect 19883 5920 19987 6020
rect 19987 5829 20021 5845
rect 21697 6113 21731 6129
rect 21731 5920 21835 6020
rect 21697 5829 21731 5845
rect 20055 5783 20071 5817
rect 21647 5783 21663 5817
rect 19668 5744 19883 5745
rect 19634 5683 19883 5744
rect 20080 5683 20280 5783
rect 20760 5683 20960 5783
rect 21420 5683 21620 5783
rect 21869 6130 22236 6213
rect 21869 6070 21930 6130
rect 21990 6070 22236 6130
rect 21869 5745 22236 6070
rect 21835 5683 22236 5745
rect 19634 5682 19945 5683
rect 1973 5649 2344 5682
rect -300 5648 2344 5649
rect 4172 5648 4544 5682
rect 6372 5648 6744 5682
rect 8572 5648 8944 5682
rect 10772 5648 11144 5682
rect 12972 5648 13344 5682
rect 15172 5648 15544 5682
rect 17372 5648 17744 5682
rect 19572 5649 19945 5682
rect 21773 5649 22236 5683
rect 19572 5648 22236 5649
rect -300 5509 22236 5648
rect -300 5475 145 5509
rect 1973 5508 19945 5509
rect 1973 5475 2344 5508
rect -300 5413 83 5475
rect -300 5330 49 5413
rect -300 5270 -70 5330
rect -10 5270 49 5330
rect -300 4945 49 5270
rect 300 5375 500 5475
rect 960 5375 1160 5475
rect 1620 5375 1820 5475
rect 2035 5474 2344 5475
rect 4172 5474 4544 5508
rect 6372 5474 6744 5508
rect 8572 5474 8944 5508
rect 10772 5474 11144 5508
rect 12972 5474 13344 5508
rect 15172 5474 15544 5508
rect 17372 5474 17744 5508
rect 19572 5475 19945 5508
rect 21773 5475 22236 5509
rect 19572 5474 19883 5475
rect 2035 5413 2282 5474
rect 255 5341 271 5375
rect 1847 5341 1863 5375
rect 187 5313 221 5329
rect 83 5120 187 5220
rect 187 5029 221 5045
rect 1897 5313 1931 5329
rect 1931 5120 2035 5220
rect 1897 5029 1931 5045
rect 255 4983 271 5017
rect 1847 4983 1863 5017
rect -300 4883 83 4945
rect 280 4883 480 4983
rect 960 4883 1160 4983
rect 1620 4883 1820 4983
rect 2069 5412 2282 5413
rect 2069 5330 2248 5412
rect 2069 5270 2130 5330
rect 2190 5270 2248 5330
rect 2069 4945 2248 5270
rect 2035 4944 2248 4945
rect 4234 5412 4482 5474
rect 2454 5340 2470 5374
rect 4046 5340 4062 5374
rect 2386 5312 2420 5328
rect 2386 5028 2420 5044
rect 4096 5312 4130 5328
rect 4096 5028 4130 5044
rect 2454 4982 2470 5016
rect 4046 4982 4062 5016
rect 2035 4883 2282 4944
rect -300 4849 145 4883
rect 1973 4882 2282 4883
rect 4268 5330 4448 5412
rect 4268 5270 4330 5330
rect 4390 5270 4448 5330
rect 4268 4944 4448 5270
rect 6434 5412 6682 5474
rect 4654 5340 4670 5374
rect 6246 5340 6262 5374
rect 4586 5312 4620 5328
rect 4586 5028 4620 5044
rect 6296 5312 6330 5328
rect 6296 5028 6330 5044
rect 4654 4982 4670 5016
rect 6246 4982 6262 5016
rect 4234 4882 4482 4944
rect 6468 5330 6648 5412
rect 6468 5270 6530 5330
rect 6590 5270 6648 5330
rect 6468 4944 6648 5270
rect 8634 5412 8882 5474
rect 6854 5340 6870 5374
rect 8446 5340 8462 5374
rect 6786 5312 6820 5328
rect 6786 5028 6820 5044
rect 8496 5312 8530 5328
rect 8496 5028 8530 5044
rect 6854 4982 6870 5016
rect 8446 4982 8462 5016
rect 6434 4882 6682 4944
rect 8668 5330 8848 5412
rect 8668 5270 8730 5330
rect 8790 5270 8848 5330
rect 8668 4944 8848 5270
rect 10834 5412 11082 5474
rect 9054 5340 9070 5374
rect 10646 5340 10662 5374
rect 8986 5312 9020 5328
rect 8986 5028 9020 5044
rect 10696 5312 10730 5328
rect 10696 5028 10730 5044
rect 9054 4982 9070 5016
rect 10646 4982 10662 5016
rect 8634 4882 8882 4944
rect 10868 5330 11048 5412
rect 10868 5270 10930 5330
rect 10990 5270 11048 5330
rect 10868 4944 11048 5270
rect 13034 5412 13282 5474
rect 11254 5340 11270 5374
rect 12846 5340 12862 5374
rect 11186 5312 11220 5328
rect 11186 5028 11220 5044
rect 12896 5312 12930 5328
rect 12896 5028 12930 5044
rect 11254 4982 11270 5016
rect 12846 4982 12862 5016
rect 10834 4882 11082 4944
rect 13068 5330 13248 5412
rect 13068 5270 13130 5330
rect 13190 5270 13248 5330
rect 13068 4944 13248 5270
rect 15234 5412 15482 5474
rect 13454 5340 13470 5374
rect 15046 5340 15062 5374
rect 13386 5312 13420 5328
rect 13386 5028 13420 5044
rect 15096 5312 15130 5328
rect 15096 5028 15130 5044
rect 13454 4982 13470 5016
rect 15046 4982 15062 5016
rect 13034 4882 13282 4944
rect 15268 5330 15448 5412
rect 15268 5270 15330 5330
rect 15390 5270 15448 5330
rect 15268 4944 15448 5270
rect 17434 5412 17682 5474
rect 15654 5340 15670 5374
rect 17246 5340 17262 5374
rect 15586 5312 15620 5328
rect 15586 5028 15620 5044
rect 17296 5312 17330 5328
rect 17296 5028 17330 5044
rect 15654 4982 15670 5016
rect 17246 4982 17262 5016
rect 15234 4882 15482 4944
rect 17468 5330 17648 5412
rect 17468 5270 17530 5330
rect 17590 5270 17648 5330
rect 17468 4944 17648 5270
rect 19634 5413 19883 5474
rect 19634 5412 19849 5413
rect 17854 5340 17870 5374
rect 19446 5340 19462 5374
rect 17786 5312 17820 5328
rect 17786 5028 17820 5044
rect 19496 5312 19530 5328
rect 19496 5028 19530 5044
rect 17854 4982 17870 5016
rect 19446 4982 19462 5016
rect 17434 4882 17682 4944
rect 19668 5330 19849 5412
rect 19668 5270 19730 5330
rect 19790 5270 19849 5330
rect 19668 4945 19849 5270
rect 20100 5375 20300 5475
rect 20760 5375 20960 5475
rect 21420 5375 21620 5475
rect 21835 5413 22236 5475
rect 20055 5341 20071 5375
rect 21647 5341 21663 5375
rect 19987 5313 20021 5329
rect 19883 5120 19987 5220
rect 19987 5029 20021 5045
rect 21697 5313 21731 5329
rect 21731 5120 21835 5220
rect 21697 5029 21731 5045
rect 20055 4983 20071 5017
rect 21647 4983 21663 5017
rect 19668 4944 19883 4945
rect 19634 4883 19883 4944
rect 20080 4883 20280 4983
rect 20760 4883 20960 4983
rect 21420 4883 21620 4983
rect 21869 5330 22236 5413
rect 21869 5270 21930 5330
rect 21990 5270 22236 5330
rect 21869 4945 22236 5270
rect 21835 4883 22236 4945
rect 19634 4882 19945 4883
rect 1973 4849 2344 4882
rect -300 4848 2344 4849
rect 4172 4848 4544 4882
rect 6372 4848 6744 4882
rect 8572 4848 8944 4882
rect 10772 4848 11144 4882
rect 12972 4848 13344 4882
rect 15172 4848 15544 4882
rect 17372 4848 17744 4882
rect 19572 4849 19945 4882
rect 21773 4849 22236 4883
rect 19572 4848 22236 4849
rect -300 4710 22236 4848
rect 22270 11400 22366 11814
rect 26932 11400 27028 11814
rect -300 4709 8946 4710
rect -300 4675 145 4709
rect 1973 4675 2345 4709
rect 4173 4675 4545 4709
rect 6373 4675 6745 4709
rect 8573 4676 8946 4709
rect 10774 4676 11146 4710
rect 12974 4709 22236 4710
rect 12974 4676 13345 4709
rect 8573 4675 8884 4676
rect -300 4613 83 4675
rect -300 4145 49 4613
rect 300 4575 500 4675
rect 960 4575 1160 4675
rect 1620 4575 1820 4675
rect 2035 4613 2283 4675
rect 255 4541 271 4575
rect 1847 4541 1863 4575
rect 187 4513 221 4529
rect 83 4320 187 4420
rect 187 4229 221 4245
rect 1897 4513 1931 4529
rect 1931 4320 2035 4420
rect 1897 4229 1931 4245
rect 255 4183 271 4217
rect 1847 4183 1863 4217
rect -300 4083 83 4145
rect 280 4083 480 4183
rect 960 4083 1160 4183
rect 1620 4083 1820 4183
rect 2069 4145 2249 4613
rect 2500 4575 2700 4675
rect 3160 4575 3360 4675
rect 3820 4575 4020 4675
rect 4235 4613 4483 4675
rect 2455 4541 2471 4575
rect 4047 4541 4063 4575
rect 2387 4513 2421 4529
rect 2283 4320 2387 4420
rect 2387 4229 2421 4245
rect 4097 4513 4131 4529
rect 4131 4320 4235 4420
rect 4097 4229 4131 4245
rect 2455 4183 2471 4217
rect 4047 4183 4063 4217
rect 2035 4083 2283 4145
rect 2480 4083 2680 4183
rect 3160 4083 3360 4183
rect 3820 4083 4020 4183
rect 4269 4145 4449 4613
rect 4700 4575 4900 4675
rect 5360 4575 5560 4675
rect 6020 4575 6220 4675
rect 6435 4613 6683 4675
rect 4655 4541 4671 4575
rect 6247 4541 6263 4575
rect 4587 4513 4621 4529
rect 4483 4320 4587 4420
rect 4587 4229 4621 4245
rect 6297 4513 6331 4529
rect 6331 4320 6435 4420
rect 6297 4229 6331 4245
rect 4655 4183 4671 4217
rect 6247 4183 6263 4217
rect 4235 4083 4483 4145
rect 4680 4083 4880 4183
rect 5360 4083 5560 4183
rect 6020 4083 6220 4183
rect 6469 4145 6649 4613
rect 6900 4575 7100 4675
rect 7560 4575 7760 4675
rect 8220 4575 8420 4675
rect 8635 4614 8884 4675
rect 8635 4613 8850 4614
rect 6855 4541 6871 4575
rect 8447 4541 8463 4575
rect 6787 4513 6821 4529
rect 6683 4320 6787 4420
rect 6787 4229 6821 4245
rect 8497 4513 8531 4529
rect 8531 4320 8635 4420
rect 8497 4229 8531 4245
rect 6855 4183 6871 4217
rect 8447 4183 8463 4217
rect 6435 4083 6683 4145
rect 6880 4083 7080 4183
rect 7560 4083 7760 4183
rect 8220 4083 8420 4183
rect 8669 4146 8850 4613
rect 10836 4614 11084 4676
rect 9056 4542 9072 4576
rect 10648 4542 10664 4576
rect 8988 4514 9022 4530
rect 8988 4230 9022 4246
rect 10698 4514 10732 4530
rect 10698 4230 10732 4246
rect 9056 4184 9072 4218
rect 10648 4184 10664 4218
rect 8669 4145 8884 4146
rect 8635 4084 8884 4145
rect 10870 4146 11050 4614
rect 13036 4675 13345 4676
rect 15173 4675 15545 4709
rect 17373 4675 17745 4709
rect 19573 4675 19945 4709
rect 21773 4675 22236 4709
rect 13036 4614 13283 4675
rect 11256 4542 11272 4576
rect 12848 4542 12864 4576
rect 11188 4514 11222 4530
rect 11188 4230 11222 4246
rect 12898 4514 12932 4530
rect 12898 4230 12932 4246
rect 11256 4184 11272 4218
rect 12848 4184 12864 4218
rect 10836 4084 11084 4146
rect 13070 4613 13283 4614
rect 13070 4146 13249 4613
rect 13036 4145 13249 4146
rect 13500 4575 13700 4675
rect 14160 4575 14360 4675
rect 14820 4575 15020 4675
rect 15235 4613 15483 4675
rect 13455 4541 13471 4575
rect 15047 4541 15063 4575
rect 13387 4513 13421 4529
rect 13283 4320 13387 4420
rect 13387 4229 13421 4245
rect 15097 4513 15131 4529
rect 15131 4320 15235 4420
rect 15097 4229 15131 4245
rect 13455 4183 13471 4217
rect 15047 4183 15063 4217
rect 13036 4084 13283 4145
rect 8635 4083 8946 4084
rect -300 4049 145 4083
rect 1973 4049 2345 4083
rect 4173 4049 4545 4083
rect 6373 4049 6745 4083
rect 8573 4050 8946 4083
rect 10774 4050 11146 4084
rect 12974 4083 13283 4084
rect 13480 4083 13680 4183
rect 14160 4083 14360 4183
rect 14820 4083 15020 4183
rect 15269 4145 15449 4613
rect 15700 4575 15900 4675
rect 16360 4575 16560 4675
rect 17020 4575 17220 4675
rect 17435 4613 17683 4675
rect 15655 4541 15671 4575
rect 17247 4541 17263 4575
rect 15587 4513 15621 4529
rect 15483 4320 15587 4420
rect 15587 4229 15621 4245
rect 17297 4513 17331 4529
rect 17331 4320 17435 4420
rect 17297 4229 17331 4245
rect 15655 4183 15671 4217
rect 17247 4183 17263 4217
rect 15235 4083 15483 4145
rect 15680 4083 15880 4183
rect 16360 4083 16560 4183
rect 17020 4083 17220 4183
rect 17469 4145 17649 4613
rect 17900 4575 18100 4675
rect 18560 4575 18760 4675
rect 19220 4575 19420 4675
rect 19635 4613 19883 4675
rect 17855 4541 17871 4575
rect 19447 4541 19463 4575
rect 17787 4513 17821 4529
rect 17683 4320 17787 4420
rect 17787 4229 17821 4245
rect 19497 4513 19531 4529
rect 19531 4320 19635 4420
rect 19497 4229 19531 4245
rect 17855 4183 17871 4217
rect 19447 4183 19463 4217
rect 17435 4083 17683 4145
rect 17880 4083 18080 4183
rect 18560 4083 18760 4183
rect 19220 4083 19420 4183
rect 19669 4145 19849 4613
rect 20100 4575 20300 4675
rect 20760 4575 20960 4675
rect 21420 4575 21620 4675
rect 21835 4613 22236 4675
rect 20055 4541 20071 4575
rect 21647 4541 21663 4575
rect 19987 4513 20021 4529
rect 19883 4320 19987 4420
rect 19987 4229 20021 4245
rect 21697 4513 21731 4529
rect 21731 4320 21835 4420
rect 21697 4229 21731 4245
rect 20055 4183 20071 4217
rect 21647 4183 21663 4217
rect 19635 4083 19883 4145
rect 20080 4083 20280 4183
rect 20760 4083 20960 4183
rect 21420 4083 21620 4183
rect 21869 4532 22236 4613
rect 22270 4566 22366 4980
rect 26932 4566 27028 4980
rect 22270 4532 22920 4566
rect 21869 4470 22920 4532
rect 26380 4532 27028 4566
rect 27062 4532 27280 11848
rect 29968 11903 30064 11920
rect 30648 11903 30757 11937
rect 31149 11903 31236 11937
rect 31550 11903 31637 11937
rect 32029 11920 32264 11937
rect 29968 11841 30002 11903
rect 27778 11558 27874 11592
rect 28850 11570 28946 11592
rect 28850 11558 29150 11570
rect 27778 11496 27812 11558
rect 28910 11496 29150 11558
rect 27922 11424 27938 11458
rect 28714 11424 28730 11458
rect 28773 11396 28807 11412
rect 28773 11312 28807 11328
rect 27922 11266 27938 11300
rect 28714 11266 28730 11300
rect 28773 11238 28807 11254
rect 28773 11154 28807 11170
rect 27922 11108 27938 11142
rect 28714 11108 28730 11142
rect 28773 11080 28807 11096
rect 28773 10996 28807 11012
rect 27922 10950 27938 10984
rect 28714 10950 28730 10984
rect 28773 10922 28807 10938
rect 28773 10838 28807 10854
rect 27922 10792 27938 10826
rect 28714 10792 28730 10826
rect 27778 10692 27812 10754
rect 28910 10754 28912 11496
rect 28946 10754 29150 11496
rect 30710 11848 30757 11903
rect 30148 11765 30164 11799
rect 30232 11765 30248 11799
rect 30306 11765 30322 11799
rect 30390 11765 30406 11799
rect 30464 11765 30480 11799
rect 30548 11765 30564 11799
rect 30102 11715 30136 11731
rect 30102 11523 30136 11539
rect 30260 11715 30294 11731
rect 30260 11523 30294 11539
rect 30418 11715 30452 11731
rect 30418 11523 30452 11539
rect 30576 11715 30610 11731
rect 30576 11523 30610 11539
rect 30148 11455 30164 11489
rect 30232 11455 30248 11489
rect 30306 11455 30322 11489
rect 30390 11455 30406 11489
rect 30464 11455 30480 11489
rect 30548 11455 30564 11489
rect 29968 11351 30002 11413
rect 30744 11406 30757 11848
rect 30903 11765 30919 11799
rect 30987 11765 31003 11799
rect 30857 11715 30891 11731
rect 30857 11523 30891 11539
rect 31015 11715 31049 11731
rect 31015 11523 31049 11539
rect 30903 11455 30919 11489
rect 30987 11455 31003 11489
rect 30710 11351 30757 11406
rect 31149 11351 31197 11903
rect 31589 11848 31637 11903
rect 31623 11841 31637 11848
rect 31343 11765 31359 11799
rect 31427 11765 31443 11799
rect 31297 11715 31331 11731
rect 31297 11523 31331 11539
rect 31455 11715 31489 11731
rect 31455 11523 31489 11539
rect 31343 11455 31359 11489
rect 31427 11455 31443 11489
rect 32029 11841 32063 11920
rect 31783 11765 31799 11799
rect 31867 11765 31883 11799
rect 31737 11715 31771 11731
rect 31737 11523 31771 11539
rect 31895 11715 31929 11731
rect 31895 11523 31929 11539
rect 31783 11455 31799 11489
rect 31867 11455 31883 11489
rect 31623 11406 31637 11413
rect 31589 11351 31637 11406
rect 32029 11351 32063 11413
rect 29968 11317 30064 11351
rect 30648 11317 30819 11351
rect 31087 11317 31259 11351
rect 31527 11317 31699 11351
rect 31967 11317 32063 11351
rect 32168 11903 32264 11920
rect 32848 11903 32957 11937
rect 33349 11903 33436 11937
rect 33750 11903 33837 11937
rect 34229 11920 34464 11937
rect 32168 11841 32202 11903
rect 32910 11848 32957 11903
rect 32348 11765 32364 11799
rect 32432 11765 32448 11799
rect 32506 11765 32522 11799
rect 32590 11765 32606 11799
rect 32664 11765 32680 11799
rect 32748 11765 32764 11799
rect 32302 11715 32336 11731
rect 32302 11523 32336 11539
rect 32460 11715 32494 11731
rect 32460 11523 32494 11539
rect 32618 11715 32652 11731
rect 32618 11523 32652 11539
rect 32776 11715 32810 11731
rect 32776 11523 32810 11539
rect 32348 11455 32364 11489
rect 32432 11455 32448 11489
rect 32506 11455 32522 11489
rect 32590 11455 32606 11489
rect 32664 11455 32680 11489
rect 32748 11455 32764 11489
rect 32168 11351 32202 11413
rect 32944 11406 32957 11848
rect 33103 11765 33119 11799
rect 33187 11765 33203 11799
rect 33057 11715 33091 11731
rect 33057 11523 33091 11539
rect 33215 11715 33249 11731
rect 33215 11523 33249 11539
rect 33103 11455 33119 11489
rect 33187 11455 33203 11489
rect 32910 11351 32957 11406
rect 33349 11351 33397 11903
rect 33789 11848 33837 11903
rect 33823 11841 33837 11848
rect 33543 11765 33559 11799
rect 33627 11765 33643 11799
rect 33497 11715 33531 11731
rect 33497 11523 33531 11539
rect 33655 11715 33689 11731
rect 33655 11523 33689 11539
rect 33543 11455 33559 11489
rect 33627 11455 33643 11489
rect 34229 11841 34263 11920
rect 33983 11765 33999 11799
rect 34067 11765 34083 11799
rect 33937 11715 33971 11731
rect 33937 11523 33971 11539
rect 34095 11715 34129 11731
rect 34095 11523 34129 11539
rect 33983 11455 33999 11489
rect 34067 11455 34083 11489
rect 33823 11406 33837 11413
rect 33789 11351 33837 11406
rect 34229 11351 34263 11413
rect 32168 11317 32264 11351
rect 32848 11317 33019 11351
rect 33287 11317 33459 11351
rect 33727 11317 33899 11351
rect 34167 11317 34263 11351
rect 34368 11903 34464 11920
rect 35048 11903 35157 11937
rect 35549 11903 35636 11937
rect 35950 11903 36037 11937
rect 34368 11841 34402 11903
rect 35110 11848 35157 11903
rect 34548 11765 34564 11799
rect 34632 11765 34648 11799
rect 34706 11765 34722 11799
rect 34790 11765 34806 11799
rect 34864 11765 34880 11799
rect 34948 11765 34964 11799
rect 34502 11715 34536 11731
rect 34502 11523 34536 11539
rect 34660 11715 34694 11731
rect 34660 11523 34694 11539
rect 34818 11715 34852 11731
rect 34818 11523 34852 11539
rect 34976 11715 35010 11731
rect 34976 11523 35010 11539
rect 34548 11455 34564 11489
rect 34632 11455 34648 11489
rect 34706 11455 34722 11489
rect 34790 11455 34806 11489
rect 34864 11455 34880 11489
rect 34948 11455 34964 11489
rect 34368 11351 34402 11413
rect 35144 11406 35157 11848
rect 35303 11765 35319 11799
rect 35387 11765 35403 11799
rect 35257 11715 35291 11731
rect 35257 11523 35291 11539
rect 35415 11715 35449 11731
rect 35415 11523 35449 11539
rect 35303 11455 35319 11489
rect 35387 11455 35403 11489
rect 35110 11351 35157 11406
rect 35549 11351 35597 11903
rect 35989 11848 36037 11903
rect 36023 11841 36037 11848
rect 35743 11765 35759 11799
rect 35827 11765 35843 11799
rect 35697 11715 35731 11731
rect 35697 11523 35731 11539
rect 35855 11715 35889 11731
rect 35855 11523 35889 11539
rect 35743 11455 35759 11489
rect 35827 11455 35843 11489
rect 36429 11841 36840 11937
rect 36183 11765 36199 11799
rect 36267 11765 36283 11799
rect 36137 11715 36171 11731
rect 36137 11523 36171 11539
rect 36295 11715 36329 11731
rect 36295 11523 36329 11539
rect 36183 11455 36199 11489
rect 36267 11455 36283 11489
rect 36023 11406 36037 11413
rect 35989 11351 36037 11406
rect 36463 11413 36840 11841
rect 36429 11351 36840 11413
rect 34368 11317 34464 11351
rect 35048 11317 35219 11351
rect 35487 11317 35659 11351
rect 35927 11317 36099 11351
rect 36367 11320 36840 11351
rect 36367 11317 36463 11320
rect 28910 10692 29150 10754
rect 27778 10658 27874 10692
rect 28850 10658 29150 10692
rect 28910 10552 29150 10658
rect 30010 11092 30106 11126
rect 30674 11092 30820 11126
rect 31088 11092 31260 11126
rect 31528 11092 31700 11126
rect 31968 11092 32064 11126
rect 30010 11030 30044 11092
rect 30724 11045 30770 11092
rect 30190 10954 30206 10988
rect 30574 10954 30590 10988
rect 30144 10895 30178 10911
rect 30144 10803 30178 10819
rect 30602 10895 30636 10911
rect 30602 10803 30636 10819
rect 30190 10726 30206 10760
rect 30574 10726 30590 10760
rect 30010 10622 30044 10684
rect 30724 10669 30736 11045
rect 30904 10954 30920 10988
rect 30988 10954 31004 10988
rect 30724 10622 30770 10669
rect 30010 10588 30106 10622
rect 30674 10588 30770 10622
rect 30858 10895 30892 10911
rect 27778 10518 27874 10552
rect 28850 10518 29150 10552
rect 27778 10456 27812 10518
rect 28910 10456 29150 10518
rect 27922 10384 27938 10418
rect 28714 10384 28730 10418
rect 28773 10356 28807 10372
rect 28773 10272 28807 10288
rect 27922 10226 27938 10260
rect 28714 10226 28730 10260
rect 28773 10198 28807 10214
rect 28773 10114 28807 10130
rect 27922 10068 27938 10102
rect 28714 10068 28730 10102
rect 28773 10040 28807 10056
rect 28773 9956 28807 9972
rect 27922 9910 27938 9944
rect 28714 9910 28730 9944
rect 28773 9882 28807 9898
rect 28773 9798 28807 9814
rect 27922 9752 27938 9786
rect 28714 9752 28730 9786
rect 27778 9652 27812 9714
rect 28910 9714 28912 10456
rect 28946 9790 29150 10456
rect 30724 10288 30758 10588
rect 30858 10503 30892 10519
rect 31016 10895 31050 10911
rect 31016 10503 31050 10519
rect 30904 10426 30920 10460
rect 30988 10426 31004 10460
rect 31150 10288 31198 11092
rect 31590 11030 31638 11092
rect 31344 10954 31360 10988
rect 31428 10954 31444 10988
rect 31298 10895 31332 10911
rect 31298 10503 31332 10519
rect 31456 10895 31490 10911
rect 31456 10503 31490 10519
rect 31344 10426 31360 10460
rect 31428 10426 31444 10460
rect 31590 10384 31604 11030
rect 32030 11030 32064 11092
rect 31784 10954 31800 10988
rect 31868 10954 31884 10988
rect 31738 10895 31772 10911
rect 31738 10503 31772 10519
rect 31896 10895 31930 10911
rect 31896 10503 31930 10519
rect 31784 10426 31800 10460
rect 31868 10426 31884 10460
rect 31590 10288 31638 10384
rect 32210 11092 32306 11126
rect 32874 11092 33020 11126
rect 33288 11092 33460 11126
rect 33728 11092 33900 11126
rect 34168 11092 34264 11126
rect 32210 11030 32244 11092
rect 32924 11045 32970 11092
rect 32390 10954 32406 10988
rect 32774 10954 32790 10988
rect 32344 10895 32378 10911
rect 32344 10803 32378 10819
rect 32802 10895 32836 10911
rect 32802 10803 32836 10819
rect 32390 10726 32406 10760
rect 32774 10726 32790 10760
rect 32210 10622 32244 10684
rect 32924 10669 32936 11045
rect 33104 10954 33120 10988
rect 33188 10954 33204 10988
rect 32924 10622 32970 10669
rect 32210 10588 32306 10622
rect 32874 10588 32970 10622
rect 33058 10895 33092 10911
rect 32030 10288 32064 10384
rect 32924 10288 32958 10588
rect 33058 10503 33092 10519
rect 33216 10895 33250 10911
rect 33216 10503 33250 10519
rect 33104 10426 33120 10460
rect 33188 10426 33204 10460
rect 33350 10288 33398 11092
rect 33790 11030 33838 11092
rect 33544 10954 33560 10988
rect 33628 10954 33644 10988
rect 33498 10895 33532 10911
rect 33498 10503 33532 10519
rect 33656 10895 33690 10911
rect 33656 10503 33690 10519
rect 33544 10426 33560 10460
rect 33628 10426 33644 10460
rect 33790 10384 33804 11030
rect 34230 11030 34264 11092
rect 33984 10954 34000 10988
rect 34068 10954 34084 10988
rect 33938 10895 33972 10911
rect 33938 10503 33972 10519
rect 34096 10895 34130 10911
rect 34096 10503 34130 10519
rect 33984 10426 34000 10460
rect 34068 10426 34084 10460
rect 33790 10288 33838 10384
rect 34410 11092 34506 11126
rect 35074 11092 35220 11126
rect 35488 11092 35660 11126
rect 35928 11092 36100 11126
rect 36368 11092 36464 11126
rect 34410 11030 34444 11092
rect 35124 11045 35170 11092
rect 34590 10954 34606 10988
rect 34974 10954 34990 10988
rect 34544 10895 34578 10911
rect 34544 10803 34578 10819
rect 35002 10895 35036 10911
rect 35002 10803 35036 10819
rect 34590 10726 34606 10760
rect 34974 10726 34990 10760
rect 34410 10622 34444 10684
rect 35124 10669 35136 11045
rect 35304 10954 35320 10988
rect 35388 10954 35404 10988
rect 35124 10622 35170 10669
rect 34410 10588 34506 10622
rect 35074 10588 35170 10622
rect 35258 10895 35292 10911
rect 34230 10288 34264 10384
rect 35124 10288 35158 10588
rect 35258 10503 35292 10519
rect 35416 10895 35450 10911
rect 35416 10503 35450 10519
rect 35304 10426 35320 10460
rect 35388 10426 35404 10460
rect 35550 10288 35598 11092
rect 35990 11030 36038 11092
rect 35744 10954 35760 10988
rect 35828 10954 35844 10988
rect 35698 10895 35732 10911
rect 35698 10503 35732 10519
rect 35856 10895 35890 10911
rect 35856 10503 35890 10519
rect 35744 10426 35760 10460
rect 35828 10426 35844 10460
rect 35990 10384 36004 11030
rect 36430 11030 36464 11092
rect 36184 10954 36200 10988
rect 36268 10954 36284 10988
rect 36138 10895 36172 10911
rect 36138 10503 36172 10519
rect 36296 10895 36330 10911
rect 36296 10503 36330 10519
rect 36184 10426 36200 10460
rect 36268 10426 36284 10460
rect 35990 10288 36038 10384
rect 36430 10288 36464 10384
rect 29598 9790 29694 9816
rect 28946 9782 29694 9790
rect 31520 9782 31616 9816
rect 28946 9720 29632 9782
rect 28946 9714 29598 9720
rect 28910 9652 29598 9714
rect 27778 9618 27874 9652
rect 28850 9618 29598 9652
rect 28910 9512 29598 9618
rect 31582 9720 31616 9782
rect 29778 9644 29794 9678
rect 30562 9644 30578 9678
rect 30636 9644 30652 9678
rect 31420 9644 31436 9678
rect 27778 9478 27874 9512
rect 28850 9478 29598 9512
rect 27778 9416 27812 9478
rect 28910 9416 29598 9478
rect 27922 9344 27938 9378
rect 28714 9344 28730 9378
rect 28773 9316 28807 9332
rect 28773 9232 28807 9248
rect 27922 9186 27938 9220
rect 28714 9186 28730 9220
rect 28773 9158 28807 9174
rect 28773 9074 28807 9090
rect 27922 9028 27938 9062
rect 28714 9028 28730 9062
rect 28773 9000 28807 9016
rect 28773 8916 28807 8932
rect 27922 8870 27938 8904
rect 28714 8870 28730 8904
rect 28773 8842 28807 8858
rect 28773 8758 28807 8774
rect 27922 8712 27938 8746
rect 28714 8712 28730 8746
rect 27778 8612 27812 8674
rect 28910 8674 28912 9416
rect 28946 9074 29598 9416
rect 29732 9585 29766 9601
rect 29732 9193 29766 9209
rect 30590 9585 30624 9601
rect 30590 9193 30624 9209
rect 31448 9585 31482 9601
rect 31448 9193 31482 9209
rect 29778 9116 29794 9150
rect 30562 9116 30578 9150
rect 30636 9116 30652 9150
rect 31420 9116 31436 9150
rect 28946 9012 29632 9074
rect 31582 9012 31616 9074
rect 28946 8978 29694 9012
rect 31520 8978 31616 9012
rect 28946 8812 31350 8978
rect 32796 8946 32830 9042
rect 28946 8778 29694 8812
rect 31520 8778 31616 8812
rect 28946 8716 29632 8778
rect 28946 8674 29598 8716
rect 28910 8612 29598 8674
rect 31582 8716 31616 8778
rect 29778 8640 29794 8674
rect 30562 8640 30578 8674
rect 30636 8640 30652 8674
rect 31420 8640 31436 8674
rect 27778 8578 27874 8612
rect 28850 8578 29598 8612
rect 28910 8472 29598 8578
rect 27778 8438 27874 8472
rect 28850 8438 29598 8472
rect 27778 8376 27812 8438
rect 28910 8376 29598 8438
rect 27922 8304 27938 8338
rect 28714 8304 28730 8338
rect 28773 8276 28807 8292
rect 28773 8192 28807 8208
rect 27922 8146 27938 8180
rect 28714 8146 28730 8180
rect 28773 8118 28807 8134
rect 28773 8034 28807 8050
rect 27922 7988 27938 8022
rect 28714 7988 28730 8022
rect 28773 7960 28807 7976
rect 28773 7876 28807 7892
rect 27922 7830 27938 7864
rect 28714 7830 28730 7864
rect 28773 7802 28807 7818
rect 28773 7718 28807 7734
rect 27922 7672 27938 7706
rect 28714 7672 28730 7706
rect 27778 7572 27812 7634
rect 28910 7634 28912 8376
rect 28946 7634 29598 8376
rect 28910 7572 29598 7634
rect 27778 7538 27874 7572
rect 28850 7538 29598 7572
rect 28910 7434 29598 7538
rect 29732 8581 29766 8597
rect 29732 8189 29766 8205
rect 30590 8581 30624 8597
rect 30590 8189 30624 8205
rect 31448 8581 31482 8597
rect 31448 8189 31482 8205
rect 29778 8112 29794 8146
rect 30562 8112 30578 8146
rect 30636 8112 30652 8146
rect 31420 8112 31436 8146
rect 29778 8004 29794 8038
rect 30562 8004 30578 8038
rect 30636 8004 30652 8038
rect 31420 8004 31436 8038
rect 29732 7945 29766 7961
rect 29732 7553 29766 7569
rect 30590 7945 30624 7961
rect 30590 7553 30624 7569
rect 31448 7945 31482 7961
rect 31448 7553 31482 7569
rect 33540 8946 33574 9042
rect 32956 8906 32972 8940
rect 33140 8906 33156 8940
rect 33214 8906 33230 8940
rect 33398 8906 33414 8940
rect 32910 8847 32944 8863
rect 32910 8055 32944 8071
rect 33168 8847 33202 8863
rect 33168 8055 33202 8071
rect 33426 8847 33460 8863
rect 33426 8055 33460 8071
rect 32956 7978 32972 8012
rect 33140 7978 33156 8012
rect 33214 7978 33230 8012
rect 33398 7978 33414 8012
rect 32796 7910 32830 7972
rect 33540 7910 33574 7972
rect 32796 7876 32892 7910
rect 33478 7876 33574 7910
rect 33636 8946 33670 9042
rect 34380 8946 34414 9042
rect 33796 8906 33812 8940
rect 33980 8906 33996 8940
rect 34054 8906 34070 8940
rect 34238 8906 34254 8940
rect 33750 8847 33784 8863
rect 33750 8055 33784 8071
rect 34008 8847 34042 8863
rect 34008 8055 34042 8071
rect 34266 8847 34300 8863
rect 34266 8055 34300 8071
rect 33796 7978 33812 8012
rect 33980 7978 33996 8012
rect 34054 7978 34070 8012
rect 34238 7978 34254 8012
rect 33636 7910 33670 7972
rect 34476 8726 34510 8822
rect 34792 8726 34826 8822
rect 34618 8686 34634 8720
rect 34668 8686 34684 8720
rect 34590 8627 34624 8643
rect 34590 8235 34624 8251
rect 34678 8627 34712 8643
rect 34678 8235 34712 8251
rect 34618 8158 34634 8192
rect 34668 8158 34684 8192
rect 34476 8090 34510 8152
rect 34792 8090 34826 8152
rect 34476 8056 34572 8090
rect 34730 8056 34826 8090
rect 34896 8726 34930 8822
rect 35212 8726 35246 8822
rect 35038 8686 35054 8720
rect 35088 8686 35104 8720
rect 35010 8627 35044 8643
rect 35010 8235 35044 8251
rect 35098 8627 35132 8643
rect 35098 8235 35132 8251
rect 35038 8158 35054 8192
rect 35088 8158 35104 8192
rect 34896 8090 34930 8152
rect 35212 8090 35246 8152
rect 34896 8056 34992 8090
rect 35150 8056 35246 8090
rect 35316 8726 35350 8822
rect 35632 8726 35666 8822
rect 35458 8686 35474 8720
rect 35508 8686 35524 8720
rect 35430 8627 35464 8643
rect 35430 8235 35464 8251
rect 35518 8627 35552 8643
rect 35518 8235 35552 8251
rect 35458 8158 35474 8192
rect 35508 8158 35524 8192
rect 35316 8090 35350 8152
rect 35632 8090 35666 8152
rect 35316 8056 35412 8090
rect 35570 8056 35666 8090
rect 34380 7910 34414 7972
rect 33636 7876 33732 7910
rect 34318 7876 34414 7910
rect 34250 7648 34490 7670
rect 29778 7476 29794 7510
rect 30562 7476 30578 7510
rect 30636 7476 30652 7510
rect 31420 7476 31436 7510
rect 28910 7432 29632 7434
rect 27778 7398 27874 7432
rect 28850 7398 29632 7432
rect 27778 7336 27812 7398
rect 28910 7372 29632 7398
rect 31582 7372 31616 7434
rect 28910 7338 29694 7372
rect 31520 7360 31616 7372
rect 33338 7614 33434 7648
rect 34176 7614 34490 7648
rect 33338 7552 33372 7614
rect 31520 7338 31800 7360
rect 28910 7336 31800 7338
rect 27922 7264 27938 7298
rect 28714 7264 28730 7298
rect 28773 7236 28807 7252
rect 28773 7152 28807 7168
rect 27922 7106 27938 7140
rect 28714 7106 28730 7140
rect 28773 7078 28807 7094
rect 28773 6994 28807 7010
rect 27922 6948 27938 6982
rect 28714 6948 28730 6982
rect 28773 6920 28807 6936
rect 28773 6836 28807 6852
rect 27922 6790 27938 6824
rect 28714 6790 28730 6824
rect 28773 6762 28807 6778
rect 28773 6678 28807 6694
rect 27922 6632 27938 6666
rect 28714 6632 28730 6666
rect 27778 6532 27812 6594
rect 28910 6594 28912 7336
rect 28946 7220 31800 7336
rect 28946 6594 29150 7220
rect 29470 7198 31800 7220
rect 29470 7180 32116 7198
rect 29538 7164 30776 7180
rect 29538 7115 29572 7164
rect 30742 7102 30776 7164
rect 29753 7030 29769 7064
rect 30545 7030 30561 7064
rect 29676 7002 29710 7018
rect 29676 6818 29710 6834
rect 30604 7002 30638 7018
rect 30604 6818 30638 6834
rect 29753 6772 29769 6806
rect 30545 6772 30561 6806
rect 29538 6672 29572 6721
rect 30742 6672 30776 6734
rect 29538 6638 30776 6672
rect 30878 7164 32116 7180
rect 30878 7102 30912 7164
rect 32082 7102 32116 7164
rect 31093 7030 31109 7064
rect 31885 7030 31901 7064
rect 31016 7002 31050 7018
rect 31016 6818 31050 6834
rect 31944 7002 31978 7018
rect 31944 6818 31978 6834
rect 31093 6772 31109 6806
rect 31885 6772 31901 6806
rect 30878 6672 30912 6734
rect 34238 7552 34490 7614
rect 33518 7476 33534 7510
rect 33602 7476 33618 7510
rect 33676 7476 33692 7510
rect 33760 7476 33776 7510
rect 33834 7476 33850 7510
rect 33918 7476 33934 7510
rect 33992 7476 34008 7510
rect 34076 7476 34092 7510
rect 33472 7426 33506 7442
rect 33472 7034 33506 7050
rect 33630 7426 33664 7442
rect 33630 7034 33664 7050
rect 33788 7426 33822 7442
rect 33788 7034 33822 7050
rect 33946 7426 33980 7442
rect 33946 7034 33980 7050
rect 34104 7426 34138 7442
rect 34104 7034 34138 7050
rect 33518 6966 33534 7000
rect 33602 6966 33618 7000
rect 33676 6966 33692 7000
rect 33760 6966 33776 7000
rect 33834 6966 33850 7000
rect 33918 6966 33934 7000
rect 33992 6966 34008 7000
rect 34076 6966 34092 7000
rect 33338 6860 33372 6924
rect 34272 7504 34490 7552
rect 34272 7470 34572 7504
rect 34730 7470 34826 7504
rect 34272 7408 34510 7470
rect 34272 7052 34476 7408
rect 34792 7408 34826 7470
rect 34618 7368 34634 7402
rect 34668 7368 34684 7402
rect 34590 7318 34624 7334
rect 34590 7126 34624 7142
rect 34678 7318 34712 7334
rect 34678 7126 34712 7142
rect 34618 7058 34634 7092
rect 34668 7058 34684 7092
rect 34272 6956 34510 7052
rect 34792 6980 34826 7052
rect 34896 7470 34992 7504
rect 35150 7470 35246 7504
rect 34896 7408 34930 7470
rect 35212 7408 35246 7470
rect 35038 7368 35054 7402
rect 35088 7368 35104 7402
rect 35010 7318 35044 7334
rect 35010 7126 35044 7142
rect 35098 7318 35132 7334
rect 35098 7126 35132 7142
rect 35038 7058 35054 7092
rect 35088 7058 35104 7092
rect 34896 6980 34930 7052
rect 34792 6956 34930 6980
rect 35212 6980 35246 7052
rect 35316 7470 35412 7504
rect 35570 7470 35666 7504
rect 35316 7408 35350 7470
rect 35632 7408 35666 7470
rect 35458 7368 35474 7402
rect 35508 7368 35524 7402
rect 35430 7318 35464 7334
rect 35430 7126 35464 7142
rect 35518 7318 35552 7334
rect 35518 7126 35552 7142
rect 35458 7058 35474 7092
rect 35508 7058 35524 7092
rect 35316 6980 35350 7052
rect 35212 6956 35350 6980
rect 35632 6956 35666 7052
rect 34272 6924 35660 6956
rect 32082 6672 32116 6734
rect 30878 6638 32116 6672
rect 33230 6828 33372 6860
rect 34238 6828 35660 6924
rect 33230 6740 35660 6828
rect 28910 6532 29150 6594
rect 27778 6498 27874 6532
rect 28850 6498 29150 6532
rect 28910 6392 29150 6498
rect 33230 6440 35130 6740
rect 27778 6358 27874 6392
rect 28850 6358 29150 6392
rect 27778 6296 27812 6358
rect 28910 6296 29150 6358
rect 27922 6224 27938 6258
rect 28714 6224 28730 6258
rect 28773 6196 28807 6212
rect 28773 6112 28807 6128
rect 27922 6066 27938 6100
rect 28714 6066 28730 6100
rect 28773 6038 28807 6054
rect 28773 5954 28807 5970
rect 27922 5908 27938 5942
rect 28714 5908 28730 5942
rect 28773 5880 28807 5896
rect 28773 5796 28807 5812
rect 27922 5750 27938 5784
rect 28714 5750 28730 5784
rect 28773 5722 28807 5738
rect 28773 5638 28807 5654
rect 27922 5592 27938 5626
rect 28714 5592 28730 5626
rect 27778 5492 27812 5554
rect 28910 5554 28912 6296
rect 28946 5554 29150 6296
rect 28910 5492 29150 5554
rect 27778 5458 27874 5492
rect 28850 5458 29150 5492
rect 28910 5376 29150 5458
rect 26380 4470 27280 4532
rect 21869 4436 22332 4470
rect 26966 4436 27280 4470
rect 21869 4145 27280 4436
rect 21835 4083 27280 4145
rect 27778 5342 27874 5376
rect 28842 5342 29150 5376
rect 27778 5280 27812 5342
rect 28904 5280 29150 5342
rect 27958 5204 27974 5238
rect 28742 5204 28758 5238
rect 27912 5145 27946 5161
rect 27912 4353 27946 4369
rect 28770 5145 28804 5161
rect 28770 4353 28804 4369
rect 27958 4276 27974 4310
rect 28742 4276 28758 4310
rect 27778 4172 27812 4234
rect 28938 4234 29150 5280
rect 29360 6368 35140 6440
rect 29360 6334 29644 6368
rect 30672 6334 30984 6368
rect 32012 6334 35140 6368
rect 29360 6272 29582 6334
rect 29360 5904 29548 6272
rect 30734 6272 30922 6334
rect 29754 6200 29770 6234
rect 30546 6200 30562 6234
rect 29686 6172 29720 6188
rect 29686 5988 29720 6004
rect 30596 6172 30630 6188
rect 30596 5988 30630 6004
rect 29754 5942 29770 5976
rect 30546 5942 30562 5976
rect 29360 5842 29582 5904
rect 30768 5904 30888 6272
rect 32074 6272 35140 6334
rect 31094 6200 31110 6234
rect 31886 6200 31902 6234
rect 31026 6172 31060 6188
rect 31026 5988 31060 6004
rect 31936 6172 31970 6188
rect 31936 5988 31970 6004
rect 31094 5942 31110 5976
rect 31886 5942 31902 5976
rect 30734 5842 30922 5904
rect 32108 5904 35140 6272
rect 32074 5842 35140 5904
rect 29360 5808 29644 5842
rect 30672 5808 30984 5842
rect 32012 5808 35140 5842
rect 29360 5718 35140 5808
rect 29360 5684 29884 5718
rect 30452 5684 31194 5718
rect 31762 5684 35140 5718
rect 29360 5622 29822 5684
rect 29360 5294 29788 5622
rect 30514 5622 31132 5684
rect 29968 5546 29984 5580
rect 30352 5546 30368 5580
rect 29922 5496 29956 5512
rect 29922 5404 29956 5420
rect 30380 5496 30414 5512
rect 30380 5404 30414 5420
rect 29968 5336 29984 5370
rect 30352 5336 30368 5370
rect 29360 5232 29822 5294
rect 30548 5294 31098 5622
rect 31824 5622 35140 5684
rect 31278 5546 31294 5580
rect 31662 5546 31678 5580
rect 31232 5496 31266 5512
rect 31232 5404 31266 5420
rect 31690 5496 31724 5512
rect 31690 5404 31724 5420
rect 31278 5336 31294 5370
rect 31662 5336 31678 5370
rect 30514 5232 31132 5294
rect 31858 5294 35140 5622
rect 31824 5232 35140 5294
rect 29360 5198 29884 5232
rect 30452 5198 31194 5232
rect 31762 5198 35140 5232
rect 29360 5108 35140 5198
rect 29360 5074 29644 5108
rect 30672 5074 30984 5108
rect 32012 5074 35140 5108
rect 29360 5012 29582 5074
rect 29360 4644 29548 5012
rect 30734 5012 30922 5074
rect 29754 4940 29770 4974
rect 30546 4940 30562 4974
rect 29686 4912 29720 4928
rect 29686 4728 29720 4744
rect 30596 4912 30630 4928
rect 30596 4728 30630 4744
rect 29754 4682 29770 4716
rect 30546 4682 30562 4716
rect 29360 4582 29582 4644
rect 30768 4644 30888 5012
rect 32074 5012 35140 5074
rect 31094 4940 31110 4974
rect 31886 4940 31902 4974
rect 31026 4912 31060 4928
rect 31026 4728 31060 4744
rect 31936 4912 31970 4928
rect 31936 4728 31970 4744
rect 31094 4682 31110 4716
rect 31886 4682 31902 4716
rect 30734 4582 30922 4644
rect 32108 4644 35140 5012
rect 32074 4582 35140 4644
rect 29360 4548 29644 4582
rect 30672 4548 30984 4582
rect 32012 4548 35140 4582
rect 29360 4500 35140 4548
rect 35380 6134 38400 6440
rect 35380 6100 36334 6134
rect 36962 6100 37120 6134
rect 37748 6100 38400 6134
rect 35380 6038 36272 6100
rect 35380 4330 36238 6038
rect 35340 4310 36238 4330
rect 28904 4172 29150 4234
rect 27778 4138 27874 4172
rect 28842 4138 29150 4172
rect 28910 4110 29150 4138
rect 29360 4168 36238 4310
rect 29360 4134 32684 4168
rect 34058 4134 34874 4168
rect 35458 4134 36238 4168
rect 12974 4050 13345 4083
rect 8573 4049 13345 4050
rect 15173 4049 15545 4083
rect 17373 4049 17745 4083
rect 19573 4049 19945 4083
rect 21773 4049 27280 4083
rect -300 3640 27280 4049
rect 29360 4072 32622 4134
rect 29360 3640 32588 4072
rect -300 3526 32588 3640
rect -300 3492 17064 3526
rect 17806 3492 32588 3526
rect -300 3430 17002 3492
rect -300 2464 16968 3430
rect 17868 3444 32588 3492
rect 34120 4072 34812 4134
rect 32768 3996 32784 4030
rect 32852 3996 32868 4030
rect 32926 3996 32942 4030
rect 33010 3996 33026 4030
rect 33084 3996 33100 4030
rect 33168 3996 33184 4030
rect 33242 3996 33258 4030
rect 33326 3996 33342 4030
rect 33400 3996 33416 4030
rect 33484 3996 33500 4030
rect 33558 3996 33574 4030
rect 33642 3996 33658 4030
rect 33716 3996 33732 4030
rect 33800 3996 33816 4030
rect 33874 3996 33890 4030
rect 33958 3996 33974 4030
rect 32722 3946 32756 3962
rect 32722 3554 32756 3570
rect 32880 3946 32914 3962
rect 32880 3554 32914 3570
rect 33038 3946 33072 3962
rect 33038 3554 33072 3570
rect 33196 3946 33230 3962
rect 33196 3554 33230 3570
rect 33354 3946 33388 3962
rect 33354 3554 33388 3570
rect 33512 3946 33546 3962
rect 33512 3554 33546 3570
rect 33670 3946 33704 3962
rect 33670 3554 33704 3570
rect 33828 3946 33862 3962
rect 33828 3554 33862 3570
rect 33986 3946 34020 3962
rect 33986 3554 34020 3570
rect 32768 3486 32784 3520
rect 32852 3486 32868 3520
rect 32926 3486 32942 3520
rect 33010 3486 33026 3520
rect 33084 3486 33100 3520
rect 33168 3486 33184 3520
rect 33242 3486 33258 3520
rect 33326 3486 33342 3520
rect 33400 3486 33416 3520
rect 33484 3486 33500 3520
rect 33558 3486 33574 3520
rect 33642 3486 33658 3520
rect 33716 3486 33732 3520
rect 33800 3486 33816 3520
rect 33874 3486 33890 3520
rect 33958 3486 33974 3520
rect 17868 3430 32622 3444
rect 17148 3354 17164 3388
rect 17232 3354 17248 3388
rect 17306 3354 17322 3388
rect 17390 3354 17406 3388
rect 17464 3354 17480 3388
rect 17548 3354 17564 3388
rect 17622 3354 17638 3388
rect 17706 3354 17722 3388
rect 17102 3304 17136 3320
rect 17102 2512 17136 2528
rect 17260 3304 17294 3320
rect 17260 2512 17294 2528
rect 17418 3304 17452 3320
rect 17418 2512 17452 2528
rect 17576 3304 17610 3320
rect 17576 2512 17610 2528
rect 17734 3304 17768 3320
rect 17734 2512 17768 2528
rect -300 2430 17002 2464
rect 17902 3382 32622 3430
rect 34154 3444 34778 4072
rect 35520 4072 36238 4134
rect 34958 3996 34974 4030
rect 35042 3996 35058 4030
rect 35116 3996 35132 4030
rect 35200 3996 35216 4030
rect 35274 3996 35290 4030
rect 35358 3996 35374 4030
rect 34912 3946 34946 3962
rect 34912 3554 34946 3570
rect 35070 3946 35104 3962
rect 35070 3554 35104 3570
rect 35228 3946 35262 3962
rect 35228 3554 35262 3570
rect 35386 3946 35420 3962
rect 35386 3554 35420 3570
rect 34958 3486 34974 3520
rect 35042 3486 35058 3520
rect 35116 3486 35132 3520
rect 35200 3486 35216 3520
rect 35274 3486 35290 3520
rect 35358 3486 35374 3520
rect 34120 3382 34812 3444
rect 35554 3864 36238 4072
rect 37024 6038 37058 6100
rect 36444 5966 36460 6000
rect 36836 5966 36852 6000
rect 36376 5938 36410 5954
rect 36376 5754 36410 5770
rect 36886 5938 36920 5954
rect 36886 5754 36920 5770
rect 36444 5708 36460 5742
rect 36836 5708 36852 5742
rect 36376 5680 36410 5696
rect 36376 5496 36410 5512
rect 36886 5680 36920 5696
rect 36886 5496 36920 5512
rect 36444 5450 36460 5484
rect 36836 5450 36852 5484
rect 36376 5422 36410 5438
rect 36376 5238 36410 5254
rect 36886 5422 36920 5438
rect 36886 5238 36920 5254
rect 36444 5192 36460 5226
rect 36836 5192 36852 5226
rect 36376 5164 36410 5180
rect 36376 4980 36410 4996
rect 36886 5164 36920 5180
rect 36886 4980 36920 4996
rect 36444 4934 36460 4968
rect 36836 4934 36852 4968
rect 36376 4906 36410 4922
rect 36376 4722 36410 4738
rect 36886 4906 36920 4922
rect 36886 4722 36920 4738
rect 36444 4676 36460 4710
rect 36836 4676 36852 4710
rect 36376 4648 36410 4664
rect 36376 4464 36410 4480
rect 36886 4648 36920 4664
rect 36886 4464 36920 4480
rect 36444 4418 36460 4452
rect 36836 4418 36852 4452
rect 36376 4390 36410 4406
rect 36376 4206 36410 4222
rect 36886 4390 36920 4406
rect 36886 4206 36920 4222
rect 36444 4160 36460 4194
rect 36836 4160 36852 4194
rect 36376 4132 36410 4148
rect 36376 3948 36410 3964
rect 36886 4132 36920 4148
rect 36886 3948 36920 3964
rect 36444 3902 36460 3936
rect 36836 3902 36852 3936
rect 35554 3802 36272 3864
rect 37810 6038 38400 6100
rect 37230 5966 37246 6000
rect 37622 5966 37638 6000
rect 37162 5938 37196 5954
rect 37162 5754 37196 5770
rect 37672 5938 37706 5954
rect 37672 5754 37706 5770
rect 37230 5708 37246 5742
rect 37622 5708 37638 5742
rect 37162 5680 37196 5696
rect 37162 5496 37196 5512
rect 37672 5680 37706 5696
rect 37672 5496 37706 5512
rect 37230 5450 37246 5484
rect 37622 5450 37638 5484
rect 37162 5422 37196 5438
rect 37162 5238 37196 5254
rect 37672 5422 37706 5438
rect 37672 5238 37706 5254
rect 37230 5192 37246 5226
rect 37622 5192 37638 5226
rect 37162 5164 37196 5180
rect 37162 4980 37196 4996
rect 37672 5164 37706 5180
rect 37672 4980 37706 4996
rect 37230 4934 37246 4968
rect 37622 4934 37638 4968
rect 37162 4906 37196 4922
rect 37162 4722 37196 4738
rect 37672 4906 37706 4922
rect 37672 4722 37706 4738
rect 37230 4676 37246 4710
rect 37622 4676 37638 4710
rect 37162 4648 37196 4664
rect 37162 4464 37196 4480
rect 37672 4648 37706 4664
rect 37672 4464 37706 4480
rect 37230 4418 37246 4452
rect 37622 4418 37638 4452
rect 37162 4390 37196 4406
rect 37162 4206 37196 4222
rect 37672 4390 37706 4406
rect 37672 4206 37706 4222
rect 37230 4160 37246 4194
rect 37622 4160 37638 4194
rect 37162 4132 37196 4148
rect 37162 3948 37196 3964
rect 37672 4132 37706 4148
rect 37672 3948 37706 3964
rect 37230 3902 37246 3936
rect 37622 3902 37638 3936
rect 37024 3802 37058 3864
rect 37844 3864 38400 6038
rect 37810 3802 38400 3864
rect 35554 3768 36334 3802
rect 36962 3768 37120 3802
rect 37748 3768 38400 3802
rect 35554 3444 38400 3768
rect 35520 3382 38400 3444
rect 17902 3348 32684 3382
rect 34058 3348 34874 3382
rect 35458 3348 38400 3382
rect 17902 3238 38400 3348
rect 17902 3204 32347 3238
rect 32787 3204 33947 3238
rect 34387 3204 35547 3238
rect 35987 3204 38400 3238
rect 17902 3142 32292 3204
rect 17902 2514 32258 3142
rect 32842 3142 33892 3204
rect 32438 3066 32454 3100
rect 32522 3066 32538 3100
rect 32596 3066 32612 3100
rect 32680 3066 32696 3100
rect 32392 3016 32426 3032
rect 32392 2624 32426 2640
rect 32550 3016 32584 3032
rect 32550 2624 32584 2640
rect 32708 3016 32742 3032
rect 32708 2624 32742 2640
rect 32438 2556 32454 2590
rect 32522 2556 32538 2590
rect 32596 2556 32612 2590
rect 32680 2556 32696 2590
rect 17902 2464 32292 2514
rect 17868 2452 32292 2464
rect 32876 2514 33858 3142
rect 34426 3142 35492 3204
rect 34038 3066 34054 3100
rect 34122 3066 34138 3100
rect 34196 3066 34212 3100
rect 34280 3066 34296 3100
rect 33992 3016 34026 3032
rect 33992 2624 34026 2640
rect 34150 3016 34184 3032
rect 34150 2624 34184 2640
rect 34308 3016 34342 3032
rect 34308 2624 34342 2640
rect 34038 2556 34054 2590
rect 34122 2556 34138 2590
rect 34196 2556 34212 2590
rect 34280 2556 34296 2590
rect 32842 2452 33892 2514
rect 34426 2514 34442 3142
rect 34476 2514 35458 3142
rect 36042 3142 38400 3204
rect 35638 3066 35654 3100
rect 35722 3066 35738 3100
rect 35796 3066 35812 3100
rect 35880 3066 35896 3100
rect 35592 3016 35626 3032
rect 35592 2624 35626 2640
rect 35750 3016 35784 3032
rect 35750 2624 35784 2640
rect 35908 3016 35942 3032
rect 35908 2624 35942 2640
rect 35638 2556 35654 2590
rect 35722 2556 35738 2590
rect 35796 2556 35812 2590
rect 35880 2556 35896 2590
rect 34426 2452 35492 2514
rect 36076 2514 38400 3142
rect 36042 2452 38400 2514
rect 17868 2430 32354 2452
rect -300 2418 32354 2430
rect 32780 2418 33954 2452
rect 34380 2418 35554 2452
rect 35980 2418 38400 2452
rect -300 2402 38400 2418
rect -300 2368 17064 2402
rect 17806 2368 38400 2402
rect -300 2229 38400 2368
rect -300 2195 -117 2229
rect 1253 2195 1483 2229
rect -300 2133 0 2195
rect -300 1165 -151 2133
rect -117 2049 0 2133
rect 180 2095 340 2195
rect 55 2061 71 2095
rect 447 2061 463 2095
rect 520 2049 620 2195
rect 800 2095 960 2195
rect 1140 2133 1483 2195
rect 673 2061 689 2095
rect 1065 2061 1081 2095
rect 1140 2049 1253 2133
rect -117 2033 21 2049
rect -117 1265 -13 2033
rect -117 1249 21 1265
rect 497 2033 639 2049
rect 531 1265 605 2033
rect 497 1249 639 1265
rect 1115 2033 1253 2049
rect 1149 1265 1253 2033
rect 1115 1249 1253 1265
rect -117 1165 0 1249
rect 55 1203 71 1237
rect 447 1203 463 1237
rect -300 1120 0 1165
rect 180 1120 340 1203
rect 520 1120 620 1249
rect 673 1203 689 1237
rect 1065 1203 1081 1237
rect 800 1120 960 1203
rect 1140 1165 1253 1249
rect 1287 1165 1449 2133
rect 2853 2133 3083 2229
rect 1655 2061 1671 2095
rect 2047 2061 2063 2095
rect 2273 2061 2289 2095
rect 2665 2061 2681 2095
rect 1587 2033 1621 2049
rect 1587 1249 1621 1265
rect 2097 2033 2131 2049
rect 2097 1249 2131 1265
rect 2205 2033 2239 2049
rect 2205 1249 2239 1265
rect 2715 2033 2749 2049
rect 2715 1249 2749 1265
rect 1655 1203 1671 1237
rect 2047 1203 2063 1237
rect 2273 1203 2289 1237
rect 2665 1203 2681 1237
rect 1140 1120 1483 1165
rect -300 1103 1483 1120
rect 2887 1165 3049 2133
rect 4453 2133 4683 2229
rect 3255 2061 3271 2095
rect 3647 2061 3663 2095
rect 3873 2061 3889 2095
rect 4265 2061 4281 2095
rect 3187 2033 3221 2049
rect 3187 1249 3221 1265
rect 3697 2033 3731 2049
rect 3697 1249 3731 1265
rect 3805 2033 3839 2049
rect 3805 1249 3839 1265
rect 4315 2033 4349 2049
rect 4315 1249 4349 1265
rect 3255 1203 3271 1237
rect 3647 1203 3663 1237
rect 3873 1203 3889 1237
rect 4265 1203 4281 1237
rect 2853 1103 3083 1165
rect 4487 1165 4649 2133
rect 6053 2133 6283 2229
rect 4855 2061 4871 2095
rect 5247 2061 5263 2095
rect 5473 2061 5489 2095
rect 5865 2061 5881 2095
rect 4787 2033 4821 2049
rect 4787 1249 4821 1265
rect 5297 2033 5331 2049
rect 5297 1249 5331 1265
rect 5405 2033 5439 2049
rect 5405 1249 5439 1265
rect 5915 2033 5949 2049
rect 5915 1249 5949 1265
rect 4855 1203 4871 1237
rect 5247 1203 5263 1237
rect 5473 1203 5489 1237
rect 5865 1203 5881 1237
rect 4453 1103 4683 1165
rect 6087 1165 6249 2133
rect 7653 2133 7883 2229
rect 6455 2061 6471 2095
rect 6847 2061 6863 2095
rect 7073 2061 7089 2095
rect 7465 2061 7481 2095
rect 6387 2033 6421 2049
rect 6387 1249 6421 1265
rect 6897 2033 6931 2049
rect 6897 1249 6931 1265
rect 7005 2033 7039 2049
rect 7005 1249 7039 1265
rect 7515 2033 7549 2049
rect 7515 1249 7549 1265
rect 6455 1203 6471 1237
rect 6847 1203 6863 1237
rect 7073 1203 7089 1237
rect 7465 1203 7481 1237
rect 6053 1103 6283 1165
rect 7687 1165 7849 2133
rect 9253 2133 9483 2229
rect 8055 2061 8071 2095
rect 8447 2061 8463 2095
rect 8673 2061 8689 2095
rect 9065 2061 9081 2095
rect 7987 2033 8021 2049
rect 7987 1249 8021 1265
rect 8497 2033 8531 2049
rect 8497 1249 8531 1265
rect 8605 2033 8639 2049
rect 8605 1249 8639 1265
rect 9115 2033 9149 2049
rect 9115 1249 9149 1265
rect 8055 1203 8071 1237
rect 8447 1203 8463 1237
rect 8673 1203 8689 1237
rect 9065 1203 9081 1237
rect 7653 1103 7883 1165
rect 9287 1165 9449 2133
rect 10853 2133 11083 2229
rect 9655 2061 9671 2095
rect 10047 2061 10063 2095
rect 10273 2061 10289 2095
rect 10665 2061 10681 2095
rect 9587 2033 9621 2049
rect 9587 1249 9621 1265
rect 10097 2033 10131 2049
rect 10097 1249 10131 1265
rect 10205 2033 10239 2049
rect 10205 1249 10239 1265
rect 10715 2033 10749 2049
rect 10715 1249 10749 1265
rect 9655 1203 9671 1237
rect 10047 1203 10063 1237
rect 10273 1203 10289 1237
rect 10665 1203 10681 1237
rect 9253 1103 9483 1165
rect 10887 1165 11049 2133
rect 12453 2133 12683 2229
rect 11255 2061 11271 2095
rect 11647 2061 11663 2095
rect 11873 2061 11889 2095
rect 12265 2061 12281 2095
rect 11187 2033 11221 2049
rect 11187 1249 11221 1265
rect 11697 2033 11731 2049
rect 11697 1249 11731 1265
rect 11805 2033 11839 2049
rect 11805 1249 11839 1265
rect 12315 2033 12349 2049
rect 12315 1249 12349 1265
rect 11255 1203 11271 1237
rect 11647 1203 11663 1237
rect 11873 1203 11889 1237
rect 12265 1203 12281 1237
rect 10853 1103 11083 1165
rect 12487 1165 12649 2133
rect 14053 2133 14283 2229
rect 12855 2061 12871 2095
rect 13247 2061 13263 2095
rect 13473 2061 13489 2095
rect 13865 2061 13881 2095
rect 12787 2033 12821 2049
rect 12787 1249 12821 1265
rect 13297 2033 13331 2049
rect 13297 1249 13331 1265
rect 13405 2033 13439 2049
rect 13405 1249 13439 1265
rect 13915 2033 13949 2049
rect 13915 1249 13949 1265
rect 12855 1203 12871 1237
rect 13247 1203 13263 1237
rect 13473 1203 13489 1237
rect 13865 1203 13881 1237
rect 12453 1103 12683 1165
rect 14087 1165 14249 2133
rect 15653 2133 15883 2229
rect 14455 2061 14471 2095
rect 14847 2061 14863 2095
rect 15073 2061 15089 2095
rect 15465 2061 15481 2095
rect 14387 2033 14421 2049
rect 14387 1249 14421 1265
rect 14897 2033 14931 2049
rect 14897 1249 14931 1265
rect 15005 2033 15039 2049
rect 15005 1249 15039 1265
rect 15515 2033 15549 2049
rect 15515 1249 15549 1265
rect 14455 1203 14471 1237
rect 14847 1203 14863 1237
rect 15073 1203 15089 1237
rect 15465 1203 15481 1237
rect 14053 1103 14283 1165
rect 15687 1165 15849 2133
rect 17253 2133 17483 2229
rect 16055 2061 16071 2095
rect 16447 2061 16463 2095
rect 16673 2061 16689 2095
rect 17065 2061 17081 2095
rect 15987 2033 16021 2049
rect 15987 1249 16021 1265
rect 16497 2033 16531 2049
rect 16497 1249 16531 1265
rect 16605 2033 16639 2049
rect 16605 1249 16639 1265
rect 17115 2033 17149 2049
rect 17115 1249 17149 1265
rect 16055 1203 16071 1237
rect 16447 1203 16463 1237
rect 16673 1203 16689 1237
rect 17065 1203 17081 1237
rect 15653 1103 15883 1165
rect 17287 1165 17449 2133
rect 18853 2133 19083 2229
rect 17655 2061 17671 2095
rect 18047 2061 18063 2095
rect 18273 2061 18289 2095
rect 18665 2061 18681 2095
rect 17587 2033 17621 2049
rect 17587 1249 17621 1265
rect 18097 2033 18131 2049
rect 18097 1249 18131 1265
rect 18205 2033 18239 2049
rect 18205 1249 18239 1265
rect 18715 2033 18749 2049
rect 18715 1249 18749 1265
rect 17655 1203 17671 1237
rect 18047 1203 18063 1237
rect 18273 1203 18289 1237
rect 18665 1203 18681 1237
rect 17253 1103 17483 1165
rect 18887 1165 19049 2133
rect 20453 2133 20683 2229
rect 19255 2061 19271 2095
rect 19647 2061 19663 2095
rect 19873 2061 19889 2095
rect 20265 2061 20281 2095
rect 19187 2033 19221 2049
rect 19187 1249 19221 1265
rect 19697 2033 19731 2049
rect 19697 1249 19731 1265
rect 19805 2033 19839 2049
rect 19805 1249 19839 1265
rect 20315 2033 20349 2049
rect 20315 1249 20349 1265
rect 19255 1203 19271 1237
rect 19647 1203 19663 1237
rect 19873 1203 19889 1237
rect 20265 1203 20281 1237
rect 18853 1103 19083 1165
rect 20487 1165 20649 2133
rect 22053 2133 22283 2229
rect 20855 2061 20871 2095
rect 21247 2061 21263 2095
rect 21473 2061 21489 2095
rect 21865 2061 21881 2095
rect 20787 2033 20821 2049
rect 20787 1249 20821 1265
rect 21297 2033 21331 2049
rect 21297 1249 21331 1265
rect 21405 2033 21439 2049
rect 21405 1249 21439 1265
rect 21915 2033 21949 2049
rect 21915 1249 21949 1265
rect 20855 1203 20871 1237
rect 21247 1203 21263 1237
rect 21473 1203 21489 1237
rect 21865 1203 21881 1237
rect 20453 1103 20683 1165
rect 22087 1165 22249 2133
rect 23653 2133 23883 2229
rect 22455 2061 22471 2095
rect 22847 2061 22863 2095
rect 23073 2061 23089 2095
rect 23465 2061 23481 2095
rect 22387 2033 22421 2049
rect 22387 1249 22421 1265
rect 22897 2033 22931 2049
rect 22897 1249 22931 1265
rect 23005 2033 23039 2049
rect 23005 1249 23039 1265
rect 23515 2033 23549 2049
rect 23515 1249 23549 1265
rect 22455 1203 22471 1237
rect 22847 1203 22863 1237
rect 23073 1203 23089 1237
rect 23465 1203 23481 1237
rect 22053 1103 22283 1165
rect 23687 1165 23849 2133
rect 25253 2133 25483 2229
rect 24055 2061 24071 2095
rect 24447 2061 24463 2095
rect 24673 2061 24689 2095
rect 25065 2061 25081 2095
rect 23987 2033 24021 2049
rect 23987 1249 24021 1265
rect 24497 2033 24531 2049
rect 24497 1249 24531 1265
rect 24605 2033 24639 2049
rect 24605 1249 24639 1265
rect 25115 2033 25149 2049
rect 25115 1249 25149 1265
rect 24055 1203 24071 1237
rect 24447 1203 24463 1237
rect 24673 1203 24689 1237
rect 25065 1203 25081 1237
rect 23653 1103 23883 1165
rect 25287 1165 25449 2133
rect 26853 2133 27083 2229
rect 25655 2061 25671 2095
rect 26047 2061 26063 2095
rect 26273 2061 26289 2095
rect 26665 2061 26681 2095
rect 25587 2033 25621 2049
rect 25587 1249 25621 1265
rect 26097 2033 26131 2049
rect 26097 1249 26131 1265
rect 26205 2033 26239 2049
rect 26205 1249 26239 1265
rect 26715 2033 26749 2049
rect 26715 1249 26749 1265
rect 25655 1203 25671 1237
rect 26047 1203 26063 1237
rect 26273 1203 26289 1237
rect 26665 1203 26681 1237
rect 25253 1103 25483 1165
rect 26887 1165 27049 2133
rect 28453 2133 28683 2229
rect 27255 2061 27271 2095
rect 27647 2061 27663 2095
rect 27873 2061 27889 2095
rect 28265 2061 28281 2095
rect 27187 2033 27221 2049
rect 27187 1249 27221 1265
rect 27697 2033 27731 2049
rect 27697 1249 27731 1265
rect 27805 2033 27839 2049
rect 27805 1249 27839 1265
rect 28315 2033 28349 2049
rect 28315 1249 28349 1265
rect 27255 1203 27271 1237
rect 27647 1203 27663 1237
rect 27873 1203 27889 1237
rect 28265 1203 28281 1237
rect 26853 1103 27083 1165
rect 28487 1165 28649 2133
rect 30053 2133 30283 2229
rect 28855 2061 28871 2095
rect 29247 2061 29263 2095
rect 29473 2061 29489 2095
rect 29865 2061 29881 2095
rect 28787 2033 28821 2049
rect 28787 1249 28821 1265
rect 29297 2033 29331 2049
rect 29297 1249 29331 1265
rect 29405 2033 29439 2049
rect 29405 1249 29439 1265
rect 29915 2033 29949 2049
rect 29915 1249 29949 1265
rect 28855 1203 28871 1237
rect 29247 1203 29263 1237
rect 29473 1203 29489 1237
rect 29865 1203 29881 1237
rect 28453 1103 28683 1165
rect 30087 1165 30249 2133
rect 31653 2133 31883 2229
rect 30455 2061 30471 2095
rect 30847 2061 30863 2095
rect 31073 2061 31089 2095
rect 31465 2061 31481 2095
rect 30387 2033 30421 2049
rect 30387 1249 30421 1265
rect 30897 2033 30931 2049
rect 30897 1249 30931 1265
rect 31005 2033 31039 2049
rect 31005 1249 31039 1265
rect 31515 2033 31549 2049
rect 31515 1249 31549 1265
rect 30455 1203 30471 1237
rect 30847 1203 30863 1237
rect 31073 1203 31089 1237
rect 31465 1203 31481 1237
rect 30053 1103 30283 1165
rect 31687 1165 31849 2133
rect 33253 2133 33483 2229
rect 32055 2061 32071 2095
rect 32447 2061 32463 2095
rect 32673 2061 32689 2095
rect 33065 2061 33081 2095
rect 31987 2033 32021 2049
rect 31987 1249 32021 1265
rect 32497 2033 32531 2049
rect 32497 1249 32531 1265
rect 32605 2033 32639 2049
rect 32605 1249 32639 1265
rect 33115 2033 33149 2049
rect 33115 1249 33149 1265
rect 32055 1203 32071 1237
rect 32447 1203 32463 1237
rect 32673 1203 32689 1237
rect 33065 1203 33081 1237
rect 31653 1103 31883 1165
rect 33287 1165 33449 2133
rect 34853 2133 35083 2229
rect 33655 2061 33671 2095
rect 34047 2061 34063 2095
rect 34273 2061 34289 2095
rect 34665 2061 34681 2095
rect 33587 2033 33621 2049
rect 33587 1249 33621 1265
rect 34097 2033 34131 2049
rect 34097 1249 34131 1265
rect 34205 2033 34239 2049
rect 34205 1249 34239 1265
rect 34715 2033 34749 2049
rect 34715 1249 34749 1265
rect 33655 1203 33671 1237
rect 34047 1203 34063 1237
rect 34273 1203 34289 1237
rect 34665 1203 34681 1237
rect 33253 1103 33483 1165
rect 34887 1165 35049 2133
rect 36453 2133 36683 2229
rect 35255 2061 35271 2095
rect 35647 2061 35663 2095
rect 35873 2061 35889 2095
rect 36265 2061 36281 2095
rect 35187 2033 35221 2049
rect 35187 1249 35221 1265
rect 35697 2033 35731 2049
rect 35697 1249 35731 1265
rect 35805 2033 35839 2049
rect 35805 1249 35839 1265
rect 36315 2033 36349 2049
rect 36315 1249 36349 1265
rect 35255 1203 35271 1237
rect 35647 1203 35663 1237
rect 35873 1203 35889 1237
rect 36265 1203 36281 1237
rect 34853 1103 35083 1165
rect 36487 1165 36649 2133
rect 38053 2133 38400 2229
rect 36855 2061 36871 2095
rect 37247 2061 37263 2095
rect 37473 2061 37489 2095
rect 37865 2061 37881 2095
rect 36787 2033 36821 2049
rect 36787 1249 36821 1265
rect 37297 2033 37331 2049
rect 37297 1249 37331 1265
rect 37405 2033 37439 2049
rect 37405 1249 37439 1265
rect 37915 2033 37949 2049
rect 37915 1249 37949 1265
rect 36855 1203 36871 1237
rect 37247 1203 37263 1237
rect 37473 1203 37489 1237
rect 37865 1203 37881 1237
rect 36453 1103 36683 1165
rect 38087 1165 38400 2133
rect 38053 1103 38400 1165
rect -300 1069 -55 1103
rect 1191 1069 1545 1103
rect 2791 1069 3145 1103
rect 4391 1069 4745 1103
rect 5991 1069 6345 1103
rect 7591 1069 7945 1103
rect 9191 1069 9545 1103
rect 10791 1069 11145 1103
rect 12391 1069 12745 1103
rect 13991 1069 14345 1103
rect 15591 1069 15945 1103
rect 17191 1069 17545 1103
rect 18791 1069 19145 1103
rect 20391 1069 20745 1103
rect 21991 1069 22345 1103
rect 23591 1069 23945 1103
rect 25191 1069 25545 1103
rect 26791 1069 27145 1103
rect 28391 1069 28745 1103
rect 29991 1069 30345 1103
rect 31591 1069 31945 1103
rect 33191 1069 33545 1103
rect 34791 1069 35145 1103
rect 36391 1069 36745 1103
rect 37991 1069 38400 1103
rect -300 1049 38400 1069
rect -300 1020 1483 1049
rect -300 987 0 1020
rect -300 619 -151 987
rect -117 903 0 987
rect 180 949 340 1020
rect 55 915 71 949
rect 447 915 463 949
rect 520 903 620 1020
rect 800 949 960 1020
rect 1140 987 1483 1020
rect 673 915 689 949
rect 1065 915 1081 949
rect 1140 903 1253 987
rect -117 887 21 903
rect -117 719 -13 887
rect -117 703 21 719
rect 497 887 639 903
rect 531 719 605 887
rect 497 703 639 719
rect 1115 887 1253 903
rect 1149 719 1253 887
rect 1115 703 1253 719
rect -117 619 0 703
rect 55 657 71 691
rect 447 657 463 691
rect -300 557 0 619
rect 180 557 340 657
rect 520 557 620 703
rect 673 657 689 691
rect 1065 657 1081 691
rect 800 557 960 657
rect 1140 619 1253 703
rect 1287 619 1449 987
rect 2853 987 3083 1049
rect 1655 915 1671 949
rect 2047 915 2063 949
rect 2273 915 2289 949
rect 2665 915 2681 949
rect 1587 887 1621 903
rect 1587 703 1621 719
rect 2097 887 2131 903
rect 2097 703 2131 719
rect 2205 887 2239 903
rect 2205 703 2239 719
rect 2715 887 2749 903
rect 2715 703 2749 719
rect 1655 657 1671 691
rect 2047 657 2063 691
rect 2273 657 2289 691
rect 2665 657 2681 691
rect 1140 557 1483 619
rect 2887 619 3049 987
rect 4453 987 4683 1049
rect 3255 915 3271 949
rect 3647 915 3663 949
rect 3873 915 3889 949
rect 4265 915 4281 949
rect 3187 887 3221 903
rect 3187 703 3221 719
rect 3697 887 3731 903
rect 3697 703 3731 719
rect 3805 887 3839 903
rect 3805 703 3839 719
rect 4315 887 4349 903
rect 4315 703 4349 719
rect 3255 657 3271 691
rect 3647 657 3663 691
rect 3873 657 3889 691
rect 4265 657 4281 691
rect 2853 557 3083 619
rect 4487 619 4649 987
rect 6053 987 6283 1049
rect 4855 915 4871 949
rect 5247 915 5263 949
rect 5473 915 5489 949
rect 5865 915 5881 949
rect 4787 887 4821 903
rect 4787 703 4821 719
rect 5297 887 5331 903
rect 5297 703 5331 719
rect 5405 887 5439 903
rect 5405 703 5439 719
rect 5915 887 5949 903
rect 5915 703 5949 719
rect 4855 657 4871 691
rect 5247 657 5263 691
rect 5473 657 5489 691
rect 5865 657 5881 691
rect 4453 557 4683 619
rect 6087 619 6249 987
rect 7653 987 7883 1049
rect 6455 915 6471 949
rect 6847 915 6863 949
rect 7073 915 7089 949
rect 7465 915 7481 949
rect 6387 887 6421 903
rect 6387 703 6421 719
rect 6897 887 6931 903
rect 6897 703 6931 719
rect 7005 887 7039 903
rect 7005 703 7039 719
rect 7515 887 7549 903
rect 7515 703 7549 719
rect 6455 657 6471 691
rect 6847 657 6863 691
rect 7073 657 7089 691
rect 7465 657 7481 691
rect 6053 557 6283 619
rect 7687 619 7849 987
rect 9253 987 9483 1049
rect 8055 915 8071 949
rect 8447 915 8463 949
rect 8673 915 8689 949
rect 9065 915 9081 949
rect 7987 887 8021 903
rect 7987 703 8021 719
rect 8497 887 8531 903
rect 8497 703 8531 719
rect 8605 887 8639 903
rect 8605 703 8639 719
rect 9115 887 9149 903
rect 9115 703 9149 719
rect 8055 657 8071 691
rect 8447 657 8463 691
rect 8673 657 8689 691
rect 9065 657 9081 691
rect 7653 557 7883 619
rect 9287 619 9449 987
rect 10853 987 11083 1049
rect 9655 915 9671 949
rect 10047 915 10063 949
rect 10273 915 10289 949
rect 10665 915 10681 949
rect 9587 887 9621 903
rect 9587 703 9621 719
rect 10097 887 10131 903
rect 10097 703 10131 719
rect 10205 887 10239 903
rect 10205 703 10239 719
rect 10715 887 10749 903
rect 10715 703 10749 719
rect 9655 657 9671 691
rect 10047 657 10063 691
rect 10273 657 10289 691
rect 10665 657 10681 691
rect 9253 557 9483 619
rect 10887 619 11049 987
rect 12453 987 12683 1049
rect 11255 915 11271 949
rect 11647 915 11663 949
rect 11873 915 11889 949
rect 12265 915 12281 949
rect 11187 887 11221 903
rect 11187 703 11221 719
rect 11697 887 11731 903
rect 11697 703 11731 719
rect 11805 887 11839 903
rect 11805 703 11839 719
rect 12315 887 12349 903
rect 12315 703 12349 719
rect 11255 657 11271 691
rect 11647 657 11663 691
rect 11873 657 11889 691
rect 12265 657 12281 691
rect 10853 557 11083 619
rect 12487 619 12649 987
rect 14053 987 14283 1049
rect 12855 915 12871 949
rect 13247 915 13263 949
rect 13473 915 13489 949
rect 13865 915 13881 949
rect 12787 887 12821 903
rect 12787 703 12821 719
rect 13297 887 13331 903
rect 13297 703 13331 719
rect 13405 887 13439 903
rect 13405 703 13439 719
rect 13915 887 13949 903
rect 13915 703 13949 719
rect 12855 657 12871 691
rect 13247 657 13263 691
rect 13473 657 13489 691
rect 13865 657 13881 691
rect 12453 557 12683 619
rect 14087 619 14249 987
rect 15653 987 15883 1049
rect 14455 915 14471 949
rect 14847 915 14863 949
rect 15073 915 15089 949
rect 15465 915 15481 949
rect 14387 887 14421 903
rect 14387 703 14421 719
rect 14897 887 14931 903
rect 14897 703 14931 719
rect 15005 887 15039 903
rect 15005 703 15039 719
rect 15515 887 15549 903
rect 15515 703 15549 719
rect 14455 657 14471 691
rect 14847 657 14863 691
rect 15073 657 15089 691
rect 15465 657 15481 691
rect 14053 557 14283 619
rect 15687 619 15849 987
rect 17253 987 17483 1049
rect 16055 915 16071 949
rect 16447 915 16463 949
rect 16673 915 16689 949
rect 17065 915 17081 949
rect 15987 887 16021 903
rect 15987 703 16021 719
rect 16497 887 16531 903
rect 16497 703 16531 719
rect 16605 887 16639 903
rect 16605 703 16639 719
rect 17115 887 17149 903
rect 17115 703 17149 719
rect 16055 657 16071 691
rect 16447 657 16463 691
rect 16673 657 16689 691
rect 17065 657 17081 691
rect 15653 557 15883 619
rect 17287 619 17449 987
rect 18853 987 19083 1049
rect 17655 915 17671 949
rect 18047 915 18063 949
rect 18273 915 18289 949
rect 18665 915 18681 949
rect 17587 887 17621 903
rect 17587 703 17621 719
rect 18097 887 18131 903
rect 18097 703 18131 719
rect 18205 887 18239 903
rect 18205 703 18239 719
rect 18715 887 18749 903
rect 18715 703 18749 719
rect 17655 657 17671 691
rect 18047 657 18063 691
rect 18273 657 18289 691
rect 18665 657 18681 691
rect 17253 557 17483 619
rect 18887 619 19049 987
rect 20453 987 20683 1049
rect 19255 915 19271 949
rect 19647 915 19663 949
rect 19873 915 19889 949
rect 20265 915 20281 949
rect 19187 887 19221 903
rect 19187 703 19221 719
rect 19697 887 19731 903
rect 19697 703 19731 719
rect 19805 887 19839 903
rect 19805 703 19839 719
rect 20315 887 20349 903
rect 20315 703 20349 719
rect 19255 657 19271 691
rect 19647 657 19663 691
rect 19873 657 19889 691
rect 20265 657 20281 691
rect 18853 557 19083 619
rect 20487 619 20649 987
rect 22053 987 22283 1049
rect 20855 915 20871 949
rect 21247 915 21263 949
rect 21473 915 21489 949
rect 21865 915 21881 949
rect 20787 887 20821 903
rect 20787 703 20821 719
rect 21297 887 21331 903
rect 21297 703 21331 719
rect 21405 887 21439 903
rect 21405 703 21439 719
rect 21915 887 21949 903
rect 21915 703 21949 719
rect 20855 657 20871 691
rect 21247 657 21263 691
rect 21473 657 21489 691
rect 21865 657 21881 691
rect 20453 557 20683 619
rect 22087 619 22249 987
rect 23653 987 23883 1049
rect 22455 915 22471 949
rect 22847 915 22863 949
rect 23073 915 23089 949
rect 23465 915 23481 949
rect 22387 887 22421 903
rect 22387 703 22421 719
rect 22897 887 22931 903
rect 22897 703 22931 719
rect 23005 887 23039 903
rect 23005 703 23039 719
rect 23515 887 23549 903
rect 23515 703 23549 719
rect 22455 657 22471 691
rect 22847 657 22863 691
rect 23073 657 23089 691
rect 23465 657 23481 691
rect 22053 557 22283 619
rect 23687 619 23849 987
rect 25253 987 25483 1049
rect 24055 915 24071 949
rect 24447 915 24463 949
rect 24673 915 24689 949
rect 25065 915 25081 949
rect 23987 887 24021 903
rect 23987 703 24021 719
rect 24497 887 24531 903
rect 24497 703 24531 719
rect 24605 887 24639 903
rect 24605 703 24639 719
rect 25115 887 25149 903
rect 25115 703 25149 719
rect 24055 657 24071 691
rect 24447 657 24463 691
rect 24673 657 24689 691
rect 25065 657 25081 691
rect 23653 557 23883 619
rect 25287 619 25449 987
rect 26853 987 27083 1049
rect 25655 915 25671 949
rect 26047 915 26063 949
rect 26273 915 26289 949
rect 26665 915 26681 949
rect 25587 887 25621 903
rect 25587 703 25621 719
rect 26097 887 26131 903
rect 26097 703 26131 719
rect 26205 887 26239 903
rect 26205 703 26239 719
rect 26715 887 26749 903
rect 26715 703 26749 719
rect 25655 657 25671 691
rect 26047 657 26063 691
rect 26273 657 26289 691
rect 26665 657 26681 691
rect 25253 557 25483 619
rect 26887 619 27049 987
rect 28453 987 28683 1049
rect 27255 915 27271 949
rect 27647 915 27663 949
rect 27873 915 27889 949
rect 28265 915 28281 949
rect 27187 887 27221 903
rect 27187 703 27221 719
rect 27697 887 27731 903
rect 27697 703 27731 719
rect 27805 887 27839 903
rect 27805 703 27839 719
rect 28315 887 28349 903
rect 28315 703 28349 719
rect 27255 657 27271 691
rect 27647 657 27663 691
rect 27873 657 27889 691
rect 28265 657 28281 691
rect 26853 557 27083 619
rect 28487 619 28649 987
rect 30053 987 30283 1049
rect 28855 915 28871 949
rect 29247 915 29263 949
rect 29473 915 29489 949
rect 29865 915 29881 949
rect 28787 887 28821 903
rect 28787 703 28821 719
rect 29297 887 29331 903
rect 29297 703 29331 719
rect 29405 887 29439 903
rect 29405 703 29439 719
rect 29915 887 29949 903
rect 29915 703 29949 719
rect 28855 657 28871 691
rect 29247 657 29263 691
rect 29473 657 29489 691
rect 29865 657 29881 691
rect 28453 557 28683 619
rect 30087 619 30249 987
rect 31653 987 31883 1049
rect 30455 915 30471 949
rect 30847 915 30863 949
rect 31073 915 31089 949
rect 31465 915 31481 949
rect 30387 887 30421 903
rect 30387 703 30421 719
rect 30897 887 30931 903
rect 30897 703 30931 719
rect 31005 887 31039 903
rect 31005 703 31039 719
rect 31515 887 31549 903
rect 31515 703 31549 719
rect 30455 657 30471 691
rect 30847 657 30863 691
rect 31073 657 31089 691
rect 31465 657 31481 691
rect 30053 557 30283 619
rect 31687 619 31849 987
rect 33253 987 33483 1049
rect 32055 915 32071 949
rect 32447 915 32463 949
rect 32673 915 32689 949
rect 33065 915 33081 949
rect 31987 887 32021 903
rect 31987 703 32021 719
rect 32497 887 32531 903
rect 32497 703 32531 719
rect 32605 887 32639 903
rect 32605 703 32639 719
rect 33115 887 33149 903
rect 33115 703 33149 719
rect 32055 657 32071 691
rect 32447 657 32463 691
rect 32673 657 32689 691
rect 33065 657 33081 691
rect 31653 557 31883 619
rect 33287 619 33449 987
rect 34853 987 35083 1049
rect 33655 915 33671 949
rect 34047 915 34063 949
rect 34273 915 34289 949
rect 34665 915 34681 949
rect 33587 887 33621 903
rect 33587 703 33621 719
rect 34097 887 34131 903
rect 34097 703 34131 719
rect 34205 887 34239 903
rect 34205 703 34239 719
rect 34715 887 34749 903
rect 34715 703 34749 719
rect 33655 657 33671 691
rect 34047 657 34063 691
rect 34273 657 34289 691
rect 34665 657 34681 691
rect 33253 557 33483 619
rect 34887 619 35049 987
rect 36453 987 36683 1049
rect 35255 915 35271 949
rect 35647 915 35663 949
rect 35873 915 35889 949
rect 36265 915 36281 949
rect 35187 887 35221 903
rect 35187 703 35221 719
rect 35697 887 35731 903
rect 35697 703 35731 719
rect 35805 887 35839 903
rect 35805 703 35839 719
rect 36315 887 36349 903
rect 36315 703 36349 719
rect 35255 657 35271 691
rect 35647 657 35663 691
rect 35873 657 35889 691
rect 36265 657 36281 691
rect 34853 557 35083 619
rect 36487 619 36649 987
rect 38053 987 38400 1049
rect 36855 915 36871 949
rect 37247 915 37263 949
rect 37473 915 37489 949
rect 37865 915 37881 949
rect 36787 887 36821 903
rect 36787 703 36821 719
rect 37297 887 37331 903
rect 37297 703 37331 719
rect 37405 887 37439 903
rect 37405 703 37439 719
rect 37915 887 37949 903
rect 37915 703 37949 719
rect 36855 657 36871 691
rect 37247 657 37263 691
rect 37473 657 37489 691
rect 37865 657 37881 691
rect 36453 557 36683 619
rect 38087 619 38400 987
rect 38053 557 38400 619
rect -300 429 38400 557
rect -300 395 -117 429
rect 1253 395 1483 429
rect -300 333 0 395
rect -300 -635 -151 333
rect -117 249 0 333
rect 180 295 340 395
rect 55 261 71 295
rect 447 261 463 295
rect 520 249 620 395
rect 800 295 960 395
rect 1140 333 1483 395
rect 673 261 689 295
rect 1065 261 1081 295
rect 1140 249 1253 333
rect -117 233 21 249
rect -117 -535 -13 233
rect -117 -551 21 -535
rect 497 233 639 249
rect 531 -535 605 233
rect 497 -551 639 -535
rect 1115 233 1253 249
rect 1149 -535 1253 233
rect 1115 -551 1253 -535
rect -117 -635 0 -551
rect 55 -597 71 -563
rect 447 -597 463 -563
rect -300 -680 0 -635
rect 180 -680 340 -597
rect 520 -680 620 -551
rect 673 -597 689 -563
rect 1065 -597 1081 -563
rect 800 -680 960 -597
rect 1140 -635 1253 -551
rect 1287 -635 1449 333
rect 2853 333 3083 429
rect 1655 261 1671 295
rect 2047 261 2063 295
rect 2273 261 2289 295
rect 2665 261 2681 295
rect 1587 233 1621 249
rect 1587 -551 1621 -535
rect 2097 233 2131 249
rect 2097 -551 2131 -535
rect 2205 233 2239 249
rect 2205 -551 2239 -535
rect 2715 233 2749 249
rect 2715 -551 2749 -535
rect 1655 -597 1671 -563
rect 2047 -597 2063 -563
rect 2273 -597 2289 -563
rect 2665 -597 2681 -563
rect 1140 -680 1483 -635
rect -300 -697 1483 -680
rect 2887 -635 3049 333
rect 4453 333 4683 429
rect 3255 261 3271 295
rect 3647 261 3663 295
rect 3873 261 3889 295
rect 4265 261 4281 295
rect 3187 233 3221 249
rect 3187 -551 3221 -535
rect 3697 233 3731 249
rect 3697 -551 3731 -535
rect 3805 233 3839 249
rect 3805 -551 3839 -535
rect 4315 233 4349 249
rect 4315 -551 4349 -535
rect 3255 -597 3271 -563
rect 3647 -597 3663 -563
rect 3873 -597 3889 -563
rect 4265 -597 4281 -563
rect 2853 -697 3083 -635
rect 4487 -635 4649 333
rect 6053 333 6283 429
rect 4855 261 4871 295
rect 5247 261 5263 295
rect 5473 261 5489 295
rect 5865 261 5881 295
rect 4787 233 4821 249
rect 4787 -551 4821 -535
rect 5297 233 5331 249
rect 5297 -551 5331 -535
rect 5405 233 5439 249
rect 5405 -551 5439 -535
rect 5915 233 5949 249
rect 5915 -551 5949 -535
rect 4855 -597 4871 -563
rect 5247 -597 5263 -563
rect 5473 -597 5489 -563
rect 5865 -597 5881 -563
rect 4453 -697 4683 -635
rect 6087 -635 6249 333
rect 7653 333 7883 429
rect 6455 261 6471 295
rect 6847 261 6863 295
rect 7073 261 7089 295
rect 7465 261 7481 295
rect 6387 233 6421 249
rect 6387 -551 6421 -535
rect 6897 233 6931 249
rect 6897 -551 6931 -535
rect 7005 233 7039 249
rect 7005 -551 7039 -535
rect 7515 233 7549 249
rect 7515 -551 7549 -535
rect 6455 -597 6471 -563
rect 6847 -597 6863 -563
rect 7073 -597 7089 -563
rect 7465 -597 7481 -563
rect 6053 -697 6283 -635
rect 7687 -635 7849 333
rect 9253 333 9483 429
rect 8055 261 8071 295
rect 8447 261 8463 295
rect 8673 261 8689 295
rect 9065 261 9081 295
rect 7987 233 8021 249
rect 7987 -551 8021 -535
rect 8497 233 8531 249
rect 8497 -551 8531 -535
rect 8605 233 8639 249
rect 8605 -551 8639 -535
rect 9115 233 9149 249
rect 9115 -551 9149 -535
rect 8055 -597 8071 -563
rect 8447 -597 8463 -563
rect 8673 -597 8689 -563
rect 9065 -597 9081 -563
rect 7653 -697 7883 -635
rect 9287 -635 9449 333
rect 10853 333 11083 429
rect 9655 261 9671 295
rect 10047 261 10063 295
rect 10273 261 10289 295
rect 10665 261 10681 295
rect 9587 233 9621 249
rect 9587 -551 9621 -535
rect 10097 233 10131 249
rect 10097 -551 10131 -535
rect 10205 233 10239 249
rect 10205 -551 10239 -535
rect 10715 233 10749 249
rect 10715 -551 10749 -535
rect 9655 -597 9671 -563
rect 10047 -597 10063 -563
rect 10273 -597 10289 -563
rect 10665 -597 10681 -563
rect 9253 -697 9483 -635
rect 10887 -635 11049 333
rect 12453 333 12683 429
rect 11255 261 11271 295
rect 11647 261 11663 295
rect 11873 261 11889 295
rect 12265 261 12281 295
rect 11187 233 11221 249
rect 11187 -551 11221 -535
rect 11697 233 11731 249
rect 11697 -551 11731 -535
rect 11805 233 11839 249
rect 11805 -551 11839 -535
rect 12315 233 12349 249
rect 12315 -551 12349 -535
rect 11255 -597 11271 -563
rect 11647 -597 11663 -563
rect 11873 -597 11889 -563
rect 12265 -597 12281 -563
rect 10853 -697 11083 -635
rect 12487 -635 12649 333
rect 14053 333 14283 429
rect 12855 261 12871 295
rect 13247 261 13263 295
rect 13473 261 13489 295
rect 13865 261 13881 295
rect 12787 233 12821 249
rect 12787 -551 12821 -535
rect 13297 233 13331 249
rect 13297 -551 13331 -535
rect 13405 233 13439 249
rect 13405 -551 13439 -535
rect 13915 233 13949 249
rect 13915 -551 13949 -535
rect 12855 -597 12871 -563
rect 13247 -597 13263 -563
rect 13473 -597 13489 -563
rect 13865 -597 13881 -563
rect 12453 -697 12683 -635
rect 14087 -635 14249 333
rect 15653 333 15883 429
rect 14455 261 14471 295
rect 14847 261 14863 295
rect 15073 261 15089 295
rect 15465 261 15481 295
rect 14387 233 14421 249
rect 14387 -551 14421 -535
rect 14897 233 14931 249
rect 14897 -551 14931 -535
rect 15005 233 15039 249
rect 15005 -551 15039 -535
rect 15515 233 15549 249
rect 15515 -551 15549 -535
rect 14455 -597 14471 -563
rect 14847 -597 14863 -563
rect 15073 -597 15089 -563
rect 15465 -597 15481 -563
rect 14053 -697 14283 -635
rect 15687 -635 15849 333
rect 17253 333 17483 429
rect 16055 261 16071 295
rect 16447 261 16463 295
rect 16673 261 16689 295
rect 17065 261 17081 295
rect 15987 233 16021 249
rect 15987 -551 16021 -535
rect 16497 233 16531 249
rect 16497 -551 16531 -535
rect 16605 233 16639 249
rect 16605 -551 16639 -535
rect 17115 233 17149 249
rect 17115 -551 17149 -535
rect 16055 -597 16071 -563
rect 16447 -597 16463 -563
rect 16673 -597 16689 -563
rect 17065 -597 17081 -563
rect 15653 -697 15883 -635
rect 17287 -635 17449 333
rect 18853 333 19083 429
rect 17655 261 17671 295
rect 18047 261 18063 295
rect 18273 261 18289 295
rect 18665 261 18681 295
rect 17587 233 17621 249
rect 17587 -551 17621 -535
rect 18097 233 18131 249
rect 18097 -551 18131 -535
rect 18205 233 18239 249
rect 18205 -551 18239 -535
rect 18715 233 18749 249
rect 18715 -551 18749 -535
rect 17655 -597 17671 -563
rect 18047 -597 18063 -563
rect 18273 -597 18289 -563
rect 18665 -597 18681 -563
rect 17253 -697 17483 -635
rect 18887 -635 19049 333
rect 20453 333 20683 429
rect 19255 261 19271 295
rect 19647 261 19663 295
rect 19873 261 19889 295
rect 20265 261 20281 295
rect 19187 233 19221 249
rect 19187 -551 19221 -535
rect 19697 233 19731 249
rect 19697 -551 19731 -535
rect 19805 233 19839 249
rect 19805 -551 19839 -535
rect 20315 233 20349 249
rect 20315 -551 20349 -535
rect 19255 -597 19271 -563
rect 19647 -597 19663 -563
rect 19873 -597 19889 -563
rect 20265 -597 20281 -563
rect 18853 -697 19083 -635
rect 20487 -635 20649 333
rect 22053 333 22283 429
rect 20855 261 20871 295
rect 21247 261 21263 295
rect 21473 261 21489 295
rect 21865 261 21881 295
rect 20787 233 20821 249
rect 20787 -551 20821 -535
rect 21297 233 21331 249
rect 21297 -551 21331 -535
rect 21405 233 21439 249
rect 21405 -551 21439 -535
rect 21915 233 21949 249
rect 21915 -551 21949 -535
rect 20855 -597 20871 -563
rect 21247 -597 21263 -563
rect 21473 -597 21489 -563
rect 21865 -597 21881 -563
rect 20453 -697 20683 -635
rect 22087 -635 22249 333
rect 23653 333 23883 429
rect 22455 261 22471 295
rect 22847 261 22863 295
rect 23073 261 23089 295
rect 23465 261 23481 295
rect 22387 233 22421 249
rect 22387 -551 22421 -535
rect 22897 233 22931 249
rect 22897 -551 22931 -535
rect 23005 233 23039 249
rect 23005 -551 23039 -535
rect 23515 233 23549 249
rect 23515 -551 23549 -535
rect 22455 -597 22471 -563
rect 22847 -597 22863 -563
rect 23073 -597 23089 -563
rect 23465 -597 23481 -563
rect 22053 -697 22283 -635
rect 23687 -635 23849 333
rect 25253 333 25483 429
rect 24055 261 24071 295
rect 24447 261 24463 295
rect 24673 261 24689 295
rect 25065 261 25081 295
rect 23987 233 24021 249
rect 23987 -551 24021 -535
rect 24497 233 24531 249
rect 24497 -551 24531 -535
rect 24605 233 24639 249
rect 24605 -551 24639 -535
rect 25115 233 25149 249
rect 25115 -551 25149 -535
rect 24055 -597 24071 -563
rect 24447 -597 24463 -563
rect 24673 -597 24689 -563
rect 25065 -597 25081 -563
rect 23653 -697 23883 -635
rect 25287 -635 25449 333
rect 26853 333 27083 429
rect 25655 261 25671 295
rect 26047 261 26063 295
rect 26273 261 26289 295
rect 26665 261 26681 295
rect 25587 233 25621 249
rect 25587 -551 25621 -535
rect 26097 233 26131 249
rect 26097 -551 26131 -535
rect 26205 233 26239 249
rect 26205 -551 26239 -535
rect 26715 233 26749 249
rect 26715 -551 26749 -535
rect 25655 -597 25671 -563
rect 26047 -597 26063 -563
rect 26273 -597 26289 -563
rect 26665 -597 26681 -563
rect 25253 -697 25483 -635
rect 26887 -635 27049 333
rect 28453 333 28683 429
rect 27255 261 27271 295
rect 27647 261 27663 295
rect 27873 261 27889 295
rect 28265 261 28281 295
rect 27187 233 27221 249
rect 27187 -551 27221 -535
rect 27697 233 27731 249
rect 27697 -551 27731 -535
rect 27805 233 27839 249
rect 27805 -551 27839 -535
rect 28315 233 28349 249
rect 28315 -551 28349 -535
rect 27255 -597 27271 -563
rect 27647 -597 27663 -563
rect 27873 -597 27889 -563
rect 28265 -597 28281 -563
rect 26853 -697 27083 -635
rect 28487 -635 28649 333
rect 30053 333 30283 429
rect 28855 261 28871 295
rect 29247 261 29263 295
rect 29473 261 29489 295
rect 29865 261 29881 295
rect 28787 233 28821 249
rect 28787 -551 28821 -535
rect 29297 233 29331 249
rect 29297 -551 29331 -535
rect 29405 233 29439 249
rect 29405 -551 29439 -535
rect 29915 233 29949 249
rect 29915 -551 29949 -535
rect 28855 -597 28871 -563
rect 29247 -597 29263 -563
rect 29473 -597 29489 -563
rect 29865 -597 29881 -563
rect 28453 -697 28683 -635
rect 30087 -635 30249 333
rect 31653 333 31883 429
rect 30455 261 30471 295
rect 30847 261 30863 295
rect 31073 261 31089 295
rect 31465 261 31481 295
rect 30387 233 30421 249
rect 30387 -551 30421 -535
rect 30897 233 30931 249
rect 30897 -551 30931 -535
rect 31005 233 31039 249
rect 31005 -551 31039 -535
rect 31515 233 31549 249
rect 31515 -551 31549 -535
rect 30455 -597 30471 -563
rect 30847 -597 30863 -563
rect 31073 -597 31089 -563
rect 31465 -597 31481 -563
rect 30053 -697 30283 -635
rect 31687 -635 31849 333
rect 33253 333 33483 429
rect 32055 261 32071 295
rect 32447 261 32463 295
rect 32673 261 32689 295
rect 33065 261 33081 295
rect 31987 233 32021 249
rect 31987 -551 32021 -535
rect 32497 233 32531 249
rect 32497 -551 32531 -535
rect 32605 233 32639 249
rect 32605 -551 32639 -535
rect 33115 233 33149 249
rect 33115 -551 33149 -535
rect 32055 -597 32071 -563
rect 32447 -597 32463 -563
rect 32673 -597 32689 -563
rect 33065 -597 33081 -563
rect 31653 -697 31883 -635
rect 33287 -635 33449 333
rect 34853 333 35083 429
rect 36453 395 36683 429
rect 38053 395 38400 429
rect 33655 261 33671 295
rect 34047 261 34063 295
rect 34273 261 34289 295
rect 34665 261 34681 295
rect 33587 233 33621 249
rect 33587 -551 33621 -535
rect 34097 233 34131 249
rect 34097 -551 34131 -535
rect 34205 233 34239 249
rect 34205 -551 34239 -535
rect 34715 233 34749 249
rect 34715 -551 34749 -535
rect 33655 -597 33671 -563
rect 34047 -597 34063 -563
rect 34273 -597 34289 -563
rect 34665 -597 34681 -563
rect 33253 -697 33483 -635
rect 34887 -635 35049 333
rect 36453 333 36800 395
rect 35255 261 35271 295
rect 35647 261 35663 295
rect 35873 261 35889 295
rect 36265 261 36281 295
rect 35187 233 35221 249
rect 35187 -551 35221 -535
rect 35697 233 35731 249
rect 35697 -551 35731 -535
rect 35805 233 35839 249
rect 35805 -551 35839 -535
rect 36315 233 36349 249
rect 36315 -551 36349 -535
rect 35255 -597 35271 -563
rect 35647 -597 35663 -563
rect 35873 -597 35889 -563
rect 36265 -597 36281 -563
rect 34853 -697 35083 -635
rect 36487 -635 36649 333
rect 36683 249 36800 333
rect 36980 295 37140 395
rect 36855 261 36871 295
rect 37247 261 37263 295
rect 37320 249 37420 395
rect 37600 295 37760 395
rect 37940 333 38400 395
rect 37473 261 37489 295
rect 37865 261 37881 295
rect 37940 249 38053 333
rect 36683 233 36821 249
rect 36683 -535 36787 233
rect 36683 -551 36821 -535
rect 37297 233 37439 249
rect 37331 -535 37405 233
rect 37297 -551 37439 -535
rect 37915 233 38053 249
rect 37949 -535 38053 233
rect 37915 -551 38053 -535
rect 36683 -635 36800 -551
rect 36855 -597 36871 -563
rect 37247 -597 37263 -563
rect 36453 -680 36800 -635
rect 36980 -680 37140 -597
rect 37320 -680 37420 -551
rect 37473 -597 37489 -563
rect 37865 -597 37881 -563
rect 37600 -680 37760 -597
rect 37940 -635 38053 -551
rect 38087 -635 38400 333
rect 37940 -680 38400 -635
rect 36453 -697 38400 -680
rect -300 -731 -55 -697
rect 1191 -731 1545 -697
rect 2791 -731 3145 -697
rect 4391 -731 4745 -697
rect 5991 -731 6345 -697
rect 7591 -731 7945 -697
rect 9191 -731 9545 -697
rect 10791 -731 11145 -697
rect 12391 -731 12745 -697
rect 13991 -731 14345 -697
rect 15591 -731 15945 -697
rect 17191 -731 17545 -697
rect 18791 -731 19145 -697
rect 20391 -731 20745 -697
rect 21991 -731 22345 -697
rect 23591 -731 23945 -697
rect 25191 -731 25545 -697
rect 26791 -731 27145 -697
rect 28391 -731 28745 -697
rect 29991 -731 30345 -697
rect 31591 -731 31945 -697
rect 33191 -731 33545 -697
rect 34791 -731 35145 -697
rect 36391 -731 36745 -697
rect 37991 -731 38400 -697
rect -300 -751 38400 -731
rect -300 -780 1483 -751
rect -300 -813 0 -780
rect -300 -1181 -151 -813
rect -117 -897 0 -813
rect 180 -851 340 -780
rect 55 -885 71 -851
rect 447 -885 463 -851
rect 520 -897 620 -780
rect 800 -851 960 -780
rect 1140 -813 1483 -780
rect 673 -885 689 -851
rect 1065 -885 1081 -851
rect 1140 -897 1253 -813
rect -117 -913 21 -897
rect -117 -1081 -13 -913
rect -117 -1097 21 -1081
rect 497 -913 639 -897
rect 531 -1081 605 -913
rect 497 -1097 639 -1081
rect 1115 -913 1253 -897
rect 1149 -1081 1253 -913
rect 1115 -1097 1253 -1081
rect -117 -1181 0 -1097
rect 55 -1143 71 -1109
rect 447 -1143 463 -1109
rect -300 -1243 0 -1181
rect 180 -1243 340 -1143
rect 520 -1243 620 -1097
rect 673 -1143 689 -1109
rect 1065 -1143 1081 -1109
rect 800 -1243 960 -1143
rect 1140 -1181 1253 -1097
rect 1287 -1181 1449 -813
rect 2853 -813 3083 -751
rect 1655 -885 1671 -851
rect 2047 -885 2063 -851
rect 2273 -885 2289 -851
rect 2665 -885 2681 -851
rect 1587 -913 1621 -897
rect 1587 -1097 1621 -1081
rect 2097 -913 2131 -897
rect 2097 -1097 2131 -1081
rect 2205 -913 2239 -897
rect 2205 -1097 2239 -1081
rect 2715 -913 2749 -897
rect 2715 -1097 2749 -1081
rect 1655 -1143 1671 -1109
rect 2047 -1143 2063 -1109
rect 2273 -1143 2289 -1109
rect 2665 -1143 2681 -1109
rect 1140 -1243 1483 -1181
rect 2887 -1181 3049 -813
rect 4453 -813 4683 -751
rect 3255 -885 3271 -851
rect 3647 -885 3663 -851
rect 3873 -885 3889 -851
rect 4265 -885 4281 -851
rect 3187 -913 3221 -897
rect 3187 -1097 3221 -1081
rect 3697 -913 3731 -897
rect 3697 -1097 3731 -1081
rect 3805 -913 3839 -897
rect 3805 -1097 3839 -1081
rect 4315 -913 4349 -897
rect 4315 -1097 4349 -1081
rect 3255 -1143 3271 -1109
rect 3647 -1143 3663 -1109
rect 3873 -1143 3889 -1109
rect 4265 -1143 4281 -1109
rect 2853 -1243 3083 -1181
rect 4487 -1181 4649 -813
rect 6053 -813 6283 -751
rect 4855 -885 4871 -851
rect 5247 -885 5263 -851
rect 5473 -885 5489 -851
rect 5865 -885 5881 -851
rect 4787 -913 4821 -897
rect 4787 -1097 4821 -1081
rect 5297 -913 5331 -897
rect 5297 -1097 5331 -1081
rect 5405 -913 5439 -897
rect 5405 -1097 5439 -1081
rect 5915 -913 5949 -897
rect 5915 -1097 5949 -1081
rect 4855 -1143 4871 -1109
rect 5247 -1143 5263 -1109
rect 5473 -1143 5489 -1109
rect 5865 -1143 5881 -1109
rect 4453 -1243 4683 -1181
rect 6087 -1181 6249 -813
rect 7653 -813 7883 -751
rect 6455 -885 6471 -851
rect 6847 -885 6863 -851
rect 7073 -885 7089 -851
rect 7465 -885 7481 -851
rect 6387 -913 6421 -897
rect 6387 -1097 6421 -1081
rect 6897 -913 6931 -897
rect 6897 -1097 6931 -1081
rect 7005 -913 7039 -897
rect 7005 -1097 7039 -1081
rect 7515 -913 7549 -897
rect 7515 -1097 7549 -1081
rect 6455 -1143 6471 -1109
rect 6847 -1143 6863 -1109
rect 7073 -1143 7089 -1109
rect 7465 -1143 7481 -1109
rect 6053 -1243 6283 -1181
rect 7687 -1181 7849 -813
rect 9253 -813 9483 -751
rect 8055 -885 8071 -851
rect 8447 -885 8463 -851
rect 8673 -885 8689 -851
rect 9065 -885 9081 -851
rect 7987 -913 8021 -897
rect 7987 -1097 8021 -1081
rect 8497 -913 8531 -897
rect 8497 -1097 8531 -1081
rect 8605 -913 8639 -897
rect 8605 -1097 8639 -1081
rect 9115 -913 9149 -897
rect 9115 -1097 9149 -1081
rect 8055 -1143 8071 -1109
rect 8447 -1143 8463 -1109
rect 8673 -1143 8689 -1109
rect 9065 -1143 9081 -1109
rect 7653 -1243 7883 -1181
rect 9287 -1181 9449 -813
rect 10853 -813 11083 -751
rect 9655 -885 9671 -851
rect 10047 -885 10063 -851
rect 10273 -885 10289 -851
rect 10665 -885 10681 -851
rect 9587 -913 9621 -897
rect 9587 -1097 9621 -1081
rect 10097 -913 10131 -897
rect 10097 -1097 10131 -1081
rect 10205 -913 10239 -897
rect 10205 -1097 10239 -1081
rect 10715 -913 10749 -897
rect 10715 -1097 10749 -1081
rect 9655 -1143 9671 -1109
rect 10047 -1143 10063 -1109
rect 10273 -1143 10289 -1109
rect 10665 -1143 10681 -1109
rect 9253 -1243 9483 -1181
rect 10887 -1181 11049 -813
rect 12453 -813 12683 -751
rect 11255 -885 11271 -851
rect 11647 -885 11663 -851
rect 11873 -885 11889 -851
rect 12265 -885 12281 -851
rect 11187 -913 11221 -897
rect 11187 -1097 11221 -1081
rect 11697 -913 11731 -897
rect 11697 -1097 11731 -1081
rect 11805 -913 11839 -897
rect 11805 -1097 11839 -1081
rect 12315 -913 12349 -897
rect 12315 -1097 12349 -1081
rect 11255 -1143 11271 -1109
rect 11647 -1143 11663 -1109
rect 11873 -1143 11889 -1109
rect 12265 -1143 12281 -1109
rect 10853 -1243 11083 -1181
rect 12487 -1181 12649 -813
rect 14053 -813 14283 -751
rect 12855 -885 12871 -851
rect 13247 -885 13263 -851
rect 13473 -885 13489 -851
rect 13865 -885 13881 -851
rect 12787 -913 12821 -897
rect 12787 -1097 12821 -1081
rect 13297 -913 13331 -897
rect 13297 -1097 13331 -1081
rect 13405 -913 13439 -897
rect 13405 -1097 13439 -1081
rect 13915 -913 13949 -897
rect 13915 -1097 13949 -1081
rect 12855 -1143 12871 -1109
rect 13247 -1143 13263 -1109
rect 13473 -1143 13489 -1109
rect 13865 -1143 13881 -1109
rect 12453 -1243 12683 -1181
rect 14087 -1181 14249 -813
rect 15653 -813 15883 -751
rect 14455 -885 14471 -851
rect 14847 -885 14863 -851
rect 15073 -885 15089 -851
rect 15465 -885 15481 -851
rect 14387 -913 14421 -897
rect 14387 -1097 14421 -1081
rect 14897 -913 14931 -897
rect 14897 -1097 14931 -1081
rect 15005 -913 15039 -897
rect 15005 -1097 15039 -1081
rect 15515 -913 15549 -897
rect 15515 -1097 15549 -1081
rect 14455 -1143 14471 -1109
rect 14847 -1143 14863 -1109
rect 15073 -1143 15089 -1109
rect 15465 -1143 15481 -1109
rect 14053 -1243 14283 -1181
rect 15687 -1181 15849 -813
rect 17253 -813 17483 -751
rect 16055 -885 16071 -851
rect 16447 -885 16463 -851
rect 16673 -885 16689 -851
rect 17065 -885 17081 -851
rect 15987 -913 16021 -897
rect 15987 -1097 16021 -1081
rect 16497 -913 16531 -897
rect 16497 -1097 16531 -1081
rect 16605 -913 16639 -897
rect 16605 -1097 16639 -1081
rect 17115 -913 17149 -897
rect 17115 -1097 17149 -1081
rect 16055 -1143 16071 -1109
rect 16447 -1143 16463 -1109
rect 16673 -1143 16689 -1109
rect 17065 -1143 17081 -1109
rect 15653 -1243 15883 -1181
rect 17287 -1181 17449 -813
rect 18853 -813 19083 -751
rect 17655 -885 17671 -851
rect 18047 -885 18063 -851
rect 18273 -885 18289 -851
rect 18665 -885 18681 -851
rect 17587 -913 17621 -897
rect 17587 -1097 17621 -1081
rect 18097 -913 18131 -897
rect 18097 -1097 18131 -1081
rect 18205 -913 18239 -897
rect 18205 -1097 18239 -1081
rect 18715 -913 18749 -897
rect 18715 -1097 18749 -1081
rect 17655 -1143 17671 -1109
rect 18047 -1143 18063 -1109
rect 18273 -1143 18289 -1109
rect 18665 -1143 18681 -1109
rect 17253 -1243 17483 -1181
rect 18887 -1181 19049 -813
rect 20453 -813 20683 -751
rect 19255 -885 19271 -851
rect 19647 -885 19663 -851
rect 19873 -885 19889 -851
rect 20265 -885 20281 -851
rect 19187 -913 19221 -897
rect 19187 -1097 19221 -1081
rect 19697 -913 19731 -897
rect 19697 -1097 19731 -1081
rect 19805 -913 19839 -897
rect 19805 -1097 19839 -1081
rect 20315 -913 20349 -897
rect 20315 -1097 20349 -1081
rect 19255 -1143 19271 -1109
rect 19647 -1143 19663 -1109
rect 19873 -1143 19889 -1109
rect 20265 -1143 20281 -1109
rect 18853 -1243 19083 -1181
rect 20487 -1181 20649 -813
rect 22053 -813 22283 -751
rect 20855 -885 20871 -851
rect 21247 -885 21263 -851
rect 21473 -885 21489 -851
rect 21865 -885 21881 -851
rect 20787 -913 20821 -897
rect 20787 -1097 20821 -1081
rect 21297 -913 21331 -897
rect 21297 -1097 21331 -1081
rect 21405 -913 21439 -897
rect 21405 -1097 21439 -1081
rect 21915 -913 21949 -897
rect 21915 -1097 21949 -1081
rect 20855 -1143 20871 -1109
rect 21247 -1143 21263 -1109
rect 21473 -1143 21489 -1109
rect 21865 -1143 21881 -1109
rect 20453 -1243 20683 -1181
rect 22087 -1181 22249 -813
rect 23653 -813 23883 -751
rect 22455 -885 22471 -851
rect 22847 -885 22863 -851
rect 23073 -885 23089 -851
rect 23465 -885 23481 -851
rect 22387 -913 22421 -897
rect 22387 -1097 22421 -1081
rect 22897 -913 22931 -897
rect 22897 -1097 22931 -1081
rect 23005 -913 23039 -897
rect 23005 -1097 23039 -1081
rect 23515 -913 23549 -897
rect 23515 -1097 23549 -1081
rect 22455 -1143 22471 -1109
rect 22847 -1143 22863 -1109
rect 23073 -1143 23089 -1109
rect 23465 -1143 23481 -1109
rect 22053 -1243 22283 -1181
rect 23687 -1181 23849 -813
rect 25253 -813 25483 -751
rect 24055 -885 24071 -851
rect 24447 -885 24463 -851
rect 24673 -885 24689 -851
rect 25065 -885 25081 -851
rect 23987 -913 24021 -897
rect 23987 -1097 24021 -1081
rect 24497 -913 24531 -897
rect 24497 -1097 24531 -1081
rect 24605 -913 24639 -897
rect 24605 -1097 24639 -1081
rect 25115 -913 25149 -897
rect 25115 -1097 25149 -1081
rect 24055 -1143 24071 -1109
rect 24447 -1143 24463 -1109
rect 24673 -1143 24689 -1109
rect 25065 -1143 25081 -1109
rect 23653 -1243 23883 -1181
rect 25287 -1181 25449 -813
rect 26853 -813 27083 -751
rect 25655 -885 25671 -851
rect 26047 -885 26063 -851
rect 26273 -885 26289 -851
rect 26665 -885 26681 -851
rect 25587 -913 25621 -897
rect 25587 -1097 25621 -1081
rect 26097 -913 26131 -897
rect 26097 -1097 26131 -1081
rect 26205 -913 26239 -897
rect 26205 -1097 26239 -1081
rect 26715 -913 26749 -897
rect 26715 -1097 26749 -1081
rect 25655 -1143 25671 -1109
rect 26047 -1143 26063 -1109
rect 26273 -1143 26289 -1109
rect 26665 -1143 26681 -1109
rect 25253 -1243 25483 -1181
rect 26887 -1181 27049 -813
rect 28453 -813 28683 -751
rect 27255 -885 27271 -851
rect 27647 -885 27663 -851
rect 27873 -885 27889 -851
rect 28265 -885 28281 -851
rect 27187 -913 27221 -897
rect 27187 -1097 27221 -1081
rect 27697 -913 27731 -897
rect 27697 -1097 27731 -1081
rect 27805 -913 27839 -897
rect 27805 -1097 27839 -1081
rect 28315 -913 28349 -897
rect 28315 -1097 28349 -1081
rect 27255 -1143 27271 -1109
rect 27647 -1143 27663 -1109
rect 27873 -1143 27889 -1109
rect 28265 -1143 28281 -1109
rect 26853 -1243 27083 -1181
rect 28487 -1181 28649 -813
rect 30053 -813 30283 -751
rect 28855 -885 28871 -851
rect 29247 -885 29263 -851
rect 29473 -885 29489 -851
rect 29865 -885 29881 -851
rect 28787 -913 28821 -897
rect 28787 -1097 28821 -1081
rect 29297 -913 29331 -897
rect 29297 -1097 29331 -1081
rect 29405 -913 29439 -897
rect 29405 -1097 29439 -1081
rect 29915 -913 29949 -897
rect 29915 -1097 29949 -1081
rect 28855 -1143 28871 -1109
rect 29247 -1143 29263 -1109
rect 29473 -1143 29489 -1109
rect 29865 -1143 29881 -1109
rect 28453 -1243 28683 -1181
rect 30087 -1181 30249 -813
rect 31653 -813 31883 -751
rect 30455 -885 30471 -851
rect 30847 -885 30863 -851
rect 31073 -885 31089 -851
rect 31465 -885 31481 -851
rect 30387 -913 30421 -897
rect 30387 -1097 30421 -1081
rect 30897 -913 30931 -897
rect 30897 -1097 30931 -1081
rect 31005 -913 31039 -897
rect 31005 -1097 31039 -1081
rect 31515 -913 31549 -897
rect 31515 -1097 31549 -1081
rect 30455 -1143 30471 -1109
rect 30847 -1143 30863 -1109
rect 31073 -1143 31089 -1109
rect 31465 -1143 31481 -1109
rect 30053 -1243 30283 -1181
rect 31687 -1181 31849 -813
rect 33253 -813 33483 -751
rect 32055 -885 32071 -851
rect 32447 -885 32463 -851
rect 32673 -885 32689 -851
rect 33065 -885 33081 -851
rect 31987 -913 32021 -897
rect 31987 -1097 32021 -1081
rect 32497 -913 32531 -897
rect 32497 -1097 32531 -1081
rect 32605 -913 32639 -897
rect 32605 -1097 32639 -1081
rect 33115 -913 33149 -897
rect 33115 -1097 33149 -1081
rect 32055 -1143 32071 -1109
rect 32447 -1143 32463 -1109
rect 32673 -1143 32689 -1109
rect 33065 -1143 33081 -1109
rect 31653 -1243 31883 -1181
rect 33287 -1181 33449 -813
rect 34853 -813 35083 -751
rect 33655 -885 33671 -851
rect 34047 -885 34063 -851
rect 34273 -885 34289 -851
rect 34665 -885 34681 -851
rect 33587 -913 33621 -897
rect 33587 -1097 33621 -1081
rect 34097 -913 34131 -897
rect 34097 -1097 34131 -1081
rect 34205 -913 34239 -897
rect 34205 -1097 34239 -1081
rect 34715 -913 34749 -897
rect 34715 -1097 34749 -1081
rect 33655 -1143 33671 -1109
rect 34047 -1143 34063 -1109
rect 34273 -1143 34289 -1109
rect 34665 -1143 34681 -1109
rect 33253 -1243 33483 -1181
rect 34887 -1181 35049 -813
rect 36453 -780 38400 -751
rect 36453 -813 36800 -780
rect 35255 -885 35271 -851
rect 35647 -885 35663 -851
rect 35873 -885 35889 -851
rect 36265 -885 36281 -851
rect 35187 -913 35221 -897
rect 35187 -1097 35221 -1081
rect 35697 -913 35731 -897
rect 35697 -1097 35731 -1081
rect 35805 -913 35839 -897
rect 35805 -1097 35839 -1081
rect 36315 -913 36349 -897
rect 36315 -1097 36349 -1081
rect 35255 -1143 35271 -1109
rect 35647 -1143 35663 -1109
rect 35873 -1143 35889 -1109
rect 36265 -1143 36281 -1109
rect 34853 -1243 35083 -1181
rect 36487 -1181 36649 -813
rect 36683 -897 36800 -813
rect 36980 -851 37140 -780
rect 36855 -885 36871 -851
rect 37247 -885 37263 -851
rect 37320 -897 37420 -780
rect 37600 -851 37760 -780
rect 37940 -813 38400 -780
rect 37473 -885 37489 -851
rect 37865 -885 37881 -851
rect 37940 -897 38053 -813
rect 36683 -913 36821 -897
rect 36683 -1081 36787 -913
rect 36683 -1097 36821 -1081
rect 37297 -913 37439 -897
rect 37331 -1081 37405 -913
rect 37297 -1097 37439 -1081
rect 37915 -913 38053 -897
rect 37949 -1081 38053 -913
rect 37915 -1097 38053 -1081
rect 36683 -1181 36800 -1097
rect 36855 -1143 36871 -1109
rect 37247 -1143 37263 -1109
rect 36453 -1243 36800 -1181
rect 36980 -1243 37140 -1143
rect 37320 -1243 37420 -1097
rect 37473 -1143 37489 -1109
rect 37865 -1143 37881 -1109
rect 37600 -1243 37760 -1143
rect 37940 -1181 38053 -1097
rect 38087 -1181 38400 -813
rect 37940 -1243 38400 -1181
rect -300 -1371 38400 -1243
rect -300 -1405 -117 -1371
rect 1253 -1405 1483 -1371
rect -300 -1467 0 -1405
rect -300 -2435 -151 -1467
rect -117 -1551 0 -1467
rect 180 -1505 340 -1405
rect 55 -1539 71 -1505
rect 447 -1539 463 -1505
rect 520 -1551 620 -1405
rect 800 -1505 960 -1405
rect 1140 -1467 1483 -1405
rect 673 -1539 689 -1505
rect 1065 -1539 1081 -1505
rect 1140 -1551 1253 -1467
rect -117 -1567 21 -1551
rect -117 -2335 -13 -1567
rect -117 -2351 21 -2335
rect 497 -1567 639 -1551
rect 531 -2335 605 -1567
rect 497 -2351 639 -2335
rect 1115 -1567 1253 -1551
rect 1149 -2335 1253 -1567
rect 1115 -2351 1253 -2335
rect -117 -2435 0 -2351
rect 55 -2397 71 -2363
rect 447 -2397 463 -2363
rect -300 -2480 0 -2435
rect 180 -2480 340 -2397
rect 520 -2480 620 -2351
rect 673 -2397 689 -2363
rect 1065 -2397 1081 -2363
rect 800 -2480 960 -2397
rect 1140 -2435 1253 -2351
rect 1287 -2435 1449 -1467
rect 2853 -1467 3083 -1371
rect 1655 -1539 1671 -1505
rect 2047 -1539 2063 -1505
rect 2273 -1539 2289 -1505
rect 2665 -1539 2681 -1505
rect 1587 -1567 1621 -1551
rect 1587 -2351 1621 -2335
rect 2097 -1567 2131 -1551
rect 2097 -2351 2131 -2335
rect 2205 -1567 2239 -1551
rect 2205 -2351 2239 -2335
rect 2715 -1567 2749 -1551
rect 2715 -2351 2749 -2335
rect 1655 -2397 1671 -2363
rect 2047 -2397 2063 -2363
rect 2273 -2397 2289 -2363
rect 2665 -2397 2681 -2363
rect 1140 -2480 1483 -2435
rect -300 -2497 1483 -2480
rect 2887 -2435 3049 -1467
rect 4453 -1467 4683 -1371
rect 3255 -1539 3271 -1505
rect 3647 -1539 3663 -1505
rect 3873 -1539 3889 -1505
rect 4265 -1539 4281 -1505
rect 3187 -1567 3221 -1551
rect 3187 -2351 3221 -2335
rect 3697 -1567 3731 -1551
rect 3697 -2351 3731 -2335
rect 3805 -1567 3839 -1551
rect 3805 -2351 3839 -2335
rect 4315 -1567 4349 -1551
rect 4315 -2351 4349 -2335
rect 3255 -2397 3271 -2363
rect 3647 -2397 3663 -2363
rect 3873 -2397 3889 -2363
rect 4265 -2397 4281 -2363
rect 2853 -2497 3083 -2435
rect 4487 -2435 4649 -1467
rect 6053 -1467 6283 -1371
rect 4855 -1539 4871 -1505
rect 5247 -1539 5263 -1505
rect 5473 -1539 5489 -1505
rect 5865 -1539 5881 -1505
rect 4787 -1567 4821 -1551
rect 4787 -2351 4821 -2335
rect 5297 -1567 5331 -1551
rect 5297 -2351 5331 -2335
rect 5405 -1567 5439 -1551
rect 5405 -2351 5439 -2335
rect 5915 -1567 5949 -1551
rect 5915 -2351 5949 -2335
rect 4855 -2397 4871 -2363
rect 5247 -2397 5263 -2363
rect 5473 -2397 5489 -2363
rect 5865 -2397 5881 -2363
rect 4453 -2497 4683 -2435
rect 6087 -2435 6249 -1467
rect 7653 -1467 7883 -1371
rect 6455 -1539 6471 -1505
rect 6847 -1539 6863 -1505
rect 7073 -1539 7089 -1505
rect 7465 -1539 7481 -1505
rect 6387 -1567 6421 -1551
rect 6387 -2351 6421 -2335
rect 6897 -1567 6931 -1551
rect 6897 -2351 6931 -2335
rect 7005 -1567 7039 -1551
rect 7005 -2351 7039 -2335
rect 7515 -1567 7549 -1551
rect 7515 -2351 7549 -2335
rect 6455 -2397 6471 -2363
rect 6847 -2397 6863 -2363
rect 7073 -2397 7089 -2363
rect 7465 -2397 7481 -2363
rect 6053 -2497 6283 -2435
rect 7687 -2435 7849 -1467
rect 9253 -1467 9483 -1371
rect 8055 -1539 8071 -1505
rect 8447 -1539 8463 -1505
rect 8673 -1539 8689 -1505
rect 9065 -1539 9081 -1505
rect 7987 -1567 8021 -1551
rect 7987 -2351 8021 -2335
rect 8497 -1567 8531 -1551
rect 8497 -2351 8531 -2335
rect 8605 -1567 8639 -1551
rect 8605 -2351 8639 -2335
rect 9115 -1567 9149 -1551
rect 9115 -2351 9149 -2335
rect 8055 -2397 8071 -2363
rect 8447 -2397 8463 -2363
rect 8673 -2397 8689 -2363
rect 9065 -2397 9081 -2363
rect 7653 -2497 7883 -2435
rect 9287 -2435 9449 -1467
rect 10853 -1467 11083 -1371
rect 9655 -1539 9671 -1505
rect 10047 -1539 10063 -1505
rect 10273 -1539 10289 -1505
rect 10665 -1539 10681 -1505
rect 9587 -1567 9621 -1551
rect 9587 -2351 9621 -2335
rect 10097 -1567 10131 -1551
rect 10097 -2351 10131 -2335
rect 10205 -1567 10239 -1551
rect 10205 -2351 10239 -2335
rect 10715 -1567 10749 -1551
rect 10715 -2351 10749 -2335
rect 9655 -2397 9671 -2363
rect 10047 -2397 10063 -2363
rect 10273 -2397 10289 -2363
rect 10665 -2397 10681 -2363
rect 9253 -2497 9483 -2435
rect 10887 -2435 11049 -1467
rect 12453 -1467 12683 -1371
rect 11255 -1539 11271 -1505
rect 11647 -1539 11663 -1505
rect 11873 -1539 11889 -1505
rect 12265 -1539 12281 -1505
rect 11187 -1567 11221 -1551
rect 11187 -2351 11221 -2335
rect 11697 -1567 11731 -1551
rect 11697 -2351 11731 -2335
rect 11805 -1567 11839 -1551
rect 11805 -2351 11839 -2335
rect 12315 -1567 12349 -1551
rect 12315 -2351 12349 -2335
rect 11255 -2397 11271 -2363
rect 11647 -2397 11663 -2363
rect 11873 -2397 11889 -2363
rect 12265 -2397 12281 -2363
rect 10853 -2497 11083 -2435
rect 12487 -2435 12649 -1467
rect 14053 -1467 14283 -1371
rect 12855 -1539 12871 -1505
rect 13247 -1539 13263 -1505
rect 13473 -1539 13489 -1505
rect 13865 -1539 13881 -1505
rect 12787 -1567 12821 -1551
rect 12787 -2351 12821 -2335
rect 13297 -1567 13331 -1551
rect 13297 -2351 13331 -2335
rect 13405 -1567 13439 -1551
rect 13405 -2351 13439 -2335
rect 13915 -1567 13949 -1551
rect 13915 -2351 13949 -2335
rect 12855 -2397 12871 -2363
rect 13247 -2397 13263 -2363
rect 13473 -2397 13489 -2363
rect 13865 -2397 13881 -2363
rect 12453 -2497 12683 -2435
rect 14087 -2435 14249 -1467
rect 15653 -1467 15883 -1371
rect 14455 -1539 14471 -1505
rect 14847 -1539 14863 -1505
rect 15073 -1539 15089 -1505
rect 15465 -1539 15481 -1505
rect 14387 -1567 14421 -1551
rect 14387 -2351 14421 -2335
rect 14897 -1567 14931 -1551
rect 14897 -2351 14931 -2335
rect 15005 -1567 15039 -1551
rect 15005 -2351 15039 -2335
rect 15515 -1567 15549 -1551
rect 15515 -2351 15549 -2335
rect 14455 -2397 14471 -2363
rect 14847 -2397 14863 -2363
rect 15073 -2397 15089 -2363
rect 15465 -2397 15481 -2363
rect 14053 -2497 14283 -2435
rect 15687 -2435 15849 -1467
rect 17253 -1467 17483 -1371
rect 16055 -1539 16071 -1505
rect 16447 -1539 16463 -1505
rect 16673 -1539 16689 -1505
rect 17065 -1539 17081 -1505
rect 15987 -1567 16021 -1551
rect 15987 -2351 16021 -2335
rect 16497 -1567 16531 -1551
rect 16497 -2351 16531 -2335
rect 16605 -1567 16639 -1551
rect 16605 -2351 16639 -2335
rect 17115 -1567 17149 -1551
rect 17115 -2351 17149 -2335
rect 16055 -2397 16071 -2363
rect 16447 -2397 16463 -2363
rect 16673 -2397 16689 -2363
rect 17065 -2397 17081 -2363
rect 15653 -2497 15883 -2435
rect 17287 -2435 17449 -1467
rect 18853 -1467 19083 -1371
rect 17655 -1539 17671 -1505
rect 18047 -1539 18063 -1505
rect 18273 -1539 18289 -1505
rect 18665 -1539 18681 -1505
rect 17587 -1567 17621 -1551
rect 17587 -2351 17621 -2335
rect 18097 -1567 18131 -1551
rect 18097 -2351 18131 -2335
rect 18205 -1567 18239 -1551
rect 18205 -2351 18239 -2335
rect 18715 -1567 18749 -1551
rect 18715 -2351 18749 -2335
rect 17655 -2397 17671 -2363
rect 18047 -2397 18063 -2363
rect 18273 -2397 18289 -2363
rect 18665 -2397 18681 -2363
rect 17253 -2497 17483 -2435
rect 18887 -2435 19049 -1467
rect 20453 -1467 20683 -1371
rect 19255 -1539 19271 -1505
rect 19647 -1539 19663 -1505
rect 19873 -1539 19889 -1505
rect 20265 -1539 20281 -1505
rect 19187 -1567 19221 -1551
rect 19187 -2351 19221 -2335
rect 19697 -1567 19731 -1551
rect 19697 -2351 19731 -2335
rect 19805 -1567 19839 -1551
rect 19805 -2351 19839 -2335
rect 20315 -1567 20349 -1551
rect 20315 -2351 20349 -2335
rect 19255 -2397 19271 -2363
rect 19647 -2397 19663 -2363
rect 19873 -2397 19889 -2363
rect 20265 -2397 20281 -2363
rect 18853 -2497 19083 -2435
rect 20487 -2435 20649 -1467
rect 22053 -1467 22283 -1371
rect 20855 -1539 20871 -1505
rect 21247 -1539 21263 -1505
rect 21473 -1539 21489 -1505
rect 21865 -1539 21881 -1505
rect 20787 -1567 20821 -1551
rect 20787 -2351 20821 -2335
rect 21297 -1567 21331 -1551
rect 21297 -2351 21331 -2335
rect 21405 -1567 21439 -1551
rect 21405 -2351 21439 -2335
rect 21915 -1567 21949 -1551
rect 21915 -2351 21949 -2335
rect 20855 -2397 20871 -2363
rect 21247 -2397 21263 -2363
rect 21473 -2397 21489 -2363
rect 21865 -2397 21881 -2363
rect 20453 -2497 20683 -2435
rect 22087 -2435 22249 -1467
rect 23653 -1467 23883 -1371
rect 22455 -1539 22471 -1505
rect 22847 -1539 22863 -1505
rect 23073 -1539 23089 -1505
rect 23465 -1539 23481 -1505
rect 22387 -1567 22421 -1551
rect 22387 -2351 22421 -2335
rect 22897 -1567 22931 -1551
rect 22897 -2351 22931 -2335
rect 23005 -1567 23039 -1551
rect 23005 -2351 23039 -2335
rect 23515 -1567 23549 -1551
rect 23515 -2351 23549 -2335
rect 22455 -2397 22471 -2363
rect 22847 -2397 22863 -2363
rect 23073 -2397 23089 -2363
rect 23465 -2397 23481 -2363
rect 22053 -2497 22283 -2435
rect 23687 -2435 23849 -1467
rect 25253 -1467 25483 -1371
rect 24055 -1539 24071 -1505
rect 24447 -1539 24463 -1505
rect 24673 -1539 24689 -1505
rect 25065 -1539 25081 -1505
rect 23987 -1567 24021 -1551
rect 23987 -2351 24021 -2335
rect 24497 -1567 24531 -1551
rect 24497 -2351 24531 -2335
rect 24605 -1567 24639 -1551
rect 24605 -2351 24639 -2335
rect 25115 -1567 25149 -1551
rect 25115 -2351 25149 -2335
rect 24055 -2397 24071 -2363
rect 24447 -2397 24463 -2363
rect 24673 -2397 24689 -2363
rect 25065 -2397 25081 -2363
rect 23653 -2497 23883 -2435
rect 25287 -2435 25449 -1467
rect 26853 -1467 27083 -1371
rect 25655 -1539 25671 -1505
rect 26047 -1539 26063 -1505
rect 26273 -1539 26289 -1505
rect 26665 -1539 26681 -1505
rect 25587 -1567 25621 -1551
rect 25587 -2351 25621 -2335
rect 26097 -1567 26131 -1551
rect 26097 -2351 26131 -2335
rect 26205 -1567 26239 -1551
rect 26205 -2351 26239 -2335
rect 26715 -1567 26749 -1551
rect 26715 -2351 26749 -2335
rect 25655 -2397 25671 -2363
rect 26047 -2397 26063 -2363
rect 26273 -2397 26289 -2363
rect 26665 -2397 26681 -2363
rect 25253 -2497 25483 -2435
rect 26887 -2435 27049 -1467
rect 28453 -1467 28683 -1371
rect 27255 -1539 27271 -1505
rect 27647 -1539 27663 -1505
rect 27873 -1539 27889 -1505
rect 28265 -1539 28281 -1505
rect 27187 -1567 27221 -1551
rect 27187 -2351 27221 -2335
rect 27697 -1567 27731 -1551
rect 27697 -2351 27731 -2335
rect 27805 -1567 27839 -1551
rect 27805 -2351 27839 -2335
rect 28315 -1567 28349 -1551
rect 28315 -2351 28349 -2335
rect 27255 -2397 27271 -2363
rect 27647 -2397 27663 -2363
rect 27873 -2397 27889 -2363
rect 28265 -2397 28281 -2363
rect 26853 -2497 27083 -2435
rect 28487 -2435 28649 -1467
rect 30053 -1467 30283 -1371
rect 28855 -1539 28871 -1505
rect 29247 -1539 29263 -1505
rect 29473 -1539 29489 -1505
rect 29865 -1539 29881 -1505
rect 28787 -1567 28821 -1551
rect 28787 -2351 28821 -2335
rect 29297 -1567 29331 -1551
rect 29297 -2351 29331 -2335
rect 29405 -1567 29439 -1551
rect 29405 -2351 29439 -2335
rect 29915 -1567 29949 -1551
rect 29915 -2351 29949 -2335
rect 28855 -2397 28871 -2363
rect 29247 -2397 29263 -2363
rect 29473 -2397 29489 -2363
rect 29865 -2397 29881 -2363
rect 28453 -2497 28683 -2435
rect 30087 -2435 30249 -1467
rect 31653 -1467 31883 -1371
rect 30455 -1539 30471 -1505
rect 30847 -1539 30863 -1505
rect 31073 -1539 31089 -1505
rect 31465 -1539 31481 -1505
rect 30387 -1567 30421 -1551
rect 30387 -2351 30421 -2335
rect 30897 -1567 30931 -1551
rect 30897 -2351 30931 -2335
rect 31005 -1567 31039 -1551
rect 31005 -2351 31039 -2335
rect 31515 -1567 31549 -1551
rect 31515 -2351 31549 -2335
rect 30455 -2397 30471 -2363
rect 30847 -2397 30863 -2363
rect 31073 -2397 31089 -2363
rect 31465 -2397 31481 -2363
rect 30053 -2497 30283 -2435
rect 31687 -2435 31849 -1467
rect 33253 -1467 33483 -1371
rect 32055 -1539 32071 -1505
rect 32447 -1539 32463 -1505
rect 32673 -1539 32689 -1505
rect 33065 -1539 33081 -1505
rect 31987 -1567 32021 -1551
rect 31987 -2351 32021 -2335
rect 32497 -1567 32531 -1551
rect 32497 -2351 32531 -2335
rect 32605 -1567 32639 -1551
rect 32605 -2351 32639 -2335
rect 33115 -1567 33149 -1551
rect 33115 -2351 33149 -2335
rect 32055 -2397 32071 -2363
rect 32447 -2397 32463 -2363
rect 32673 -2397 32689 -2363
rect 33065 -2397 33081 -2363
rect 31653 -2497 31883 -2435
rect 33287 -2435 33449 -1467
rect 34853 -1467 35083 -1371
rect 36453 -1405 36683 -1371
rect 38053 -1405 38400 -1371
rect 33655 -1539 33671 -1505
rect 34047 -1539 34063 -1505
rect 34273 -1539 34289 -1505
rect 34665 -1539 34681 -1505
rect 33587 -1567 33621 -1551
rect 33587 -2351 33621 -2335
rect 34097 -1567 34131 -1551
rect 34097 -2351 34131 -2335
rect 34205 -1567 34239 -1551
rect 34205 -2351 34239 -2335
rect 34715 -1567 34749 -1551
rect 34715 -2351 34749 -2335
rect 33655 -2397 33671 -2363
rect 34047 -2397 34063 -2363
rect 34273 -2397 34289 -2363
rect 34665 -2397 34681 -2363
rect 33253 -2497 33483 -2435
rect 34887 -2435 35049 -1467
rect 36453 -1467 36800 -1405
rect 35255 -1539 35271 -1505
rect 35647 -1539 35663 -1505
rect 35873 -1539 35889 -1505
rect 36265 -1539 36281 -1505
rect 35187 -1567 35221 -1551
rect 35187 -2351 35221 -2335
rect 35697 -1567 35731 -1551
rect 35697 -2351 35731 -2335
rect 35805 -1567 35839 -1551
rect 35805 -2351 35839 -2335
rect 36315 -1567 36349 -1551
rect 36315 -2351 36349 -2335
rect 35255 -2397 35271 -2363
rect 35647 -2397 35663 -2363
rect 35873 -2397 35889 -2363
rect 36265 -2397 36281 -2363
rect 34853 -2497 35083 -2435
rect 36487 -2435 36649 -1467
rect 36683 -1551 36800 -1467
rect 36980 -1505 37140 -1405
rect 36855 -1539 36871 -1505
rect 37247 -1539 37263 -1505
rect 37320 -1551 37420 -1405
rect 37600 -1505 37760 -1405
rect 37940 -1467 38400 -1405
rect 37473 -1539 37489 -1505
rect 37865 -1539 37881 -1505
rect 37940 -1551 38053 -1467
rect 36683 -1567 36821 -1551
rect 36683 -2335 36787 -1567
rect 36683 -2351 36821 -2335
rect 37297 -1567 37439 -1551
rect 37331 -2335 37405 -1567
rect 37297 -2351 37439 -2335
rect 37915 -1567 38053 -1551
rect 37949 -2335 38053 -1567
rect 37915 -2351 38053 -2335
rect 36683 -2435 36800 -2351
rect 36855 -2397 36871 -2363
rect 37247 -2397 37263 -2363
rect 36453 -2480 36800 -2435
rect 36980 -2480 37140 -2397
rect 37320 -2480 37420 -2351
rect 37473 -2397 37489 -2363
rect 37865 -2397 37881 -2363
rect 37600 -2480 37760 -2397
rect 37940 -2435 38053 -2351
rect 38087 -2435 38400 -1467
rect 37940 -2480 38400 -2435
rect 36453 -2497 38400 -2480
rect -300 -2531 -55 -2497
rect 1191 -2531 1545 -2497
rect 2791 -2531 3145 -2497
rect 4391 -2531 4745 -2497
rect 5991 -2531 6345 -2497
rect 7591 -2531 7945 -2497
rect 9191 -2531 9545 -2497
rect 10791 -2531 11145 -2497
rect 12391 -2531 12745 -2497
rect 13991 -2531 14345 -2497
rect 15591 -2531 15945 -2497
rect 17191 -2531 17545 -2497
rect 18791 -2531 19145 -2497
rect 20391 -2531 20745 -2497
rect 21991 -2531 22345 -2497
rect 23591 -2531 23945 -2497
rect 25191 -2531 25545 -2497
rect 26791 -2531 27145 -2497
rect 28391 -2531 28745 -2497
rect 29991 -2531 30345 -2497
rect 31591 -2531 31945 -2497
rect 33191 -2531 33545 -2497
rect 34791 -2531 35145 -2497
rect 36391 -2531 36745 -2497
rect 37991 -2531 38400 -2497
rect -300 -2551 38400 -2531
rect -300 -2580 1483 -2551
rect -300 -2613 0 -2580
rect -300 -2981 -151 -2613
rect -117 -2697 0 -2613
rect 180 -2651 340 -2580
rect 55 -2685 71 -2651
rect 447 -2685 463 -2651
rect 520 -2697 620 -2580
rect 800 -2651 960 -2580
rect 1140 -2613 1483 -2580
rect 673 -2685 689 -2651
rect 1065 -2685 1081 -2651
rect 1140 -2697 1253 -2613
rect -117 -2713 21 -2697
rect -117 -2881 -13 -2713
rect -117 -2897 21 -2881
rect 497 -2713 639 -2697
rect 531 -2881 605 -2713
rect 497 -2897 639 -2881
rect 1115 -2713 1253 -2697
rect 1149 -2881 1253 -2713
rect 1115 -2897 1253 -2881
rect -117 -2981 0 -2897
rect 55 -2943 71 -2909
rect 447 -2943 463 -2909
rect -300 -3043 0 -2981
rect 180 -3043 340 -2943
rect 520 -3043 620 -2897
rect 673 -2943 689 -2909
rect 1065 -2943 1081 -2909
rect 800 -3043 960 -2943
rect 1140 -2981 1253 -2897
rect 1287 -2981 1449 -2613
rect 2853 -2613 3083 -2551
rect 1655 -2685 1671 -2651
rect 2047 -2685 2063 -2651
rect 2273 -2685 2289 -2651
rect 2665 -2685 2681 -2651
rect 1587 -2713 1621 -2697
rect 1587 -2897 1621 -2881
rect 2097 -2713 2131 -2697
rect 2097 -2897 2131 -2881
rect 2205 -2713 2239 -2697
rect 2205 -2897 2239 -2881
rect 2715 -2713 2749 -2697
rect 2715 -2897 2749 -2881
rect 1655 -2943 1671 -2909
rect 2047 -2943 2063 -2909
rect 2273 -2943 2289 -2909
rect 2665 -2943 2681 -2909
rect 1140 -3043 1483 -2981
rect 2887 -2981 3049 -2613
rect 4453 -2613 4683 -2551
rect 3255 -2685 3271 -2651
rect 3647 -2685 3663 -2651
rect 3873 -2685 3889 -2651
rect 4265 -2685 4281 -2651
rect 3187 -2713 3221 -2697
rect 3187 -2897 3221 -2881
rect 3697 -2713 3731 -2697
rect 3697 -2897 3731 -2881
rect 3805 -2713 3839 -2697
rect 3805 -2897 3839 -2881
rect 4315 -2713 4349 -2697
rect 4315 -2897 4349 -2881
rect 3255 -2943 3271 -2909
rect 3647 -2943 3663 -2909
rect 3873 -2943 3889 -2909
rect 4265 -2943 4281 -2909
rect 2853 -3043 3083 -2981
rect 4487 -2981 4649 -2613
rect 6053 -2613 6283 -2551
rect 4855 -2685 4871 -2651
rect 5247 -2685 5263 -2651
rect 5473 -2685 5489 -2651
rect 5865 -2685 5881 -2651
rect 4787 -2713 4821 -2697
rect 4787 -2897 4821 -2881
rect 5297 -2713 5331 -2697
rect 5297 -2897 5331 -2881
rect 5405 -2713 5439 -2697
rect 5405 -2897 5439 -2881
rect 5915 -2713 5949 -2697
rect 5915 -2897 5949 -2881
rect 4855 -2943 4871 -2909
rect 5247 -2943 5263 -2909
rect 5473 -2943 5489 -2909
rect 5865 -2943 5881 -2909
rect 4453 -3043 4683 -2981
rect 6087 -2981 6249 -2613
rect 7653 -2613 7883 -2551
rect 6455 -2685 6471 -2651
rect 6847 -2685 6863 -2651
rect 7073 -2685 7089 -2651
rect 7465 -2685 7481 -2651
rect 6387 -2713 6421 -2697
rect 6387 -2897 6421 -2881
rect 6897 -2713 6931 -2697
rect 6897 -2897 6931 -2881
rect 7005 -2713 7039 -2697
rect 7005 -2897 7039 -2881
rect 7515 -2713 7549 -2697
rect 7515 -2897 7549 -2881
rect 6455 -2943 6471 -2909
rect 6847 -2943 6863 -2909
rect 7073 -2943 7089 -2909
rect 7465 -2943 7481 -2909
rect 6053 -3043 6283 -2981
rect 7687 -2981 7849 -2613
rect 9253 -2613 9483 -2551
rect 8055 -2685 8071 -2651
rect 8447 -2685 8463 -2651
rect 8673 -2685 8689 -2651
rect 9065 -2685 9081 -2651
rect 7987 -2713 8021 -2697
rect 7987 -2897 8021 -2881
rect 8497 -2713 8531 -2697
rect 8497 -2897 8531 -2881
rect 8605 -2713 8639 -2697
rect 8605 -2897 8639 -2881
rect 9115 -2713 9149 -2697
rect 9115 -2897 9149 -2881
rect 8055 -2943 8071 -2909
rect 8447 -2943 8463 -2909
rect 8673 -2943 8689 -2909
rect 9065 -2943 9081 -2909
rect 7653 -3043 7883 -2981
rect 9287 -2981 9449 -2613
rect 10853 -2613 11083 -2551
rect 9655 -2685 9671 -2651
rect 10047 -2685 10063 -2651
rect 10273 -2685 10289 -2651
rect 10665 -2685 10681 -2651
rect 9587 -2713 9621 -2697
rect 9587 -2897 9621 -2881
rect 10097 -2713 10131 -2697
rect 10097 -2897 10131 -2881
rect 10205 -2713 10239 -2697
rect 10205 -2897 10239 -2881
rect 10715 -2713 10749 -2697
rect 10715 -2897 10749 -2881
rect 9655 -2943 9671 -2909
rect 10047 -2943 10063 -2909
rect 10273 -2943 10289 -2909
rect 10665 -2943 10681 -2909
rect 9253 -3043 9483 -2981
rect 10887 -2981 11049 -2613
rect 12453 -2613 12683 -2551
rect 11255 -2685 11271 -2651
rect 11647 -2685 11663 -2651
rect 11873 -2685 11889 -2651
rect 12265 -2685 12281 -2651
rect 11187 -2713 11221 -2697
rect 11187 -2897 11221 -2881
rect 11697 -2713 11731 -2697
rect 11697 -2897 11731 -2881
rect 11805 -2713 11839 -2697
rect 11805 -2897 11839 -2881
rect 12315 -2713 12349 -2697
rect 12315 -2897 12349 -2881
rect 11255 -2943 11271 -2909
rect 11647 -2943 11663 -2909
rect 11873 -2943 11889 -2909
rect 12265 -2943 12281 -2909
rect 10853 -3043 11083 -2981
rect 12487 -2981 12649 -2613
rect 14053 -2613 14283 -2551
rect 12855 -2685 12871 -2651
rect 13247 -2685 13263 -2651
rect 13473 -2685 13489 -2651
rect 13865 -2685 13881 -2651
rect 12787 -2713 12821 -2697
rect 12787 -2897 12821 -2881
rect 13297 -2713 13331 -2697
rect 13297 -2897 13331 -2881
rect 13405 -2713 13439 -2697
rect 13405 -2897 13439 -2881
rect 13915 -2713 13949 -2697
rect 13915 -2897 13949 -2881
rect 12855 -2943 12871 -2909
rect 13247 -2943 13263 -2909
rect 13473 -2943 13489 -2909
rect 13865 -2943 13881 -2909
rect 12453 -3043 12683 -2981
rect 14087 -2981 14249 -2613
rect 15653 -2613 15883 -2551
rect 14455 -2685 14471 -2651
rect 14847 -2685 14863 -2651
rect 15073 -2685 15089 -2651
rect 15465 -2685 15481 -2651
rect 14387 -2713 14421 -2697
rect 14387 -2897 14421 -2881
rect 14897 -2713 14931 -2697
rect 14897 -2897 14931 -2881
rect 15005 -2713 15039 -2697
rect 15005 -2897 15039 -2881
rect 15515 -2713 15549 -2697
rect 15515 -2897 15549 -2881
rect 14455 -2943 14471 -2909
rect 14847 -2943 14863 -2909
rect 15073 -2943 15089 -2909
rect 15465 -2943 15481 -2909
rect 14053 -3043 14283 -2981
rect 15687 -2981 15849 -2613
rect 17253 -2613 17483 -2551
rect 16055 -2685 16071 -2651
rect 16447 -2685 16463 -2651
rect 16673 -2685 16689 -2651
rect 17065 -2685 17081 -2651
rect 15987 -2713 16021 -2697
rect 15987 -2897 16021 -2881
rect 16497 -2713 16531 -2697
rect 16497 -2897 16531 -2881
rect 16605 -2713 16639 -2697
rect 16605 -2897 16639 -2881
rect 17115 -2713 17149 -2697
rect 17115 -2897 17149 -2881
rect 16055 -2943 16071 -2909
rect 16447 -2943 16463 -2909
rect 16673 -2943 16689 -2909
rect 17065 -2943 17081 -2909
rect 15653 -3043 15883 -2981
rect 17287 -2981 17449 -2613
rect 18853 -2613 19083 -2551
rect 17655 -2685 17671 -2651
rect 18047 -2685 18063 -2651
rect 18273 -2685 18289 -2651
rect 18665 -2685 18681 -2651
rect 17587 -2713 17621 -2697
rect 17587 -2897 17621 -2881
rect 18097 -2713 18131 -2697
rect 18097 -2897 18131 -2881
rect 18205 -2713 18239 -2697
rect 18205 -2897 18239 -2881
rect 18715 -2713 18749 -2697
rect 18715 -2897 18749 -2881
rect 17655 -2943 17671 -2909
rect 18047 -2943 18063 -2909
rect 18273 -2943 18289 -2909
rect 18665 -2943 18681 -2909
rect 17253 -3043 17483 -2981
rect 18887 -2981 19049 -2613
rect 20453 -2613 20683 -2551
rect 19255 -2685 19271 -2651
rect 19647 -2685 19663 -2651
rect 19873 -2685 19889 -2651
rect 20265 -2685 20281 -2651
rect 19187 -2713 19221 -2697
rect 19187 -2897 19221 -2881
rect 19697 -2713 19731 -2697
rect 19697 -2897 19731 -2881
rect 19805 -2713 19839 -2697
rect 19805 -2897 19839 -2881
rect 20315 -2713 20349 -2697
rect 20315 -2897 20349 -2881
rect 19255 -2943 19271 -2909
rect 19647 -2943 19663 -2909
rect 19873 -2943 19889 -2909
rect 20265 -2943 20281 -2909
rect 18853 -3043 19083 -2981
rect 20487 -2981 20649 -2613
rect 22053 -2613 22283 -2551
rect 20855 -2685 20871 -2651
rect 21247 -2685 21263 -2651
rect 21473 -2685 21489 -2651
rect 21865 -2685 21881 -2651
rect 20787 -2713 20821 -2697
rect 20787 -2897 20821 -2881
rect 21297 -2713 21331 -2697
rect 21297 -2897 21331 -2881
rect 21405 -2713 21439 -2697
rect 21405 -2897 21439 -2881
rect 21915 -2713 21949 -2697
rect 21915 -2897 21949 -2881
rect 20855 -2943 20871 -2909
rect 21247 -2943 21263 -2909
rect 21473 -2943 21489 -2909
rect 21865 -2943 21881 -2909
rect 20453 -3043 20683 -2981
rect 22087 -2981 22249 -2613
rect 23653 -2613 23883 -2551
rect 22455 -2685 22471 -2651
rect 22847 -2685 22863 -2651
rect 23073 -2685 23089 -2651
rect 23465 -2685 23481 -2651
rect 22387 -2713 22421 -2697
rect 22387 -2897 22421 -2881
rect 22897 -2713 22931 -2697
rect 22897 -2897 22931 -2881
rect 23005 -2713 23039 -2697
rect 23005 -2897 23039 -2881
rect 23515 -2713 23549 -2697
rect 23515 -2897 23549 -2881
rect 22455 -2943 22471 -2909
rect 22847 -2943 22863 -2909
rect 23073 -2943 23089 -2909
rect 23465 -2943 23481 -2909
rect 22053 -3043 22283 -2981
rect 23687 -2981 23849 -2613
rect 25253 -2613 25483 -2551
rect 24055 -2685 24071 -2651
rect 24447 -2685 24463 -2651
rect 24673 -2685 24689 -2651
rect 25065 -2685 25081 -2651
rect 23987 -2713 24021 -2697
rect 23987 -2897 24021 -2881
rect 24497 -2713 24531 -2697
rect 24497 -2897 24531 -2881
rect 24605 -2713 24639 -2697
rect 24605 -2897 24639 -2881
rect 25115 -2713 25149 -2697
rect 25115 -2897 25149 -2881
rect 24055 -2943 24071 -2909
rect 24447 -2943 24463 -2909
rect 24673 -2943 24689 -2909
rect 25065 -2943 25081 -2909
rect 23653 -3043 23883 -2981
rect 25287 -2981 25449 -2613
rect 26853 -2613 27083 -2551
rect 25655 -2685 25671 -2651
rect 26047 -2685 26063 -2651
rect 26273 -2685 26289 -2651
rect 26665 -2685 26681 -2651
rect 25587 -2713 25621 -2697
rect 25587 -2897 25621 -2881
rect 26097 -2713 26131 -2697
rect 26097 -2897 26131 -2881
rect 26205 -2713 26239 -2697
rect 26205 -2897 26239 -2881
rect 26715 -2713 26749 -2697
rect 26715 -2897 26749 -2881
rect 25655 -2943 25671 -2909
rect 26047 -2943 26063 -2909
rect 26273 -2943 26289 -2909
rect 26665 -2943 26681 -2909
rect 25253 -3043 25483 -2981
rect 26887 -2981 27049 -2613
rect 28453 -2613 28683 -2551
rect 27255 -2685 27271 -2651
rect 27647 -2685 27663 -2651
rect 27873 -2685 27889 -2651
rect 28265 -2685 28281 -2651
rect 27187 -2713 27221 -2697
rect 27187 -2897 27221 -2881
rect 27697 -2713 27731 -2697
rect 27697 -2897 27731 -2881
rect 27805 -2713 27839 -2697
rect 27805 -2897 27839 -2881
rect 28315 -2713 28349 -2697
rect 28315 -2897 28349 -2881
rect 27255 -2943 27271 -2909
rect 27647 -2943 27663 -2909
rect 27873 -2943 27889 -2909
rect 28265 -2943 28281 -2909
rect 26853 -3043 27083 -2981
rect 28487 -2981 28649 -2613
rect 30053 -2613 30283 -2551
rect 28855 -2685 28871 -2651
rect 29247 -2685 29263 -2651
rect 29473 -2685 29489 -2651
rect 29865 -2685 29881 -2651
rect 28787 -2713 28821 -2697
rect 28787 -2897 28821 -2881
rect 29297 -2713 29331 -2697
rect 29297 -2897 29331 -2881
rect 29405 -2713 29439 -2697
rect 29405 -2897 29439 -2881
rect 29915 -2713 29949 -2697
rect 29915 -2897 29949 -2881
rect 28855 -2943 28871 -2909
rect 29247 -2943 29263 -2909
rect 29473 -2943 29489 -2909
rect 29865 -2943 29881 -2909
rect 28453 -3043 28683 -2981
rect 30087 -2981 30249 -2613
rect 31653 -2613 31883 -2551
rect 30455 -2685 30471 -2651
rect 30847 -2685 30863 -2651
rect 31073 -2685 31089 -2651
rect 31465 -2685 31481 -2651
rect 30387 -2713 30421 -2697
rect 30387 -2897 30421 -2881
rect 30897 -2713 30931 -2697
rect 30897 -2897 30931 -2881
rect 31005 -2713 31039 -2697
rect 31005 -2897 31039 -2881
rect 31515 -2713 31549 -2697
rect 31515 -2897 31549 -2881
rect 30455 -2943 30471 -2909
rect 30847 -2943 30863 -2909
rect 31073 -2943 31089 -2909
rect 31465 -2943 31481 -2909
rect 30053 -3043 30283 -2981
rect 31687 -2981 31849 -2613
rect 33253 -2613 33483 -2551
rect 32055 -2685 32071 -2651
rect 32447 -2685 32463 -2651
rect 32673 -2685 32689 -2651
rect 33065 -2685 33081 -2651
rect 31987 -2713 32021 -2697
rect 31987 -2897 32021 -2881
rect 32497 -2713 32531 -2697
rect 32497 -2897 32531 -2881
rect 32605 -2713 32639 -2697
rect 32605 -2897 32639 -2881
rect 33115 -2713 33149 -2697
rect 33115 -2897 33149 -2881
rect 32055 -2943 32071 -2909
rect 32447 -2943 32463 -2909
rect 32673 -2943 32689 -2909
rect 33065 -2943 33081 -2909
rect 31653 -3043 31883 -2981
rect 33287 -2981 33449 -2613
rect 34853 -2613 35083 -2551
rect 33655 -2685 33671 -2651
rect 34047 -2685 34063 -2651
rect 34273 -2685 34289 -2651
rect 34665 -2685 34681 -2651
rect 33587 -2713 33621 -2697
rect 33587 -2897 33621 -2881
rect 34097 -2713 34131 -2697
rect 34097 -2897 34131 -2881
rect 34205 -2713 34239 -2697
rect 34205 -2897 34239 -2881
rect 34715 -2713 34749 -2697
rect 34715 -2897 34749 -2881
rect 33655 -2943 33671 -2909
rect 34047 -2943 34063 -2909
rect 34273 -2943 34289 -2909
rect 34665 -2943 34681 -2909
rect 33253 -3043 33483 -2981
rect 34887 -2981 35049 -2613
rect 36453 -2580 38400 -2551
rect 36453 -2613 36800 -2580
rect 35255 -2685 35271 -2651
rect 35647 -2685 35663 -2651
rect 35873 -2685 35889 -2651
rect 36265 -2685 36281 -2651
rect 35187 -2713 35221 -2697
rect 35187 -2897 35221 -2881
rect 35697 -2713 35731 -2697
rect 35697 -2897 35731 -2881
rect 35805 -2713 35839 -2697
rect 35805 -2897 35839 -2881
rect 36315 -2713 36349 -2697
rect 36315 -2897 36349 -2881
rect 35255 -2943 35271 -2909
rect 35647 -2943 35663 -2909
rect 35873 -2943 35889 -2909
rect 36265 -2943 36281 -2909
rect 34853 -3043 35083 -2981
rect 36487 -2981 36649 -2613
rect 36683 -2697 36800 -2613
rect 36980 -2651 37140 -2580
rect 36855 -2685 36871 -2651
rect 37247 -2685 37263 -2651
rect 37320 -2697 37420 -2580
rect 37600 -2651 37760 -2580
rect 37940 -2613 38400 -2580
rect 37473 -2685 37489 -2651
rect 37865 -2685 37881 -2651
rect 37940 -2697 38053 -2613
rect 36683 -2713 36821 -2697
rect 36683 -2881 36787 -2713
rect 36683 -2897 36821 -2881
rect 37297 -2713 37439 -2697
rect 37331 -2881 37405 -2713
rect 37297 -2897 37439 -2881
rect 37915 -2713 38053 -2697
rect 37949 -2881 38053 -2713
rect 37915 -2897 38053 -2881
rect 36683 -2981 36800 -2897
rect 36855 -2943 36871 -2909
rect 37247 -2943 37263 -2909
rect 36453 -3043 36800 -2981
rect 36980 -3043 37140 -2943
rect 37320 -3043 37420 -2897
rect 37473 -2943 37489 -2909
rect 37865 -2943 37881 -2909
rect 37600 -3043 37760 -2943
rect 37940 -2981 38053 -2897
rect 38087 -2981 38400 -2613
rect 37940 -3043 38400 -2981
rect -300 -3171 38400 -3043
rect -300 -3205 -117 -3171
rect 1253 -3205 1483 -3171
rect -300 -3267 0 -3205
rect -300 -4235 -151 -3267
rect -117 -3351 0 -3267
rect 180 -3305 340 -3205
rect 55 -3339 71 -3305
rect 447 -3339 463 -3305
rect 520 -3351 620 -3205
rect 800 -3305 960 -3205
rect 1140 -3267 1483 -3205
rect 673 -3339 689 -3305
rect 1065 -3339 1081 -3305
rect 1140 -3351 1253 -3267
rect -117 -3367 21 -3351
rect -117 -4135 -13 -3367
rect -117 -4151 21 -4135
rect 497 -3367 639 -3351
rect 531 -4135 605 -3367
rect 497 -4151 639 -4135
rect 1115 -3367 1253 -3351
rect 1149 -4135 1253 -3367
rect 1115 -4151 1253 -4135
rect -117 -4235 0 -4151
rect 55 -4197 71 -4163
rect 447 -4197 463 -4163
rect -300 -4280 0 -4235
rect 180 -4280 340 -4197
rect 520 -4280 620 -4151
rect 673 -4197 689 -4163
rect 1065 -4197 1081 -4163
rect 800 -4280 960 -4197
rect 1140 -4235 1253 -4151
rect 1287 -4235 1449 -3267
rect 2853 -3267 3083 -3171
rect 1655 -3339 1671 -3305
rect 2047 -3339 2063 -3305
rect 2273 -3339 2289 -3305
rect 2665 -3339 2681 -3305
rect 1587 -3367 1621 -3351
rect 1587 -4151 1621 -4135
rect 2097 -3367 2131 -3351
rect 2097 -4151 2131 -4135
rect 2205 -3367 2239 -3351
rect 2205 -4151 2239 -4135
rect 2715 -3367 2749 -3351
rect 2715 -4151 2749 -4135
rect 1655 -4197 1671 -4163
rect 2047 -4197 2063 -4163
rect 2273 -4197 2289 -4163
rect 2665 -4197 2681 -4163
rect 1140 -4280 1483 -4235
rect -300 -4297 1483 -4280
rect 2887 -4235 3049 -3267
rect 4453 -3267 4683 -3171
rect 3255 -3339 3271 -3305
rect 3647 -3339 3663 -3305
rect 3873 -3339 3889 -3305
rect 4265 -3339 4281 -3305
rect 3187 -3367 3221 -3351
rect 3187 -4151 3221 -4135
rect 3697 -3367 3731 -3351
rect 3697 -4151 3731 -4135
rect 3805 -3367 3839 -3351
rect 3805 -4151 3839 -4135
rect 4315 -3367 4349 -3351
rect 4315 -4151 4349 -4135
rect 3255 -4197 3271 -4163
rect 3647 -4197 3663 -4163
rect 3873 -4197 3889 -4163
rect 4265 -4197 4281 -4163
rect 2853 -4297 3083 -4235
rect 4487 -4235 4649 -3267
rect 6053 -3267 6283 -3171
rect 4855 -3339 4871 -3305
rect 5247 -3339 5263 -3305
rect 5473 -3339 5489 -3305
rect 5865 -3339 5881 -3305
rect 4787 -3367 4821 -3351
rect 4787 -4151 4821 -4135
rect 5297 -3367 5331 -3351
rect 5297 -4151 5331 -4135
rect 5405 -3367 5439 -3351
rect 5405 -4151 5439 -4135
rect 5915 -3367 5949 -3351
rect 5915 -4151 5949 -4135
rect 4855 -4197 4871 -4163
rect 5247 -4197 5263 -4163
rect 5473 -4197 5489 -4163
rect 5865 -4197 5881 -4163
rect 4453 -4297 4683 -4235
rect 6087 -4235 6249 -3267
rect 7653 -3267 7883 -3171
rect 6455 -3339 6471 -3305
rect 6847 -3339 6863 -3305
rect 7073 -3339 7089 -3305
rect 7465 -3339 7481 -3305
rect 6387 -3367 6421 -3351
rect 6387 -4151 6421 -4135
rect 6897 -3367 6931 -3351
rect 6897 -4151 6931 -4135
rect 7005 -3367 7039 -3351
rect 7005 -4151 7039 -4135
rect 7515 -3367 7549 -3351
rect 7515 -4151 7549 -4135
rect 6455 -4197 6471 -4163
rect 6847 -4197 6863 -4163
rect 7073 -4197 7089 -4163
rect 7465 -4197 7481 -4163
rect 6053 -4297 6283 -4235
rect 7687 -4235 7849 -3267
rect 9253 -3267 9483 -3171
rect 8055 -3339 8071 -3305
rect 8447 -3339 8463 -3305
rect 8673 -3339 8689 -3305
rect 9065 -3339 9081 -3305
rect 7987 -3367 8021 -3351
rect 7987 -4151 8021 -4135
rect 8497 -3367 8531 -3351
rect 8497 -4151 8531 -4135
rect 8605 -3367 8639 -3351
rect 8605 -4151 8639 -4135
rect 9115 -3367 9149 -3351
rect 9115 -4151 9149 -4135
rect 8055 -4197 8071 -4163
rect 8447 -4197 8463 -4163
rect 8673 -4197 8689 -4163
rect 9065 -4197 9081 -4163
rect 7653 -4297 7883 -4235
rect 9287 -4235 9449 -3267
rect 10853 -3267 11083 -3171
rect 9655 -3339 9671 -3305
rect 10047 -3339 10063 -3305
rect 10273 -3339 10289 -3305
rect 10665 -3339 10681 -3305
rect 9587 -3367 9621 -3351
rect 9587 -4151 9621 -4135
rect 10097 -3367 10131 -3351
rect 10097 -4151 10131 -4135
rect 10205 -3367 10239 -3351
rect 10205 -4151 10239 -4135
rect 10715 -3367 10749 -3351
rect 10715 -4151 10749 -4135
rect 9655 -4197 9671 -4163
rect 10047 -4197 10063 -4163
rect 10273 -4197 10289 -4163
rect 10665 -4197 10681 -4163
rect 9253 -4297 9483 -4235
rect 10887 -4235 11049 -3267
rect 12453 -3267 12683 -3171
rect 11255 -3339 11271 -3305
rect 11647 -3339 11663 -3305
rect 11873 -3339 11889 -3305
rect 12265 -3339 12281 -3305
rect 11187 -3367 11221 -3351
rect 11187 -4151 11221 -4135
rect 11697 -3367 11731 -3351
rect 11697 -4151 11731 -4135
rect 11805 -3367 11839 -3351
rect 11805 -4151 11839 -4135
rect 12315 -3367 12349 -3351
rect 12315 -4151 12349 -4135
rect 11255 -4197 11271 -4163
rect 11647 -4197 11663 -4163
rect 11873 -4197 11889 -4163
rect 12265 -4197 12281 -4163
rect 10853 -4297 11083 -4235
rect 12487 -4235 12649 -3267
rect 14053 -3267 14283 -3171
rect 12855 -3339 12871 -3305
rect 13247 -3339 13263 -3305
rect 13473 -3339 13489 -3305
rect 13865 -3339 13881 -3305
rect 12787 -3367 12821 -3351
rect 12787 -4151 12821 -4135
rect 13297 -3367 13331 -3351
rect 13297 -4151 13331 -4135
rect 13405 -3367 13439 -3351
rect 13405 -4151 13439 -4135
rect 13915 -3367 13949 -3351
rect 13915 -4151 13949 -4135
rect 12855 -4197 12871 -4163
rect 13247 -4197 13263 -4163
rect 13473 -4197 13489 -4163
rect 13865 -4197 13881 -4163
rect 12453 -4297 12683 -4235
rect 14087 -4235 14249 -3267
rect 15653 -3267 15883 -3171
rect 14455 -3339 14471 -3305
rect 14847 -3339 14863 -3305
rect 15073 -3339 15089 -3305
rect 15465 -3339 15481 -3305
rect 14387 -3367 14421 -3351
rect 14387 -4151 14421 -4135
rect 14897 -3367 14931 -3351
rect 14897 -4151 14931 -4135
rect 15005 -3367 15039 -3351
rect 15005 -4151 15039 -4135
rect 15515 -3367 15549 -3351
rect 15515 -4151 15549 -4135
rect 14455 -4197 14471 -4163
rect 14847 -4197 14863 -4163
rect 15073 -4197 15089 -4163
rect 15465 -4197 15481 -4163
rect 14053 -4297 14283 -4235
rect 15687 -4235 15849 -3267
rect 17253 -3267 17483 -3171
rect 16055 -3339 16071 -3305
rect 16447 -3339 16463 -3305
rect 16673 -3339 16689 -3305
rect 17065 -3339 17081 -3305
rect 15987 -3367 16021 -3351
rect 15987 -4151 16021 -4135
rect 16497 -3367 16531 -3351
rect 16497 -4151 16531 -4135
rect 16605 -3367 16639 -3351
rect 16605 -4151 16639 -4135
rect 17115 -3367 17149 -3351
rect 17115 -4151 17149 -4135
rect 16055 -4197 16071 -4163
rect 16447 -4197 16463 -4163
rect 16673 -4197 16689 -4163
rect 17065 -4197 17081 -4163
rect 15653 -4297 15883 -4235
rect 17287 -4235 17449 -3267
rect 18853 -3267 19083 -3171
rect 17655 -3339 17671 -3305
rect 18047 -3339 18063 -3305
rect 18273 -3339 18289 -3305
rect 18665 -3339 18681 -3305
rect 17587 -3367 17621 -3351
rect 17587 -4151 17621 -4135
rect 18097 -3367 18131 -3351
rect 18097 -4151 18131 -4135
rect 18205 -3367 18239 -3351
rect 18205 -4151 18239 -4135
rect 18715 -3367 18749 -3351
rect 18715 -4151 18749 -4135
rect 17655 -4197 17671 -4163
rect 18047 -4197 18063 -4163
rect 18273 -4197 18289 -4163
rect 18665 -4197 18681 -4163
rect 17253 -4297 17483 -4235
rect 18887 -4235 19049 -3267
rect 20453 -3267 20683 -3171
rect 19255 -3339 19271 -3305
rect 19647 -3339 19663 -3305
rect 19873 -3339 19889 -3305
rect 20265 -3339 20281 -3305
rect 19187 -3367 19221 -3351
rect 19187 -4151 19221 -4135
rect 19697 -3367 19731 -3351
rect 19697 -4151 19731 -4135
rect 19805 -3367 19839 -3351
rect 19805 -4151 19839 -4135
rect 20315 -3367 20349 -3351
rect 20315 -4151 20349 -4135
rect 19255 -4197 19271 -4163
rect 19647 -4197 19663 -4163
rect 19873 -4197 19889 -4163
rect 20265 -4197 20281 -4163
rect 18853 -4297 19083 -4235
rect 20487 -4235 20649 -3267
rect 22053 -3267 22283 -3171
rect 20855 -3339 20871 -3305
rect 21247 -3339 21263 -3305
rect 21473 -3339 21489 -3305
rect 21865 -3339 21881 -3305
rect 20787 -3367 20821 -3351
rect 20787 -4151 20821 -4135
rect 21297 -3367 21331 -3351
rect 21297 -4151 21331 -4135
rect 21405 -3367 21439 -3351
rect 21405 -4151 21439 -4135
rect 21915 -3367 21949 -3351
rect 21915 -4151 21949 -4135
rect 20855 -4197 20871 -4163
rect 21247 -4197 21263 -4163
rect 21473 -4197 21489 -4163
rect 21865 -4197 21881 -4163
rect 20453 -4297 20683 -4235
rect 22087 -4235 22249 -3267
rect 23653 -3267 23883 -3171
rect 22455 -3339 22471 -3305
rect 22847 -3339 22863 -3305
rect 23073 -3339 23089 -3305
rect 23465 -3339 23481 -3305
rect 22387 -3367 22421 -3351
rect 22387 -4151 22421 -4135
rect 22897 -3367 22931 -3351
rect 22897 -4151 22931 -4135
rect 23005 -3367 23039 -3351
rect 23005 -4151 23039 -4135
rect 23515 -3367 23549 -3351
rect 23515 -4151 23549 -4135
rect 22455 -4197 22471 -4163
rect 22847 -4197 22863 -4163
rect 23073 -4197 23089 -4163
rect 23465 -4197 23481 -4163
rect 22053 -4297 22283 -4235
rect 23687 -4235 23849 -3267
rect 25253 -3267 25483 -3171
rect 24055 -3339 24071 -3305
rect 24447 -3339 24463 -3305
rect 24673 -3339 24689 -3305
rect 25065 -3339 25081 -3305
rect 23987 -3367 24021 -3351
rect 23987 -4151 24021 -4135
rect 24497 -3367 24531 -3351
rect 24497 -4151 24531 -4135
rect 24605 -3367 24639 -3351
rect 24605 -4151 24639 -4135
rect 25115 -3367 25149 -3351
rect 25115 -4151 25149 -4135
rect 24055 -4197 24071 -4163
rect 24447 -4197 24463 -4163
rect 24673 -4197 24689 -4163
rect 25065 -4197 25081 -4163
rect 23653 -4297 23883 -4235
rect 25287 -4235 25449 -3267
rect 26853 -3267 27083 -3171
rect 25655 -3339 25671 -3305
rect 26047 -3339 26063 -3305
rect 26273 -3339 26289 -3305
rect 26665 -3339 26681 -3305
rect 25587 -3367 25621 -3351
rect 25587 -4151 25621 -4135
rect 26097 -3367 26131 -3351
rect 26097 -4151 26131 -4135
rect 26205 -3367 26239 -3351
rect 26205 -4151 26239 -4135
rect 26715 -3367 26749 -3351
rect 26715 -4151 26749 -4135
rect 25655 -4197 25671 -4163
rect 26047 -4197 26063 -4163
rect 26273 -4197 26289 -4163
rect 26665 -4197 26681 -4163
rect 25253 -4297 25483 -4235
rect 26887 -4235 27049 -3267
rect 28453 -3267 28683 -3171
rect 27255 -3339 27271 -3305
rect 27647 -3339 27663 -3305
rect 27873 -3339 27889 -3305
rect 28265 -3339 28281 -3305
rect 27187 -3367 27221 -3351
rect 27187 -4151 27221 -4135
rect 27697 -3367 27731 -3351
rect 27697 -4151 27731 -4135
rect 27805 -3367 27839 -3351
rect 27805 -4151 27839 -4135
rect 28315 -3367 28349 -3351
rect 28315 -4151 28349 -4135
rect 27255 -4197 27271 -4163
rect 27647 -4197 27663 -4163
rect 27873 -4197 27889 -4163
rect 28265 -4197 28281 -4163
rect 26853 -4297 27083 -4235
rect 28487 -4235 28649 -3267
rect 30053 -3267 30283 -3171
rect 28855 -3339 28871 -3305
rect 29247 -3339 29263 -3305
rect 29473 -3339 29489 -3305
rect 29865 -3339 29881 -3305
rect 28787 -3367 28821 -3351
rect 28787 -4151 28821 -4135
rect 29297 -3367 29331 -3351
rect 29297 -4151 29331 -4135
rect 29405 -3367 29439 -3351
rect 29405 -4151 29439 -4135
rect 29915 -3367 29949 -3351
rect 29915 -4151 29949 -4135
rect 28855 -4197 28871 -4163
rect 29247 -4197 29263 -4163
rect 29473 -4197 29489 -4163
rect 29865 -4197 29881 -4163
rect 28453 -4297 28683 -4235
rect 30087 -4235 30249 -3267
rect 31653 -3267 31883 -3171
rect 30455 -3339 30471 -3305
rect 30847 -3339 30863 -3305
rect 31073 -3339 31089 -3305
rect 31465 -3339 31481 -3305
rect 30387 -3367 30421 -3351
rect 30387 -4151 30421 -4135
rect 30897 -3367 30931 -3351
rect 30897 -4151 30931 -4135
rect 31005 -3367 31039 -3351
rect 31005 -4151 31039 -4135
rect 31515 -3367 31549 -3351
rect 31515 -4151 31549 -4135
rect 30455 -4197 30471 -4163
rect 30847 -4197 30863 -4163
rect 31073 -4197 31089 -4163
rect 31465 -4197 31481 -4163
rect 30053 -4297 30283 -4235
rect 31687 -4235 31849 -3267
rect 33253 -3267 33483 -3171
rect 32055 -3339 32071 -3305
rect 32447 -3339 32463 -3305
rect 32673 -3339 32689 -3305
rect 33065 -3339 33081 -3305
rect 31987 -3367 32021 -3351
rect 31987 -4151 32021 -4135
rect 32497 -3367 32531 -3351
rect 32497 -4151 32531 -4135
rect 32605 -3367 32639 -3351
rect 32605 -4151 32639 -4135
rect 33115 -3367 33149 -3351
rect 33115 -4151 33149 -4135
rect 32055 -4197 32071 -4163
rect 32447 -4197 32463 -4163
rect 32673 -4197 32689 -4163
rect 33065 -4197 33081 -4163
rect 31653 -4297 31883 -4235
rect 33287 -4235 33449 -3267
rect 34853 -3267 35083 -3171
rect 36453 -3205 36683 -3171
rect 38053 -3205 38400 -3171
rect 33655 -3339 33671 -3305
rect 34047 -3339 34063 -3305
rect 34273 -3339 34289 -3305
rect 34665 -3339 34681 -3305
rect 33587 -3367 33621 -3351
rect 33587 -4151 33621 -4135
rect 34097 -3367 34131 -3351
rect 34097 -4151 34131 -4135
rect 34205 -3367 34239 -3351
rect 34205 -4151 34239 -4135
rect 34715 -3367 34749 -3351
rect 34715 -4151 34749 -4135
rect 33655 -4197 33671 -4163
rect 34047 -4197 34063 -4163
rect 34273 -4197 34289 -4163
rect 34665 -4197 34681 -4163
rect 33253 -4297 33483 -4235
rect 34887 -4235 35049 -3267
rect 36453 -3267 36800 -3205
rect 35255 -3339 35271 -3305
rect 35647 -3339 35663 -3305
rect 35873 -3339 35889 -3305
rect 36265 -3339 36281 -3305
rect 35187 -3367 35221 -3351
rect 35187 -4151 35221 -4135
rect 35697 -3367 35731 -3351
rect 35697 -4151 35731 -4135
rect 35805 -3367 35839 -3351
rect 35805 -4151 35839 -4135
rect 36315 -3367 36349 -3351
rect 36315 -4151 36349 -4135
rect 35255 -4197 35271 -4163
rect 35647 -4197 35663 -4163
rect 35873 -4197 35889 -4163
rect 36265 -4197 36281 -4163
rect 34853 -4297 35083 -4235
rect 36487 -4235 36649 -3267
rect 36683 -3351 36800 -3267
rect 36980 -3305 37140 -3205
rect 36855 -3339 36871 -3305
rect 37247 -3339 37263 -3305
rect 37320 -3351 37420 -3205
rect 37600 -3305 37760 -3205
rect 37940 -3267 38400 -3205
rect 37473 -3339 37489 -3305
rect 37865 -3339 37881 -3305
rect 37940 -3351 38053 -3267
rect 36683 -3367 36821 -3351
rect 36683 -4135 36787 -3367
rect 36683 -4151 36821 -4135
rect 37297 -3367 37439 -3351
rect 37331 -4135 37405 -3367
rect 37297 -4151 37439 -4135
rect 37915 -3367 38053 -3351
rect 37949 -4135 38053 -3367
rect 37915 -4151 38053 -4135
rect 36683 -4235 36800 -4151
rect 36855 -4197 36871 -4163
rect 37247 -4197 37263 -4163
rect 36453 -4280 36800 -4235
rect 36980 -4280 37140 -4197
rect 37320 -4280 37420 -4151
rect 37473 -4197 37489 -4163
rect 37865 -4197 37881 -4163
rect 37600 -4280 37760 -4197
rect 37940 -4235 38053 -4151
rect 38087 -4235 38400 -3267
rect 37940 -4280 38400 -4235
rect 36453 -4297 38400 -4280
rect -300 -4331 -55 -4297
rect 1191 -4331 1545 -4297
rect 2791 -4331 3145 -4297
rect 4391 -4331 4745 -4297
rect 5991 -4331 6345 -4297
rect 7591 -4331 7945 -4297
rect 9191 -4331 9545 -4297
rect 10791 -4331 11145 -4297
rect 12391 -4331 12745 -4297
rect 13991 -4331 14345 -4297
rect 15591 -4331 15945 -4297
rect 17191 -4331 17545 -4297
rect 18791 -4331 19145 -4297
rect 20391 -4331 20745 -4297
rect 21991 -4331 22345 -4297
rect 23591 -4331 23945 -4297
rect 25191 -4331 25545 -4297
rect 26791 -4331 27145 -4297
rect 28391 -4331 28745 -4297
rect 29991 -4331 30345 -4297
rect 31591 -4331 31945 -4297
rect 33191 -4331 33545 -4297
rect 34791 -4331 35145 -4297
rect 36391 -4331 36745 -4297
rect 37991 -4331 38400 -4297
rect -300 -4351 38400 -4331
rect -300 -4380 1483 -4351
rect -300 -4413 0 -4380
rect -300 -4781 -151 -4413
rect -117 -4497 0 -4413
rect 180 -4451 340 -4380
rect 55 -4485 71 -4451
rect 447 -4485 463 -4451
rect 520 -4497 620 -4380
rect 800 -4451 960 -4380
rect 1140 -4413 1483 -4380
rect 673 -4485 689 -4451
rect 1065 -4485 1081 -4451
rect 1140 -4497 1253 -4413
rect -117 -4513 21 -4497
rect -117 -4681 -13 -4513
rect -117 -4697 21 -4681
rect 497 -4513 639 -4497
rect 531 -4681 605 -4513
rect 497 -4697 639 -4681
rect 1115 -4513 1253 -4497
rect 1149 -4681 1253 -4513
rect 1115 -4697 1253 -4681
rect -117 -4781 0 -4697
rect 55 -4743 71 -4709
rect 447 -4743 463 -4709
rect -300 -4843 0 -4781
rect 180 -4843 340 -4743
rect 520 -4843 620 -4697
rect 673 -4743 689 -4709
rect 1065 -4743 1081 -4709
rect 800 -4843 960 -4743
rect 1140 -4781 1253 -4697
rect 1287 -4781 1449 -4413
rect 2853 -4413 3083 -4351
rect 1655 -4485 1671 -4451
rect 2047 -4485 2063 -4451
rect 2273 -4485 2289 -4451
rect 2665 -4485 2681 -4451
rect 1587 -4513 1621 -4497
rect 1587 -4697 1621 -4681
rect 2097 -4513 2131 -4497
rect 2097 -4697 2131 -4681
rect 2205 -4513 2239 -4497
rect 2205 -4697 2239 -4681
rect 2715 -4513 2749 -4497
rect 2715 -4697 2749 -4681
rect 1655 -4743 1671 -4709
rect 2047 -4743 2063 -4709
rect 2273 -4743 2289 -4709
rect 2665 -4743 2681 -4709
rect 1140 -4843 1483 -4781
rect 2887 -4781 3049 -4413
rect 4453 -4413 4683 -4351
rect 3255 -4485 3271 -4451
rect 3647 -4485 3663 -4451
rect 3873 -4485 3889 -4451
rect 4265 -4485 4281 -4451
rect 3187 -4513 3221 -4497
rect 3187 -4697 3221 -4681
rect 3697 -4513 3731 -4497
rect 3697 -4697 3731 -4681
rect 3805 -4513 3839 -4497
rect 3805 -4697 3839 -4681
rect 4315 -4513 4349 -4497
rect 4315 -4697 4349 -4681
rect 3255 -4743 3271 -4709
rect 3647 -4743 3663 -4709
rect 3873 -4743 3889 -4709
rect 4265 -4743 4281 -4709
rect 2853 -4843 3083 -4781
rect 4487 -4781 4649 -4413
rect 6053 -4413 6283 -4351
rect 4855 -4485 4871 -4451
rect 5247 -4485 5263 -4451
rect 5473 -4485 5489 -4451
rect 5865 -4485 5881 -4451
rect 4787 -4513 4821 -4497
rect 4787 -4697 4821 -4681
rect 5297 -4513 5331 -4497
rect 5297 -4697 5331 -4681
rect 5405 -4513 5439 -4497
rect 5405 -4697 5439 -4681
rect 5915 -4513 5949 -4497
rect 5915 -4697 5949 -4681
rect 4855 -4743 4871 -4709
rect 5247 -4743 5263 -4709
rect 5473 -4743 5489 -4709
rect 5865 -4743 5881 -4709
rect 4453 -4843 4683 -4781
rect 6087 -4781 6249 -4413
rect 7653 -4413 7883 -4351
rect 6455 -4485 6471 -4451
rect 6847 -4485 6863 -4451
rect 7073 -4485 7089 -4451
rect 7465 -4485 7481 -4451
rect 6387 -4513 6421 -4497
rect 6387 -4697 6421 -4681
rect 6897 -4513 6931 -4497
rect 6897 -4697 6931 -4681
rect 7005 -4513 7039 -4497
rect 7005 -4697 7039 -4681
rect 7515 -4513 7549 -4497
rect 7515 -4697 7549 -4681
rect 6455 -4743 6471 -4709
rect 6847 -4743 6863 -4709
rect 7073 -4743 7089 -4709
rect 7465 -4743 7481 -4709
rect 6053 -4843 6283 -4781
rect 7687 -4781 7849 -4413
rect 9253 -4413 9483 -4351
rect 8055 -4485 8071 -4451
rect 8447 -4485 8463 -4451
rect 8673 -4485 8689 -4451
rect 9065 -4485 9081 -4451
rect 7987 -4513 8021 -4497
rect 7987 -4697 8021 -4681
rect 8497 -4513 8531 -4497
rect 8497 -4697 8531 -4681
rect 8605 -4513 8639 -4497
rect 8605 -4697 8639 -4681
rect 9115 -4513 9149 -4497
rect 9115 -4697 9149 -4681
rect 8055 -4743 8071 -4709
rect 8447 -4743 8463 -4709
rect 8673 -4743 8689 -4709
rect 9065 -4743 9081 -4709
rect 7653 -4843 7883 -4781
rect 9287 -4781 9449 -4413
rect 10853 -4413 11083 -4351
rect 9655 -4485 9671 -4451
rect 10047 -4485 10063 -4451
rect 10273 -4485 10289 -4451
rect 10665 -4485 10681 -4451
rect 9587 -4513 9621 -4497
rect 9587 -4697 9621 -4681
rect 10097 -4513 10131 -4497
rect 10097 -4697 10131 -4681
rect 10205 -4513 10239 -4497
rect 10205 -4697 10239 -4681
rect 10715 -4513 10749 -4497
rect 10715 -4697 10749 -4681
rect 9655 -4743 9671 -4709
rect 10047 -4743 10063 -4709
rect 10273 -4743 10289 -4709
rect 10665 -4743 10681 -4709
rect 9253 -4843 9483 -4781
rect 10887 -4781 11049 -4413
rect 12453 -4413 12683 -4351
rect 11255 -4485 11271 -4451
rect 11647 -4485 11663 -4451
rect 11873 -4485 11889 -4451
rect 12265 -4485 12281 -4451
rect 11187 -4513 11221 -4497
rect 11187 -4697 11221 -4681
rect 11697 -4513 11731 -4497
rect 11697 -4697 11731 -4681
rect 11805 -4513 11839 -4497
rect 11805 -4697 11839 -4681
rect 12315 -4513 12349 -4497
rect 12315 -4697 12349 -4681
rect 11255 -4743 11271 -4709
rect 11647 -4743 11663 -4709
rect 11873 -4743 11889 -4709
rect 12265 -4743 12281 -4709
rect 10853 -4843 11083 -4781
rect 12487 -4781 12649 -4413
rect 14053 -4413 14283 -4351
rect 12855 -4485 12871 -4451
rect 13247 -4485 13263 -4451
rect 13473 -4485 13489 -4451
rect 13865 -4485 13881 -4451
rect 12787 -4513 12821 -4497
rect 12787 -4697 12821 -4681
rect 13297 -4513 13331 -4497
rect 13297 -4697 13331 -4681
rect 13405 -4513 13439 -4497
rect 13405 -4697 13439 -4681
rect 13915 -4513 13949 -4497
rect 13915 -4697 13949 -4681
rect 12855 -4743 12871 -4709
rect 13247 -4743 13263 -4709
rect 13473 -4743 13489 -4709
rect 13865 -4743 13881 -4709
rect 12453 -4843 12683 -4781
rect 14087 -4781 14249 -4413
rect 15653 -4413 15883 -4351
rect 14455 -4485 14471 -4451
rect 14847 -4485 14863 -4451
rect 15073 -4485 15089 -4451
rect 15465 -4485 15481 -4451
rect 14387 -4513 14421 -4497
rect 14387 -4697 14421 -4681
rect 14897 -4513 14931 -4497
rect 14897 -4697 14931 -4681
rect 15005 -4513 15039 -4497
rect 15005 -4697 15039 -4681
rect 15515 -4513 15549 -4497
rect 15515 -4697 15549 -4681
rect 14455 -4743 14471 -4709
rect 14847 -4743 14863 -4709
rect 15073 -4743 15089 -4709
rect 15465 -4743 15481 -4709
rect 14053 -4843 14283 -4781
rect 15687 -4781 15849 -4413
rect 17253 -4413 17483 -4351
rect 16055 -4485 16071 -4451
rect 16447 -4485 16463 -4451
rect 16673 -4485 16689 -4451
rect 17065 -4485 17081 -4451
rect 15987 -4513 16021 -4497
rect 15987 -4697 16021 -4681
rect 16497 -4513 16531 -4497
rect 16497 -4697 16531 -4681
rect 16605 -4513 16639 -4497
rect 16605 -4697 16639 -4681
rect 17115 -4513 17149 -4497
rect 17115 -4697 17149 -4681
rect 16055 -4743 16071 -4709
rect 16447 -4743 16463 -4709
rect 16673 -4743 16689 -4709
rect 17065 -4743 17081 -4709
rect 15653 -4843 15883 -4781
rect 17287 -4781 17449 -4413
rect 18853 -4413 19083 -4351
rect 17655 -4485 17671 -4451
rect 18047 -4485 18063 -4451
rect 18273 -4485 18289 -4451
rect 18665 -4485 18681 -4451
rect 17587 -4513 17621 -4497
rect 17587 -4697 17621 -4681
rect 18097 -4513 18131 -4497
rect 18097 -4697 18131 -4681
rect 18205 -4513 18239 -4497
rect 18205 -4697 18239 -4681
rect 18715 -4513 18749 -4497
rect 18715 -4697 18749 -4681
rect 17655 -4743 17671 -4709
rect 18047 -4743 18063 -4709
rect 18273 -4743 18289 -4709
rect 18665 -4743 18681 -4709
rect 17253 -4843 17483 -4781
rect 18887 -4781 19049 -4413
rect 20453 -4413 20683 -4351
rect 19255 -4485 19271 -4451
rect 19647 -4485 19663 -4451
rect 19873 -4485 19889 -4451
rect 20265 -4485 20281 -4451
rect 19187 -4513 19221 -4497
rect 19187 -4697 19221 -4681
rect 19697 -4513 19731 -4497
rect 19697 -4697 19731 -4681
rect 19805 -4513 19839 -4497
rect 19805 -4697 19839 -4681
rect 20315 -4513 20349 -4497
rect 20315 -4697 20349 -4681
rect 19255 -4743 19271 -4709
rect 19647 -4743 19663 -4709
rect 19873 -4743 19889 -4709
rect 20265 -4743 20281 -4709
rect 18853 -4843 19083 -4781
rect 20487 -4781 20649 -4413
rect 22053 -4413 22283 -4351
rect 20855 -4485 20871 -4451
rect 21247 -4485 21263 -4451
rect 21473 -4485 21489 -4451
rect 21865 -4485 21881 -4451
rect 20787 -4513 20821 -4497
rect 20787 -4697 20821 -4681
rect 21297 -4513 21331 -4497
rect 21297 -4697 21331 -4681
rect 21405 -4513 21439 -4497
rect 21405 -4697 21439 -4681
rect 21915 -4513 21949 -4497
rect 21915 -4697 21949 -4681
rect 20855 -4743 20871 -4709
rect 21247 -4743 21263 -4709
rect 21473 -4743 21489 -4709
rect 21865 -4743 21881 -4709
rect 20453 -4843 20683 -4781
rect 22087 -4781 22249 -4413
rect 23653 -4413 23883 -4351
rect 22455 -4485 22471 -4451
rect 22847 -4485 22863 -4451
rect 23073 -4485 23089 -4451
rect 23465 -4485 23481 -4451
rect 22387 -4513 22421 -4497
rect 22387 -4697 22421 -4681
rect 22897 -4513 22931 -4497
rect 22897 -4697 22931 -4681
rect 23005 -4513 23039 -4497
rect 23005 -4697 23039 -4681
rect 23515 -4513 23549 -4497
rect 23515 -4697 23549 -4681
rect 22455 -4743 22471 -4709
rect 22847 -4743 22863 -4709
rect 23073 -4743 23089 -4709
rect 23465 -4743 23481 -4709
rect 22053 -4843 22283 -4781
rect 23687 -4781 23849 -4413
rect 25253 -4413 25483 -4351
rect 24055 -4485 24071 -4451
rect 24447 -4485 24463 -4451
rect 24673 -4485 24689 -4451
rect 25065 -4485 25081 -4451
rect 23987 -4513 24021 -4497
rect 23987 -4697 24021 -4681
rect 24497 -4513 24531 -4497
rect 24497 -4697 24531 -4681
rect 24605 -4513 24639 -4497
rect 24605 -4697 24639 -4681
rect 25115 -4513 25149 -4497
rect 25115 -4697 25149 -4681
rect 24055 -4743 24071 -4709
rect 24447 -4743 24463 -4709
rect 24673 -4743 24689 -4709
rect 25065 -4743 25081 -4709
rect 23653 -4843 23883 -4781
rect 25287 -4781 25449 -4413
rect 26853 -4413 27083 -4351
rect 25655 -4485 25671 -4451
rect 26047 -4485 26063 -4451
rect 26273 -4485 26289 -4451
rect 26665 -4485 26681 -4451
rect 25587 -4513 25621 -4497
rect 25587 -4697 25621 -4681
rect 26097 -4513 26131 -4497
rect 26097 -4697 26131 -4681
rect 26205 -4513 26239 -4497
rect 26205 -4697 26239 -4681
rect 26715 -4513 26749 -4497
rect 26715 -4697 26749 -4681
rect 25655 -4743 25671 -4709
rect 26047 -4743 26063 -4709
rect 26273 -4743 26289 -4709
rect 26665 -4743 26681 -4709
rect 25253 -4843 25483 -4781
rect 26887 -4781 27049 -4413
rect 28453 -4413 28683 -4351
rect 27255 -4485 27271 -4451
rect 27647 -4485 27663 -4451
rect 27873 -4485 27889 -4451
rect 28265 -4485 28281 -4451
rect 27187 -4513 27221 -4497
rect 27187 -4697 27221 -4681
rect 27697 -4513 27731 -4497
rect 27697 -4697 27731 -4681
rect 27805 -4513 27839 -4497
rect 27805 -4697 27839 -4681
rect 28315 -4513 28349 -4497
rect 28315 -4697 28349 -4681
rect 27255 -4743 27271 -4709
rect 27647 -4743 27663 -4709
rect 27873 -4743 27889 -4709
rect 28265 -4743 28281 -4709
rect 26853 -4843 27083 -4781
rect 28487 -4781 28649 -4413
rect 30053 -4413 30283 -4351
rect 28855 -4485 28871 -4451
rect 29247 -4485 29263 -4451
rect 29473 -4485 29489 -4451
rect 29865 -4485 29881 -4451
rect 28787 -4513 28821 -4497
rect 28787 -4697 28821 -4681
rect 29297 -4513 29331 -4497
rect 29297 -4697 29331 -4681
rect 29405 -4513 29439 -4497
rect 29405 -4697 29439 -4681
rect 29915 -4513 29949 -4497
rect 29915 -4697 29949 -4681
rect 28855 -4743 28871 -4709
rect 29247 -4743 29263 -4709
rect 29473 -4743 29489 -4709
rect 29865 -4743 29881 -4709
rect 28453 -4843 28683 -4781
rect 30087 -4781 30249 -4413
rect 31653 -4413 31883 -4351
rect 30455 -4485 30471 -4451
rect 30847 -4485 30863 -4451
rect 31073 -4485 31089 -4451
rect 31465 -4485 31481 -4451
rect 30387 -4513 30421 -4497
rect 30387 -4697 30421 -4681
rect 30897 -4513 30931 -4497
rect 30897 -4697 30931 -4681
rect 31005 -4513 31039 -4497
rect 31005 -4697 31039 -4681
rect 31515 -4513 31549 -4497
rect 31515 -4697 31549 -4681
rect 30455 -4743 30471 -4709
rect 30847 -4743 30863 -4709
rect 31073 -4743 31089 -4709
rect 31465 -4743 31481 -4709
rect 30053 -4843 30283 -4781
rect 31687 -4781 31849 -4413
rect 33253 -4413 33483 -4351
rect 32055 -4485 32071 -4451
rect 32447 -4485 32463 -4451
rect 32673 -4485 32689 -4451
rect 33065 -4485 33081 -4451
rect 31987 -4513 32021 -4497
rect 31987 -4697 32021 -4681
rect 32497 -4513 32531 -4497
rect 32497 -4697 32531 -4681
rect 32605 -4513 32639 -4497
rect 32605 -4697 32639 -4681
rect 33115 -4513 33149 -4497
rect 33115 -4697 33149 -4681
rect 32055 -4743 32071 -4709
rect 32447 -4743 32463 -4709
rect 32673 -4743 32689 -4709
rect 33065 -4743 33081 -4709
rect 31653 -4843 31883 -4781
rect 33287 -4781 33449 -4413
rect 34853 -4413 35083 -4351
rect 33655 -4485 33671 -4451
rect 34047 -4485 34063 -4451
rect 34273 -4485 34289 -4451
rect 34665 -4485 34681 -4451
rect 33587 -4513 33621 -4497
rect 33587 -4697 33621 -4681
rect 34097 -4513 34131 -4497
rect 34097 -4697 34131 -4681
rect 34205 -4513 34239 -4497
rect 34205 -4697 34239 -4681
rect 34715 -4513 34749 -4497
rect 34715 -4697 34749 -4681
rect 33655 -4743 33671 -4709
rect 34047 -4743 34063 -4709
rect 34273 -4743 34289 -4709
rect 34665 -4743 34681 -4709
rect 33253 -4843 33483 -4781
rect 34887 -4781 35049 -4413
rect 36453 -4380 38400 -4351
rect 36453 -4413 36800 -4380
rect 35255 -4485 35271 -4451
rect 35647 -4485 35663 -4451
rect 35873 -4485 35889 -4451
rect 36265 -4485 36281 -4451
rect 35187 -4513 35221 -4497
rect 35187 -4697 35221 -4681
rect 35697 -4513 35731 -4497
rect 35697 -4697 35731 -4681
rect 35805 -4513 35839 -4497
rect 35805 -4697 35839 -4681
rect 36315 -4513 36349 -4497
rect 36315 -4697 36349 -4681
rect 35255 -4743 35271 -4709
rect 35647 -4743 35663 -4709
rect 35873 -4743 35889 -4709
rect 36265 -4743 36281 -4709
rect 34853 -4843 35083 -4781
rect 36487 -4781 36649 -4413
rect 36683 -4497 36800 -4413
rect 36980 -4451 37140 -4380
rect 36855 -4485 36871 -4451
rect 37247 -4485 37263 -4451
rect 37320 -4497 37420 -4380
rect 37600 -4451 37760 -4380
rect 37940 -4413 38400 -4380
rect 37473 -4485 37489 -4451
rect 37865 -4485 37881 -4451
rect 37940 -4497 38053 -4413
rect 36683 -4513 36821 -4497
rect 36683 -4681 36787 -4513
rect 36683 -4697 36821 -4681
rect 37297 -4513 37439 -4497
rect 37331 -4681 37405 -4513
rect 37297 -4697 37439 -4681
rect 37915 -4513 38053 -4497
rect 37949 -4681 38053 -4513
rect 37915 -4697 38053 -4681
rect 36683 -4781 36800 -4697
rect 36855 -4743 36871 -4709
rect 37247 -4743 37263 -4709
rect 36453 -4843 36800 -4781
rect 36980 -4843 37140 -4743
rect 37320 -4843 37420 -4697
rect 37473 -4743 37489 -4709
rect 37865 -4743 37881 -4709
rect 37600 -4843 37760 -4743
rect 37940 -4781 38053 -4697
rect 38087 -4781 38400 -4413
rect 37940 -4843 38400 -4781
rect -300 -5600 38400 -4843
rect -140 -8036 38100 -7840
rect -162 -8070 -66 -8036
rect 1216 -8070 1534 -8036
rect 2816 -8060 3134 -8036
rect 2816 -8070 2912 -8060
rect -162 -8132 1472 -8070
rect -128 -8170 1278 -8132
rect -128 -8204 69 -8170
rect 445 -8204 705 -8170
rect 1081 -8204 1278 -8170
rect -128 -8232 1278 -8204
rect -128 -8400 -24 -8232
rect 10 -8400 504 -8232
rect 538 -8400 612 -8232
rect 646 -8400 1140 -8232
rect 1174 -8400 1278 -8232
rect -128 -8428 1278 -8400
rect -128 -8462 69 -8428
rect 445 -8462 705 -8428
rect 1081 -8462 1278 -8428
rect -128 -8500 1278 -8462
rect 1312 -8500 1438 -8132
rect 2878 -8132 2912 -8070
rect 1653 -8204 1669 -8170
rect 2045 -8204 2061 -8170
rect 2289 -8204 2305 -8170
rect 2681 -8204 2697 -8170
rect 1576 -8232 1610 -8216
rect 1576 -8416 1610 -8400
rect 2104 -8232 2138 -8216
rect 2104 -8416 2138 -8400
rect 2212 -8232 2246 -8216
rect 2212 -8416 2246 -8400
rect 2740 -8232 2774 -8216
rect 2740 -8416 2774 -8400
rect 1653 -8462 1669 -8428
rect 2045 -8462 2061 -8428
rect 2289 -8462 2305 -8428
rect 2681 -8462 2697 -8428
rect -162 -8562 1472 -8500
rect 2878 -8562 2912 -8500
rect -162 -8596 -66 -8562
rect 1216 -8596 1534 -8562
rect 2816 -8596 2912 -8562
rect -162 -8658 1472 -8596
rect -128 -8696 1278 -8658
rect -128 -8730 69 -8696
rect 445 -8730 705 -8696
rect 1081 -8730 1278 -8696
rect -128 -8758 1278 -8730
rect -128 -9526 -24 -8758
rect 10 -9526 504 -8758
rect 538 -9526 612 -8758
rect 646 -9526 1140 -8758
rect 1174 -9526 1278 -8758
rect -128 -9554 1278 -9526
rect -128 -9588 69 -9554
rect 445 -9588 705 -9554
rect 1081 -9588 1278 -9554
rect -128 -9626 1278 -9588
rect 1312 -9626 1438 -8658
rect 2878 -8658 2912 -8596
rect 1653 -8730 1669 -8696
rect 2045 -8730 2061 -8696
rect 2289 -8730 2305 -8696
rect 2681 -8730 2697 -8696
rect 1576 -8758 1610 -8742
rect 1576 -9542 1610 -9526
rect 2104 -8758 2138 -8742
rect 2104 -9542 2138 -9526
rect 2212 -8758 2246 -8742
rect 2212 -9542 2246 -9526
rect 2740 -8758 2774 -8742
rect 2740 -9542 2774 -9526
rect 1653 -9588 1669 -9554
rect 2045 -9588 2061 -9554
rect 2289 -9588 2305 -9554
rect 2681 -9588 2697 -9554
rect -162 -9688 1472 -9626
rect 2878 -9688 2912 -9626
rect -162 -9722 -66 -9688
rect 1216 -9722 1534 -9688
rect 2816 -9722 2912 -9688
rect 3038 -8070 3134 -8060
rect 4416 -8060 4734 -8036
rect 4416 -8070 4512 -8060
rect 3038 -8132 3072 -8070
rect 4478 -8132 4512 -8070
rect 3253 -8204 3269 -8170
rect 3645 -8204 3661 -8170
rect 3889 -8204 3905 -8170
rect 4281 -8204 4297 -8170
rect 3176 -8232 3210 -8216
rect 3176 -8416 3210 -8400
rect 3704 -8232 3738 -8216
rect 3704 -8416 3738 -8400
rect 3812 -8232 3846 -8216
rect 3812 -8416 3846 -8400
rect 4340 -8232 4374 -8216
rect 4340 -8416 4374 -8400
rect 3253 -8462 3269 -8428
rect 3645 -8462 3661 -8428
rect 3889 -8462 3905 -8428
rect 4281 -8462 4297 -8428
rect 3038 -8562 3072 -8500
rect 4478 -8562 4512 -8500
rect 3038 -8596 3134 -8562
rect 4416 -8596 4512 -8562
rect 3038 -8658 3072 -8596
rect 4478 -8658 4512 -8596
rect 3253 -8730 3269 -8696
rect 3645 -8730 3661 -8696
rect 3889 -8730 3905 -8696
rect 4281 -8730 4297 -8696
rect 3176 -8758 3210 -8742
rect 3176 -9542 3210 -9526
rect 3704 -8758 3738 -8742
rect 3704 -9542 3738 -9526
rect 3812 -8758 3846 -8742
rect 3812 -9542 3846 -9526
rect 4340 -8758 4374 -8742
rect 4340 -9542 4374 -9526
rect 3253 -9588 3269 -9554
rect 3645 -9588 3661 -9554
rect 3889 -9588 3905 -9554
rect 4281 -9588 4297 -9554
rect 3038 -9688 3072 -9626
rect 4478 -9688 4512 -9626
rect 3038 -9722 3134 -9688
rect 4416 -9722 4512 -9688
rect 4638 -8070 4734 -8060
rect 6016 -8060 6334 -8036
rect 6016 -8070 6112 -8060
rect 4638 -8132 4672 -8070
rect 6078 -8132 6112 -8070
rect 4853 -8204 4869 -8170
rect 5245 -8204 5261 -8170
rect 5489 -8204 5505 -8170
rect 5881 -8204 5897 -8170
rect 4776 -8232 4810 -8216
rect 4776 -8416 4810 -8400
rect 5304 -8232 5338 -8216
rect 5304 -8416 5338 -8400
rect 5412 -8232 5446 -8216
rect 5412 -8416 5446 -8400
rect 5940 -8232 5974 -8216
rect 5940 -8416 5974 -8400
rect 4853 -8462 4869 -8428
rect 5245 -8462 5261 -8428
rect 5489 -8462 5505 -8428
rect 5881 -8462 5897 -8428
rect 4638 -8562 4672 -8500
rect 6078 -8562 6112 -8500
rect 4638 -8596 4734 -8562
rect 6016 -8596 6112 -8562
rect 4638 -8658 4672 -8596
rect 6078 -8658 6112 -8596
rect 4853 -8730 4869 -8696
rect 5245 -8730 5261 -8696
rect 5489 -8730 5505 -8696
rect 5881 -8730 5897 -8696
rect 4776 -8758 4810 -8742
rect 4776 -9542 4810 -9526
rect 5304 -8758 5338 -8742
rect 5304 -9542 5338 -9526
rect 5412 -8758 5446 -8742
rect 5412 -9542 5446 -9526
rect 5940 -8758 5974 -8742
rect 5940 -9542 5974 -9526
rect 4853 -9588 4869 -9554
rect 5245 -9588 5261 -9554
rect 5489 -9588 5505 -9554
rect 5881 -9588 5897 -9554
rect 4638 -9688 4672 -9626
rect 6078 -9688 6112 -9626
rect 4638 -9722 4734 -9688
rect 6016 -9722 6112 -9688
rect 6238 -8070 6334 -8060
rect 7616 -8060 7934 -8036
rect 7616 -8070 7712 -8060
rect 6238 -8132 6272 -8070
rect 7678 -8132 7712 -8070
rect 6453 -8204 6469 -8170
rect 6845 -8204 6861 -8170
rect 7089 -8204 7105 -8170
rect 7481 -8204 7497 -8170
rect 6376 -8232 6410 -8216
rect 6376 -8416 6410 -8400
rect 6904 -8232 6938 -8216
rect 6904 -8416 6938 -8400
rect 7012 -8232 7046 -8216
rect 7012 -8416 7046 -8400
rect 7540 -8232 7574 -8216
rect 7540 -8416 7574 -8400
rect 6453 -8462 6469 -8428
rect 6845 -8462 6861 -8428
rect 7089 -8462 7105 -8428
rect 7481 -8462 7497 -8428
rect 6238 -8562 6272 -8500
rect 7678 -8562 7712 -8500
rect 6238 -8596 6334 -8562
rect 7616 -8596 7712 -8562
rect 6238 -8658 6272 -8596
rect 7678 -8658 7712 -8596
rect 6453 -8730 6469 -8696
rect 6845 -8730 6861 -8696
rect 7089 -8730 7105 -8696
rect 7481 -8730 7497 -8696
rect 6376 -8758 6410 -8742
rect 6376 -9542 6410 -9526
rect 6904 -8758 6938 -8742
rect 6904 -9542 6938 -9526
rect 7012 -8758 7046 -8742
rect 7012 -9542 7046 -9526
rect 7540 -8758 7574 -8742
rect 7540 -9542 7574 -9526
rect 6453 -9588 6469 -9554
rect 6845 -9588 6861 -9554
rect 7089 -9588 7105 -9554
rect 7481 -9588 7497 -9554
rect 6238 -9688 6272 -9626
rect 7678 -9688 7712 -9626
rect 6238 -9722 6334 -9688
rect 7616 -9722 7712 -9688
rect 7838 -8070 7934 -8060
rect 9216 -8060 9534 -8036
rect 9216 -8070 9312 -8060
rect 7838 -8132 7872 -8070
rect 9278 -8132 9312 -8070
rect 8053 -8204 8069 -8170
rect 8445 -8204 8461 -8170
rect 8689 -8204 8705 -8170
rect 9081 -8204 9097 -8170
rect 7976 -8232 8010 -8216
rect 7976 -8416 8010 -8400
rect 8504 -8232 8538 -8216
rect 8504 -8416 8538 -8400
rect 8612 -8232 8646 -8216
rect 8612 -8416 8646 -8400
rect 9140 -8232 9174 -8216
rect 9140 -8416 9174 -8400
rect 8053 -8462 8069 -8428
rect 8445 -8462 8461 -8428
rect 8689 -8462 8705 -8428
rect 9081 -8462 9097 -8428
rect 7838 -8562 7872 -8500
rect 9278 -8562 9312 -8500
rect 7838 -8596 7934 -8562
rect 9216 -8596 9312 -8562
rect 7838 -8658 7872 -8596
rect 9278 -8658 9312 -8596
rect 8053 -8730 8069 -8696
rect 8445 -8730 8461 -8696
rect 8689 -8730 8705 -8696
rect 9081 -8730 9097 -8696
rect 7976 -8758 8010 -8742
rect 7976 -9542 8010 -9526
rect 8504 -8758 8538 -8742
rect 8504 -9542 8538 -9526
rect 8612 -8758 8646 -8742
rect 8612 -9542 8646 -9526
rect 9140 -8758 9174 -8742
rect 9140 -9542 9174 -9526
rect 8053 -9588 8069 -9554
rect 8445 -9588 8461 -9554
rect 8689 -9588 8705 -9554
rect 9081 -9588 9097 -9554
rect 7838 -9688 7872 -9626
rect 9278 -9688 9312 -9626
rect 7838 -9722 7934 -9688
rect 9216 -9722 9312 -9688
rect 9438 -8070 9534 -8060
rect 10816 -8060 11134 -8036
rect 10816 -8070 10912 -8060
rect 9438 -8132 9472 -8070
rect 10878 -8132 10912 -8070
rect 9653 -8204 9669 -8170
rect 10045 -8204 10061 -8170
rect 10289 -8204 10305 -8170
rect 10681 -8204 10697 -8170
rect 9576 -8232 9610 -8216
rect 9576 -8416 9610 -8400
rect 10104 -8232 10138 -8216
rect 10104 -8416 10138 -8400
rect 10212 -8232 10246 -8216
rect 10212 -8416 10246 -8400
rect 10740 -8232 10774 -8216
rect 10740 -8416 10774 -8400
rect 9653 -8462 9669 -8428
rect 10045 -8462 10061 -8428
rect 10289 -8462 10305 -8428
rect 10681 -8462 10697 -8428
rect 9438 -8562 9472 -8500
rect 10878 -8562 10912 -8500
rect 9438 -8596 9534 -8562
rect 10816 -8596 10912 -8562
rect 9438 -8658 9472 -8596
rect 10878 -8658 10912 -8596
rect 9653 -8730 9669 -8696
rect 10045 -8730 10061 -8696
rect 10289 -8730 10305 -8696
rect 10681 -8730 10697 -8696
rect 9576 -8758 9610 -8742
rect 9576 -9542 9610 -9526
rect 10104 -8758 10138 -8742
rect 10104 -9542 10138 -9526
rect 10212 -8758 10246 -8742
rect 10212 -9542 10246 -9526
rect 10740 -8758 10774 -8742
rect 10740 -9542 10774 -9526
rect 9653 -9588 9669 -9554
rect 10045 -9588 10061 -9554
rect 10289 -9588 10305 -9554
rect 10681 -9588 10697 -9554
rect 9438 -9688 9472 -9626
rect 10878 -9688 10912 -9626
rect 9438 -9722 9534 -9688
rect 10816 -9722 10912 -9688
rect 11038 -8070 11134 -8060
rect 12416 -8060 12734 -8036
rect 12416 -8070 12512 -8060
rect 11038 -8132 11072 -8070
rect 12478 -8132 12512 -8070
rect 11253 -8204 11269 -8170
rect 11645 -8204 11661 -8170
rect 11889 -8204 11905 -8170
rect 12281 -8204 12297 -8170
rect 11176 -8232 11210 -8216
rect 11176 -8416 11210 -8400
rect 11704 -8232 11738 -8216
rect 11704 -8416 11738 -8400
rect 11812 -8232 11846 -8216
rect 11812 -8416 11846 -8400
rect 12340 -8232 12374 -8216
rect 12340 -8416 12374 -8400
rect 11253 -8462 11269 -8428
rect 11645 -8462 11661 -8428
rect 11889 -8462 11905 -8428
rect 12281 -8462 12297 -8428
rect 11038 -8562 11072 -8500
rect 12478 -8562 12512 -8500
rect 11038 -8596 11134 -8562
rect 12416 -8596 12512 -8562
rect 11038 -8658 11072 -8596
rect 12478 -8658 12512 -8596
rect 11253 -8730 11269 -8696
rect 11645 -8730 11661 -8696
rect 11889 -8730 11905 -8696
rect 12281 -8730 12297 -8696
rect 11176 -8758 11210 -8742
rect 11176 -9542 11210 -9526
rect 11704 -8758 11738 -8742
rect 11704 -9542 11738 -9526
rect 11812 -8758 11846 -8742
rect 11812 -9542 11846 -9526
rect 12340 -8758 12374 -8742
rect 12340 -9542 12374 -9526
rect 11253 -9588 11269 -9554
rect 11645 -9588 11661 -9554
rect 11889 -9588 11905 -9554
rect 12281 -9588 12297 -9554
rect 11038 -9688 11072 -9626
rect 12478 -9688 12512 -9626
rect 11038 -9722 11134 -9688
rect 12416 -9722 12512 -9688
rect 12638 -8070 12734 -8060
rect 14016 -8060 14334 -8036
rect 14016 -8070 14112 -8060
rect 12638 -8132 12672 -8070
rect 14078 -8132 14112 -8070
rect 12853 -8204 12869 -8170
rect 13245 -8204 13261 -8170
rect 13489 -8204 13505 -8170
rect 13881 -8204 13897 -8170
rect 12776 -8232 12810 -8216
rect 12776 -8416 12810 -8400
rect 13304 -8232 13338 -8216
rect 13304 -8416 13338 -8400
rect 13412 -8232 13446 -8216
rect 13412 -8416 13446 -8400
rect 13940 -8232 13974 -8216
rect 13940 -8416 13974 -8400
rect 12853 -8462 12869 -8428
rect 13245 -8462 13261 -8428
rect 13489 -8462 13505 -8428
rect 13881 -8462 13897 -8428
rect 12638 -8562 12672 -8500
rect 14078 -8562 14112 -8500
rect 12638 -8596 12734 -8562
rect 14016 -8596 14112 -8562
rect 12638 -8658 12672 -8596
rect 14078 -8658 14112 -8596
rect 12853 -8730 12869 -8696
rect 13245 -8730 13261 -8696
rect 13489 -8730 13505 -8696
rect 13881 -8730 13897 -8696
rect 12776 -8758 12810 -8742
rect 12776 -9542 12810 -9526
rect 13304 -8758 13338 -8742
rect 13304 -9542 13338 -9526
rect 13412 -8758 13446 -8742
rect 13412 -9542 13446 -9526
rect 13940 -8758 13974 -8742
rect 13940 -9542 13974 -9526
rect 12853 -9588 12869 -9554
rect 13245 -9588 13261 -9554
rect 13489 -9588 13505 -9554
rect 13881 -9588 13897 -9554
rect 12638 -9688 12672 -9626
rect 14078 -9688 14112 -9626
rect 12638 -9722 12734 -9688
rect 14016 -9722 14112 -9688
rect 14238 -8070 14334 -8060
rect 15616 -8060 15934 -8036
rect 15616 -8070 15712 -8060
rect 14238 -8132 14272 -8070
rect 15678 -8132 15712 -8070
rect 14453 -8204 14469 -8170
rect 14845 -8204 14861 -8170
rect 15089 -8204 15105 -8170
rect 15481 -8204 15497 -8170
rect 14376 -8232 14410 -8216
rect 14376 -8416 14410 -8400
rect 14904 -8232 14938 -8216
rect 14904 -8416 14938 -8400
rect 15012 -8232 15046 -8216
rect 15012 -8416 15046 -8400
rect 15540 -8232 15574 -8216
rect 15540 -8416 15574 -8400
rect 14453 -8462 14469 -8428
rect 14845 -8462 14861 -8428
rect 15089 -8462 15105 -8428
rect 15481 -8462 15497 -8428
rect 14238 -8562 14272 -8500
rect 15678 -8562 15712 -8500
rect 14238 -8596 14334 -8562
rect 15616 -8596 15712 -8562
rect 14238 -8658 14272 -8596
rect 15678 -8658 15712 -8596
rect 14453 -8730 14469 -8696
rect 14845 -8730 14861 -8696
rect 15089 -8730 15105 -8696
rect 15481 -8730 15497 -8696
rect 14376 -8758 14410 -8742
rect 14376 -9542 14410 -9526
rect 14904 -8758 14938 -8742
rect 14904 -9542 14938 -9526
rect 15012 -8758 15046 -8742
rect 15012 -9542 15046 -9526
rect 15540 -8758 15574 -8742
rect 15540 -9542 15574 -9526
rect 14453 -9588 14469 -9554
rect 14845 -9588 14861 -9554
rect 15089 -9588 15105 -9554
rect 15481 -9588 15497 -9554
rect 14238 -9688 14272 -9626
rect 15678 -9688 15712 -9626
rect 14238 -9722 14334 -9688
rect 15616 -9722 15712 -9688
rect 15838 -8070 15934 -8060
rect 17216 -8060 17534 -8036
rect 17216 -8070 17312 -8060
rect 15838 -8132 15872 -8070
rect 17278 -8132 17312 -8070
rect 16053 -8204 16069 -8170
rect 16445 -8204 16461 -8170
rect 16689 -8204 16705 -8170
rect 17081 -8204 17097 -8170
rect 15976 -8232 16010 -8216
rect 15976 -8416 16010 -8400
rect 16504 -8232 16538 -8216
rect 16504 -8416 16538 -8400
rect 16612 -8232 16646 -8216
rect 16612 -8416 16646 -8400
rect 17140 -8232 17174 -8216
rect 17140 -8416 17174 -8400
rect 16053 -8462 16069 -8428
rect 16445 -8462 16461 -8428
rect 16689 -8462 16705 -8428
rect 17081 -8462 17097 -8428
rect 15838 -8562 15872 -8500
rect 17278 -8562 17312 -8500
rect 15838 -8596 15934 -8562
rect 17216 -8596 17312 -8562
rect 15838 -8658 15872 -8596
rect 17278 -8658 17312 -8596
rect 16053 -8730 16069 -8696
rect 16445 -8730 16461 -8696
rect 16689 -8730 16705 -8696
rect 17081 -8730 17097 -8696
rect 15976 -8758 16010 -8742
rect 15976 -9542 16010 -9526
rect 16504 -8758 16538 -8742
rect 16504 -9542 16538 -9526
rect 16612 -8758 16646 -8742
rect 16612 -9542 16646 -9526
rect 17140 -8758 17174 -8742
rect 17140 -9542 17174 -9526
rect 16053 -9588 16069 -9554
rect 16445 -9588 16461 -9554
rect 16689 -9588 16705 -9554
rect 17081 -9588 17097 -9554
rect 15838 -9688 15872 -9626
rect 17278 -9688 17312 -9626
rect 15838 -9722 15934 -9688
rect 17216 -9722 17312 -9688
rect 17438 -8070 17534 -8060
rect 18816 -8060 19134 -8036
rect 18816 -8070 18912 -8060
rect 17438 -8132 17472 -8070
rect 18878 -8132 18912 -8070
rect 17653 -8204 17669 -8170
rect 18045 -8204 18061 -8170
rect 18289 -8204 18305 -8170
rect 18681 -8204 18697 -8170
rect 17576 -8232 17610 -8216
rect 17576 -8416 17610 -8400
rect 18104 -8232 18138 -8216
rect 18104 -8416 18138 -8400
rect 18212 -8232 18246 -8216
rect 18212 -8416 18246 -8400
rect 18740 -8232 18774 -8216
rect 18740 -8416 18774 -8400
rect 17653 -8462 17669 -8428
rect 18045 -8462 18061 -8428
rect 18289 -8462 18305 -8428
rect 18681 -8462 18697 -8428
rect 17438 -8562 17472 -8500
rect 18878 -8562 18912 -8500
rect 17438 -8596 17534 -8562
rect 18816 -8596 18912 -8562
rect 17438 -8658 17472 -8596
rect 18878 -8658 18912 -8596
rect 17653 -8730 17669 -8696
rect 18045 -8730 18061 -8696
rect 18289 -8730 18305 -8696
rect 18681 -8730 18697 -8696
rect 17576 -8758 17610 -8742
rect 17576 -9542 17610 -9526
rect 18104 -8758 18138 -8742
rect 18104 -9542 18138 -9526
rect 18212 -8758 18246 -8742
rect 18212 -9542 18246 -9526
rect 18740 -8758 18774 -8742
rect 18740 -9542 18774 -9526
rect 17653 -9588 17669 -9554
rect 18045 -9588 18061 -9554
rect 18289 -9588 18305 -9554
rect 18681 -9588 18697 -9554
rect 17438 -9688 17472 -9626
rect 18878 -9688 18912 -9626
rect 17438 -9722 17534 -9688
rect 18816 -9722 18912 -9688
rect 19038 -8070 19134 -8060
rect 20416 -8060 20734 -8036
rect 20416 -8070 20512 -8060
rect 19038 -8132 19072 -8070
rect 20478 -8132 20512 -8070
rect 19253 -8204 19269 -8170
rect 19645 -8204 19661 -8170
rect 19889 -8204 19905 -8170
rect 20281 -8204 20297 -8170
rect 19176 -8232 19210 -8216
rect 19176 -8416 19210 -8400
rect 19704 -8232 19738 -8216
rect 19704 -8416 19738 -8400
rect 19812 -8232 19846 -8216
rect 19812 -8416 19846 -8400
rect 20340 -8232 20374 -8216
rect 20340 -8416 20374 -8400
rect 19253 -8462 19269 -8428
rect 19645 -8462 19661 -8428
rect 19889 -8462 19905 -8428
rect 20281 -8462 20297 -8428
rect 19038 -8562 19072 -8500
rect 20478 -8562 20512 -8500
rect 19038 -8596 19134 -8562
rect 20416 -8596 20512 -8562
rect 19038 -8658 19072 -8596
rect 20478 -8658 20512 -8596
rect 19253 -8730 19269 -8696
rect 19645 -8730 19661 -8696
rect 19889 -8730 19905 -8696
rect 20281 -8730 20297 -8696
rect 19176 -8758 19210 -8742
rect 19176 -9542 19210 -9526
rect 19704 -8758 19738 -8742
rect 19704 -9542 19738 -9526
rect 19812 -8758 19846 -8742
rect 19812 -9542 19846 -9526
rect 20340 -8758 20374 -8742
rect 20340 -9542 20374 -9526
rect 19253 -9588 19269 -9554
rect 19645 -9588 19661 -9554
rect 19889 -9588 19905 -9554
rect 20281 -9588 20297 -9554
rect 19038 -9688 19072 -9626
rect 20478 -9688 20512 -9626
rect 19038 -9722 19134 -9688
rect 20416 -9722 20512 -9688
rect 20638 -8070 20734 -8060
rect 22016 -8060 22334 -8036
rect 22016 -8070 22112 -8060
rect 20638 -8132 20672 -8070
rect 22078 -8132 22112 -8070
rect 20853 -8204 20869 -8170
rect 21245 -8204 21261 -8170
rect 21489 -8204 21505 -8170
rect 21881 -8204 21897 -8170
rect 20776 -8232 20810 -8216
rect 20776 -8416 20810 -8400
rect 21304 -8232 21338 -8216
rect 21304 -8416 21338 -8400
rect 21412 -8232 21446 -8216
rect 21412 -8416 21446 -8400
rect 21940 -8232 21974 -8216
rect 21940 -8416 21974 -8400
rect 20853 -8462 20869 -8428
rect 21245 -8462 21261 -8428
rect 21489 -8462 21505 -8428
rect 21881 -8462 21897 -8428
rect 20638 -8562 20672 -8500
rect 22078 -8562 22112 -8500
rect 20638 -8596 20734 -8562
rect 22016 -8596 22112 -8562
rect 20638 -8658 20672 -8596
rect 22078 -8658 22112 -8596
rect 20853 -8730 20869 -8696
rect 21245 -8730 21261 -8696
rect 21489 -8730 21505 -8696
rect 21881 -8730 21897 -8696
rect 20776 -8758 20810 -8742
rect 20776 -9542 20810 -9526
rect 21304 -8758 21338 -8742
rect 21304 -9542 21338 -9526
rect 21412 -8758 21446 -8742
rect 21412 -9542 21446 -9526
rect 21940 -8758 21974 -8742
rect 21940 -9542 21974 -9526
rect 20853 -9588 20869 -9554
rect 21245 -9588 21261 -9554
rect 21489 -9588 21505 -9554
rect 21881 -9588 21897 -9554
rect 20638 -9688 20672 -9626
rect 22078 -9688 22112 -9626
rect 20638 -9722 20734 -9688
rect 22016 -9722 22112 -9688
rect 22238 -8070 22334 -8060
rect 23616 -8060 23934 -8036
rect 23616 -8070 23712 -8060
rect 22238 -8132 22272 -8070
rect 23678 -8132 23712 -8070
rect 22453 -8204 22469 -8170
rect 22845 -8204 22861 -8170
rect 23089 -8204 23105 -8170
rect 23481 -8204 23497 -8170
rect 22376 -8232 22410 -8216
rect 22376 -8416 22410 -8400
rect 22904 -8232 22938 -8216
rect 22904 -8416 22938 -8400
rect 23012 -8232 23046 -8216
rect 23012 -8416 23046 -8400
rect 23540 -8232 23574 -8216
rect 23540 -8416 23574 -8400
rect 22453 -8462 22469 -8428
rect 22845 -8462 22861 -8428
rect 23089 -8462 23105 -8428
rect 23481 -8462 23497 -8428
rect 22238 -8562 22272 -8500
rect 23678 -8562 23712 -8500
rect 22238 -8596 22334 -8562
rect 23616 -8596 23712 -8562
rect 22238 -8658 22272 -8596
rect 23678 -8658 23712 -8596
rect 22453 -8730 22469 -8696
rect 22845 -8730 22861 -8696
rect 23089 -8730 23105 -8696
rect 23481 -8730 23497 -8696
rect 22376 -8758 22410 -8742
rect 22376 -9542 22410 -9526
rect 22904 -8758 22938 -8742
rect 22904 -9542 22938 -9526
rect 23012 -8758 23046 -8742
rect 23012 -9542 23046 -9526
rect 23540 -8758 23574 -8742
rect 23540 -9542 23574 -9526
rect 22453 -9588 22469 -9554
rect 22845 -9588 22861 -9554
rect 23089 -9588 23105 -9554
rect 23481 -9588 23497 -9554
rect 22238 -9688 22272 -9626
rect 23678 -9688 23712 -9626
rect 22238 -9722 22334 -9688
rect 23616 -9722 23712 -9688
rect 23838 -8070 23934 -8060
rect 25216 -8060 25534 -8036
rect 25216 -8070 25312 -8060
rect 23838 -8132 23872 -8070
rect 25278 -8132 25312 -8070
rect 24053 -8204 24069 -8170
rect 24445 -8204 24461 -8170
rect 24689 -8204 24705 -8170
rect 25081 -8204 25097 -8170
rect 23976 -8232 24010 -8216
rect 23976 -8416 24010 -8400
rect 24504 -8232 24538 -8216
rect 24504 -8416 24538 -8400
rect 24612 -8232 24646 -8216
rect 24612 -8416 24646 -8400
rect 25140 -8232 25174 -8216
rect 25140 -8416 25174 -8400
rect 24053 -8462 24069 -8428
rect 24445 -8462 24461 -8428
rect 24689 -8462 24705 -8428
rect 25081 -8462 25097 -8428
rect 23838 -8562 23872 -8500
rect 25278 -8562 25312 -8500
rect 23838 -8596 23934 -8562
rect 25216 -8596 25312 -8562
rect 23838 -8658 23872 -8596
rect 25278 -8658 25312 -8596
rect 24053 -8730 24069 -8696
rect 24445 -8730 24461 -8696
rect 24689 -8730 24705 -8696
rect 25081 -8730 25097 -8696
rect 23976 -8758 24010 -8742
rect 23976 -9542 24010 -9526
rect 24504 -8758 24538 -8742
rect 24504 -9542 24538 -9526
rect 24612 -8758 24646 -8742
rect 24612 -9542 24646 -9526
rect 25140 -8758 25174 -8742
rect 25140 -9542 25174 -9526
rect 24053 -9588 24069 -9554
rect 24445 -9588 24461 -9554
rect 24689 -9588 24705 -9554
rect 25081 -9588 25097 -9554
rect 23838 -9688 23872 -9626
rect 25278 -9688 25312 -9626
rect 23838 -9722 23934 -9688
rect 25216 -9722 25312 -9688
rect 25438 -8070 25534 -8060
rect 26816 -8060 27134 -8036
rect 26816 -8070 26912 -8060
rect 25438 -8132 25472 -8070
rect 26878 -8132 26912 -8070
rect 25653 -8204 25669 -8170
rect 26045 -8204 26061 -8170
rect 26289 -8204 26305 -8170
rect 26681 -8204 26697 -8170
rect 25576 -8232 25610 -8216
rect 25576 -8416 25610 -8400
rect 26104 -8232 26138 -8216
rect 26104 -8416 26138 -8400
rect 26212 -8232 26246 -8216
rect 26212 -8416 26246 -8400
rect 26740 -8232 26774 -8216
rect 26740 -8416 26774 -8400
rect 25653 -8462 25669 -8428
rect 26045 -8462 26061 -8428
rect 26289 -8462 26305 -8428
rect 26681 -8462 26697 -8428
rect 25438 -8562 25472 -8500
rect 26878 -8562 26912 -8500
rect 25438 -8596 25534 -8562
rect 26816 -8596 26912 -8562
rect 25438 -8658 25472 -8596
rect 26878 -8658 26912 -8596
rect 25653 -8730 25669 -8696
rect 26045 -8730 26061 -8696
rect 26289 -8730 26305 -8696
rect 26681 -8730 26697 -8696
rect 25576 -8758 25610 -8742
rect 25576 -9542 25610 -9526
rect 26104 -8758 26138 -8742
rect 26104 -9542 26138 -9526
rect 26212 -8758 26246 -8742
rect 26212 -9542 26246 -9526
rect 26740 -8758 26774 -8742
rect 26740 -9542 26774 -9526
rect 25653 -9588 25669 -9554
rect 26045 -9588 26061 -9554
rect 26289 -9588 26305 -9554
rect 26681 -9588 26697 -9554
rect 25438 -9688 25472 -9626
rect 26878 -9688 26912 -9626
rect 25438 -9722 25534 -9688
rect 26816 -9722 26912 -9688
rect 27038 -8070 27134 -8060
rect 28416 -8060 28734 -8036
rect 28416 -8070 28512 -8060
rect 27038 -8132 27072 -8070
rect 28478 -8132 28512 -8070
rect 27253 -8204 27269 -8170
rect 27645 -8204 27661 -8170
rect 27889 -8204 27905 -8170
rect 28281 -8204 28297 -8170
rect 27176 -8232 27210 -8216
rect 27176 -8416 27210 -8400
rect 27704 -8232 27738 -8216
rect 27704 -8416 27738 -8400
rect 27812 -8232 27846 -8216
rect 27812 -8416 27846 -8400
rect 28340 -8232 28374 -8216
rect 28340 -8416 28374 -8400
rect 27253 -8462 27269 -8428
rect 27645 -8462 27661 -8428
rect 27889 -8462 27905 -8428
rect 28281 -8462 28297 -8428
rect 27038 -8562 27072 -8500
rect 28478 -8562 28512 -8500
rect 27038 -8596 27134 -8562
rect 28416 -8596 28512 -8562
rect 27038 -8658 27072 -8596
rect 28478 -8658 28512 -8596
rect 27253 -8730 27269 -8696
rect 27645 -8730 27661 -8696
rect 27889 -8730 27905 -8696
rect 28281 -8730 28297 -8696
rect 27176 -8758 27210 -8742
rect 27176 -9542 27210 -9526
rect 27704 -8758 27738 -8742
rect 27704 -9542 27738 -9526
rect 27812 -8758 27846 -8742
rect 27812 -9542 27846 -9526
rect 28340 -8758 28374 -8742
rect 28340 -9542 28374 -9526
rect 27253 -9588 27269 -9554
rect 27645 -9588 27661 -9554
rect 27889 -9588 27905 -9554
rect 28281 -9588 28297 -9554
rect 27038 -9688 27072 -9626
rect 28478 -9688 28512 -9626
rect 27038 -9722 27134 -9688
rect 28416 -9722 28512 -9688
rect 28638 -8070 28734 -8060
rect 30016 -8060 30334 -8036
rect 30016 -8070 30112 -8060
rect 28638 -8132 28672 -8070
rect 30078 -8132 30112 -8070
rect 28853 -8204 28869 -8170
rect 29245 -8204 29261 -8170
rect 29489 -8204 29505 -8170
rect 29881 -8204 29897 -8170
rect 28776 -8232 28810 -8216
rect 28776 -8416 28810 -8400
rect 29304 -8232 29338 -8216
rect 29304 -8416 29338 -8400
rect 29412 -8232 29446 -8216
rect 29412 -8416 29446 -8400
rect 29940 -8232 29974 -8216
rect 29940 -8416 29974 -8400
rect 28853 -8462 28869 -8428
rect 29245 -8462 29261 -8428
rect 29489 -8462 29505 -8428
rect 29881 -8462 29897 -8428
rect 28638 -8562 28672 -8500
rect 30078 -8562 30112 -8500
rect 28638 -8596 28734 -8562
rect 30016 -8596 30112 -8562
rect 28638 -8658 28672 -8596
rect 30078 -8658 30112 -8596
rect 28853 -8730 28869 -8696
rect 29245 -8730 29261 -8696
rect 29489 -8730 29505 -8696
rect 29881 -8730 29897 -8696
rect 28776 -8758 28810 -8742
rect 28776 -9542 28810 -9526
rect 29304 -8758 29338 -8742
rect 29304 -9542 29338 -9526
rect 29412 -8758 29446 -8742
rect 29412 -9542 29446 -9526
rect 29940 -8758 29974 -8742
rect 29940 -9542 29974 -9526
rect 28853 -9588 28869 -9554
rect 29245 -9588 29261 -9554
rect 29489 -9588 29505 -9554
rect 29881 -9588 29897 -9554
rect 28638 -9688 28672 -9626
rect 30078 -9688 30112 -9626
rect 28638 -9722 28734 -9688
rect 30016 -9722 30112 -9688
rect 30238 -8070 30334 -8060
rect 31616 -8060 31934 -8036
rect 31616 -8070 31712 -8060
rect 30238 -8132 30272 -8070
rect 31678 -8132 31712 -8070
rect 30453 -8204 30469 -8170
rect 30845 -8204 30861 -8170
rect 31089 -8204 31105 -8170
rect 31481 -8204 31497 -8170
rect 30376 -8232 30410 -8216
rect 30376 -8416 30410 -8400
rect 30904 -8232 30938 -8216
rect 30904 -8416 30938 -8400
rect 31012 -8232 31046 -8216
rect 31012 -8416 31046 -8400
rect 31540 -8232 31574 -8216
rect 31540 -8416 31574 -8400
rect 30453 -8462 30469 -8428
rect 30845 -8462 30861 -8428
rect 31089 -8462 31105 -8428
rect 31481 -8462 31497 -8428
rect 30238 -8562 30272 -8500
rect 31678 -8562 31712 -8500
rect 30238 -8596 30334 -8562
rect 31616 -8596 31712 -8562
rect 30238 -8658 30272 -8596
rect 31678 -8658 31712 -8596
rect 30453 -8730 30469 -8696
rect 30845 -8730 30861 -8696
rect 31089 -8730 31105 -8696
rect 31481 -8730 31497 -8696
rect 30376 -8758 30410 -8742
rect 30376 -9542 30410 -9526
rect 30904 -8758 30938 -8742
rect 30904 -9542 30938 -9526
rect 31012 -8758 31046 -8742
rect 31012 -9542 31046 -9526
rect 31540 -8758 31574 -8742
rect 31540 -9542 31574 -9526
rect 30453 -9588 30469 -9554
rect 30845 -9588 30861 -9554
rect 31089 -9588 31105 -9554
rect 31481 -9588 31497 -9554
rect 30238 -9688 30272 -9626
rect 31678 -9688 31712 -9626
rect 30238 -9722 30334 -9688
rect 31616 -9722 31712 -9688
rect 31838 -8070 31934 -8060
rect 33216 -8060 33534 -8036
rect 33216 -8070 33312 -8060
rect 31838 -8132 31872 -8070
rect 33278 -8132 33312 -8070
rect 32053 -8204 32069 -8170
rect 32445 -8204 32461 -8170
rect 32689 -8204 32705 -8170
rect 33081 -8204 33097 -8170
rect 31976 -8232 32010 -8216
rect 31976 -8416 32010 -8400
rect 32504 -8232 32538 -8216
rect 32504 -8416 32538 -8400
rect 32612 -8232 32646 -8216
rect 32612 -8416 32646 -8400
rect 33140 -8232 33174 -8216
rect 33140 -8416 33174 -8400
rect 32053 -8462 32069 -8428
rect 32445 -8462 32461 -8428
rect 32689 -8462 32705 -8428
rect 33081 -8462 33097 -8428
rect 31838 -8562 31872 -8500
rect 33278 -8562 33312 -8500
rect 31838 -8596 31934 -8562
rect 33216 -8596 33312 -8562
rect 31838 -8658 31872 -8596
rect 33278 -8658 33312 -8596
rect 32053 -8730 32069 -8696
rect 32445 -8730 32461 -8696
rect 32689 -8730 32705 -8696
rect 33081 -8730 33097 -8696
rect 31976 -8758 32010 -8742
rect 31976 -9542 32010 -9526
rect 32504 -8758 32538 -8742
rect 32504 -9542 32538 -9526
rect 32612 -8758 32646 -8742
rect 32612 -9542 32646 -9526
rect 33140 -8758 33174 -8742
rect 33140 -9542 33174 -9526
rect 32053 -9588 32069 -9554
rect 32445 -9588 32461 -9554
rect 32689 -9588 32705 -9554
rect 33081 -9588 33097 -9554
rect 31838 -9688 31872 -9626
rect 33278 -9688 33312 -9626
rect 31838 -9722 31934 -9688
rect 33216 -9722 33312 -9688
rect 33438 -8070 33534 -8060
rect 34816 -8060 35134 -8036
rect 34816 -8070 34912 -8060
rect 33438 -8132 33472 -8070
rect 34878 -8132 34912 -8070
rect 33653 -8204 33669 -8170
rect 34045 -8204 34061 -8170
rect 34289 -8204 34305 -8170
rect 34681 -8204 34697 -8170
rect 33576 -8232 33610 -8216
rect 33576 -8416 33610 -8400
rect 34104 -8232 34138 -8216
rect 34104 -8416 34138 -8400
rect 34212 -8232 34246 -8216
rect 34212 -8416 34246 -8400
rect 34740 -8232 34774 -8216
rect 34740 -8416 34774 -8400
rect 33653 -8462 33669 -8428
rect 34045 -8462 34061 -8428
rect 34289 -8462 34305 -8428
rect 34681 -8462 34697 -8428
rect 33438 -8562 33472 -8500
rect 34878 -8562 34912 -8500
rect 33438 -8596 33534 -8562
rect 34816 -8596 34912 -8562
rect 33438 -8658 33472 -8596
rect 34878 -8658 34912 -8596
rect 33653 -8730 33669 -8696
rect 34045 -8730 34061 -8696
rect 34289 -8730 34305 -8696
rect 34681 -8730 34697 -8696
rect 33576 -8758 33610 -8742
rect 33576 -9542 33610 -9526
rect 34104 -8758 34138 -8742
rect 34104 -9542 34138 -9526
rect 34212 -8758 34246 -8742
rect 34212 -9542 34246 -9526
rect 34740 -8758 34774 -8742
rect 34740 -9542 34774 -9526
rect 33653 -9588 33669 -9554
rect 34045 -9588 34061 -9554
rect 34289 -9588 34305 -9554
rect 34681 -9588 34697 -9554
rect 33438 -9688 33472 -9626
rect 34878 -9688 34912 -9626
rect 33438 -9722 33534 -9688
rect 34816 -9722 34912 -9688
rect 35038 -8070 35134 -8060
rect 36416 -8070 36734 -8036
rect 38016 -8070 38112 -8036
rect 35038 -8132 35072 -8070
rect 36478 -8132 38112 -8070
rect 35253 -8204 35269 -8170
rect 35645 -8204 35661 -8170
rect 35889 -8204 35905 -8170
rect 36281 -8204 36297 -8170
rect 35176 -8232 35210 -8216
rect 35176 -8416 35210 -8400
rect 35704 -8232 35738 -8216
rect 35704 -8416 35738 -8400
rect 35812 -8232 35846 -8216
rect 35812 -8416 35846 -8400
rect 36340 -8232 36374 -8216
rect 36340 -8416 36374 -8400
rect 35253 -8462 35269 -8428
rect 35645 -8462 35661 -8428
rect 35889 -8462 35905 -8428
rect 36281 -8462 36297 -8428
rect 35038 -8562 35072 -8500
rect 36512 -8500 36638 -8132
rect 36672 -8170 38078 -8132
rect 36672 -8204 36869 -8170
rect 37245 -8204 37505 -8170
rect 37881 -8204 38078 -8170
rect 36672 -8232 38078 -8204
rect 36672 -8400 36776 -8232
rect 36810 -8400 37304 -8232
rect 37338 -8400 37412 -8232
rect 37446 -8400 37940 -8232
rect 37974 -8400 38078 -8232
rect 36672 -8428 38078 -8400
rect 36672 -8462 36869 -8428
rect 37245 -8462 37505 -8428
rect 37881 -8462 38078 -8428
rect 36672 -8500 38078 -8462
rect 36478 -8562 38112 -8500
rect 35038 -8596 35134 -8562
rect 36416 -8596 36734 -8562
rect 38016 -8596 38112 -8562
rect 35038 -8658 35072 -8596
rect 36478 -8658 38112 -8596
rect 35253 -8730 35269 -8696
rect 35645 -8730 35661 -8696
rect 35889 -8730 35905 -8696
rect 36281 -8730 36297 -8696
rect 35176 -8758 35210 -8742
rect 35176 -9542 35210 -9526
rect 35704 -8758 35738 -8742
rect 35704 -9542 35738 -9526
rect 35812 -8758 35846 -8742
rect 35812 -9542 35846 -9526
rect 36340 -8758 36374 -8742
rect 36340 -9542 36374 -9526
rect 35253 -9588 35269 -9554
rect 35645 -9588 35661 -9554
rect 35889 -9588 35905 -9554
rect 36281 -9588 36297 -9554
rect 35038 -9688 35072 -9626
rect 36512 -9626 36638 -8658
rect 36672 -8696 38078 -8658
rect 36672 -8730 36869 -8696
rect 37245 -8730 37505 -8696
rect 37881 -8730 38078 -8696
rect 36672 -8758 38078 -8730
rect 36672 -9526 36776 -8758
rect 36810 -9526 37304 -8758
rect 37338 -9526 37412 -8758
rect 37446 -9526 37940 -8758
rect 37974 -9526 38078 -8758
rect 36672 -9554 38078 -9526
rect 36672 -9588 36869 -9554
rect 37245 -9588 37505 -9554
rect 37881 -9588 38078 -9554
rect 36672 -9626 38078 -9588
rect 36478 -9688 38112 -9626
rect 35038 -9722 35134 -9688
rect 36416 -9722 36734 -9688
rect 38016 -9722 38112 -9688
rect -140 -9836 1460 -9722
rect 36500 -9836 38100 -9722
rect -162 -9870 -66 -9836
rect 1216 -9870 1534 -9836
rect 2816 -9870 2912 -9836
rect -162 -9932 1472 -9870
rect -128 -9970 1278 -9932
rect -128 -10004 69 -9970
rect 445 -10004 705 -9970
rect 1081 -10004 1278 -9970
rect -128 -10032 1278 -10004
rect -128 -10200 -24 -10032
rect 10 -10200 504 -10032
rect 538 -10200 612 -10032
rect 646 -10200 1140 -10032
rect 1174 -10200 1278 -10032
rect -128 -10228 1278 -10200
rect -128 -10262 69 -10228
rect 445 -10262 705 -10228
rect 1081 -10262 1278 -10228
rect -128 -10300 1278 -10262
rect 1312 -10300 1438 -9932
rect 2878 -9932 2912 -9870
rect 1653 -10004 1669 -9970
rect 2045 -10004 2061 -9970
rect 2289 -10004 2305 -9970
rect 2681 -10004 2697 -9970
rect 1576 -10032 1610 -10016
rect 1576 -10216 1610 -10200
rect 2104 -10032 2138 -10016
rect 2104 -10216 2138 -10200
rect 2212 -10032 2246 -10016
rect 2212 -10216 2246 -10200
rect 2740 -10032 2774 -10016
rect 2740 -10216 2774 -10200
rect 1653 -10262 1669 -10228
rect 2045 -10262 2061 -10228
rect 2289 -10262 2305 -10228
rect 2681 -10262 2697 -10228
rect -162 -10362 1472 -10300
rect 2878 -10362 2912 -10300
rect -162 -10396 -66 -10362
rect 1216 -10396 1534 -10362
rect 2816 -10396 2912 -10362
rect -162 -10458 1472 -10396
rect -128 -10496 1278 -10458
rect -128 -10530 69 -10496
rect 445 -10530 705 -10496
rect 1081 -10530 1278 -10496
rect -128 -10558 1278 -10530
rect -128 -11326 -24 -10558
rect 10 -11326 504 -10558
rect 538 -11326 612 -10558
rect 646 -11326 1140 -10558
rect 1174 -11326 1278 -10558
rect -128 -11354 1278 -11326
rect -128 -11388 69 -11354
rect 445 -11388 705 -11354
rect 1081 -11388 1278 -11354
rect -128 -11426 1278 -11388
rect 1312 -11426 1438 -10458
rect 2878 -10458 2912 -10396
rect 1653 -10530 1669 -10496
rect 2045 -10530 2061 -10496
rect 2289 -10530 2305 -10496
rect 2681 -10530 2697 -10496
rect 1576 -10558 1610 -10542
rect 1576 -11342 1610 -11326
rect 2104 -10558 2138 -10542
rect 2104 -11342 2138 -11326
rect 2212 -10558 2246 -10542
rect 2212 -11342 2246 -11326
rect 2740 -10558 2774 -10542
rect 2740 -11342 2774 -11326
rect 1653 -11388 1669 -11354
rect 2045 -11388 2061 -11354
rect 2289 -11388 2305 -11354
rect 2681 -11388 2697 -11354
rect -162 -11488 1472 -11426
rect 2878 -11488 2912 -11426
rect -162 -11522 -66 -11488
rect 1216 -11522 1534 -11488
rect 2816 -11522 2912 -11488
rect 3038 -9870 3134 -9836
rect 4416 -9870 4512 -9836
rect 3038 -9932 3072 -9870
rect 4478 -9932 4512 -9870
rect 3253 -10004 3269 -9970
rect 3645 -10004 3661 -9970
rect 3889 -10004 3905 -9970
rect 4281 -10004 4297 -9970
rect 3176 -10032 3210 -10016
rect 3176 -10216 3210 -10200
rect 3704 -10032 3738 -10016
rect 3704 -10216 3738 -10200
rect 3812 -10032 3846 -10016
rect 3812 -10216 3846 -10200
rect 4340 -10032 4374 -10016
rect 4340 -10216 4374 -10200
rect 3253 -10262 3269 -10228
rect 3645 -10262 3661 -10228
rect 3889 -10262 3905 -10228
rect 4281 -10262 4297 -10228
rect 3038 -10362 3072 -10300
rect 4478 -10362 4512 -10300
rect 3038 -10396 3134 -10362
rect 4416 -10396 4512 -10362
rect 3038 -10458 3072 -10396
rect 4478 -10458 4512 -10396
rect 3253 -10530 3269 -10496
rect 3645 -10530 3661 -10496
rect 3889 -10530 3905 -10496
rect 4281 -10530 4297 -10496
rect 3176 -10558 3210 -10542
rect 3176 -11342 3210 -11326
rect 3704 -10558 3738 -10542
rect 3704 -11342 3738 -11326
rect 3812 -10558 3846 -10542
rect 3812 -11342 3846 -11326
rect 4340 -10558 4374 -10542
rect 4340 -11342 4374 -11326
rect 3253 -11388 3269 -11354
rect 3645 -11388 3661 -11354
rect 3889 -11388 3905 -11354
rect 4281 -11388 4297 -11354
rect 3038 -11488 3072 -11426
rect 4478 -11488 4512 -11426
rect 3038 -11522 3134 -11488
rect 4416 -11522 4512 -11488
rect 4638 -9870 4734 -9836
rect 6016 -9870 6112 -9836
rect 4638 -9932 4672 -9870
rect 6078 -9932 6112 -9870
rect 4853 -10004 4869 -9970
rect 5245 -10004 5261 -9970
rect 5489 -10004 5505 -9970
rect 5881 -10004 5897 -9970
rect 4776 -10032 4810 -10016
rect 4776 -10216 4810 -10200
rect 5304 -10032 5338 -10016
rect 5304 -10216 5338 -10200
rect 5412 -10032 5446 -10016
rect 5412 -10216 5446 -10200
rect 5940 -10032 5974 -10016
rect 5940 -10216 5974 -10200
rect 4853 -10262 4869 -10228
rect 5245 -10262 5261 -10228
rect 5489 -10262 5505 -10228
rect 5881 -10262 5897 -10228
rect 4638 -10362 4672 -10300
rect 6078 -10362 6112 -10300
rect 4638 -10396 4734 -10362
rect 6016 -10396 6112 -10362
rect 4638 -10458 4672 -10396
rect 6078 -10458 6112 -10396
rect 4853 -10530 4869 -10496
rect 5245 -10530 5261 -10496
rect 5489 -10530 5505 -10496
rect 5881 -10530 5897 -10496
rect 4776 -10558 4810 -10542
rect 4776 -11342 4810 -11326
rect 5304 -10558 5338 -10542
rect 5304 -11342 5338 -11326
rect 5412 -10558 5446 -10542
rect 5412 -11342 5446 -11326
rect 5940 -10558 5974 -10542
rect 5940 -11342 5974 -11326
rect 4853 -11388 4869 -11354
rect 5245 -11388 5261 -11354
rect 5489 -11388 5505 -11354
rect 5881 -11388 5897 -11354
rect 4638 -11488 4672 -11426
rect 6078 -11488 6112 -11426
rect 4638 -11522 4734 -11488
rect 6016 -11522 6112 -11488
rect 6238 -9870 6334 -9836
rect 7616 -9870 7712 -9836
rect 6238 -9932 6272 -9870
rect 7678 -9932 7712 -9870
rect 6453 -10004 6469 -9970
rect 6845 -10004 6861 -9970
rect 7089 -10004 7105 -9970
rect 7481 -10004 7497 -9970
rect 6376 -10032 6410 -10016
rect 6376 -10216 6410 -10200
rect 6904 -10032 6938 -10016
rect 6904 -10216 6938 -10200
rect 7012 -10032 7046 -10016
rect 7012 -10216 7046 -10200
rect 7540 -10032 7574 -10016
rect 7540 -10216 7574 -10200
rect 6453 -10262 6469 -10228
rect 6845 -10262 6861 -10228
rect 7089 -10262 7105 -10228
rect 7481 -10262 7497 -10228
rect 6238 -10362 6272 -10300
rect 7678 -10362 7712 -10300
rect 6238 -10396 6334 -10362
rect 7616 -10396 7712 -10362
rect 6238 -10458 6272 -10396
rect 7678 -10458 7712 -10396
rect 6453 -10530 6469 -10496
rect 6845 -10530 6861 -10496
rect 7089 -10530 7105 -10496
rect 7481 -10530 7497 -10496
rect 6376 -10558 6410 -10542
rect 6376 -11342 6410 -11326
rect 6904 -10558 6938 -10542
rect 6904 -11342 6938 -11326
rect 7012 -10558 7046 -10542
rect 7012 -11342 7046 -11326
rect 7540 -10558 7574 -10542
rect 7540 -11342 7574 -11326
rect 6453 -11388 6469 -11354
rect 6845 -11388 6861 -11354
rect 7089 -11388 7105 -11354
rect 7481 -11388 7497 -11354
rect 6238 -11488 6272 -11426
rect 7678 -11488 7712 -11426
rect 6238 -11522 6334 -11488
rect 7616 -11522 7712 -11488
rect 7838 -9870 7934 -9836
rect 9216 -9870 9312 -9836
rect 7838 -9932 7872 -9870
rect 9278 -9932 9312 -9870
rect 8053 -10004 8069 -9970
rect 8445 -10004 8461 -9970
rect 8689 -10004 8705 -9970
rect 9081 -10004 9097 -9970
rect 7976 -10032 8010 -10016
rect 7976 -10216 8010 -10200
rect 8504 -10032 8538 -10016
rect 8504 -10216 8538 -10200
rect 8612 -10032 8646 -10016
rect 8612 -10216 8646 -10200
rect 9140 -10032 9174 -10016
rect 9140 -10216 9174 -10200
rect 8053 -10262 8069 -10228
rect 8445 -10262 8461 -10228
rect 8689 -10262 8705 -10228
rect 9081 -10262 9097 -10228
rect 7838 -10362 7872 -10300
rect 9278 -10362 9312 -10300
rect 7838 -10396 7934 -10362
rect 9216 -10396 9312 -10362
rect 7838 -10458 7872 -10396
rect 9278 -10458 9312 -10396
rect 8053 -10530 8069 -10496
rect 8445 -10530 8461 -10496
rect 8689 -10530 8705 -10496
rect 9081 -10530 9097 -10496
rect 7976 -10558 8010 -10542
rect 7976 -11342 8010 -11326
rect 8504 -10558 8538 -10542
rect 8504 -11342 8538 -11326
rect 8612 -10558 8646 -10542
rect 8612 -11342 8646 -11326
rect 9140 -10558 9174 -10542
rect 9140 -11342 9174 -11326
rect 8053 -11388 8069 -11354
rect 8445 -11388 8461 -11354
rect 8689 -11388 8705 -11354
rect 9081 -11388 9097 -11354
rect 7838 -11488 7872 -11426
rect 9278 -11488 9312 -11426
rect 7838 -11522 7934 -11488
rect 9216 -11522 9312 -11488
rect 9438 -9870 9534 -9836
rect 10816 -9870 10912 -9836
rect 9438 -9932 9472 -9870
rect 10878 -9932 10912 -9870
rect 9653 -10004 9669 -9970
rect 10045 -10004 10061 -9970
rect 10289 -10004 10305 -9970
rect 10681 -10004 10697 -9970
rect 9576 -10032 9610 -10016
rect 9576 -10216 9610 -10200
rect 10104 -10032 10138 -10016
rect 10104 -10216 10138 -10200
rect 10212 -10032 10246 -10016
rect 10212 -10216 10246 -10200
rect 10740 -10032 10774 -10016
rect 10740 -10216 10774 -10200
rect 9653 -10262 9669 -10228
rect 10045 -10262 10061 -10228
rect 10289 -10262 10305 -10228
rect 10681 -10262 10697 -10228
rect 9438 -10362 9472 -10300
rect 10878 -10362 10912 -10300
rect 9438 -10396 9534 -10362
rect 10816 -10396 10912 -10362
rect 9438 -10458 9472 -10396
rect 10878 -10458 10912 -10396
rect 9653 -10530 9669 -10496
rect 10045 -10530 10061 -10496
rect 10289 -10530 10305 -10496
rect 10681 -10530 10697 -10496
rect 9576 -10558 9610 -10542
rect 9576 -11342 9610 -11326
rect 10104 -10558 10138 -10542
rect 10104 -11342 10138 -11326
rect 10212 -10558 10246 -10542
rect 10212 -11342 10246 -11326
rect 10740 -10558 10774 -10542
rect 10740 -11342 10774 -11326
rect 9653 -11388 9669 -11354
rect 10045 -11388 10061 -11354
rect 10289 -11388 10305 -11354
rect 10681 -11388 10697 -11354
rect 9438 -11488 9472 -11426
rect 10878 -11488 10912 -11426
rect 9438 -11522 9534 -11488
rect 10816 -11522 10912 -11488
rect 11038 -9870 11134 -9836
rect 12416 -9870 12512 -9836
rect 11038 -9932 11072 -9870
rect 12478 -9932 12512 -9870
rect 11253 -10004 11269 -9970
rect 11645 -10004 11661 -9970
rect 11889 -10004 11905 -9970
rect 12281 -10004 12297 -9970
rect 11176 -10032 11210 -10016
rect 11176 -10216 11210 -10200
rect 11704 -10032 11738 -10016
rect 11704 -10216 11738 -10200
rect 11812 -10032 11846 -10016
rect 11812 -10216 11846 -10200
rect 12340 -10032 12374 -10016
rect 12340 -10216 12374 -10200
rect 11253 -10262 11269 -10228
rect 11645 -10262 11661 -10228
rect 11889 -10262 11905 -10228
rect 12281 -10262 12297 -10228
rect 11038 -10362 11072 -10300
rect 12478 -10362 12512 -10300
rect 11038 -10396 11134 -10362
rect 12416 -10396 12512 -10362
rect 11038 -10458 11072 -10396
rect 12478 -10458 12512 -10396
rect 11253 -10530 11269 -10496
rect 11645 -10530 11661 -10496
rect 11889 -10530 11905 -10496
rect 12281 -10530 12297 -10496
rect 11176 -10558 11210 -10542
rect 11176 -11342 11210 -11326
rect 11704 -10558 11738 -10542
rect 11704 -11342 11738 -11326
rect 11812 -10558 11846 -10542
rect 11812 -11342 11846 -11326
rect 12340 -10558 12374 -10542
rect 12340 -11342 12374 -11326
rect 11253 -11388 11269 -11354
rect 11645 -11388 11661 -11354
rect 11889 -11388 11905 -11354
rect 12281 -11388 12297 -11354
rect 11038 -11488 11072 -11426
rect 12478 -11488 12512 -11426
rect 11038 -11522 11134 -11488
rect 12416 -11522 12512 -11488
rect 12638 -9870 12734 -9836
rect 14016 -9870 14112 -9836
rect 12638 -9932 12672 -9870
rect 14078 -9932 14112 -9870
rect 12853 -10004 12869 -9970
rect 13245 -10004 13261 -9970
rect 13489 -10004 13505 -9970
rect 13881 -10004 13897 -9970
rect 12776 -10032 12810 -10016
rect 12776 -10216 12810 -10200
rect 13304 -10032 13338 -10016
rect 13304 -10216 13338 -10200
rect 13412 -10032 13446 -10016
rect 13412 -10216 13446 -10200
rect 13940 -10032 13974 -10016
rect 13940 -10216 13974 -10200
rect 12853 -10262 12869 -10228
rect 13245 -10262 13261 -10228
rect 13489 -10262 13505 -10228
rect 13881 -10262 13897 -10228
rect 12638 -10362 12672 -10300
rect 14078 -10362 14112 -10300
rect 12638 -10396 12734 -10362
rect 14016 -10396 14112 -10362
rect 12638 -10458 12672 -10396
rect 14078 -10458 14112 -10396
rect 12853 -10530 12869 -10496
rect 13245 -10530 13261 -10496
rect 13489 -10530 13505 -10496
rect 13881 -10530 13897 -10496
rect 12776 -10558 12810 -10542
rect 12776 -11342 12810 -11326
rect 13304 -10558 13338 -10542
rect 13304 -11342 13338 -11326
rect 13412 -10558 13446 -10542
rect 13412 -11342 13446 -11326
rect 13940 -10558 13974 -10542
rect 13940 -11342 13974 -11326
rect 12853 -11388 12869 -11354
rect 13245 -11388 13261 -11354
rect 13489 -11388 13505 -11354
rect 13881 -11388 13897 -11354
rect 12638 -11488 12672 -11426
rect 14078 -11488 14112 -11426
rect 12638 -11522 12734 -11488
rect 14016 -11522 14112 -11488
rect 14238 -9870 14334 -9836
rect 15616 -9870 15712 -9836
rect 14238 -9932 14272 -9870
rect 15678 -9932 15712 -9870
rect 14453 -10004 14469 -9970
rect 14845 -10004 14861 -9970
rect 15089 -10004 15105 -9970
rect 15481 -10004 15497 -9970
rect 14376 -10032 14410 -10016
rect 14376 -10216 14410 -10200
rect 14904 -10032 14938 -10016
rect 14904 -10216 14938 -10200
rect 15012 -10032 15046 -10016
rect 15012 -10216 15046 -10200
rect 15540 -10032 15574 -10016
rect 15540 -10216 15574 -10200
rect 14453 -10262 14469 -10228
rect 14845 -10262 14861 -10228
rect 15089 -10262 15105 -10228
rect 15481 -10262 15497 -10228
rect 14238 -10362 14272 -10300
rect 15678 -10362 15712 -10300
rect 14238 -10396 14334 -10362
rect 15616 -10396 15712 -10362
rect 14238 -10458 14272 -10396
rect 15678 -10458 15712 -10396
rect 14453 -10530 14469 -10496
rect 14845 -10530 14861 -10496
rect 15089 -10530 15105 -10496
rect 15481 -10530 15497 -10496
rect 14376 -10558 14410 -10542
rect 14376 -11342 14410 -11326
rect 14904 -10558 14938 -10542
rect 14904 -11342 14938 -11326
rect 15012 -10558 15046 -10542
rect 15012 -11342 15046 -11326
rect 15540 -10558 15574 -10542
rect 15540 -11342 15574 -11326
rect 14453 -11388 14469 -11354
rect 14845 -11388 14861 -11354
rect 15089 -11388 15105 -11354
rect 15481 -11388 15497 -11354
rect 14238 -11488 14272 -11426
rect 15678 -11488 15712 -11426
rect 14238 -11522 14334 -11488
rect 15616 -11522 15712 -11488
rect 15838 -9870 15934 -9836
rect 17216 -9870 17312 -9836
rect 15838 -9932 15872 -9870
rect 17278 -9932 17312 -9870
rect 16053 -10004 16069 -9970
rect 16445 -10004 16461 -9970
rect 16689 -10004 16705 -9970
rect 17081 -10004 17097 -9970
rect 15976 -10032 16010 -10016
rect 15976 -10216 16010 -10200
rect 16504 -10032 16538 -10016
rect 16504 -10216 16538 -10200
rect 16612 -10032 16646 -10016
rect 16612 -10216 16646 -10200
rect 17140 -10032 17174 -10016
rect 17140 -10216 17174 -10200
rect 16053 -10262 16069 -10228
rect 16445 -10262 16461 -10228
rect 16689 -10262 16705 -10228
rect 17081 -10262 17097 -10228
rect 15838 -10362 15872 -10300
rect 17278 -10362 17312 -10300
rect 15838 -10396 15934 -10362
rect 17216 -10396 17312 -10362
rect 15838 -10458 15872 -10396
rect 17278 -10458 17312 -10396
rect 16053 -10530 16069 -10496
rect 16445 -10530 16461 -10496
rect 16689 -10530 16705 -10496
rect 17081 -10530 17097 -10496
rect 15976 -10558 16010 -10542
rect 15976 -11342 16010 -11326
rect 16504 -10558 16538 -10542
rect 16504 -11342 16538 -11326
rect 16612 -10558 16646 -10542
rect 16612 -11342 16646 -11326
rect 17140 -10558 17174 -10542
rect 17140 -11342 17174 -11326
rect 16053 -11388 16069 -11354
rect 16445 -11388 16461 -11354
rect 16689 -11388 16705 -11354
rect 17081 -11388 17097 -11354
rect 15838 -11488 15872 -11426
rect 17278 -11488 17312 -11426
rect 15838 -11522 15934 -11488
rect 17216 -11522 17312 -11488
rect 17438 -9870 17534 -9836
rect 18816 -9870 18912 -9836
rect 17438 -9932 17472 -9870
rect 18878 -9932 18912 -9870
rect 17653 -10004 17669 -9970
rect 18045 -10004 18061 -9970
rect 18289 -10004 18305 -9970
rect 18681 -10004 18697 -9970
rect 17576 -10032 17610 -10016
rect 17576 -10216 17610 -10200
rect 18104 -10032 18138 -10016
rect 18104 -10216 18138 -10200
rect 18212 -10032 18246 -10016
rect 18212 -10216 18246 -10200
rect 18740 -10032 18774 -10016
rect 18740 -10216 18774 -10200
rect 17653 -10262 17669 -10228
rect 18045 -10262 18061 -10228
rect 18289 -10262 18305 -10228
rect 18681 -10262 18697 -10228
rect 17438 -10362 17472 -10300
rect 18878 -10362 18912 -10300
rect 17438 -10396 17534 -10362
rect 18816 -10396 18912 -10362
rect 17438 -10458 17472 -10396
rect 18878 -10458 18912 -10396
rect 17653 -10530 17669 -10496
rect 18045 -10530 18061 -10496
rect 18289 -10530 18305 -10496
rect 18681 -10530 18697 -10496
rect 17576 -10558 17610 -10542
rect 17576 -11342 17610 -11326
rect 18104 -10558 18138 -10542
rect 18104 -11342 18138 -11326
rect 18212 -10558 18246 -10542
rect 18212 -11342 18246 -11326
rect 18740 -10558 18774 -10542
rect 18740 -11342 18774 -11326
rect 17653 -11388 17669 -11354
rect 18045 -11388 18061 -11354
rect 18289 -11388 18305 -11354
rect 18681 -11388 18697 -11354
rect 17438 -11488 17472 -11426
rect 18878 -11488 18912 -11426
rect 17438 -11522 17534 -11488
rect 18816 -11522 18912 -11488
rect 19038 -9870 19134 -9836
rect 20416 -9870 20512 -9836
rect 19038 -9932 19072 -9870
rect 20478 -9932 20512 -9870
rect 19253 -10004 19269 -9970
rect 19645 -10004 19661 -9970
rect 19889 -10004 19905 -9970
rect 20281 -10004 20297 -9970
rect 19176 -10032 19210 -10016
rect 19176 -10216 19210 -10200
rect 19704 -10032 19738 -10016
rect 19704 -10216 19738 -10200
rect 19812 -10032 19846 -10016
rect 19812 -10216 19846 -10200
rect 20340 -10032 20374 -10016
rect 20340 -10216 20374 -10200
rect 19253 -10262 19269 -10228
rect 19645 -10262 19661 -10228
rect 19889 -10262 19905 -10228
rect 20281 -10262 20297 -10228
rect 19038 -10362 19072 -10300
rect 20478 -10362 20512 -10300
rect 19038 -10396 19134 -10362
rect 20416 -10396 20512 -10362
rect 19038 -10458 19072 -10396
rect 20478 -10458 20512 -10396
rect 19253 -10530 19269 -10496
rect 19645 -10530 19661 -10496
rect 19889 -10530 19905 -10496
rect 20281 -10530 20297 -10496
rect 19176 -10558 19210 -10542
rect 19176 -11342 19210 -11326
rect 19704 -10558 19738 -10542
rect 19704 -11342 19738 -11326
rect 19812 -10558 19846 -10542
rect 19812 -11342 19846 -11326
rect 20340 -10558 20374 -10542
rect 20340 -11342 20374 -11326
rect 19253 -11388 19269 -11354
rect 19645 -11388 19661 -11354
rect 19889 -11388 19905 -11354
rect 20281 -11388 20297 -11354
rect 19038 -11488 19072 -11426
rect 20478 -11488 20512 -11426
rect 19038 -11522 19134 -11488
rect 20416 -11522 20512 -11488
rect 20638 -9870 20734 -9836
rect 22016 -9870 22112 -9836
rect 20638 -9932 20672 -9870
rect 22078 -9932 22112 -9870
rect 20853 -10004 20869 -9970
rect 21245 -10004 21261 -9970
rect 21489 -10004 21505 -9970
rect 21881 -10004 21897 -9970
rect 20776 -10032 20810 -10016
rect 20776 -10216 20810 -10200
rect 21304 -10032 21338 -10016
rect 21304 -10216 21338 -10200
rect 21412 -10032 21446 -10016
rect 21412 -10216 21446 -10200
rect 21940 -10032 21974 -10016
rect 21940 -10216 21974 -10200
rect 20853 -10262 20869 -10228
rect 21245 -10262 21261 -10228
rect 21489 -10262 21505 -10228
rect 21881 -10262 21897 -10228
rect 20638 -10362 20672 -10300
rect 22078 -10362 22112 -10300
rect 20638 -10396 20734 -10362
rect 22016 -10396 22112 -10362
rect 20638 -10458 20672 -10396
rect 22078 -10458 22112 -10396
rect 20853 -10530 20869 -10496
rect 21245 -10530 21261 -10496
rect 21489 -10530 21505 -10496
rect 21881 -10530 21897 -10496
rect 20776 -10558 20810 -10542
rect 20776 -11342 20810 -11326
rect 21304 -10558 21338 -10542
rect 21304 -11342 21338 -11326
rect 21412 -10558 21446 -10542
rect 21412 -11342 21446 -11326
rect 21940 -10558 21974 -10542
rect 21940 -11342 21974 -11326
rect 20853 -11388 20869 -11354
rect 21245 -11388 21261 -11354
rect 21489 -11388 21505 -11354
rect 21881 -11388 21897 -11354
rect 20638 -11488 20672 -11426
rect 22078 -11488 22112 -11426
rect 20638 -11522 20734 -11488
rect 22016 -11522 22112 -11488
rect 22238 -9870 22334 -9836
rect 23616 -9870 23712 -9836
rect 22238 -9932 22272 -9870
rect 23678 -9932 23712 -9870
rect 22453 -10004 22469 -9970
rect 22845 -10004 22861 -9970
rect 23089 -10004 23105 -9970
rect 23481 -10004 23497 -9970
rect 22376 -10032 22410 -10016
rect 22376 -10216 22410 -10200
rect 22904 -10032 22938 -10016
rect 22904 -10216 22938 -10200
rect 23012 -10032 23046 -10016
rect 23012 -10216 23046 -10200
rect 23540 -10032 23574 -10016
rect 23540 -10216 23574 -10200
rect 22453 -10262 22469 -10228
rect 22845 -10262 22861 -10228
rect 23089 -10262 23105 -10228
rect 23481 -10262 23497 -10228
rect 22238 -10362 22272 -10300
rect 23678 -10362 23712 -10300
rect 22238 -10396 22334 -10362
rect 23616 -10396 23712 -10362
rect 22238 -10458 22272 -10396
rect 23678 -10458 23712 -10396
rect 22453 -10530 22469 -10496
rect 22845 -10530 22861 -10496
rect 23089 -10530 23105 -10496
rect 23481 -10530 23497 -10496
rect 22376 -10558 22410 -10542
rect 22376 -11342 22410 -11326
rect 22904 -10558 22938 -10542
rect 22904 -11342 22938 -11326
rect 23012 -10558 23046 -10542
rect 23012 -11342 23046 -11326
rect 23540 -10558 23574 -10542
rect 23540 -11342 23574 -11326
rect 22453 -11388 22469 -11354
rect 22845 -11388 22861 -11354
rect 23089 -11388 23105 -11354
rect 23481 -11388 23497 -11354
rect 22238 -11488 22272 -11426
rect 23678 -11488 23712 -11426
rect 22238 -11522 22334 -11488
rect 23616 -11522 23712 -11488
rect 23838 -9870 23934 -9836
rect 25216 -9870 25312 -9836
rect 23838 -9932 23872 -9870
rect 25278 -9932 25312 -9870
rect 24053 -10004 24069 -9970
rect 24445 -10004 24461 -9970
rect 24689 -10004 24705 -9970
rect 25081 -10004 25097 -9970
rect 23976 -10032 24010 -10016
rect 23976 -10216 24010 -10200
rect 24504 -10032 24538 -10016
rect 24504 -10216 24538 -10200
rect 24612 -10032 24646 -10016
rect 24612 -10216 24646 -10200
rect 25140 -10032 25174 -10016
rect 25140 -10216 25174 -10200
rect 24053 -10262 24069 -10228
rect 24445 -10262 24461 -10228
rect 24689 -10262 24705 -10228
rect 25081 -10262 25097 -10228
rect 23838 -10362 23872 -10300
rect 25278 -10362 25312 -10300
rect 23838 -10396 23934 -10362
rect 25216 -10396 25312 -10362
rect 23838 -10458 23872 -10396
rect 25278 -10458 25312 -10396
rect 24053 -10530 24069 -10496
rect 24445 -10530 24461 -10496
rect 24689 -10530 24705 -10496
rect 25081 -10530 25097 -10496
rect 23976 -10558 24010 -10542
rect 23976 -11342 24010 -11326
rect 24504 -10558 24538 -10542
rect 24504 -11342 24538 -11326
rect 24612 -10558 24646 -10542
rect 24612 -11342 24646 -11326
rect 25140 -10558 25174 -10542
rect 25140 -11342 25174 -11326
rect 24053 -11388 24069 -11354
rect 24445 -11388 24461 -11354
rect 24689 -11388 24705 -11354
rect 25081 -11388 25097 -11354
rect 23838 -11488 23872 -11426
rect 25278 -11488 25312 -11426
rect 23838 -11522 23934 -11488
rect 25216 -11522 25312 -11488
rect 25438 -9870 25534 -9836
rect 26816 -9870 26912 -9836
rect 25438 -9932 25472 -9870
rect 26878 -9932 26912 -9870
rect 25653 -10004 25669 -9970
rect 26045 -10004 26061 -9970
rect 26289 -10004 26305 -9970
rect 26681 -10004 26697 -9970
rect 25576 -10032 25610 -10016
rect 25576 -10216 25610 -10200
rect 26104 -10032 26138 -10016
rect 26104 -10216 26138 -10200
rect 26212 -10032 26246 -10016
rect 26212 -10216 26246 -10200
rect 26740 -10032 26774 -10016
rect 26740 -10216 26774 -10200
rect 25653 -10262 25669 -10228
rect 26045 -10262 26061 -10228
rect 26289 -10262 26305 -10228
rect 26681 -10262 26697 -10228
rect 25438 -10362 25472 -10300
rect 26878 -10362 26912 -10300
rect 25438 -10396 25534 -10362
rect 26816 -10396 26912 -10362
rect 25438 -10458 25472 -10396
rect 26878 -10458 26912 -10396
rect 25653 -10530 25669 -10496
rect 26045 -10530 26061 -10496
rect 26289 -10530 26305 -10496
rect 26681 -10530 26697 -10496
rect 25576 -10558 25610 -10542
rect 25576 -11342 25610 -11326
rect 26104 -10558 26138 -10542
rect 26104 -11342 26138 -11326
rect 26212 -10558 26246 -10542
rect 26212 -11342 26246 -11326
rect 26740 -10558 26774 -10542
rect 26740 -11342 26774 -11326
rect 25653 -11388 25669 -11354
rect 26045 -11388 26061 -11354
rect 26289 -11388 26305 -11354
rect 26681 -11388 26697 -11354
rect 25438 -11488 25472 -11426
rect 26878 -11488 26912 -11426
rect 25438 -11522 25534 -11488
rect 26816 -11522 26912 -11488
rect 27038 -9870 27134 -9836
rect 28416 -9870 28512 -9836
rect 27038 -9932 27072 -9870
rect 28478 -9932 28512 -9870
rect 27253 -10004 27269 -9970
rect 27645 -10004 27661 -9970
rect 27889 -10004 27905 -9970
rect 28281 -10004 28297 -9970
rect 27176 -10032 27210 -10016
rect 27176 -10216 27210 -10200
rect 27704 -10032 27738 -10016
rect 27704 -10216 27738 -10200
rect 27812 -10032 27846 -10016
rect 27812 -10216 27846 -10200
rect 28340 -10032 28374 -10016
rect 28340 -10216 28374 -10200
rect 27253 -10262 27269 -10228
rect 27645 -10262 27661 -10228
rect 27889 -10262 27905 -10228
rect 28281 -10262 28297 -10228
rect 27038 -10362 27072 -10300
rect 28478 -10362 28512 -10300
rect 27038 -10396 27134 -10362
rect 28416 -10396 28512 -10362
rect 27038 -10458 27072 -10396
rect 28478 -10458 28512 -10396
rect 27253 -10530 27269 -10496
rect 27645 -10530 27661 -10496
rect 27889 -10530 27905 -10496
rect 28281 -10530 28297 -10496
rect 27176 -10558 27210 -10542
rect 27176 -11342 27210 -11326
rect 27704 -10558 27738 -10542
rect 27704 -11342 27738 -11326
rect 27812 -10558 27846 -10542
rect 27812 -11342 27846 -11326
rect 28340 -10558 28374 -10542
rect 28340 -11342 28374 -11326
rect 27253 -11388 27269 -11354
rect 27645 -11388 27661 -11354
rect 27889 -11388 27905 -11354
rect 28281 -11388 28297 -11354
rect 27038 -11488 27072 -11426
rect 28478 -11488 28512 -11426
rect 27038 -11522 27134 -11488
rect 28416 -11522 28512 -11488
rect 28638 -9870 28734 -9836
rect 30016 -9870 30112 -9836
rect 28638 -9932 28672 -9870
rect 30078 -9932 30112 -9870
rect 28853 -10004 28869 -9970
rect 29245 -10004 29261 -9970
rect 29489 -10004 29505 -9970
rect 29881 -10004 29897 -9970
rect 28776 -10032 28810 -10016
rect 28776 -10216 28810 -10200
rect 29304 -10032 29338 -10016
rect 29304 -10216 29338 -10200
rect 29412 -10032 29446 -10016
rect 29412 -10216 29446 -10200
rect 29940 -10032 29974 -10016
rect 29940 -10216 29974 -10200
rect 28853 -10262 28869 -10228
rect 29245 -10262 29261 -10228
rect 29489 -10262 29505 -10228
rect 29881 -10262 29897 -10228
rect 28638 -10362 28672 -10300
rect 30078 -10362 30112 -10300
rect 28638 -10396 28734 -10362
rect 30016 -10396 30112 -10362
rect 28638 -10458 28672 -10396
rect 30078 -10458 30112 -10396
rect 28853 -10530 28869 -10496
rect 29245 -10530 29261 -10496
rect 29489 -10530 29505 -10496
rect 29881 -10530 29897 -10496
rect 28776 -10558 28810 -10542
rect 28776 -11342 28810 -11326
rect 29304 -10558 29338 -10542
rect 29304 -11342 29338 -11326
rect 29412 -10558 29446 -10542
rect 29412 -11342 29446 -11326
rect 29940 -10558 29974 -10542
rect 29940 -11342 29974 -11326
rect 28853 -11388 28869 -11354
rect 29245 -11388 29261 -11354
rect 29489 -11388 29505 -11354
rect 29881 -11388 29897 -11354
rect 28638 -11488 28672 -11426
rect 30078 -11488 30112 -11426
rect 28638 -11522 28734 -11488
rect 30016 -11522 30112 -11488
rect 30238 -9870 30334 -9836
rect 31616 -9870 31712 -9836
rect 30238 -9932 30272 -9870
rect 31678 -9932 31712 -9870
rect 30453 -10004 30469 -9970
rect 30845 -10004 30861 -9970
rect 31089 -10004 31105 -9970
rect 31481 -10004 31497 -9970
rect 30376 -10032 30410 -10016
rect 30376 -10216 30410 -10200
rect 30904 -10032 30938 -10016
rect 30904 -10216 30938 -10200
rect 31012 -10032 31046 -10016
rect 31012 -10216 31046 -10200
rect 31540 -10032 31574 -10016
rect 31540 -10216 31574 -10200
rect 30453 -10262 30469 -10228
rect 30845 -10262 30861 -10228
rect 31089 -10262 31105 -10228
rect 31481 -10262 31497 -10228
rect 30238 -10362 30272 -10300
rect 31678 -10362 31712 -10300
rect 30238 -10396 30334 -10362
rect 31616 -10396 31712 -10362
rect 30238 -10458 30272 -10396
rect 31678 -10458 31712 -10396
rect 30453 -10530 30469 -10496
rect 30845 -10530 30861 -10496
rect 31089 -10530 31105 -10496
rect 31481 -10530 31497 -10496
rect 30376 -10558 30410 -10542
rect 30376 -11342 30410 -11326
rect 30904 -10558 30938 -10542
rect 30904 -11342 30938 -11326
rect 31012 -10558 31046 -10542
rect 31012 -11342 31046 -11326
rect 31540 -10558 31574 -10542
rect 31540 -11342 31574 -11326
rect 30453 -11388 30469 -11354
rect 30845 -11388 30861 -11354
rect 31089 -11388 31105 -11354
rect 31481 -11388 31497 -11354
rect 30238 -11488 30272 -11426
rect 31678 -11488 31712 -11426
rect 30238 -11522 30334 -11488
rect 31616 -11522 31712 -11488
rect 31838 -9870 31934 -9836
rect 33216 -9870 33312 -9836
rect 31838 -9932 31872 -9870
rect 33278 -9932 33312 -9870
rect 32053 -10004 32069 -9970
rect 32445 -10004 32461 -9970
rect 32689 -10004 32705 -9970
rect 33081 -10004 33097 -9970
rect 31976 -10032 32010 -10016
rect 31976 -10216 32010 -10200
rect 32504 -10032 32538 -10016
rect 32504 -10216 32538 -10200
rect 32612 -10032 32646 -10016
rect 32612 -10216 32646 -10200
rect 33140 -10032 33174 -10016
rect 33140 -10216 33174 -10200
rect 32053 -10262 32069 -10228
rect 32445 -10262 32461 -10228
rect 32689 -10262 32705 -10228
rect 33081 -10262 33097 -10228
rect 31838 -10362 31872 -10300
rect 33278 -10362 33312 -10300
rect 31838 -10396 31934 -10362
rect 33216 -10396 33312 -10362
rect 31838 -10458 31872 -10396
rect 33278 -10458 33312 -10396
rect 32053 -10530 32069 -10496
rect 32445 -10530 32461 -10496
rect 32689 -10530 32705 -10496
rect 33081 -10530 33097 -10496
rect 31976 -10558 32010 -10542
rect 31976 -11342 32010 -11326
rect 32504 -10558 32538 -10542
rect 32504 -11342 32538 -11326
rect 32612 -10558 32646 -10542
rect 32612 -11342 32646 -11326
rect 33140 -10558 33174 -10542
rect 33140 -11342 33174 -11326
rect 32053 -11388 32069 -11354
rect 32445 -11388 32461 -11354
rect 32689 -11388 32705 -11354
rect 33081 -11388 33097 -11354
rect 31838 -11488 31872 -11426
rect 33278 -11488 33312 -11426
rect 31838 -11522 31934 -11488
rect 33216 -11522 33312 -11488
rect 33438 -9870 33534 -9836
rect 34816 -9870 34912 -9836
rect 33438 -9932 33472 -9870
rect 34878 -9932 34912 -9870
rect 33653 -10004 33669 -9970
rect 34045 -10004 34061 -9970
rect 34289 -10004 34305 -9970
rect 34681 -10004 34697 -9970
rect 33576 -10032 33610 -10016
rect 33576 -10216 33610 -10200
rect 34104 -10032 34138 -10016
rect 34104 -10216 34138 -10200
rect 34212 -10032 34246 -10016
rect 34212 -10216 34246 -10200
rect 34740 -10032 34774 -10016
rect 34740 -10216 34774 -10200
rect 33653 -10262 33669 -10228
rect 34045 -10262 34061 -10228
rect 34289 -10262 34305 -10228
rect 34681 -10262 34697 -10228
rect 33438 -10362 33472 -10300
rect 34878 -10362 34912 -10300
rect 33438 -10396 33534 -10362
rect 34816 -10396 34912 -10362
rect 33438 -10458 33472 -10396
rect 34878 -10458 34912 -10396
rect 33653 -10530 33669 -10496
rect 34045 -10530 34061 -10496
rect 34289 -10530 34305 -10496
rect 34681 -10530 34697 -10496
rect 33576 -10558 33610 -10542
rect 33576 -11342 33610 -11326
rect 34104 -10558 34138 -10542
rect 34104 -11342 34138 -11326
rect 34212 -10558 34246 -10542
rect 34212 -11342 34246 -11326
rect 34740 -10558 34774 -10542
rect 34740 -11342 34774 -11326
rect 33653 -11388 33669 -11354
rect 34045 -11388 34061 -11354
rect 34289 -11388 34305 -11354
rect 34681 -11388 34697 -11354
rect 33438 -11488 33472 -11426
rect 34878 -11488 34912 -11426
rect 33438 -11522 33534 -11488
rect 34816 -11522 34912 -11488
rect 35038 -9870 35134 -9836
rect 36416 -9870 36734 -9836
rect 38016 -9870 38112 -9836
rect 35038 -9932 35072 -9870
rect 36478 -9932 38112 -9870
rect 35253 -10004 35269 -9970
rect 35645 -10004 35661 -9970
rect 35889 -10004 35905 -9970
rect 36281 -10004 36297 -9970
rect 35176 -10032 35210 -10016
rect 35176 -10216 35210 -10200
rect 35704 -10032 35738 -10016
rect 35704 -10216 35738 -10200
rect 35812 -10032 35846 -10016
rect 35812 -10216 35846 -10200
rect 36340 -10032 36374 -10016
rect 36340 -10216 36374 -10200
rect 35253 -10262 35269 -10228
rect 35645 -10262 35661 -10228
rect 35889 -10262 35905 -10228
rect 36281 -10262 36297 -10228
rect 35038 -10362 35072 -10300
rect 36512 -10300 36638 -9932
rect 36672 -9970 38078 -9932
rect 36672 -10004 36869 -9970
rect 37245 -10004 37505 -9970
rect 37881 -10004 38078 -9970
rect 36672 -10032 38078 -10004
rect 36672 -10200 36776 -10032
rect 36810 -10200 37304 -10032
rect 37338 -10200 37412 -10032
rect 37446 -10200 37940 -10032
rect 37974 -10200 38078 -10032
rect 36672 -10228 38078 -10200
rect 36672 -10262 36869 -10228
rect 37245 -10262 37505 -10228
rect 37881 -10262 38078 -10228
rect 36672 -10300 38078 -10262
rect 36478 -10362 38112 -10300
rect 35038 -10396 35134 -10362
rect 36416 -10396 36734 -10362
rect 38016 -10396 38112 -10362
rect 35038 -10458 35072 -10396
rect 36478 -10458 38112 -10396
rect 35253 -10530 35269 -10496
rect 35645 -10530 35661 -10496
rect 35889 -10530 35905 -10496
rect 36281 -10530 36297 -10496
rect 35176 -10558 35210 -10542
rect 35176 -11342 35210 -11326
rect 35704 -10558 35738 -10542
rect 35704 -11342 35738 -11326
rect 35812 -10558 35846 -10542
rect 35812 -11342 35846 -11326
rect 36340 -10558 36374 -10542
rect 36340 -11342 36374 -11326
rect 35253 -11388 35269 -11354
rect 35645 -11388 35661 -11354
rect 35889 -11388 35905 -11354
rect 36281 -11388 36297 -11354
rect 35038 -11488 35072 -11426
rect 36512 -11426 36638 -10458
rect 36672 -10496 38078 -10458
rect 36672 -10530 36869 -10496
rect 37245 -10530 37505 -10496
rect 37881 -10530 38078 -10496
rect 36672 -10558 38078 -10530
rect 36672 -11326 36776 -10558
rect 36810 -11326 37304 -10558
rect 37338 -11326 37412 -10558
rect 37446 -11326 37940 -10558
rect 37974 -11326 38078 -10558
rect 36672 -11354 38078 -11326
rect 36672 -11388 36869 -11354
rect 37245 -11388 37505 -11354
rect 37881 -11388 38078 -11354
rect 36672 -11426 38078 -11388
rect 36478 -11488 38112 -11426
rect 35038 -11522 35134 -11488
rect 36416 -11522 36734 -11488
rect 38016 -11522 38112 -11488
rect -140 -11636 1460 -11522
rect 36500 -11636 38100 -11522
rect -162 -11670 -66 -11636
rect 1216 -11670 1534 -11636
rect 2816 -11670 2912 -11636
rect -162 -11732 1472 -11670
rect -128 -11770 1278 -11732
rect -128 -11804 69 -11770
rect 445 -11804 705 -11770
rect 1081 -11804 1278 -11770
rect -128 -11832 1278 -11804
rect -128 -12000 -24 -11832
rect 10 -12000 504 -11832
rect 538 -12000 612 -11832
rect 646 -12000 1140 -11832
rect 1174 -12000 1278 -11832
rect -128 -12028 1278 -12000
rect -128 -12062 69 -12028
rect 445 -12062 705 -12028
rect 1081 -12062 1278 -12028
rect -128 -12100 1278 -12062
rect 1312 -12100 1438 -11732
rect 2878 -11732 2912 -11670
rect 1653 -11804 1669 -11770
rect 2045 -11804 2061 -11770
rect 2289 -11804 2305 -11770
rect 2681 -11804 2697 -11770
rect 1576 -11832 1610 -11816
rect 1576 -12016 1610 -12000
rect 2104 -11832 2138 -11816
rect 2104 -12016 2138 -12000
rect 2212 -11832 2246 -11816
rect 2212 -12016 2246 -12000
rect 2740 -11832 2774 -11816
rect 2740 -12016 2774 -12000
rect 1653 -12062 1669 -12028
rect 2045 -12062 2061 -12028
rect 2289 -12062 2305 -12028
rect 2681 -12062 2697 -12028
rect -162 -12162 1472 -12100
rect 2878 -12162 2912 -12100
rect -162 -12196 -66 -12162
rect 1216 -12196 1534 -12162
rect 2816 -12196 2912 -12162
rect -162 -12258 1472 -12196
rect -128 -12296 1278 -12258
rect -128 -12330 69 -12296
rect 445 -12330 705 -12296
rect 1081 -12330 1278 -12296
rect -128 -12358 1278 -12330
rect -128 -13126 -24 -12358
rect 10 -13126 504 -12358
rect 538 -13126 612 -12358
rect 646 -13126 1140 -12358
rect 1174 -13126 1278 -12358
rect -128 -13154 1278 -13126
rect -128 -13188 69 -13154
rect 445 -13188 705 -13154
rect 1081 -13188 1278 -13154
rect -128 -13226 1278 -13188
rect 1312 -13226 1438 -12258
rect 2878 -12258 2912 -12196
rect 1653 -12330 1669 -12296
rect 2045 -12330 2061 -12296
rect 2289 -12330 2305 -12296
rect 2681 -12330 2697 -12296
rect 1576 -12358 1610 -12342
rect 1576 -13142 1610 -13126
rect 2104 -12358 2138 -12342
rect 2104 -13142 2138 -13126
rect 2212 -12358 2246 -12342
rect 2212 -13142 2246 -13126
rect 2740 -12358 2774 -12342
rect 2740 -13142 2774 -13126
rect 1653 -13188 1669 -13154
rect 2045 -13188 2061 -13154
rect 2289 -13188 2305 -13154
rect 2681 -13188 2697 -13154
rect -162 -13288 1472 -13226
rect 2878 -13288 2912 -13226
rect -162 -13322 -66 -13288
rect 1216 -13322 1534 -13288
rect 2816 -13322 2912 -13288
rect 3038 -11670 3134 -11636
rect 4416 -11670 4512 -11636
rect 3038 -11732 3072 -11670
rect 4478 -11732 4512 -11670
rect 3253 -11804 3269 -11770
rect 3645 -11804 3661 -11770
rect 3889 -11804 3905 -11770
rect 4281 -11804 4297 -11770
rect 3176 -11832 3210 -11816
rect 3176 -12016 3210 -12000
rect 3704 -11832 3738 -11816
rect 3704 -12016 3738 -12000
rect 3812 -11832 3846 -11816
rect 3812 -12016 3846 -12000
rect 4340 -11832 4374 -11816
rect 4340 -12016 4374 -12000
rect 3253 -12062 3269 -12028
rect 3645 -12062 3661 -12028
rect 3889 -12062 3905 -12028
rect 4281 -12062 4297 -12028
rect 3038 -12162 3072 -12100
rect 4478 -12162 4512 -12100
rect 3038 -12196 3134 -12162
rect 4416 -12196 4512 -12162
rect 3038 -12258 3072 -12196
rect 4478 -12258 4512 -12196
rect 3253 -12330 3269 -12296
rect 3645 -12330 3661 -12296
rect 3889 -12330 3905 -12296
rect 4281 -12330 4297 -12296
rect 3176 -12358 3210 -12342
rect 3176 -13142 3210 -13126
rect 3704 -12358 3738 -12342
rect 3704 -13142 3738 -13126
rect 3812 -12358 3846 -12342
rect 3812 -13142 3846 -13126
rect 4340 -12358 4374 -12342
rect 4340 -13142 4374 -13126
rect 3253 -13188 3269 -13154
rect 3645 -13188 3661 -13154
rect 3889 -13188 3905 -13154
rect 4281 -13188 4297 -13154
rect 3038 -13288 3072 -13226
rect 4478 -13288 4512 -13226
rect 3038 -13322 3134 -13288
rect 4416 -13322 4512 -13288
rect 4638 -11670 4734 -11636
rect 6016 -11670 6112 -11636
rect 4638 -11732 4672 -11670
rect 6078 -11732 6112 -11670
rect 4853 -11804 4869 -11770
rect 5245 -11804 5261 -11770
rect 5489 -11804 5505 -11770
rect 5881 -11804 5897 -11770
rect 4776 -11832 4810 -11816
rect 4776 -12016 4810 -12000
rect 5304 -11832 5338 -11816
rect 5304 -12016 5338 -12000
rect 5412 -11832 5446 -11816
rect 5412 -12016 5446 -12000
rect 5940 -11832 5974 -11816
rect 5940 -12016 5974 -12000
rect 4853 -12062 4869 -12028
rect 5245 -12062 5261 -12028
rect 5489 -12062 5505 -12028
rect 5881 -12062 5897 -12028
rect 4638 -12162 4672 -12100
rect 6078 -12162 6112 -12100
rect 4638 -12196 4734 -12162
rect 6016 -12196 6112 -12162
rect 4638 -12258 4672 -12196
rect 6078 -12258 6112 -12196
rect 4853 -12330 4869 -12296
rect 5245 -12330 5261 -12296
rect 5489 -12330 5505 -12296
rect 5881 -12330 5897 -12296
rect 4776 -12358 4810 -12342
rect 4776 -13142 4810 -13126
rect 5304 -12358 5338 -12342
rect 5304 -13142 5338 -13126
rect 5412 -12358 5446 -12342
rect 5412 -13142 5446 -13126
rect 5940 -12358 5974 -12342
rect 5940 -13142 5974 -13126
rect 4853 -13188 4869 -13154
rect 5245 -13188 5261 -13154
rect 5489 -13188 5505 -13154
rect 5881 -13188 5897 -13154
rect 4638 -13288 4672 -13226
rect 6078 -13288 6112 -13226
rect 4638 -13322 4734 -13288
rect 6016 -13322 6112 -13288
rect 6238 -11670 6334 -11636
rect 7616 -11670 7712 -11636
rect 6238 -11732 6272 -11670
rect 7678 -11732 7712 -11670
rect 6453 -11804 6469 -11770
rect 6845 -11804 6861 -11770
rect 7089 -11804 7105 -11770
rect 7481 -11804 7497 -11770
rect 6376 -11832 6410 -11816
rect 6376 -12016 6410 -12000
rect 6904 -11832 6938 -11816
rect 6904 -12016 6938 -12000
rect 7012 -11832 7046 -11816
rect 7012 -12016 7046 -12000
rect 7540 -11832 7574 -11816
rect 7540 -12016 7574 -12000
rect 6453 -12062 6469 -12028
rect 6845 -12062 6861 -12028
rect 7089 -12062 7105 -12028
rect 7481 -12062 7497 -12028
rect 6238 -12162 6272 -12100
rect 7678 -12162 7712 -12100
rect 6238 -12196 6334 -12162
rect 7616 -12196 7712 -12162
rect 6238 -12258 6272 -12196
rect 7678 -12258 7712 -12196
rect 6453 -12330 6469 -12296
rect 6845 -12330 6861 -12296
rect 7089 -12330 7105 -12296
rect 7481 -12330 7497 -12296
rect 6376 -12358 6410 -12342
rect 6376 -13142 6410 -13126
rect 6904 -12358 6938 -12342
rect 6904 -13142 6938 -13126
rect 7012 -12358 7046 -12342
rect 7012 -13142 7046 -13126
rect 7540 -12358 7574 -12342
rect 7540 -13142 7574 -13126
rect 6453 -13188 6469 -13154
rect 6845 -13188 6861 -13154
rect 7089 -13188 7105 -13154
rect 7481 -13188 7497 -13154
rect 6238 -13288 6272 -13226
rect 7678 -13288 7712 -13226
rect 6238 -13322 6334 -13288
rect 7616 -13322 7712 -13288
rect 7838 -11670 7934 -11636
rect 9216 -11670 9312 -11636
rect 7838 -11732 7872 -11670
rect 9278 -11732 9312 -11670
rect 8053 -11804 8069 -11770
rect 8445 -11804 8461 -11770
rect 8689 -11804 8705 -11770
rect 9081 -11804 9097 -11770
rect 7976 -11832 8010 -11816
rect 7976 -12016 8010 -12000
rect 8504 -11832 8538 -11816
rect 8504 -12016 8538 -12000
rect 8612 -11832 8646 -11816
rect 8612 -12016 8646 -12000
rect 9140 -11832 9174 -11816
rect 9140 -12016 9174 -12000
rect 8053 -12062 8069 -12028
rect 8445 -12062 8461 -12028
rect 8689 -12062 8705 -12028
rect 9081 -12062 9097 -12028
rect 7838 -12162 7872 -12100
rect 9278 -12162 9312 -12100
rect 7838 -12196 7934 -12162
rect 9216 -12196 9312 -12162
rect 7838 -12258 7872 -12196
rect 9278 -12258 9312 -12196
rect 8053 -12330 8069 -12296
rect 8445 -12330 8461 -12296
rect 8689 -12330 8705 -12296
rect 9081 -12330 9097 -12296
rect 7976 -12358 8010 -12342
rect 7976 -13142 8010 -13126
rect 8504 -12358 8538 -12342
rect 8504 -13142 8538 -13126
rect 8612 -12358 8646 -12342
rect 8612 -13142 8646 -13126
rect 9140 -12358 9174 -12342
rect 9140 -13142 9174 -13126
rect 8053 -13188 8069 -13154
rect 8445 -13188 8461 -13154
rect 8689 -13188 8705 -13154
rect 9081 -13188 9097 -13154
rect 7838 -13288 7872 -13226
rect 9278 -13288 9312 -13226
rect 7838 -13322 7934 -13288
rect 9216 -13322 9312 -13288
rect 9438 -11670 9534 -11636
rect 10816 -11670 10912 -11636
rect 9438 -11732 9472 -11670
rect 10878 -11732 10912 -11670
rect 9653 -11804 9669 -11770
rect 10045 -11804 10061 -11770
rect 10289 -11804 10305 -11770
rect 10681 -11804 10697 -11770
rect 9576 -11832 9610 -11816
rect 9576 -12016 9610 -12000
rect 10104 -11832 10138 -11816
rect 10104 -12016 10138 -12000
rect 10212 -11832 10246 -11816
rect 10212 -12016 10246 -12000
rect 10740 -11832 10774 -11816
rect 10740 -12016 10774 -12000
rect 9653 -12062 9669 -12028
rect 10045 -12062 10061 -12028
rect 10289 -12062 10305 -12028
rect 10681 -12062 10697 -12028
rect 9438 -12162 9472 -12100
rect 10878 -12162 10912 -12100
rect 9438 -12196 9534 -12162
rect 10816 -12196 10912 -12162
rect 9438 -12258 9472 -12196
rect 10878 -12258 10912 -12196
rect 9653 -12330 9669 -12296
rect 10045 -12330 10061 -12296
rect 10289 -12330 10305 -12296
rect 10681 -12330 10697 -12296
rect 9576 -12358 9610 -12342
rect 9576 -13142 9610 -13126
rect 10104 -12358 10138 -12342
rect 10104 -13142 10138 -13126
rect 10212 -12358 10246 -12342
rect 10212 -13142 10246 -13126
rect 10740 -12358 10774 -12342
rect 10740 -13142 10774 -13126
rect 9653 -13188 9669 -13154
rect 10045 -13188 10061 -13154
rect 10289 -13188 10305 -13154
rect 10681 -13188 10697 -13154
rect 9438 -13288 9472 -13226
rect 10878 -13288 10912 -13226
rect 9438 -13322 9534 -13288
rect 10816 -13322 10912 -13288
rect 11038 -11670 11134 -11636
rect 12416 -11670 12512 -11636
rect 11038 -11732 11072 -11670
rect 12478 -11732 12512 -11670
rect 11253 -11804 11269 -11770
rect 11645 -11804 11661 -11770
rect 11889 -11804 11905 -11770
rect 12281 -11804 12297 -11770
rect 11176 -11832 11210 -11816
rect 11176 -12016 11210 -12000
rect 11704 -11832 11738 -11816
rect 11704 -12016 11738 -12000
rect 11812 -11832 11846 -11816
rect 11812 -12016 11846 -12000
rect 12340 -11832 12374 -11816
rect 12340 -12016 12374 -12000
rect 11253 -12062 11269 -12028
rect 11645 -12062 11661 -12028
rect 11889 -12062 11905 -12028
rect 12281 -12062 12297 -12028
rect 11038 -12162 11072 -12100
rect 12478 -12162 12512 -12100
rect 11038 -12196 11134 -12162
rect 12416 -12196 12512 -12162
rect 11038 -12258 11072 -12196
rect 12478 -12258 12512 -12196
rect 11253 -12330 11269 -12296
rect 11645 -12330 11661 -12296
rect 11889 -12330 11905 -12296
rect 12281 -12330 12297 -12296
rect 11176 -12358 11210 -12342
rect 11176 -13142 11210 -13126
rect 11704 -12358 11738 -12342
rect 11704 -13142 11738 -13126
rect 11812 -12358 11846 -12342
rect 11812 -13142 11846 -13126
rect 12340 -12358 12374 -12342
rect 12340 -13142 12374 -13126
rect 11253 -13188 11269 -13154
rect 11645 -13188 11661 -13154
rect 11889 -13188 11905 -13154
rect 12281 -13188 12297 -13154
rect 11038 -13288 11072 -13226
rect 12478 -13288 12512 -13226
rect 11038 -13322 11134 -13288
rect 12416 -13322 12512 -13288
rect 12638 -11670 12734 -11636
rect 14016 -11670 14112 -11636
rect 12638 -11732 12672 -11670
rect 14078 -11732 14112 -11670
rect 12853 -11804 12869 -11770
rect 13245 -11804 13261 -11770
rect 13489 -11804 13505 -11770
rect 13881 -11804 13897 -11770
rect 12776 -11832 12810 -11816
rect 12776 -12016 12810 -12000
rect 13304 -11832 13338 -11816
rect 13304 -12016 13338 -12000
rect 13412 -11832 13446 -11816
rect 13412 -12016 13446 -12000
rect 13940 -11832 13974 -11816
rect 13940 -12016 13974 -12000
rect 12853 -12062 12869 -12028
rect 13245 -12062 13261 -12028
rect 13489 -12062 13505 -12028
rect 13881 -12062 13897 -12028
rect 12638 -12162 12672 -12100
rect 14078 -12162 14112 -12100
rect 12638 -12196 12734 -12162
rect 14016 -12196 14112 -12162
rect 12638 -12258 12672 -12196
rect 14078 -12258 14112 -12196
rect 12853 -12330 12869 -12296
rect 13245 -12330 13261 -12296
rect 13489 -12330 13505 -12296
rect 13881 -12330 13897 -12296
rect 12776 -12358 12810 -12342
rect 12776 -13142 12810 -13126
rect 13304 -12358 13338 -12342
rect 13304 -13142 13338 -13126
rect 13412 -12358 13446 -12342
rect 13412 -13142 13446 -13126
rect 13940 -12358 13974 -12342
rect 13940 -13142 13974 -13126
rect 12853 -13188 12869 -13154
rect 13245 -13188 13261 -13154
rect 13489 -13188 13505 -13154
rect 13881 -13188 13897 -13154
rect 12638 -13288 12672 -13226
rect 14078 -13288 14112 -13226
rect 12638 -13322 12734 -13288
rect 14016 -13322 14112 -13288
rect 14238 -11670 14334 -11636
rect 15616 -11670 15712 -11636
rect 14238 -11732 14272 -11670
rect 15678 -11732 15712 -11670
rect 14453 -11804 14469 -11770
rect 14845 -11804 14861 -11770
rect 15089 -11804 15105 -11770
rect 15481 -11804 15497 -11770
rect 14376 -11832 14410 -11816
rect 14376 -12016 14410 -12000
rect 14904 -11832 14938 -11816
rect 14904 -12016 14938 -12000
rect 15012 -11832 15046 -11816
rect 15012 -12016 15046 -12000
rect 15540 -11832 15574 -11816
rect 15540 -12016 15574 -12000
rect 14453 -12062 14469 -12028
rect 14845 -12062 14861 -12028
rect 15089 -12062 15105 -12028
rect 15481 -12062 15497 -12028
rect 14238 -12162 14272 -12100
rect 15678 -12162 15712 -12100
rect 14238 -12196 14334 -12162
rect 15616 -12196 15712 -12162
rect 14238 -12258 14272 -12196
rect 15678 -12258 15712 -12196
rect 14453 -12330 14469 -12296
rect 14845 -12330 14861 -12296
rect 15089 -12330 15105 -12296
rect 15481 -12330 15497 -12296
rect 14376 -12358 14410 -12342
rect 14376 -13142 14410 -13126
rect 14904 -12358 14938 -12342
rect 14904 -13142 14938 -13126
rect 15012 -12358 15046 -12342
rect 15012 -13142 15046 -13126
rect 15540 -12358 15574 -12342
rect 15540 -13142 15574 -13126
rect 14453 -13188 14469 -13154
rect 14845 -13188 14861 -13154
rect 15089 -13188 15105 -13154
rect 15481 -13188 15497 -13154
rect 14238 -13288 14272 -13226
rect 15678 -13288 15712 -13226
rect 14238 -13322 14334 -13288
rect 15616 -13322 15712 -13288
rect 15838 -11670 15934 -11636
rect 17216 -11670 17312 -11636
rect 15838 -11732 15872 -11670
rect 17278 -11732 17312 -11670
rect 16053 -11804 16069 -11770
rect 16445 -11804 16461 -11770
rect 16689 -11804 16705 -11770
rect 17081 -11804 17097 -11770
rect 15976 -11832 16010 -11816
rect 15976 -12016 16010 -12000
rect 16504 -11832 16538 -11816
rect 16504 -12016 16538 -12000
rect 16612 -11832 16646 -11816
rect 16612 -12016 16646 -12000
rect 17140 -11832 17174 -11816
rect 17140 -12016 17174 -12000
rect 16053 -12062 16069 -12028
rect 16445 -12062 16461 -12028
rect 16689 -12062 16705 -12028
rect 17081 -12062 17097 -12028
rect 15838 -12162 15872 -12100
rect 17278 -12162 17312 -12100
rect 15838 -12196 15934 -12162
rect 17216 -12196 17312 -12162
rect 15838 -12258 15872 -12196
rect 17278 -12258 17312 -12196
rect 16053 -12330 16069 -12296
rect 16445 -12330 16461 -12296
rect 16689 -12330 16705 -12296
rect 17081 -12330 17097 -12296
rect 15976 -12358 16010 -12342
rect 15976 -13142 16010 -13126
rect 16504 -12358 16538 -12342
rect 16504 -13142 16538 -13126
rect 16612 -12358 16646 -12342
rect 16612 -13142 16646 -13126
rect 17140 -12358 17174 -12342
rect 17140 -13142 17174 -13126
rect 16053 -13188 16069 -13154
rect 16445 -13188 16461 -13154
rect 16689 -13188 16705 -13154
rect 17081 -13188 17097 -13154
rect 15838 -13288 15872 -13226
rect 17278 -13288 17312 -13226
rect 15838 -13322 15934 -13288
rect 17216 -13322 17312 -13288
rect 17438 -11670 17534 -11636
rect 18816 -11670 18912 -11636
rect 17438 -11732 17472 -11670
rect 18878 -11732 18912 -11670
rect 17653 -11804 17669 -11770
rect 18045 -11804 18061 -11770
rect 18289 -11804 18305 -11770
rect 18681 -11804 18697 -11770
rect 17576 -11832 17610 -11816
rect 17576 -12016 17610 -12000
rect 18104 -11832 18138 -11816
rect 18104 -12016 18138 -12000
rect 18212 -11832 18246 -11816
rect 18212 -12016 18246 -12000
rect 18740 -11832 18774 -11816
rect 18740 -12016 18774 -12000
rect 17653 -12062 17669 -12028
rect 18045 -12062 18061 -12028
rect 18289 -12062 18305 -12028
rect 18681 -12062 18697 -12028
rect 17438 -12162 17472 -12100
rect 18878 -12162 18912 -12100
rect 17438 -12196 17534 -12162
rect 18816 -12196 18912 -12162
rect 17438 -12258 17472 -12196
rect 18878 -12258 18912 -12196
rect 17653 -12330 17669 -12296
rect 18045 -12330 18061 -12296
rect 18289 -12330 18305 -12296
rect 18681 -12330 18697 -12296
rect 17576 -12358 17610 -12342
rect 17576 -13142 17610 -13126
rect 18104 -12358 18138 -12342
rect 18104 -13142 18138 -13126
rect 18212 -12358 18246 -12342
rect 18212 -13142 18246 -13126
rect 18740 -12358 18774 -12342
rect 18740 -13142 18774 -13126
rect 17653 -13188 17669 -13154
rect 18045 -13188 18061 -13154
rect 18289 -13188 18305 -13154
rect 18681 -13188 18697 -13154
rect 17438 -13288 17472 -13226
rect 18878 -13288 18912 -13226
rect 17438 -13322 17534 -13288
rect 18816 -13322 18912 -13288
rect 19038 -11670 19134 -11636
rect 20416 -11670 20512 -11636
rect 19038 -11732 19072 -11670
rect 20478 -11732 20512 -11670
rect 19253 -11804 19269 -11770
rect 19645 -11804 19661 -11770
rect 19889 -11804 19905 -11770
rect 20281 -11804 20297 -11770
rect 19176 -11832 19210 -11816
rect 19176 -12016 19210 -12000
rect 19704 -11832 19738 -11816
rect 19704 -12016 19738 -12000
rect 19812 -11832 19846 -11816
rect 19812 -12016 19846 -12000
rect 20340 -11832 20374 -11816
rect 20340 -12016 20374 -12000
rect 19253 -12062 19269 -12028
rect 19645 -12062 19661 -12028
rect 19889 -12062 19905 -12028
rect 20281 -12062 20297 -12028
rect 19038 -12162 19072 -12100
rect 20478 -12162 20512 -12100
rect 19038 -12196 19134 -12162
rect 20416 -12196 20512 -12162
rect 19038 -12258 19072 -12196
rect 20478 -12258 20512 -12196
rect 19253 -12330 19269 -12296
rect 19645 -12330 19661 -12296
rect 19889 -12330 19905 -12296
rect 20281 -12330 20297 -12296
rect 19176 -12358 19210 -12342
rect 19176 -13142 19210 -13126
rect 19704 -12358 19738 -12342
rect 19704 -13142 19738 -13126
rect 19812 -12358 19846 -12342
rect 19812 -13142 19846 -13126
rect 20340 -12358 20374 -12342
rect 20340 -13142 20374 -13126
rect 19253 -13188 19269 -13154
rect 19645 -13188 19661 -13154
rect 19889 -13188 19905 -13154
rect 20281 -13188 20297 -13154
rect 19038 -13288 19072 -13226
rect 20478 -13288 20512 -13226
rect 19038 -13322 19134 -13288
rect 20416 -13322 20512 -13288
rect 20638 -11670 20734 -11636
rect 22016 -11670 22112 -11636
rect 20638 -11732 20672 -11670
rect 22078 -11732 22112 -11670
rect 20853 -11804 20869 -11770
rect 21245 -11804 21261 -11770
rect 21489 -11804 21505 -11770
rect 21881 -11804 21897 -11770
rect 20776 -11832 20810 -11816
rect 20776 -12016 20810 -12000
rect 21304 -11832 21338 -11816
rect 21304 -12016 21338 -12000
rect 21412 -11832 21446 -11816
rect 21412 -12016 21446 -12000
rect 21940 -11832 21974 -11816
rect 21940 -12016 21974 -12000
rect 20853 -12062 20869 -12028
rect 21245 -12062 21261 -12028
rect 21489 -12062 21505 -12028
rect 21881 -12062 21897 -12028
rect 20638 -12162 20672 -12100
rect 22078 -12162 22112 -12100
rect 20638 -12196 20734 -12162
rect 22016 -12196 22112 -12162
rect 20638 -12258 20672 -12196
rect 22078 -12258 22112 -12196
rect 20853 -12330 20869 -12296
rect 21245 -12330 21261 -12296
rect 21489 -12330 21505 -12296
rect 21881 -12330 21897 -12296
rect 20776 -12358 20810 -12342
rect 20776 -13142 20810 -13126
rect 21304 -12358 21338 -12342
rect 21304 -13142 21338 -13126
rect 21412 -12358 21446 -12342
rect 21412 -13142 21446 -13126
rect 21940 -12358 21974 -12342
rect 21940 -13142 21974 -13126
rect 20853 -13188 20869 -13154
rect 21245 -13188 21261 -13154
rect 21489 -13188 21505 -13154
rect 21881 -13188 21897 -13154
rect 20638 -13288 20672 -13226
rect 22078 -13288 22112 -13226
rect 20638 -13322 20734 -13288
rect 22016 -13322 22112 -13288
rect 22238 -11670 22334 -11636
rect 23616 -11670 23712 -11636
rect 22238 -11732 22272 -11670
rect 23678 -11732 23712 -11670
rect 22453 -11804 22469 -11770
rect 22845 -11804 22861 -11770
rect 23089 -11804 23105 -11770
rect 23481 -11804 23497 -11770
rect 22376 -11832 22410 -11816
rect 22376 -12016 22410 -12000
rect 22904 -11832 22938 -11816
rect 22904 -12016 22938 -12000
rect 23012 -11832 23046 -11816
rect 23012 -12016 23046 -12000
rect 23540 -11832 23574 -11816
rect 23540 -12016 23574 -12000
rect 22453 -12062 22469 -12028
rect 22845 -12062 22861 -12028
rect 23089 -12062 23105 -12028
rect 23481 -12062 23497 -12028
rect 22238 -12162 22272 -12100
rect 23678 -12162 23712 -12100
rect 22238 -12196 22334 -12162
rect 23616 -12196 23712 -12162
rect 22238 -12258 22272 -12196
rect 23678 -12258 23712 -12196
rect 22453 -12330 22469 -12296
rect 22845 -12330 22861 -12296
rect 23089 -12330 23105 -12296
rect 23481 -12330 23497 -12296
rect 22376 -12358 22410 -12342
rect 22376 -13142 22410 -13126
rect 22904 -12358 22938 -12342
rect 22904 -13142 22938 -13126
rect 23012 -12358 23046 -12342
rect 23012 -13142 23046 -13126
rect 23540 -12358 23574 -12342
rect 23540 -13142 23574 -13126
rect 22453 -13188 22469 -13154
rect 22845 -13188 22861 -13154
rect 23089 -13188 23105 -13154
rect 23481 -13188 23497 -13154
rect 22238 -13288 22272 -13226
rect 23678 -13288 23712 -13226
rect 22238 -13322 22334 -13288
rect 23616 -13322 23712 -13288
rect 23838 -11670 23934 -11636
rect 25216 -11670 25312 -11636
rect 23838 -11732 23872 -11670
rect 25278 -11732 25312 -11670
rect 24053 -11804 24069 -11770
rect 24445 -11804 24461 -11770
rect 24689 -11804 24705 -11770
rect 25081 -11804 25097 -11770
rect 23976 -11832 24010 -11816
rect 23976 -12016 24010 -12000
rect 24504 -11832 24538 -11816
rect 24504 -12016 24538 -12000
rect 24612 -11832 24646 -11816
rect 24612 -12016 24646 -12000
rect 25140 -11832 25174 -11816
rect 25140 -12016 25174 -12000
rect 24053 -12062 24069 -12028
rect 24445 -12062 24461 -12028
rect 24689 -12062 24705 -12028
rect 25081 -12062 25097 -12028
rect 23838 -12162 23872 -12100
rect 25278 -12162 25312 -12100
rect 23838 -12196 23934 -12162
rect 25216 -12196 25312 -12162
rect 23838 -12258 23872 -12196
rect 25278 -12258 25312 -12196
rect 24053 -12330 24069 -12296
rect 24445 -12330 24461 -12296
rect 24689 -12330 24705 -12296
rect 25081 -12330 25097 -12296
rect 23976 -12358 24010 -12342
rect 23976 -13142 24010 -13126
rect 24504 -12358 24538 -12342
rect 24504 -13142 24538 -13126
rect 24612 -12358 24646 -12342
rect 24612 -13142 24646 -13126
rect 25140 -12358 25174 -12342
rect 25140 -13142 25174 -13126
rect 24053 -13188 24069 -13154
rect 24445 -13188 24461 -13154
rect 24689 -13188 24705 -13154
rect 25081 -13188 25097 -13154
rect 23838 -13288 23872 -13226
rect 25278 -13288 25312 -13226
rect 23838 -13322 23934 -13288
rect 25216 -13322 25312 -13288
rect 25438 -11670 25534 -11636
rect 26816 -11670 26912 -11636
rect 25438 -11732 25472 -11670
rect 26878 -11732 26912 -11670
rect 25653 -11804 25669 -11770
rect 26045 -11804 26061 -11770
rect 26289 -11804 26305 -11770
rect 26681 -11804 26697 -11770
rect 25576 -11832 25610 -11816
rect 25576 -12016 25610 -12000
rect 26104 -11832 26138 -11816
rect 26104 -12016 26138 -12000
rect 26212 -11832 26246 -11816
rect 26212 -12016 26246 -12000
rect 26740 -11832 26774 -11816
rect 26740 -12016 26774 -12000
rect 25653 -12062 25669 -12028
rect 26045 -12062 26061 -12028
rect 26289 -12062 26305 -12028
rect 26681 -12062 26697 -12028
rect 25438 -12162 25472 -12100
rect 26878 -12162 26912 -12100
rect 25438 -12196 25534 -12162
rect 26816 -12196 26912 -12162
rect 25438 -12258 25472 -12196
rect 26878 -12258 26912 -12196
rect 25653 -12330 25669 -12296
rect 26045 -12330 26061 -12296
rect 26289 -12330 26305 -12296
rect 26681 -12330 26697 -12296
rect 25576 -12358 25610 -12342
rect 25576 -13142 25610 -13126
rect 26104 -12358 26138 -12342
rect 26104 -13142 26138 -13126
rect 26212 -12358 26246 -12342
rect 26212 -13142 26246 -13126
rect 26740 -12358 26774 -12342
rect 26740 -13142 26774 -13126
rect 25653 -13188 25669 -13154
rect 26045 -13188 26061 -13154
rect 26289 -13188 26305 -13154
rect 26681 -13188 26697 -13154
rect 25438 -13288 25472 -13226
rect 26878 -13288 26912 -13226
rect 25438 -13322 25534 -13288
rect 26816 -13322 26912 -13288
rect 27038 -11670 27134 -11636
rect 28416 -11670 28512 -11636
rect 27038 -11732 27072 -11670
rect 28478 -11732 28512 -11670
rect 27253 -11804 27269 -11770
rect 27645 -11804 27661 -11770
rect 27889 -11804 27905 -11770
rect 28281 -11804 28297 -11770
rect 27176 -11832 27210 -11816
rect 27176 -12016 27210 -12000
rect 27704 -11832 27738 -11816
rect 27704 -12016 27738 -12000
rect 27812 -11832 27846 -11816
rect 27812 -12016 27846 -12000
rect 28340 -11832 28374 -11816
rect 28340 -12016 28374 -12000
rect 27253 -12062 27269 -12028
rect 27645 -12062 27661 -12028
rect 27889 -12062 27905 -12028
rect 28281 -12062 28297 -12028
rect 27038 -12162 27072 -12100
rect 28478 -12162 28512 -12100
rect 27038 -12196 27134 -12162
rect 28416 -12196 28512 -12162
rect 27038 -12258 27072 -12196
rect 28478 -12258 28512 -12196
rect 27253 -12330 27269 -12296
rect 27645 -12330 27661 -12296
rect 27889 -12330 27905 -12296
rect 28281 -12330 28297 -12296
rect 27176 -12358 27210 -12342
rect 27176 -13142 27210 -13126
rect 27704 -12358 27738 -12342
rect 27704 -13142 27738 -13126
rect 27812 -12358 27846 -12342
rect 27812 -13142 27846 -13126
rect 28340 -12358 28374 -12342
rect 28340 -13142 28374 -13126
rect 27253 -13188 27269 -13154
rect 27645 -13188 27661 -13154
rect 27889 -13188 27905 -13154
rect 28281 -13188 28297 -13154
rect 27038 -13288 27072 -13226
rect 28478 -13288 28512 -13226
rect 27038 -13322 27134 -13288
rect 28416 -13322 28512 -13288
rect 28638 -11670 28734 -11636
rect 30016 -11670 30112 -11636
rect 28638 -11732 28672 -11670
rect 30078 -11732 30112 -11670
rect 28853 -11804 28869 -11770
rect 29245 -11804 29261 -11770
rect 29489 -11804 29505 -11770
rect 29881 -11804 29897 -11770
rect 28776 -11832 28810 -11816
rect 28776 -12016 28810 -12000
rect 29304 -11832 29338 -11816
rect 29304 -12016 29338 -12000
rect 29412 -11832 29446 -11816
rect 29412 -12016 29446 -12000
rect 29940 -11832 29974 -11816
rect 29940 -12016 29974 -12000
rect 28853 -12062 28869 -12028
rect 29245 -12062 29261 -12028
rect 29489 -12062 29505 -12028
rect 29881 -12062 29897 -12028
rect 28638 -12162 28672 -12100
rect 30078 -12162 30112 -12100
rect 28638 -12196 28734 -12162
rect 30016 -12196 30112 -12162
rect 28638 -12258 28672 -12196
rect 30078 -12258 30112 -12196
rect 28853 -12330 28869 -12296
rect 29245 -12330 29261 -12296
rect 29489 -12330 29505 -12296
rect 29881 -12330 29897 -12296
rect 28776 -12358 28810 -12342
rect 28776 -13142 28810 -13126
rect 29304 -12358 29338 -12342
rect 29304 -13142 29338 -13126
rect 29412 -12358 29446 -12342
rect 29412 -13142 29446 -13126
rect 29940 -12358 29974 -12342
rect 29940 -13142 29974 -13126
rect 28853 -13188 28869 -13154
rect 29245 -13188 29261 -13154
rect 29489 -13188 29505 -13154
rect 29881 -13188 29897 -13154
rect 28638 -13288 28672 -13226
rect 30078 -13288 30112 -13226
rect 28638 -13322 28734 -13288
rect 30016 -13322 30112 -13288
rect 30238 -11670 30334 -11636
rect 31616 -11670 31712 -11636
rect 30238 -11732 30272 -11670
rect 31678 -11732 31712 -11670
rect 30453 -11804 30469 -11770
rect 30845 -11804 30861 -11770
rect 31089 -11804 31105 -11770
rect 31481 -11804 31497 -11770
rect 30376 -11832 30410 -11816
rect 30376 -12016 30410 -12000
rect 30904 -11832 30938 -11816
rect 30904 -12016 30938 -12000
rect 31012 -11832 31046 -11816
rect 31012 -12016 31046 -12000
rect 31540 -11832 31574 -11816
rect 31540 -12016 31574 -12000
rect 30453 -12062 30469 -12028
rect 30845 -12062 30861 -12028
rect 31089 -12062 31105 -12028
rect 31481 -12062 31497 -12028
rect 30238 -12162 30272 -12100
rect 31678 -12162 31712 -12100
rect 30238 -12196 30334 -12162
rect 31616 -12196 31712 -12162
rect 30238 -12258 30272 -12196
rect 31678 -12258 31712 -12196
rect 30453 -12330 30469 -12296
rect 30845 -12330 30861 -12296
rect 31089 -12330 31105 -12296
rect 31481 -12330 31497 -12296
rect 30376 -12358 30410 -12342
rect 30376 -13142 30410 -13126
rect 30904 -12358 30938 -12342
rect 30904 -13142 30938 -13126
rect 31012 -12358 31046 -12342
rect 31012 -13142 31046 -13126
rect 31540 -12358 31574 -12342
rect 31540 -13142 31574 -13126
rect 30453 -13188 30469 -13154
rect 30845 -13188 30861 -13154
rect 31089 -13188 31105 -13154
rect 31481 -13188 31497 -13154
rect 30238 -13288 30272 -13226
rect 31678 -13288 31712 -13226
rect 30238 -13322 30334 -13288
rect 31616 -13322 31712 -13288
rect 31838 -11670 31934 -11636
rect 33216 -11670 33312 -11636
rect 31838 -11732 31872 -11670
rect 33278 -11732 33312 -11670
rect 32053 -11804 32069 -11770
rect 32445 -11804 32461 -11770
rect 32689 -11804 32705 -11770
rect 33081 -11804 33097 -11770
rect 31976 -11832 32010 -11816
rect 31976 -12016 32010 -12000
rect 32504 -11832 32538 -11816
rect 32504 -12016 32538 -12000
rect 32612 -11832 32646 -11816
rect 32612 -12016 32646 -12000
rect 33140 -11832 33174 -11816
rect 33140 -12016 33174 -12000
rect 32053 -12062 32069 -12028
rect 32445 -12062 32461 -12028
rect 32689 -12062 32705 -12028
rect 33081 -12062 33097 -12028
rect 31838 -12162 31872 -12100
rect 33278 -12162 33312 -12100
rect 31838 -12196 31934 -12162
rect 33216 -12196 33312 -12162
rect 31838 -12258 31872 -12196
rect 33278 -12258 33312 -12196
rect 32053 -12330 32069 -12296
rect 32445 -12330 32461 -12296
rect 32689 -12330 32705 -12296
rect 33081 -12330 33097 -12296
rect 31976 -12358 32010 -12342
rect 31976 -13142 32010 -13126
rect 32504 -12358 32538 -12342
rect 32504 -13142 32538 -13126
rect 32612 -12358 32646 -12342
rect 32612 -13142 32646 -13126
rect 33140 -12358 33174 -12342
rect 33140 -13142 33174 -13126
rect 32053 -13188 32069 -13154
rect 32445 -13188 32461 -13154
rect 32689 -13188 32705 -13154
rect 33081 -13188 33097 -13154
rect 31838 -13288 31872 -13226
rect 33278 -13288 33312 -13226
rect 31838 -13322 31934 -13288
rect 33216 -13322 33312 -13288
rect 33438 -11670 33534 -11636
rect 34816 -11670 34912 -11636
rect 33438 -11732 33472 -11670
rect 34878 -11732 34912 -11670
rect 33653 -11804 33669 -11770
rect 34045 -11804 34061 -11770
rect 34289 -11804 34305 -11770
rect 34681 -11804 34697 -11770
rect 33576 -11832 33610 -11816
rect 33576 -12016 33610 -12000
rect 34104 -11832 34138 -11816
rect 34104 -12016 34138 -12000
rect 34212 -11832 34246 -11816
rect 34212 -12016 34246 -12000
rect 34740 -11832 34774 -11816
rect 34740 -12016 34774 -12000
rect 33653 -12062 33669 -12028
rect 34045 -12062 34061 -12028
rect 34289 -12062 34305 -12028
rect 34681 -12062 34697 -12028
rect 33438 -12162 33472 -12100
rect 34878 -12162 34912 -12100
rect 33438 -12196 33534 -12162
rect 34816 -12196 34912 -12162
rect 33438 -12258 33472 -12196
rect 34878 -12258 34912 -12196
rect 33653 -12330 33669 -12296
rect 34045 -12330 34061 -12296
rect 34289 -12330 34305 -12296
rect 34681 -12330 34697 -12296
rect 33576 -12358 33610 -12342
rect 33576 -13142 33610 -13126
rect 34104 -12358 34138 -12342
rect 34104 -13142 34138 -13126
rect 34212 -12358 34246 -12342
rect 34212 -13142 34246 -13126
rect 34740 -12358 34774 -12342
rect 34740 -13142 34774 -13126
rect 33653 -13188 33669 -13154
rect 34045 -13188 34061 -13154
rect 34289 -13188 34305 -13154
rect 34681 -13188 34697 -13154
rect 33438 -13288 33472 -13226
rect 34878 -13288 34912 -13226
rect 33438 -13322 33534 -13288
rect 34816 -13322 34912 -13288
rect 35038 -11670 35134 -11636
rect 36416 -11670 36734 -11636
rect 38016 -11670 38112 -11636
rect 35038 -11732 35072 -11670
rect 36478 -11732 38112 -11670
rect 35253 -11804 35269 -11770
rect 35645 -11804 35661 -11770
rect 35889 -11804 35905 -11770
rect 36281 -11804 36297 -11770
rect 35176 -11832 35210 -11816
rect 35176 -12016 35210 -12000
rect 35704 -11832 35738 -11816
rect 35704 -12016 35738 -12000
rect 35812 -11832 35846 -11816
rect 35812 -12016 35846 -12000
rect 36340 -11832 36374 -11816
rect 36340 -12016 36374 -12000
rect 35253 -12062 35269 -12028
rect 35645 -12062 35661 -12028
rect 35889 -12062 35905 -12028
rect 36281 -12062 36297 -12028
rect 35038 -12162 35072 -12100
rect 36512 -12100 36638 -11732
rect 36672 -11770 38078 -11732
rect 36672 -11804 36869 -11770
rect 37245 -11804 37505 -11770
rect 37881 -11804 38078 -11770
rect 36672 -11832 38078 -11804
rect 36672 -12000 36776 -11832
rect 36810 -12000 37304 -11832
rect 37338 -12000 37412 -11832
rect 37446 -12000 37940 -11832
rect 37974 -12000 38078 -11832
rect 36672 -12028 38078 -12000
rect 36672 -12062 36869 -12028
rect 37245 -12062 37505 -12028
rect 37881 -12062 38078 -12028
rect 36672 -12100 38078 -12062
rect 36478 -12162 38112 -12100
rect 35038 -12196 35134 -12162
rect 36416 -12196 36734 -12162
rect 38016 -12196 38112 -12162
rect 35038 -12258 35072 -12196
rect 36478 -12258 38112 -12196
rect 35253 -12330 35269 -12296
rect 35645 -12330 35661 -12296
rect 35889 -12330 35905 -12296
rect 36281 -12330 36297 -12296
rect 35176 -12358 35210 -12342
rect 35176 -13142 35210 -13126
rect 35704 -12358 35738 -12342
rect 35704 -13142 35738 -13126
rect 35812 -12358 35846 -12342
rect 35812 -13142 35846 -13126
rect 36340 -12358 36374 -12342
rect 36340 -13142 36374 -13126
rect 35253 -13188 35269 -13154
rect 35645 -13188 35661 -13154
rect 35889 -13188 35905 -13154
rect 36281 -13188 36297 -13154
rect 35038 -13288 35072 -13226
rect 36512 -13226 36638 -12258
rect 36672 -12296 38078 -12258
rect 36672 -12330 36869 -12296
rect 37245 -12330 37505 -12296
rect 37881 -12330 38078 -12296
rect 36672 -12358 38078 -12330
rect 36672 -13126 36776 -12358
rect 36810 -13126 37304 -12358
rect 37338 -13126 37412 -12358
rect 37446 -13126 37940 -12358
rect 37974 -13126 38078 -12358
rect 36672 -13154 38078 -13126
rect 36672 -13188 36869 -13154
rect 37245 -13188 37505 -13154
rect 37881 -13188 38078 -13154
rect 36672 -13226 38078 -13188
rect 36478 -13288 38112 -13226
rect 35038 -13322 35134 -13288
rect 36416 -13322 36734 -13288
rect 38016 -13322 38112 -13288
rect -140 -13436 1460 -13322
rect 36500 -13436 38100 -13322
rect -162 -13470 -66 -13436
rect 1216 -13470 1534 -13436
rect 2816 -13470 2912 -13436
rect -162 -13532 1472 -13470
rect -128 -13570 1278 -13532
rect -128 -13604 69 -13570
rect 445 -13604 705 -13570
rect 1081 -13604 1278 -13570
rect -128 -13632 1278 -13604
rect -128 -13800 -24 -13632
rect 10 -13800 504 -13632
rect 538 -13800 612 -13632
rect 646 -13800 1140 -13632
rect 1174 -13800 1278 -13632
rect -128 -13828 1278 -13800
rect -128 -13862 69 -13828
rect 445 -13862 705 -13828
rect 1081 -13862 1278 -13828
rect -128 -13900 1278 -13862
rect 1312 -13900 1438 -13532
rect 2878 -13532 2912 -13470
rect 1653 -13604 1669 -13570
rect 2045 -13604 2061 -13570
rect 2289 -13604 2305 -13570
rect 2681 -13604 2697 -13570
rect 1576 -13632 1610 -13616
rect 1576 -13816 1610 -13800
rect 2104 -13632 2138 -13616
rect 2104 -13816 2138 -13800
rect 2212 -13632 2246 -13616
rect 2212 -13816 2246 -13800
rect 2740 -13632 2774 -13616
rect 2740 -13816 2774 -13800
rect 1653 -13862 1669 -13828
rect 2045 -13862 2061 -13828
rect 2289 -13862 2305 -13828
rect 2681 -13862 2697 -13828
rect -162 -13962 1472 -13900
rect 2878 -13962 2912 -13900
rect -162 -13996 -66 -13962
rect 1216 -13996 1534 -13962
rect 2816 -13996 2912 -13962
rect -162 -14058 1472 -13996
rect -128 -14096 1278 -14058
rect -128 -14130 69 -14096
rect 445 -14130 705 -14096
rect 1081 -14130 1278 -14096
rect -128 -14158 1278 -14130
rect -128 -14926 -24 -14158
rect 10 -14926 504 -14158
rect 538 -14926 612 -14158
rect 646 -14926 1140 -14158
rect 1174 -14926 1278 -14158
rect -128 -14954 1278 -14926
rect -128 -14988 69 -14954
rect 445 -14988 705 -14954
rect 1081 -14988 1278 -14954
rect -128 -15026 1278 -14988
rect 1312 -15026 1438 -14058
rect 2878 -14058 2912 -13996
rect 1653 -14130 1669 -14096
rect 2045 -14130 2061 -14096
rect 2289 -14130 2305 -14096
rect 2681 -14130 2697 -14096
rect 1576 -14158 1610 -14142
rect 1576 -14942 1610 -14926
rect 2104 -14158 2138 -14142
rect 2104 -14942 2138 -14926
rect 2212 -14158 2246 -14142
rect 2212 -14942 2246 -14926
rect 2740 -14158 2774 -14142
rect 2740 -14942 2774 -14926
rect 1653 -14988 1669 -14954
rect 2045 -14988 2061 -14954
rect 2289 -14988 2305 -14954
rect 2681 -14988 2697 -14954
rect -162 -15088 1472 -15026
rect 2878 -15088 2912 -15026
rect -162 -15122 -66 -15088
rect 1216 -15122 1534 -15088
rect 2816 -15122 2912 -15088
rect 3038 -13470 3134 -13436
rect 4416 -13470 4512 -13436
rect 3038 -13532 3072 -13470
rect 4478 -13532 4512 -13470
rect 3253 -13604 3269 -13570
rect 3645 -13604 3661 -13570
rect 3889 -13604 3905 -13570
rect 4281 -13604 4297 -13570
rect 3176 -13632 3210 -13616
rect 3176 -13816 3210 -13800
rect 3704 -13632 3738 -13616
rect 3704 -13816 3738 -13800
rect 3812 -13632 3846 -13616
rect 3812 -13816 3846 -13800
rect 4340 -13632 4374 -13616
rect 4340 -13816 4374 -13800
rect 3253 -13862 3269 -13828
rect 3645 -13862 3661 -13828
rect 3889 -13862 3905 -13828
rect 4281 -13862 4297 -13828
rect 3038 -13962 3072 -13900
rect 4478 -13962 4512 -13900
rect 3038 -13996 3134 -13962
rect 4416 -13996 4512 -13962
rect 3038 -14058 3072 -13996
rect 4478 -14058 4512 -13996
rect 3253 -14130 3269 -14096
rect 3645 -14130 3661 -14096
rect 3889 -14130 3905 -14096
rect 4281 -14130 4297 -14096
rect 3176 -14158 3210 -14142
rect 3176 -14942 3210 -14926
rect 3704 -14158 3738 -14142
rect 3704 -14942 3738 -14926
rect 3812 -14158 3846 -14142
rect 3812 -14942 3846 -14926
rect 4340 -14158 4374 -14142
rect 4340 -14942 4374 -14926
rect 3253 -14988 3269 -14954
rect 3645 -14988 3661 -14954
rect 3889 -14988 3905 -14954
rect 4281 -14988 4297 -14954
rect 3038 -15088 3072 -15026
rect 4478 -15088 4512 -15026
rect 3038 -15122 3134 -15088
rect 4416 -15122 4512 -15088
rect 4638 -13470 4734 -13436
rect 6016 -13470 6112 -13436
rect 4638 -13532 4672 -13470
rect 6078 -13532 6112 -13470
rect 4853 -13604 4869 -13570
rect 5245 -13604 5261 -13570
rect 5489 -13604 5505 -13570
rect 5881 -13604 5897 -13570
rect 4776 -13632 4810 -13616
rect 4776 -13816 4810 -13800
rect 5304 -13632 5338 -13616
rect 5304 -13816 5338 -13800
rect 5412 -13632 5446 -13616
rect 5412 -13816 5446 -13800
rect 5940 -13632 5974 -13616
rect 5940 -13816 5974 -13800
rect 4853 -13862 4869 -13828
rect 5245 -13862 5261 -13828
rect 5489 -13862 5505 -13828
rect 5881 -13862 5897 -13828
rect 4638 -13962 4672 -13900
rect 6078 -13962 6112 -13900
rect 4638 -13996 4734 -13962
rect 6016 -13996 6112 -13962
rect 4638 -14058 4672 -13996
rect 6078 -14058 6112 -13996
rect 4853 -14130 4869 -14096
rect 5245 -14130 5261 -14096
rect 5489 -14130 5505 -14096
rect 5881 -14130 5897 -14096
rect 4776 -14158 4810 -14142
rect 4776 -14942 4810 -14926
rect 5304 -14158 5338 -14142
rect 5304 -14942 5338 -14926
rect 5412 -14158 5446 -14142
rect 5412 -14942 5446 -14926
rect 5940 -14158 5974 -14142
rect 5940 -14942 5974 -14926
rect 4853 -14988 4869 -14954
rect 5245 -14988 5261 -14954
rect 5489 -14988 5505 -14954
rect 5881 -14988 5897 -14954
rect 4638 -15088 4672 -15026
rect 6078 -15088 6112 -15026
rect 4638 -15122 4734 -15088
rect 6016 -15122 6112 -15088
rect 6238 -13470 6334 -13436
rect 7616 -13470 7712 -13436
rect 6238 -13532 6272 -13470
rect 7678 -13532 7712 -13470
rect 6453 -13604 6469 -13570
rect 6845 -13604 6861 -13570
rect 7089 -13604 7105 -13570
rect 7481 -13604 7497 -13570
rect 6376 -13632 6410 -13616
rect 6376 -13816 6410 -13800
rect 6904 -13632 6938 -13616
rect 6904 -13816 6938 -13800
rect 7012 -13632 7046 -13616
rect 7012 -13816 7046 -13800
rect 7540 -13632 7574 -13616
rect 7540 -13816 7574 -13800
rect 6453 -13862 6469 -13828
rect 6845 -13862 6861 -13828
rect 7089 -13862 7105 -13828
rect 7481 -13862 7497 -13828
rect 6238 -13962 6272 -13900
rect 7678 -13962 7712 -13900
rect 6238 -13996 6334 -13962
rect 7616 -13996 7712 -13962
rect 6238 -14058 6272 -13996
rect 7678 -14058 7712 -13996
rect 6453 -14130 6469 -14096
rect 6845 -14130 6861 -14096
rect 7089 -14130 7105 -14096
rect 7481 -14130 7497 -14096
rect 6376 -14158 6410 -14142
rect 6376 -14942 6410 -14926
rect 6904 -14158 6938 -14142
rect 6904 -14942 6938 -14926
rect 7012 -14158 7046 -14142
rect 7012 -14942 7046 -14926
rect 7540 -14158 7574 -14142
rect 7540 -14942 7574 -14926
rect 6453 -14988 6469 -14954
rect 6845 -14988 6861 -14954
rect 7089 -14988 7105 -14954
rect 7481 -14988 7497 -14954
rect 6238 -15088 6272 -15026
rect 7678 -15088 7712 -15026
rect 6238 -15122 6334 -15088
rect 7616 -15122 7712 -15088
rect 7838 -13470 7934 -13436
rect 9216 -13470 9312 -13436
rect 7838 -13532 7872 -13470
rect 9278 -13532 9312 -13470
rect 8053 -13604 8069 -13570
rect 8445 -13604 8461 -13570
rect 8689 -13604 8705 -13570
rect 9081 -13604 9097 -13570
rect 7976 -13632 8010 -13616
rect 7976 -13816 8010 -13800
rect 8504 -13632 8538 -13616
rect 8504 -13816 8538 -13800
rect 8612 -13632 8646 -13616
rect 8612 -13816 8646 -13800
rect 9140 -13632 9174 -13616
rect 9140 -13816 9174 -13800
rect 8053 -13862 8069 -13828
rect 8445 -13862 8461 -13828
rect 8689 -13862 8705 -13828
rect 9081 -13862 9097 -13828
rect 7838 -13962 7872 -13900
rect 9278 -13962 9312 -13900
rect 7838 -13996 7934 -13962
rect 9216 -13996 9312 -13962
rect 7838 -14058 7872 -13996
rect 9278 -14058 9312 -13996
rect 8053 -14130 8069 -14096
rect 8445 -14130 8461 -14096
rect 8689 -14130 8705 -14096
rect 9081 -14130 9097 -14096
rect 7976 -14158 8010 -14142
rect 7976 -14942 8010 -14926
rect 8504 -14158 8538 -14142
rect 8504 -14942 8538 -14926
rect 8612 -14158 8646 -14142
rect 8612 -14942 8646 -14926
rect 9140 -14158 9174 -14142
rect 9140 -14942 9174 -14926
rect 8053 -14988 8069 -14954
rect 8445 -14988 8461 -14954
rect 8689 -14988 8705 -14954
rect 9081 -14988 9097 -14954
rect 7838 -15088 7872 -15026
rect 9278 -15088 9312 -15026
rect 7838 -15122 7934 -15088
rect 9216 -15122 9312 -15088
rect 9438 -13470 9534 -13436
rect 10816 -13470 10912 -13436
rect 9438 -13532 9472 -13470
rect 10878 -13532 10912 -13470
rect 9653 -13604 9669 -13570
rect 10045 -13604 10061 -13570
rect 10289 -13604 10305 -13570
rect 10681 -13604 10697 -13570
rect 9576 -13632 9610 -13616
rect 9576 -13816 9610 -13800
rect 10104 -13632 10138 -13616
rect 10104 -13816 10138 -13800
rect 10212 -13632 10246 -13616
rect 10212 -13816 10246 -13800
rect 10740 -13632 10774 -13616
rect 10740 -13816 10774 -13800
rect 9653 -13862 9669 -13828
rect 10045 -13862 10061 -13828
rect 10289 -13862 10305 -13828
rect 10681 -13862 10697 -13828
rect 9438 -13962 9472 -13900
rect 10878 -13962 10912 -13900
rect 9438 -13996 9534 -13962
rect 10816 -13996 10912 -13962
rect 9438 -14058 9472 -13996
rect 10878 -14058 10912 -13996
rect 9653 -14130 9669 -14096
rect 10045 -14130 10061 -14096
rect 10289 -14130 10305 -14096
rect 10681 -14130 10697 -14096
rect 9576 -14158 9610 -14142
rect 9576 -14942 9610 -14926
rect 10104 -14158 10138 -14142
rect 10104 -14942 10138 -14926
rect 10212 -14158 10246 -14142
rect 10212 -14942 10246 -14926
rect 10740 -14158 10774 -14142
rect 10740 -14942 10774 -14926
rect 9653 -14988 9669 -14954
rect 10045 -14988 10061 -14954
rect 10289 -14988 10305 -14954
rect 10681 -14988 10697 -14954
rect 9438 -15088 9472 -15026
rect 10878 -15088 10912 -15026
rect 9438 -15122 9534 -15088
rect 10816 -15122 10912 -15088
rect 11038 -13470 11134 -13436
rect 12416 -13470 12512 -13436
rect 11038 -13532 11072 -13470
rect 12478 -13532 12512 -13470
rect 11253 -13604 11269 -13570
rect 11645 -13604 11661 -13570
rect 11889 -13604 11905 -13570
rect 12281 -13604 12297 -13570
rect 11176 -13632 11210 -13616
rect 11176 -13816 11210 -13800
rect 11704 -13632 11738 -13616
rect 11704 -13816 11738 -13800
rect 11812 -13632 11846 -13616
rect 11812 -13816 11846 -13800
rect 12340 -13632 12374 -13616
rect 12340 -13816 12374 -13800
rect 11253 -13862 11269 -13828
rect 11645 -13862 11661 -13828
rect 11889 -13862 11905 -13828
rect 12281 -13862 12297 -13828
rect 11038 -13962 11072 -13900
rect 12478 -13962 12512 -13900
rect 11038 -13996 11134 -13962
rect 12416 -13996 12512 -13962
rect 11038 -14058 11072 -13996
rect 12478 -14058 12512 -13996
rect 11253 -14130 11269 -14096
rect 11645 -14130 11661 -14096
rect 11889 -14130 11905 -14096
rect 12281 -14130 12297 -14096
rect 11176 -14158 11210 -14142
rect 11176 -14942 11210 -14926
rect 11704 -14158 11738 -14142
rect 11704 -14942 11738 -14926
rect 11812 -14158 11846 -14142
rect 11812 -14942 11846 -14926
rect 12340 -14158 12374 -14142
rect 12340 -14942 12374 -14926
rect 11253 -14988 11269 -14954
rect 11645 -14988 11661 -14954
rect 11889 -14988 11905 -14954
rect 12281 -14988 12297 -14954
rect 11038 -15088 11072 -15026
rect 12478 -15088 12512 -15026
rect 11038 -15122 11134 -15088
rect 12416 -15122 12512 -15088
rect 12638 -13470 12734 -13436
rect 14016 -13470 14112 -13436
rect 12638 -13532 12672 -13470
rect 14078 -13532 14112 -13470
rect 12853 -13604 12869 -13570
rect 13245 -13604 13261 -13570
rect 13489 -13604 13505 -13570
rect 13881 -13604 13897 -13570
rect 12776 -13632 12810 -13616
rect 12776 -13816 12810 -13800
rect 13304 -13632 13338 -13616
rect 13304 -13816 13338 -13800
rect 13412 -13632 13446 -13616
rect 13412 -13816 13446 -13800
rect 13940 -13632 13974 -13616
rect 13940 -13816 13974 -13800
rect 12853 -13862 12869 -13828
rect 13245 -13862 13261 -13828
rect 13489 -13862 13505 -13828
rect 13881 -13862 13897 -13828
rect 12638 -13962 12672 -13900
rect 14078 -13962 14112 -13900
rect 12638 -13996 12734 -13962
rect 14016 -13996 14112 -13962
rect 12638 -14058 12672 -13996
rect 14078 -14058 14112 -13996
rect 12853 -14130 12869 -14096
rect 13245 -14130 13261 -14096
rect 13489 -14130 13505 -14096
rect 13881 -14130 13897 -14096
rect 12776 -14158 12810 -14142
rect 12776 -14942 12810 -14926
rect 13304 -14158 13338 -14142
rect 13304 -14942 13338 -14926
rect 13412 -14158 13446 -14142
rect 13412 -14942 13446 -14926
rect 13940 -14158 13974 -14142
rect 13940 -14942 13974 -14926
rect 12853 -14988 12869 -14954
rect 13245 -14988 13261 -14954
rect 13489 -14988 13505 -14954
rect 13881 -14988 13897 -14954
rect 12638 -15088 12672 -15026
rect 14078 -15088 14112 -15026
rect 12638 -15122 12734 -15088
rect 14016 -15122 14112 -15088
rect 14238 -13470 14334 -13436
rect 15616 -13470 15712 -13436
rect 14238 -13532 14272 -13470
rect 15678 -13532 15712 -13470
rect 14453 -13604 14469 -13570
rect 14845 -13604 14861 -13570
rect 15089 -13604 15105 -13570
rect 15481 -13604 15497 -13570
rect 14376 -13632 14410 -13616
rect 14376 -13816 14410 -13800
rect 14904 -13632 14938 -13616
rect 14904 -13816 14938 -13800
rect 15012 -13632 15046 -13616
rect 15012 -13816 15046 -13800
rect 15540 -13632 15574 -13616
rect 15540 -13816 15574 -13800
rect 14453 -13862 14469 -13828
rect 14845 -13862 14861 -13828
rect 15089 -13862 15105 -13828
rect 15481 -13862 15497 -13828
rect 14238 -13962 14272 -13900
rect 15678 -13962 15712 -13900
rect 14238 -13996 14334 -13962
rect 15616 -13996 15712 -13962
rect 14238 -14058 14272 -13996
rect 15678 -14058 15712 -13996
rect 14453 -14130 14469 -14096
rect 14845 -14130 14861 -14096
rect 15089 -14130 15105 -14096
rect 15481 -14130 15497 -14096
rect 14376 -14158 14410 -14142
rect 14376 -14942 14410 -14926
rect 14904 -14158 14938 -14142
rect 14904 -14942 14938 -14926
rect 15012 -14158 15046 -14142
rect 15012 -14942 15046 -14926
rect 15540 -14158 15574 -14142
rect 15540 -14942 15574 -14926
rect 14453 -14988 14469 -14954
rect 14845 -14988 14861 -14954
rect 15089 -14988 15105 -14954
rect 15481 -14988 15497 -14954
rect 14238 -15088 14272 -15026
rect 15678 -15088 15712 -15026
rect 14238 -15122 14334 -15088
rect 15616 -15122 15712 -15088
rect 15838 -13470 15934 -13436
rect 17216 -13470 17312 -13436
rect 15838 -13532 15872 -13470
rect 17278 -13532 17312 -13470
rect 16053 -13604 16069 -13570
rect 16445 -13604 16461 -13570
rect 16689 -13604 16705 -13570
rect 17081 -13604 17097 -13570
rect 15976 -13632 16010 -13616
rect 15976 -13816 16010 -13800
rect 16504 -13632 16538 -13616
rect 16504 -13816 16538 -13800
rect 16612 -13632 16646 -13616
rect 16612 -13816 16646 -13800
rect 17140 -13632 17174 -13616
rect 17140 -13816 17174 -13800
rect 16053 -13862 16069 -13828
rect 16445 -13862 16461 -13828
rect 16689 -13862 16705 -13828
rect 17081 -13862 17097 -13828
rect 15838 -13962 15872 -13900
rect 17278 -13962 17312 -13900
rect 15838 -13996 15934 -13962
rect 17216 -13996 17312 -13962
rect 15838 -14058 15872 -13996
rect 17278 -14058 17312 -13996
rect 16053 -14130 16069 -14096
rect 16445 -14130 16461 -14096
rect 16689 -14130 16705 -14096
rect 17081 -14130 17097 -14096
rect 15976 -14158 16010 -14142
rect 15976 -14942 16010 -14926
rect 16504 -14158 16538 -14142
rect 16504 -14942 16538 -14926
rect 16612 -14158 16646 -14142
rect 16612 -14942 16646 -14926
rect 17140 -14158 17174 -14142
rect 17140 -14942 17174 -14926
rect 16053 -14988 16069 -14954
rect 16445 -14988 16461 -14954
rect 16689 -14988 16705 -14954
rect 17081 -14988 17097 -14954
rect 15838 -15088 15872 -15026
rect 17278 -15088 17312 -15026
rect 15838 -15122 15934 -15088
rect 17216 -15122 17312 -15088
rect 17438 -13470 17534 -13436
rect 18816 -13470 18912 -13436
rect 17438 -13532 17472 -13470
rect 18878 -13532 18912 -13470
rect 17653 -13604 17669 -13570
rect 18045 -13604 18061 -13570
rect 18289 -13604 18305 -13570
rect 18681 -13604 18697 -13570
rect 17576 -13632 17610 -13616
rect 17576 -13816 17610 -13800
rect 18104 -13632 18138 -13616
rect 18104 -13816 18138 -13800
rect 18212 -13632 18246 -13616
rect 18212 -13816 18246 -13800
rect 18740 -13632 18774 -13616
rect 18740 -13816 18774 -13800
rect 17653 -13862 17669 -13828
rect 18045 -13862 18061 -13828
rect 18289 -13862 18305 -13828
rect 18681 -13862 18697 -13828
rect 17438 -13962 17472 -13900
rect 18878 -13962 18912 -13900
rect 17438 -13996 17534 -13962
rect 18816 -13996 18912 -13962
rect 17438 -14058 17472 -13996
rect 18878 -14058 18912 -13996
rect 17653 -14130 17669 -14096
rect 18045 -14130 18061 -14096
rect 18289 -14130 18305 -14096
rect 18681 -14130 18697 -14096
rect 17576 -14158 17610 -14142
rect 17576 -14942 17610 -14926
rect 18104 -14158 18138 -14142
rect 18104 -14942 18138 -14926
rect 18212 -14158 18246 -14142
rect 18212 -14942 18246 -14926
rect 18740 -14158 18774 -14142
rect 18740 -14942 18774 -14926
rect 17653 -14988 17669 -14954
rect 18045 -14988 18061 -14954
rect 18289 -14988 18305 -14954
rect 18681 -14988 18697 -14954
rect 17438 -15088 17472 -15026
rect 18878 -15088 18912 -15026
rect 17438 -15122 17534 -15088
rect 18816 -15122 18912 -15088
rect 19038 -13470 19134 -13436
rect 20416 -13470 20512 -13436
rect 19038 -13532 19072 -13470
rect 20478 -13532 20512 -13470
rect 19253 -13604 19269 -13570
rect 19645 -13604 19661 -13570
rect 19889 -13604 19905 -13570
rect 20281 -13604 20297 -13570
rect 19176 -13632 19210 -13616
rect 19176 -13816 19210 -13800
rect 19704 -13632 19738 -13616
rect 19704 -13816 19738 -13800
rect 19812 -13632 19846 -13616
rect 19812 -13816 19846 -13800
rect 20340 -13632 20374 -13616
rect 20340 -13816 20374 -13800
rect 19253 -13862 19269 -13828
rect 19645 -13862 19661 -13828
rect 19889 -13862 19905 -13828
rect 20281 -13862 20297 -13828
rect 19038 -13962 19072 -13900
rect 20478 -13962 20512 -13900
rect 19038 -13996 19134 -13962
rect 20416 -13996 20512 -13962
rect 19038 -14058 19072 -13996
rect 20478 -14058 20512 -13996
rect 19253 -14130 19269 -14096
rect 19645 -14130 19661 -14096
rect 19889 -14130 19905 -14096
rect 20281 -14130 20297 -14096
rect 19176 -14158 19210 -14142
rect 19176 -14942 19210 -14926
rect 19704 -14158 19738 -14142
rect 19704 -14942 19738 -14926
rect 19812 -14158 19846 -14142
rect 19812 -14942 19846 -14926
rect 20340 -14158 20374 -14142
rect 20340 -14942 20374 -14926
rect 19253 -14988 19269 -14954
rect 19645 -14988 19661 -14954
rect 19889 -14988 19905 -14954
rect 20281 -14988 20297 -14954
rect 19038 -15088 19072 -15026
rect 20478 -15088 20512 -15026
rect 19038 -15122 19134 -15088
rect 20416 -15122 20512 -15088
rect 20638 -13470 20734 -13436
rect 22016 -13470 22112 -13436
rect 20638 -13532 20672 -13470
rect 22078 -13532 22112 -13470
rect 20853 -13604 20869 -13570
rect 21245 -13604 21261 -13570
rect 21489 -13604 21505 -13570
rect 21881 -13604 21897 -13570
rect 20776 -13632 20810 -13616
rect 20776 -13816 20810 -13800
rect 21304 -13632 21338 -13616
rect 21304 -13816 21338 -13800
rect 21412 -13632 21446 -13616
rect 21412 -13816 21446 -13800
rect 21940 -13632 21974 -13616
rect 21940 -13816 21974 -13800
rect 20853 -13862 20869 -13828
rect 21245 -13862 21261 -13828
rect 21489 -13862 21505 -13828
rect 21881 -13862 21897 -13828
rect 20638 -13962 20672 -13900
rect 22078 -13962 22112 -13900
rect 20638 -13996 20734 -13962
rect 22016 -13996 22112 -13962
rect 20638 -14058 20672 -13996
rect 22078 -14058 22112 -13996
rect 20853 -14130 20869 -14096
rect 21245 -14130 21261 -14096
rect 21489 -14130 21505 -14096
rect 21881 -14130 21897 -14096
rect 20776 -14158 20810 -14142
rect 20776 -14942 20810 -14926
rect 21304 -14158 21338 -14142
rect 21304 -14942 21338 -14926
rect 21412 -14158 21446 -14142
rect 21412 -14942 21446 -14926
rect 21940 -14158 21974 -14142
rect 21940 -14942 21974 -14926
rect 20853 -14988 20869 -14954
rect 21245 -14988 21261 -14954
rect 21489 -14988 21505 -14954
rect 21881 -14988 21897 -14954
rect 20638 -15088 20672 -15026
rect 22078 -15088 22112 -15026
rect 20638 -15122 20734 -15088
rect 22016 -15122 22112 -15088
rect 22238 -13470 22334 -13436
rect 23616 -13470 23712 -13436
rect 22238 -13532 22272 -13470
rect 23678 -13532 23712 -13470
rect 22453 -13604 22469 -13570
rect 22845 -13604 22861 -13570
rect 23089 -13604 23105 -13570
rect 23481 -13604 23497 -13570
rect 22376 -13632 22410 -13616
rect 22376 -13816 22410 -13800
rect 22904 -13632 22938 -13616
rect 22904 -13816 22938 -13800
rect 23012 -13632 23046 -13616
rect 23012 -13816 23046 -13800
rect 23540 -13632 23574 -13616
rect 23540 -13816 23574 -13800
rect 22453 -13862 22469 -13828
rect 22845 -13862 22861 -13828
rect 23089 -13862 23105 -13828
rect 23481 -13862 23497 -13828
rect 22238 -13962 22272 -13900
rect 23678 -13962 23712 -13900
rect 22238 -13996 22334 -13962
rect 23616 -13996 23712 -13962
rect 22238 -14058 22272 -13996
rect 23678 -14058 23712 -13996
rect 22453 -14130 22469 -14096
rect 22845 -14130 22861 -14096
rect 23089 -14130 23105 -14096
rect 23481 -14130 23497 -14096
rect 22376 -14158 22410 -14142
rect 22376 -14942 22410 -14926
rect 22904 -14158 22938 -14142
rect 22904 -14942 22938 -14926
rect 23012 -14158 23046 -14142
rect 23012 -14942 23046 -14926
rect 23540 -14158 23574 -14142
rect 23540 -14942 23574 -14926
rect 22453 -14988 22469 -14954
rect 22845 -14988 22861 -14954
rect 23089 -14988 23105 -14954
rect 23481 -14988 23497 -14954
rect 22238 -15088 22272 -15026
rect 23678 -15088 23712 -15026
rect 22238 -15122 22334 -15088
rect 23616 -15122 23712 -15088
rect 23838 -13470 23934 -13436
rect 25216 -13470 25312 -13436
rect 23838 -13532 23872 -13470
rect 25278 -13532 25312 -13470
rect 24053 -13604 24069 -13570
rect 24445 -13604 24461 -13570
rect 24689 -13604 24705 -13570
rect 25081 -13604 25097 -13570
rect 23976 -13632 24010 -13616
rect 23976 -13816 24010 -13800
rect 24504 -13632 24538 -13616
rect 24504 -13816 24538 -13800
rect 24612 -13632 24646 -13616
rect 24612 -13816 24646 -13800
rect 25140 -13632 25174 -13616
rect 25140 -13816 25174 -13800
rect 24053 -13862 24069 -13828
rect 24445 -13862 24461 -13828
rect 24689 -13862 24705 -13828
rect 25081 -13862 25097 -13828
rect 23838 -13962 23872 -13900
rect 25278 -13962 25312 -13900
rect 23838 -13996 23934 -13962
rect 25216 -13996 25312 -13962
rect 23838 -14058 23872 -13996
rect 25278 -14058 25312 -13996
rect 24053 -14130 24069 -14096
rect 24445 -14130 24461 -14096
rect 24689 -14130 24705 -14096
rect 25081 -14130 25097 -14096
rect 23976 -14158 24010 -14142
rect 23976 -14942 24010 -14926
rect 24504 -14158 24538 -14142
rect 24504 -14942 24538 -14926
rect 24612 -14158 24646 -14142
rect 24612 -14942 24646 -14926
rect 25140 -14158 25174 -14142
rect 25140 -14942 25174 -14926
rect 24053 -14988 24069 -14954
rect 24445 -14988 24461 -14954
rect 24689 -14988 24705 -14954
rect 25081 -14988 25097 -14954
rect 23838 -15088 23872 -15026
rect 25278 -15088 25312 -15026
rect 23838 -15122 23934 -15088
rect 25216 -15122 25312 -15088
rect 25438 -13470 25534 -13436
rect 26816 -13470 26912 -13436
rect 25438 -13532 25472 -13470
rect 26878 -13532 26912 -13470
rect 25653 -13604 25669 -13570
rect 26045 -13604 26061 -13570
rect 26289 -13604 26305 -13570
rect 26681 -13604 26697 -13570
rect 25576 -13632 25610 -13616
rect 25576 -13816 25610 -13800
rect 26104 -13632 26138 -13616
rect 26104 -13816 26138 -13800
rect 26212 -13632 26246 -13616
rect 26212 -13816 26246 -13800
rect 26740 -13632 26774 -13616
rect 26740 -13816 26774 -13800
rect 25653 -13862 25669 -13828
rect 26045 -13862 26061 -13828
rect 26289 -13862 26305 -13828
rect 26681 -13862 26697 -13828
rect 25438 -13962 25472 -13900
rect 26878 -13962 26912 -13900
rect 25438 -13996 25534 -13962
rect 26816 -13996 26912 -13962
rect 25438 -14058 25472 -13996
rect 26878 -14058 26912 -13996
rect 25653 -14130 25669 -14096
rect 26045 -14130 26061 -14096
rect 26289 -14130 26305 -14096
rect 26681 -14130 26697 -14096
rect 25576 -14158 25610 -14142
rect 25576 -14942 25610 -14926
rect 26104 -14158 26138 -14142
rect 26104 -14942 26138 -14926
rect 26212 -14158 26246 -14142
rect 26212 -14942 26246 -14926
rect 26740 -14158 26774 -14142
rect 26740 -14942 26774 -14926
rect 25653 -14988 25669 -14954
rect 26045 -14988 26061 -14954
rect 26289 -14988 26305 -14954
rect 26681 -14988 26697 -14954
rect 25438 -15088 25472 -15026
rect 26878 -15088 26912 -15026
rect 25438 -15122 25534 -15088
rect 26816 -15122 26912 -15088
rect 27038 -13470 27134 -13436
rect 28416 -13470 28512 -13436
rect 27038 -13532 27072 -13470
rect 28478 -13532 28512 -13470
rect 27253 -13604 27269 -13570
rect 27645 -13604 27661 -13570
rect 27889 -13604 27905 -13570
rect 28281 -13604 28297 -13570
rect 27176 -13632 27210 -13616
rect 27176 -13816 27210 -13800
rect 27704 -13632 27738 -13616
rect 27704 -13816 27738 -13800
rect 27812 -13632 27846 -13616
rect 27812 -13816 27846 -13800
rect 28340 -13632 28374 -13616
rect 28340 -13816 28374 -13800
rect 27253 -13862 27269 -13828
rect 27645 -13862 27661 -13828
rect 27889 -13862 27905 -13828
rect 28281 -13862 28297 -13828
rect 27038 -13962 27072 -13900
rect 28478 -13962 28512 -13900
rect 27038 -13996 27134 -13962
rect 28416 -13996 28512 -13962
rect 27038 -14058 27072 -13996
rect 28478 -14058 28512 -13996
rect 27253 -14130 27269 -14096
rect 27645 -14130 27661 -14096
rect 27889 -14130 27905 -14096
rect 28281 -14130 28297 -14096
rect 27176 -14158 27210 -14142
rect 27176 -14942 27210 -14926
rect 27704 -14158 27738 -14142
rect 27704 -14942 27738 -14926
rect 27812 -14158 27846 -14142
rect 27812 -14942 27846 -14926
rect 28340 -14158 28374 -14142
rect 28340 -14942 28374 -14926
rect 27253 -14988 27269 -14954
rect 27645 -14988 27661 -14954
rect 27889 -14988 27905 -14954
rect 28281 -14988 28297 -14954
rect 27038 -15088 27072 -15026
rect 28478 -15088 28512 -15026
rect 27038 -15122 27134 -15088
rect 28416 -15122 28512 -15088
rect 28638 -13470 28734 -13436
rect 30016 -13470 30112 -13436
rect 28638 -13532 28672 -13470
rect 30078 -13532 30112 -13470
rect 28853 -13604 28869 -13570
rect 29245 -13604 29261 -13570
rect 29489 -13604 29505 -13570
rect 29881 -13604 29897 -13570
rect 28776 -13632 28810 -13616
rect 28776 -13816 28810 -13800
rect 29304 -13632 29338 -13616
rect 29304 -13816 29338 -13800
rect 29412 -13632 29446 -13616
rect 29412 -13816 29446 -13800
rect 29940 -13632 29974 -13616
rect 29940 -13816 29974 -13800
rect 28853 -13862 28869 -13828
rect 29245 -13862 29261 -13828
rect 29489 -13862 29505 -13828
rect 29881 -13862 29897 -13828
rect 28638 -13962 28672 -13900
rect 30078 -13962 30112 -13900
rect 28638 -13996 28734 -13962
rect 30016 -13996 30112 -13962
rect 28638 -14058 28672 -13996
rect 30078 -14058 30112 -13996
rect 28853 -14130 28869 -14096
rect 29245 -14130 29261 -14096
rect 29489 -14130 29505 -14096
rect 29881 -14130 29897 -14096
rect 28776 -14158 28810 -14142
rect 28776 -14942 28810 -14926
rect 29304 -14158 29338 -14142
rect 29304 -14942 29338 -14926
rect 29412 -14158 29446 -14142
rect 29412 -14942 29446 -14926
rect 29940 -14158 29974 -14142
rect 29940 -14942 29974 -14926
rect 28853 -14988 28869 -14954
rect 29245 -14988 29261 -14954
rect 29489 -14988 29505 -14954
rect 29881 -14988 29897 -14954
rect 28638 -15088 28672 -15026
rect 30078 -15088 30112 -15026
rect 28638 -15122 28734 -15088
rect 30016 -15122 30112 -15088
rect 30238 -13470 30334 -13436
rect 31616 -13470 31712 -13436
rect 30238 -13532 30272 -13470
rect 31678 -13532 31712 -13470
rect 30453 -13604 30469 -13570
rect 30845 -13604 30861 -13570
rect 31089 -13604 31105 -13570
rect 31481 -13604 31497 -13570
rect 30376 -13632 30410 -13616
rect 30376 -13816 30410 -13800
rect 30904 -13632 30938 -13616
rect 30904 -13816 30938 -13800
rect 31012 -13632 31046 -13616
rect 31012 -13816 31046 -13800
rect 31540 -13632 31574 -13616
rect 31540 -13816 31574 -13800
rect 30453 -13862 30469 -13828
rect 30845 -13862 30861 -13828
rect 31089 -13862 31105 -13828
rect 31481 -13862 31497 -13828
rect 30238 -13962 30272 -13900
rect 31678 -13962 31712 -13900
rect 30238 -13996 30334 -13962
rect 31616 -13996 31712 -13962
rect 30238 -14058 30272 -13996
rect 31678 -14058 31712 -13996
rect 30453 -14130 30469 -14096
rect 30845 -14130 30861 -14096
rect 31089 -14130 31105 -14096
rect 31481 -14130 31497 -14096
rect 30376 -14158 30410 -14142
rect 30376 -14942 30410 -14926
rect 30904 -14158 30938 -14142
rect 30904 -14942 30938 -14926
rect 31012 -14158 31046 -14142
rect 31012 -14942 31046 -14926
rect 31540 -14158 31574 -14142
rect 31540 -14942 31574 -14926
rect 30453 -14988 30469 -14954
rect 30845 -14988 30861 -14954
rect 31089 -14988 31105 -14954
rect 31481 -14988 31497 -14954
rect 30238 -15088 30272 -15026
rect 31678 -15088 31712 -15026
rect 30238 -15122 30334 -15088
rect 31616 -15122 31712 -15088
rect 31838 -13470 31934 -13436
rect 33216 -13470 33312 -13436
rect 31838 -13532 31872 -13470
rect 33278 -13532 33312 -13470
rect 32053 -13604 32069 -13570
rect 32445 -13604 32461 -13570
rect 32689 -13604 32705 -13570
rect 33081 -13604 33097 -13570
rect 31976 -13632 32010 -13616
rect 31976 -13816 32010 -13800
rect 32504 -13632 32538 -13616
rect 32504 -13816 32538 -13800
rect 32612 -13632 32646 -13616
rect 32612 -13816 32646 -13800
rect 33140 -13632 33174 -13616
rect 33140 -13816 33174 -13800
rect 32053 -13862 32069 -13828
rect 32445 -13862 32461 -13828
rect 32689 -13862 32705 -13828
rect 33081 -13862 33097 -13828
rect 31838 -13962 31872 -13900
rect 33278 -13962 33312 -13900
rect 31838 -13996 31934 -13962
rect 33216 -13996 33312 -13962
rect 31838 -14058 31872 -13996
rect 33278 -14058 33312 -13996
rect 32053 -14130 32069 -14096
rect 32445 -14130 32461 -14096
rect 32689 -14130 32705 -14096
rect 33081 -14130 33097 -14096
rect 31976 -14158 32010 -14142
rect 31976 -14942 32010 -14926
rect 32504 -14158 32538 -14142
rect 32504 -14942 32538 -14926
rect 32612 -14158 32646 -14142
rect 32612 -14942 32646 -14926
rect 33140 -14158 33174 -14142
rect 33140 -14942 33174 -14926
rect 32053 -14988 32069 -14954
rect 32445 -14988 32461 -14954
rect 32689 -14988 32705 -14954
rect 33081 -14988 33097 -14954
rect 31838 -15088 31872 -15026
rect 33278 -15088 33312 -15026
rect 31838 -15122 31934 -15088
rect 33216 -15122 33312 -15088
rect 33438 -13470 33534 -13436
rect 34816 -13470 34912 -13436
rect 33438 -13532 33472 -13470
rect 34878 -13532 34912 -13470
rect 33653 -13604 33669 -13570
rect 34045 -13604 34061 -13570
rect 34289 -13604 34305 -13570
rect 34681 -13604 34697 -13570
rect 33576 -13632 33610 -13616
rect 33576 -13816 33610 -13800
rect 34104 -13632 34138 -13616
rect 34104 -13816 34138 -13800
rect 34212 -13632 34246 -13616
rect 34212 -13816 34246 -13800
rect 34740 -13632 34774 -13616
rect 34740 -13816 34774 -13800
rect 33653 -13862 33669 -13828
rect 34045 -13862 34061 -13828
rect 34289 -13862 34305 -13828
rect 34681 -13862 34697 -13828
rect 33438 -13962 33472 -13900
rect 34878 -13962 34912 -13900
rect 33438 -13996 33534 -13962
rect 34816 -13996 34912 -13962
rect 33438 -14058 33472 -13996
rect 34878 -14058 34912 -13996
rect 33653 -14130 33669 -14096
rect 34045 -14130 34061 -14096
rect 34289 -14130 34305 -14096
rect 34681 -14130 34697 -14096
rect 33576 -14158 33610 -14142
rect 33576 -14942 33610 -14926
rect 34104 -14158 34138 -14142
rect 34104 -14942 34138 -14926
rect 34212 -14158 34246 -14142
rect 34212 -14942 34246 -14926
rect 34740 -14158 34774 -14142
rect 34740 -14942 34774 -14926
rect 33653 -14988 33669 -14954
rect 34045 -14988 34061 -14954
rect 34289 -14988 34305 -14954
rect 34681 -14988 34697 -14954
rect 33438 -15088 33472 -15026
rect 34878 -15088 34912 -15026
rect 33438 -15122 33534 -15088
rect 34816 -15122 34912 -15088
rect 35038 -13470 35134 -13436
rect 36416 -13470 36734 -13436
rect 38016 -13470 38112 -13436
rect 35038 -13532 35072 -13470
rect 36478 -13532 38112 -13470
rect 35253 -13604 35269 -13570
rect 35645 -13604 35661 -13570
rect 35889 -13604 35905 -13570
rect 36281 -13604 36297 -13570
rect 35176 -13632 35210 -13616
rect 35176 -13816 35210 -13800
rect 35704 -13632 35738 -13616
rect 35704 -13816 35738 -13800
rect 35812 -13632 35846 -13616
rect 35812 -13816 35846 -13800
rect 36340 -13632 36374 -13616
rect 36340 -13816 36374 -13800
rect 35253 -13862 35269 -13828
rect 35645 -13862 35661 -13828
rect 35889 -13862 35905 -13828
rect 36281 -13862 36297 -13828
rect 35038 -13962 35072 -13900
rect 36512 -13900 36638 -13532
rect 36672 -13570 38078 -13532
rect 36672 -13604 36869 -13570
rect 37245 -13604 37505 -13570
rect 37881 -13604 38078 -13570
rect 36672 -13632 38078 -13604
rect 36672 -13800 36776 -13632
rect 36810 -13800 37304 -13632
rect 37338 -13800 37412 -13632
rect 37446 -13800 37940 -13632
rect 37974 -13800 38078 -13632
rect 36672 -13828 38078 -13800
rect 36672 -13862 36869 -13828
rect 37245 -13862 37505 -13828
rect 37881 -13862 38078 -13828
rect 36672 -13900 38078 -13862
rect 36478 -13962 38112 -13900
rect 35038 -13996 35134 -13962
rect 36416 -13996 36734 -13962
rect 38016 -13996 38112 -13962
rect 35038 -14058 35072 -13996
rect 36478 -14058 38112 -13996
rect 35253 -14130 35269 -14096
rect 35645 -14130 35661 -14096
rect 35889 -14130 35905 -14096
rect 36281 -14130 36297 -14096
rect 35176 -14158 35210 -14142
rect 35176 -14942 35210 -14926
rect 35704 -14158 35738 -14142
rect 35704 -14942 35738 -14926
rect 35812 -14158 35846 -14142
rect 35812 -14942 35846 -14926
rect 36340 -14158 36374 -14142
rect 36340 -14942 36374 -14926
rect 35253 -14988 35269 -14954
rect 35645 -14988 35661 -14954
rect 35889 -14988 35905 -14954
rect 36281 -14988 36297 -14954
rect 35038 -15088 35072 -15026
rect 36512 -15026 36638 -14058
rect 36672 -14096 38078 -14058
rect 36672 -14130 36869 -14096
rect 37245 -14130 37505 -14096
rect 37881 -14130 38078 -14096
rect 36672 -14158 38078 -14130
rect 36672 -14926 36776 -14158
rect 36810 -14926 37304 -14158
rect 37338 -14926 37412 -14158
rect 37446 -14926 37940 -14158
rect 37974 -14926 38078 -14158
rect 36672 -14954 38078 -14926
rect 36672 -14988 36869 -14954
rect 37245 -14988 37505 -14954
rect 37881 -14988 38078 -14954
rect 36672 -15026 38078 -14988
rect 36478 -15088 38112 -15026
rect 35038 -15122 35134 -15088
rect 36416 -15122 36734 -15088
rect 38016 -15122 38112 -15088
rect -140 -15236 1460 -15122
rect 36500 -15236 38100 -15122
rect -162 -15270 -66 -15236
rect 1216 -15270 1534 -15236
rect 2816 -15270 2912 -15236
rect -162 -15332 1472 -15270
rect -128 -15370 1278 -15332
rect -128 -15404 69 -15370
rect 445 -15404 705 -15370
rect 1081 -15404 1278 -15370
rect -128 -15432 1278 -15404
rect -128 -15600 -24 -15432
rect 10 -15600 504 -15432
rect 538 -15600 612 -15432
rect 646 -15600 1140 -15432
rect 1174 -15600 1278 -15432
rect -128 -15628 1278 -15600
rect -128 -15662 69 -15628
rect 445 -15662 705 -15628
rect 1081 -15662 1278 -15628
rect -128 -15700 1278 -15662
rect 1312 -15700 1438 -15332
rect 2878 -15332 2912 -15270
rect 1653 -15404 1669 -15370
rect 2045 -15404 2061 -15370
rect 2289 -15404 2305 -15370
rect 2681 -15404 2697 -15370
rect 1576 -15432 1610 -15416
rect 1576 -15616 1610 -15600
rect 2104 -15432 2138 -15416
rect 2104 -15616 2138 -15600
rect 2212 -15432 2246 -15416
rect 2212 -15616 2246 -15600
rect 2740 -15432 2774 -15416
rect 2740 -15616 2774 -15600
rect 1653 -15662 1669 -15628
rect 2045 -15662 2061 -15628
rect 2289 -15662 2305 -15628
rect 2681 -15662 2697 -15628
rect -162 -15762 1472 -15700
rect 2878 -15762 2912 -15700
rect -162 -15796 -66 -15762
rect 1216 -15796 1534 -15762
rect 2816 -15796 2912 -15762
rect -162 -15858 1472 -15796
rect -128 -15896 1278 -15858
rect -128 -15930 69 -15896
rect 445 -15930 705 -15896
rect 1081 -15930 1278 -15896
rect -128 -15958 1278 -15930
rect -128 -16726 -24 -15958
rect 10 -16726 504 -15958
rect 538 -16726 612 -15958
rect 646 -16726 1140 -15958
rect 1174 -16726 1278 -15958
rect -128 -16754 1278 -16726
rect -128 -16788 69 -16754
rect 445 -16788 705 -16754
rect 1081 -16788 1278 -16754
rect -128 -16826 1278 -16788
rect 1312 -16826 1438 -15858
rect 2878 -15858 2912 -15796
rect 1653 -15930 1669 -15896
rect 2045 -15930 2061 -15896
rect 2289 -15930 2305 -15896
rect 2681 -15930 2697 -15896
rect 1576 -15958 1610 -15942
rect 1576 -16742 1610 -16726
rect 2104 -15958 2138 -15942
rect 2104 -16742 2138 -16726
rect 2212 -15958 2246 -15942
rect 2212 -16742 2246 -16726
rect 2740 -15958 2774 -15942
rect 2740 -16742 2774 -16726
rect 1653 -16788 1669 -16754
rect 2045 -16788 2061 -16754
rect 2289 -16788 2305 -16754
rect 2681 -16788 2697 -16754
rect -162 -16888 1472 -16826
rect 2878 -16888 2912 -16826
rect -162 -16922 -66 -16888
rect 1216 -16922 1534 -16888
rect 2816 -16922 2912 -16888
rect 3038 -15270 3134 -15236
rect 4416 -15270 4512 -15236
rect 3038 -15332 3072 -15270
rect 4478 -15332 4512 -15270
rect 3253 -15404 3269 -15370
rect 3645 -15404 3661 -15370
rect 3889 -15404 3905 -15370
rect 4281 -15404 4297 -15370
rect 3176 -15432 3210 -15416
rect 3176 -15616 3210 -15600
rect 3704 -15432 3738 -15416
rect 3704 -15616 3738 -15600
rect 3812 -15432 3846 -15416
rect 3812 -15616 3846 -15600
rect 4340 -15432 4374 -15416
rect 4340 -15616 4374 -15600
rect 3253 -15662 3269 -15628
rect 3645 -15662 3661 -15628
rect 3889 -15662 3905 -15628
rect 4281 -15662 4297 -15628
rect 3038 -15762 3072 -15700
rect 4478 -15762 4512 -15700
rect 3038 -15796 3134 -15762
rect 4416 -15796 4512 -15762
rect 3038 -15858 3072 -15796
rect 4478 -15858 4512 -15796
rect 3253 -15930 3269 -15896
rect 3645 -15930 3661 -15896
rect 3889 -15930 3905 -15896
rect 4281 -15930 4297 -15896
rect 3176 -15958 3210 -15942
rect 3176 -16742 3210 -16726
rect 3704 -15958 3738 -15942
rect 3704 -16742 3738 -16726
rect 3812 -15958 3846 -15942
rect 3812 -16742 3846 -16726
rect 4340 -15958 4374 -15942
rect 4340 -16742 4374 -16726
rect 3253 -16788 3269 -16754
rect 3645 -16788 3661 -16754
rect 3889 -16788 3905 -16754
rect 4281 -16788 4297 -16754
rect 3038 -16888 3072 -16826
rect 4478 -16888 4512 -16826
rect 3038 -16922 3134 -16888
rect 4416 -16922 4512 -16888
rect 4638 -15270 4734 -15236
rect 6016 -15270 6112 -15236
rect 4638 -15332 4672 -15270
rect 6078 -15332 6112 -15270
rect 4853 -15404 4869 -15370
rect 5245 -15404 5261 -15370
rect 5489 -15404 5505 -15370
rect 5881 -15404 5897 -15370
rect 4776 -15432 4810 -15416
rect 4776 -15616 4810 -15600
rect 5304 -15432 5338 -15416
rect 5304 -15616 5338 -15600
rect 5412 -15432 5446 -15416
rect 5412 -15616 5446 -15600
rect 5940 -15432 5974 -15416
rect 5940 -15616 5974 -15600
rect 4853 -15662 4869 -15628
rect 5245 -15662 5261 -15628
rect 5489 -15662 5505 -15628
rect 5881 -15662 5897 -15628
rect 4638 -15762 4672 -15700
rect 6078 -15762 6112 -15700
rect 4638 -15796 4734 -15762
rect 6016 -15796 6112 -15762
rect 4638 -15858 4672 -15796
rect 6078 -15858 6112 -15796
rect 4853 -15930 4869 -15896
rect 5245 -15930 5261 -15896
rect 5489 -15930 5505 -15896
rect 5881 -15930 5897 -15896
rect 4776 -15958 4810 -15942
rect 4776 -16742 4810 -16726
rect 5304 -15958 5338 -15942
rect 5304 -16742 5338 -16726
rect 5412 -15958 5446 -15942
rect 5412 -16742 5446 -16726
rect 5940 -15958 5974 -15942
rect 5940 -16742 5974 -16726
rect 4853 -16788 4869 -16754
rect 5245 -16788 5261 -16754
rect 5489 -16788 5505 -16754
rect 5881 -16788 5897 -16754
rect 4638 -16888 4672 -16826
rect 6078 -16888 6112 -16826
rect 4638 -16922 4734 -16888
rect 6016 -16922 6112 -16888
rect 6238 -15270 6334 -15236
rect 7616 -15270 7712 -15236
rect 6238 -15332 6272 -15270
rect 7678 -15332 7712 -15270
rect 6453 -15404 6469 -15370
rect 6845 -15404 6861 -15370
rect 7089 -15404 7105 -15370
rect 7481 -15404 7497 -15370
rect 6376 -15432 6410 -15416
rect 6376 -15616 6410 -15600
rect 6904 -15432 6938 -15416
rect 6904 -15616 6938 -15600
rect 7012 -15432 7046 -15416
rect 7012 -15616 7046 -15600
rect 7540 -15432 7574 -15416
rect 7540 -15616 7574 -15600
rect 6453 -15662 6469 -15628
rect 6845 -15662 6861 -15628
rect 7089 -15662 7105 -15628
rect 7481 -15662 7497 -15628
rect 6238 -15762 6272 -15700
rect 7678 -15762 7712 -15700
rect 6238 -15796 6334 -15762
rect 7616 -15796 7712 -15762
rect 6238 -15858 6272 -15796
rect 7678 -15858 7712 -15796
rect 6453 -15930 6469 -15896
rect 6845 -15930 6861 -15896
rect 7089 -15930 7105 -15896
rect 7481 -15930 7497 -15896
rect 6376 -15958 6410 -15942
rect 6376 -16742 6410 -16726
rect 6904 -15958 6938 -15942
rect 6904 -16742 6938 -16726
rect 7012 -15958 7046 -15942
rect 7012 -16742 7046 -16726
rect 7540 -15958 7574 -15942
rect 7540 -16742 7574 -16726
rect 6453 -16788 6469 -16754
rect 6845 -16788 6861 -16754
rect 7089 -16788 7105 -16754
rect 7481 -16788 7497 -16754
rect 6238 -16888 6272 -16826
rect 7678 -16888 7712 -16826
rect 6238 -16922 6334 -16888
rect 7616 -16922 7712 -16888
rect 7838 -15270 7934 -15236
rect 9216 -15270 9312 -15236
rect 7838 -15332 7872 -15270
rect 9278 -15332 9312 -15270
rect 8053 -15404 8069 -15370
rect 8445 -15404 8461 -15370
rect 8689 -15404 8705 -15370
rect 9081 -15404 9097 -15370
rect 7976 -15432 8010 -15416
rect 7976 -15616 8010 -15600
rect 8504 -15432 8538 -15416
rect 8504 -15616 8538 -15600
rect 8612 -15432 8646 -15416
rect 8612 -15616 8646 -15600
rect 9140 -15432 9174 -15416
rect 9140 -15616 9174 -15600
rect 8053 -15662 8069 -15628
rect 8445 -15662 8461 -15628
rect 8689 -15662 8705 -15628
rect 9081 -15662 9097 -15628
rect 7838 -15762 7872 -15700
rect 9278 -15762 9312 -15700
rect 7838 -15796 7934 -15762
rect 9216 -15796 9312 -15762
rect 7838 -15858 7872 -15796
rect 9278 -15858 9312 -15796
rect 8053 -15930 8069 -15896
rect 8445 -15930 8461 -15896
rect 8689 -15930 8705 -15896
rect 9081 -15930 9097 -15896
rect 7976 -15958 8010 -15942
rect 7976 -16742 8010 -16726
rect 8504 -15958 8538 -15942
rect 8504 -16742 8538 -16726
rect 8612 -15958 8646 -15942
rect 8612 -16742 8646 -16726
rect 9140 -15958 9174 -15942
rect 9140 -16742 9174 -16726
rect 8053 -16788 8069 -16754
rect 8445 -16788 8461 -16754
rect 8689 -16788 8705 -16754
rect 9081 -16788 9097 -16754
rect 7838 -16888 7872 -16826
rect 9278 -16888 9312 -16826
rect 7838 -16922 7934 -16888
rect 9216 -16922 9312 -16888
rect 9438 -15270 9534 -15236
rect 10816 -15270 10912 -15236
rect 9438 -15332 9472 -15270
rect 10878 -15332 10912 -15270
rect 9653 -15404 9669 -15370
rect 10045 -15404 10061 -15370
rect 10289 -15404 10305 -15370
rect 10681 -15404 10697 -15370
rect 9576 -15432 9610 -15416
rect 9576 -15616 9610 -15600
rect 10104 -15432 10138 -15416
rect 10104 -15616 10138 -15600
rect 10212 -15432 10246 -15416
rect 10212 -15616 10246 -15600
rect 10740 -15432 10774 -15416
rect 10740 -15616 10774 -15600
rect 9653 -15662 9669 -15628
rect 10045 -15662 10061 -15628
rect 10289 -15662 10305 -15628
rect 10681 -15662 10697 -15628
rect 9438 -15762 9472 -15700
rect 10878 -15762 10912 -15700
rect 9438 -15796 9534 -15762
rect 10816 -15796 10912 -15762
rect 9438 -15858 9472 -15796
rect 10878 -15858 10912 -15796
rect 9653 -15930 9669 -15896
rect 10045 -15930 10061 -15896
rect 10289 -15930 10305 -15896
rect 10681 -15930 10697 -15896
rect 9576 -15958 9610 -15942
rect 9576 -16742 9610 -16726
rect 10104 -15958 10138 -15942
rect 10104 -16742 10138 -16726
rect 10212 -15958 10246 -15942
rect 10212 -16742 10246 -16726
rect 10740 -15958 10774 -15942
rect 10740 -16742 10774 -16726
rect 9653 -16788 9669 -16754
rect 10045 -16788 10061 -16754
rect 10289 -16788 10305 -16754
rect 10681 -16788 10697 -16754
rect 9438 -16888 9472 -16826
rect 10878 -16888 10912 -16826
rect 9438 -16922 9534 -16888
rect 10816 -16922 10912 -16888
rect 11038 -15270 11134 -15236
rect 12416 -15270 12512 -15236
rect 11038 -15332 11072 -15270
rect 12478 -15332 12512 -15270
rect 11253 -15404 11269 -15370
rect 11645 -15404 11661 -15370
rect 11889 -15404 11905 -15370
rect 12281 -15404 12297 -15370
rect 11176 -15432 11210 -15416
rect 11176 -15616 11210 -15600
rect 11704 -15432 11738 -15416
rect 11704 -15616 11738 -15600
rect 11812 -15432 11846 -15416
rect 11812 -15616 11846 -15600
rect 12340 -15432 12374 -15416
rect 12340 -15616 12374 -15600
rect 11253 -15662 11269 -15628
rect 11645 -15662 11661 -15628
rect 11889 -15662 11905 -15628
rect 12281 -15662 12297 -15628
rect 11038 -15762 11072 -15700
rect 12478 -15762 12512 -15700
rect 11038 -15796 11134 -15762
rect 12416 -15796 12512 -15762
rect 11038 -15858 11072 -15796
rect 12478 -15858 12512 -15796
rect 11253 -15930 11269 -15896
rect 11645 -15930 11661 -15896
rect 11889 -15930 11905 -15896
rect 12281 -15930 12297 -15896
rect 11176 -15958 11210 -15942
rect 11176 -16742 11210 -16726
rect 11704 -15958 11738 -15942
rect 11704 -16742 11738 -16726
rect 11812 -15958 11846 -15942
rect 11812 -16742 11846 -16726
rect 12340 -15958 12374 -15942
rect 12340 -16742 12374 -16726
rect 11253 -16788 11269 -16754
rect 11645 -16788 11661 -16754
rect 11889 -16788 11905 -16754
rect 12281 -16788 12297 -16754
rect 11038 -16888 11072 -16826
rect 12478 -16888 12512 -16826
rect 11038 -16922 11134 -16888
rect 12416 -16922 12512 -16888
rect 12638 -15270 12734 -15236
rect 14016 -15270 14112 -15236
rect 12638 -15332 12672 -15270
rect 14078 -15332 14112 -15270
rect 12853 -15404 12869 -15370
rect 13245 -15404 13261 -15370
rect 13489 -15404 13505 -15370
rect 13881 -15404 13897 -15370
rect 12776 -15432 12810 -15416
rect 12776 -15616 12810 -15600
rect 13304 -15432 13338 -15416
rect 13304 -15616 13338 -15600
rect 13412 -15432 13446 -15416
rect 13412 -15616 13446 -15600
rect 13940 -15432 13974 -15416
rect 13940 -15616 13974 -15600
rect 12853 -15662 12869 -15628
rect 13245 -15662 13261 -15628
rect 13489 -15662 13505 -15628
rect 13881 -15662 13897 -15628
rect 12638 -15762 12672 -15700
rect 14078 -15762 14112 -15700
rect 12638 -15796 12734 -15762
rect 14016 -15796 14112 -15762
rect 12638 -15858 12672 -15796
rect 14078 -15858 14112 -15796
rect 12853 -15930 12869 -15896
rect 13245 -15930 13261 -15896
rect 13489 -15930 13505 -15896
rect 13881 -15930 13897 -15896
rect 12776 -15958 12810 -15942
rect 12776 -16742 12810 -16726
rect 13304 -15958 13338 -15942
rect 13304 -16742 13338 -16726
rect 13412 -15958 13446 -15942
rect 13412 -16742 13446 -16726
rect 13940 -15958 13974 -15942
rect 13940 -16742 13974 -16726
rect 12853 -16788 12869 -16754
rect 13245 -16788 13261 -16754
rect 13489 -16788 13505 -16754
rect 13881 -16788 13897 -16754
rect 12638 -16888 12672 -16826
rect 14078 -16888 14112 -16826
rect 12638 -16922 12734 -16888
rect 14016 -16922 14112 -16888
rect 14238 -15270 14334 -15236
rect 15616 -15270 15712 -15236
rect 14238 -15332 14272 -15270
rect 15678 -15332 15712 -15270
rect 14453 -15404 14469 -15370
rect 14845 -15404 14861 -15370
rect 15089 -15404 15105 -15370
rect 15481 -15404 15497 -15370
rect 14376 -15432 14410 -15416
rect 14376 -15616 14410 -15600
rect 14904 -15432 14938 -15416
rect 14904 -15616 14938 -15600
rect 15012 -15432 15046 -15416
rect 15012 -15616 15046 -15600
rect 15540 -15432 15574 -15416
rect 15540 -15616 15574 -15600
rect 14453 -15662 14469 -15628
rect 14845 -15662 14861 -15628
rect 15089 -15662 15105 -15628
rect 15481 -15662 15497 -15628
rect 14238 -15762 14272 -15700
rect 15678 -15762 15712 -15700
rect 14238 -15796 14334 -15762
rect 15616 -15796 15712 -15762
rect 14238 -15858 14272 -15796
rect 15678 -15858 15712 -15796
rect 14453 -15930 14469 -15896
rect 14845 -15930 14861 -15896
rect 15089 -15930 15105 -15896
rect 15481 -15930 15497 -15896
rect 14376 -15958 14410 -15942
rect 14376 -16742 14410 -16726
rect 14904 -15958 14938 -15942
rect 14904 -16742 14938 -16726
rect 15012 -15958 15046 -15942
rect 15012 -16742 15046 -16726
rect 15540 -15958 15574 -15942
rect 15540 -16742 15574 -16726
rect 14453 -16788 14469 -16754
rect 14845 -16788 14861 -16754
rect 15089 -16788 15105 -16754
rect 15481 -16788 15497 -16754
rect 14238 -16888 14272 -16826
rect 15678 -16888 15712 -16826
rect 14238 -16922 14334 -16888
rect 15616 -16922 15712 -16888
rect 15838 -15270 15934 -15236
rect 17216 -15270 17312 -15236
rect 15838 -15332 15872 -15270
rect 17278 -15332 17312 -15270
rect 16053 -15404 16069 -15370
rect 16445 -15404 16461 -15370
rect 16689 -15404 16705 -15370
rect 17081 -15404 17097 -15370
rect 15976 -15432 16010 -15416
rect 15976 -15616 16010 -15600
rect 16504 -15432 16538 -15416
rect 16504 -15616 16538 -15600
rect 16612 -15432 16646 -15416
rect 16612 -15616 16646 -15600
rect 17140 -15432 17174 -15416
rect 17140 -15616 17174 -15600
rect 16053 -15662 16069 -15628
rect 16445 -15662 16461 -15628
rect 16689 -15662 16705 -15628
rect 17081 -15662 17097 -15628
rect 15838 -15762 15872 -15700
rect 17278 -15762 17312 -15700
rect 15838 -15796 15934 -15762
rect 17216 -15796 17312 -15762
rect 15838 -15858 15872 -15796
rect 17278 -15858 17312 -15796
rect 16053 -15930 16069 -15896
rect 16445 -15930 16461 -15896
rect 16689 -15930 16705 -15896
rect 17081 -15930 17097 -15896
rect 15976 -15958 16010 -15942
rect 15976 -16742 16010 -16726
rect 16504 -15958 16538 -15942
rect 16504 -16742 16538 -16726
rect 16612 -15958 16646 -15942
rect 16612 -16742 16646 -16726
rect 17140 -15958 17174 -15942
rect 17140 -16742 17174 -16726
rect 16053 -16788 16069 -16754
rect 16445 -16788 16461 -16754
rect 16689 -16788 16705 -16754
rect 17081 -16788 17097 -16754
rect 15838 -16888 15872 -16826
rect 17278 -16888 17312 -16826
rect 15838 -16922 15934 -16888
rect 17216 -16922 17312 -16888
rect 17438 -15270 17534 -15236
rect 18816 -15270 18912 -15236
rect 17438 -15332 17472 -15270
rect 18878 -15332 18912 -15270
rect 17653 -15404 17669 -15370
rect 18045 -15404 18061 -15370
rect 18289 -15404 18305 -15370
rect 18681 -15404 18697 -15370
rect 17576 -15432 17610 -15416
rect 17576 -15616 17610 -15600
rect 18104 -15432 18138 -15416
rect 18104 -15616 18138 -15600
rect 18212 -15432 18246 -15416
rect 18212 -15616 18246 -15600
rect 18740 -15432 18774 -15416
rect 18740 -15616 18774 -15600
rect 17653 -15662 17669 -15628
rect 18045 -15662 18061 -15628
rect 18289 -15662 18305 -15628
rect 18681 -15662 18697 -15628
rect 17438 -15762 17472 -15700
rect 18878 -15762 18912 -15700
rect 17438 -15796 17534 -15762
rect 18816 -15796 18912 -15762
rect 17438 -15858 17472 -15796
rect 18878 -15858 18912 -15796
rect 17653 -15930 17669 -15896
rect 18045 -15930 18061 -15896
rect 18289 -15930 18305 -15896
rect 18681 -15930 18697 -15896
rect 17576 -15958 17610 -15942
rect 17576 -16742 17610 -16726
rect 18104 -15958 18138 -15942
rect 18104 -16742 18138 -16726
rect 18212 -15958 18246 -15942
rect 18212 -16742 18246 -16726
rect 18740 -15958 18774 -15942
rect 18740 -16742 18774 -16726
rect 17653 -16788 17669 -16754
rect 18045 -16788 18061 -16754
rect 18289 -16788 18305 -16754
rect 18681 -16788 18697 -16754
rect 17438 -16888 17472 -16826
rect 18878 -16888 18912 -16826
rect 17438 -16922 17534 -16888
rect 18816 -16922 18912 -16888
rect 19038 -15270 19134 -15236
rect 20416 -15270 20512 -15236
rect 19038 -15332 19072 -15270
rect 20478 -15332 20512 -15270
rect 19253 -15404 19269 -15370
rect 19645 -15404 19661 -15370
rect 19889 -15404 19905 -15370
rect 20281 -15404 20297 -15370
rect 19176 -15432 19210 -15416
rect 19176 -15616 19210 -15600
rect 19704 -15432 19738 -15416
rect 19704 -15616 19738 -15600
rect 19812 -15432 19846 -15416
rect 19812 -15616 19846 -15600
rect 20340 -15432 20374 -15416
rect 20340 -15616 20374 -15600
rect 19253 -15662 19269 -15628
rect 19645 -15662 19661 -15628
rect 19889 -15662 19905 -15628
rect 20281 -15662 20297 -15628
rect 19038 -15762 19072 -15700
rect 20478 -15762 20512 -15700
rect 19038 -15796 19134 -15762
rect 20416 -15796 20512 -15762
rect 19038 -15858 19072 -15796
rect 20478 -15858 20512 -15796
rect 19253 -15930 19269 -15896
rect 19645 -15930 19661 -15896
rect 19889 -15930 19905 -15896
rect 20281 -15930 20297 -15896
rect 19176 -15958 19210 -15942
rect 19176 -16742 19210 -16726
rect 19704 -15958 19738 -15942
rect 19704 -16742 19738 -16726
rect 19812 -15958 19846 -15942
rect 19812 -16742 19846 -16726
rect 20340 -15958 20374 -15942
rect 20340 -16742 20374 -16726
rect 19253 -16788 19269 -16754
rect 19645 -16788 19661 -16754
rect 19889 -16788 19905 -16754
rect 20281 -16788 20297 -16754
rect 19038 -16888 19072 -16826
rect 20478 -16888 20512 -16826
rect 19038 -16922 19134 -16888
rect 20416 -16922 20512 -16888
rect 20638 -15270 20734 -15236
rect 22016 -15270 22112 -15236
rect 20638 -15332 20672 -15270
rect 22078 -15332 22112 -15270
rect 20853 -15404 20869 -15370
rect 21245 -15404 21261 -15370
rect 21489 -15404 21505 -15370
rect 21881 -15404 21897 -15370
rect 20776 -15432 20810 -15416
rect 20776 -15616 20810 -15600
rect 21304 -15432 21338 -15416
rect 21304 -15616 21338 -15600
rect 21412 -15432 21446 -15416
rect 21412 -15616 21446 -15600
rect 21940 -15432 21974 -15416
rect 21940 -15616 21974 -15600
rect 20853 -15662 20869 -15628
rect 21245 -15662 21261 -15628
rect 21489 -15662 21505 -15628
rect 21881 -15662 21897 -15628
rect 20638 -15762 20672 -15700
rect 22078 -15762 22112 -15700
rect 20638 -15796 20734 -15762
rect 22016 -15796 22112 -15762
rect 20638 -15858 20672 -15796
rect 22078 -15858 22112 -15796
rect 20853 -15930 20869 -15896
rect 21245 -15930 21261 -15896
rect 21489 -15930 21505 -15896
rect 21881 -15930 21897 -15896
rect 20776 -15958 20810 -15942
rect 20776 -16742 20810 -16726
rect 21304 -15958 21338 -15942
rect 21304 -16742 21338 -16726
rect 21412 -15958 21446 -15942
rect 21412 -16742 21446 -16726
rect 21940 -15958 21974 -15942
rect 21940 -16742 21974 -16726
rect 20853 -16788 20869 -16754
rect 21245 -16788 21261 -16754
rect 21489 -16788 21505 -16754
rect 21881 -16788 21897 -16754
rect 20638 -16888 20672 -16826
rect 22078 -16888 22112 -16826
rect 20638 -16922 20734 -16888
rect 22016 -16922 22112 -16888
rect 22238 -15270 22334 -15236
rect 23616 -15270 23712 -15236
rect 22238 -15332 22272 -15270
rect 23678 -15332 23712 -15270
rect 22453 -15404 22469 -15370
rect 22845 -15404 22861 -15370
rect 23089 -15404 23105 -15370
rect 23481 -15404 23497 -15370
rect 22376 -15432 22410 -15416
rect 22376 -15616 22410 -15600
rect 22904 -15432 22938 -15416
rect 22904 -15616 22938 -15600
rect 23012 -15432 23046 -15416
rect 23012 -15616 23046 -15600
rect 23540 -15432 23574 -15416
rect 23540 -15616 23574 -15600
rect 22453 -15662 22469 -15628
rect 22845 -15662 22861 -15628
rect 23089 -15662 23105 -15628
rect 23481 -15662 23497 -15628
rect 22238 -15762 22272 -15700
rect 23678 -15762 23712 -15700
rect 22238 -15796 22334 -15762
rect 23616 -15796 23712 -15762
rect 22238 -15858 22272 -15796
rect 23678 -15858 23712 -15796
rect 22453 -15930 22469 -15896
rect 22845 -15930 22861 -15896
rect 23089 -15930 23105 -15896
rect 23481 -15930 23497 -15896
rect 22376 -15958 22410 -15942
rect 22376 -16742 22410 -16726
rect 22904 -15958 22938 -15942
rect 22904 -16742 22938 -16726
rect 23012 -15958 23046 -15942
rect 23012 -16742 23046 -16726
rect 23540 -15958 23574 -15942
rect 23540 -16742 23574 -16726
rect 22453 -16788 22469 -16754
rect 22845 -16788 22861 -16754
rect 23089 -16788 23105 -16754
rect 23481 -16788 23497 -16754
rect 22238 -16888 22272 -16826
rect 23678 -16888 23712 -16826
rect 22238 -16922 22334 -16888
rect 23616 -16922 23712 -16888
rect 23838 -15270 23934 -15236
rect 25216 -15270 25312 -15236
rect 23838 -15332 23872 -15270
rect 25278 -15332 25312 -15270
rect 24053 -15404 24069 -15370
rect 24445 -15404 24461 -15370
rect 24689 -15404 24705 -15370
rect 25081 -15404 25097 -15370
rect 23976 -15432 24010 -15416
rect 23976 -15616 24010 -15600
rect 24504 -15432 24538 -15416
rect 24504 -15616 24538 -15600
rect 24612 -15432 24646 -15416
rect 24612 -15616 24646 -15600
rect 25140 -15432 25174 -15416
rect 25140 -15616 25174 -15600
rect 24053 -15662 24069 -15628
rect 24445 -15662 24461 -15628
rect 24689 -15662 24705 -15628
rect 25081 -15662 25097 -15628
rect 23838 -15762 23872 -15700
rect 25278 -15762 25312 -15700
rect 23838 -15796 23934 -15762
rect 25216 -15796 25312 -15762
rect 23838 -15858 23872 -15796
rect 25278 -15858 25312 -15796
rect 24053 -15930 24069 -15896
rect 24445 -15930 24461 -15896
rect 24689 -15930 24705 -15896
rect 25081 -15930 25097 -15896
rect 23976 -15958 24010 -15942
rect 23976 -16742 24010 -16726
rect 24504 -15958 24538 -15942
rect 24504 -16742 24538 -16726
rect 24612 -15958 24646 -15942
rect 24612 -16742 24646 -16726
rect 25140 -15958 25174 -15942
rect 25140 -16742 25174 -16726
rect 24053 -16788 24069 -16754
rect 24445 -16788 24461 -16754
rect 24689 -16788 24705 -16754
rect 25081 -16788 25097 -16754
rect 23838 -16888 23872 -16826
rect 25278 -16888 25312 -16826
rect 23838 -16922 23934 -16888
rect 25216 -16922 25312 -16888
rect 25438 -15270 25534 -15236
rect 26816 -15270 26912 -15236
rect 25438 -15332 25472 -15270
rect 26878 -15332 26912 -15270
rect 25653 -15404 25669 -15370
rect 26045 -15404 26061 -15370
rect 26289 -15404 26305 -15370
rect 26681 -15404 26697 -15370
rect 25576 -15432 25610 -15416
rect 25576 -15616 25610 -15600
rect 26104 -15432 26138 -15416
rect 26104 -15616 26138 -15600
rect 26212 -15432 26246 -15416
rect 26212 -15616 26246 -15600
rect 26740 -15432 26774 -15416
rect 26740 -15616 26774 -15600
rect 25653 -15662 25669 -15628
rect 26045 -15662 26061 -15628
rect 26289 -15662 26305 -15628
rect 26681 -15662 26697 -15628
rect 25438 -15762 25472 -15700
rect 26878 -15762 26912 -15700
rect 25438 -15796 25534 -15762
rect 26816 -15796 26912 -15762
rect 25438 -15858 25472 -15796
rect 26878 -15858 26912 -15796
rect 25653 -15930 25669 -15896
rect 26045 -15930 26061 -15896
rect 26289 -15930 26305 -15896
rect 26681 -15930 26697 -15896
rect 25576 -15958 25610 -15942
rect 25576 -16742 25610 -16726
rect 26104 -15958 26138 -15942
rect 26104 -16742 26138 -16726
rect 26212 -15958 26246 -15942
rect 26212 -16742 26246 -16726
rect 26740 -15958 26774 -15942
rect 26740 -16742 26774 -16726
rect 25653 -16788 25669 -16754
rect 26045 -16788 26061 -16754
rect 26289 -16788 26305 -16754
rect 26681 -16788 26697 -16754
rect 25438 -16888 25472 -16826
rect 26878 -16888 26912 -16826
rect 25438 -16922 25534 -16888
rect 26816 -16922 26912 -16888
rect 27038 -15270 27134 -15236
rect 28416 -15270 28512 -15236
rect 27038 -15332 27072 -15270
rect 28478 -15332 28512 -15270
rect 27253 -15404 27269 -15370
rect 27645 -15404 27661 -15370
rect 27889 -15404 27905 -15370
rect 28281 -15404 28297 -15370
rect 27176 -15432 27210 -15416
rect 27176 -15616 27210 -15600
rect 27704 -15432 27738 -15416
rect 27704 -15616 27738 -15600
rect 27812 -15432 27846 -15416
rect 27812 -15616 27846 -15600
rect 28340 -15432 28374 -15416
rect 28340 -15616 28374 -15600
rect 27253 -15662 27269 -15628
rect 27645 -15662 27661 -15628
rect 27889 -15662 27905 -15628
rect 28281 -15662 28297 -15628
rect 27038 -15762 27072 -15700
rect 28478 -15762 28512 -15700
rect 27038 -15796 27134 -15762
rect 28416 -15796 28512 -15762
rect 27038 -15858 27072 -15796
rect 28478 -15858 28512 -15796
rect 27253 -15930 27269 -15896
rect 27645 -15930 27661 -15896
rect 27889 -15930 27905 -15896
rect 28281 -15930 28297 -15896
rect 27176 -15958 27210 -15942
rect 27176 -16742 27210 -16726
rect 27704 -15958 27738 -15942
rect 27704 -16742 27738 -16726
rect 27812 -15958 27846 -15942
rect 27812 -16742 27846 -16726
rect 28340 -15958 28374 -15942
rect 28340 -16742 28374 -16726
rect 27253 -16788 27269 -16754
rect 27645 -16788 27661 -16754
rect 27889 -16788 27905 -16754
rect 28281 -16788 28297 -16754
rect 27038 -16888 27072 -16826
rect 28478 -16888 28512 -16826
rect 27038 -16922 27134 -16888
rect 28416 -16922 28512 -16888
rect 28638 -15270 28734 -15236
rect 30016 -15270 30112 -15236
rect 28638 -15332 28672 -15270
rect 30078 -15332 30112 -15270
rect 28853 -15404 28869 -15370
rect 29245 -15404 29261 -15370
rect 29489 -15404 29505 -15370
rect 29881 -15404 29897 -15370
rect 28776 -15432 28810 -15416
rect 28776 -15616 28810 -15600
rect 29304 -15432 29338 -15416
rect 29304 -15616 29338 -15600
rect 29412 -15432 29446 -15416
rect 29412 -15616 29446 -15600
rect 29940 -15432 29974 -15416
rect 29940 -15616 29974 -15600
rect 28853 -15662 28869 -15628
rect 29245 -15662 29261 -15628
rect 29489 -15662 29505 -15628
rect 29881 -15662 29897 -15628
rect 28638 -15762 28672 -15700
rect 30078 -15762 30112 -15700
rect 28638 -15796 28734 -15762
rect 30016 -15796 30112 -15762
rect 28638 -15858 28672 -15796
rect 30078 -15858 30112 -15796
rect 28853 -15930 28869 -15896
rect 29245 -15930 29261 -15896
rect 29489 -15930 29505 -15896
rect 29881 -15930 29897 -15896
rect 28776 -15958 28810 -15942
rect 28776 -16742 28810 -16726
rect 29304 -15958 29338 -15942
rect 29304 -16742 29338 -16726
rect 29412 -15958 29446 -15942
rect 29412 -16742 29446 -16726
rect 29940 -15958 29974 -15942
rect 29940 -16742 29974 -16726
rect 28853 -16788 28869 -16754
rect 29245 -16788 29261 -16754
rect 29489 -16788 29505 -16754
rect 29881 -16788 29897 -16754
rect 28638 -16888 28672 -16826
rect 30078 -16888 30112 -16826
rect 28638 -16922 28734 -16888
rect 30016 -16922 30112 -16888
rect 30238 -15270 30334 -15236
rect 31616 -15270 31712 -15236
rect 30238 -15332 30272 -15270
rect 31678 -15332 31712 -15270
rect 30453 -15404 30469 -15370
rect 30845 -15404 30861 -15370
rect 31089 -15404 31105 -15370
rect 31481 -15404 31497 -15370
rect 30376 -15432 30410 -15416
rect 30376 -15616 30410 -15600
rect 30904 -15432 30938 -15416
rect 30904 -15616 30938 -15600
rect 31012 -15432 31046 -15416
rect 31012 -15616 31046 -15600
rect 31540 -15432 31574 -15416
rect 31540 -15616 31574 -15600
rect 30453 -15662 30469 -15628
rect 30845 -15662 30861 -15628
rect 31089 -15662 31105 -15628
rect 31481 -15662 31497 -15628
rect 30238 -15762 30272 -15700
rect 31678 -15762 31712 -15700
rect 30238 -15796 30334 -15762
rect 31616 -15796 31712 -15762
rect 30238 -15858 30272 -15796
rect 31678 -15858 31712 -15796
rect 30453 -15930 30469 -15896
rect 30845 -15930 30861 -15896
rect 31089 -15930 31105 -15896
rect 31481 -15930 31497 -15896
rect 30376 -15958 30410 -15942
rect 30376 -16742 30410 -16726
rect 30904 -15958 30938 -15942
rect 30904 -16742 30938 -16726
rect 31012 -15958 31046 -15942
rect 31012 -16742 31046 -16726
rect 31540 -15958 31574 -15942
rect 31540 -16742 31574 -16726
rect 30453 -16788 30469 -16754
rect 30845 -16788 30861 -16754
rect 31089 -16788 31105 -16754
rect 31481 -16788 31497 -16754
rect 30238 -16888 30272 -16826
rect 31678 -16888 31712 -16826
rect 30238 -16922 30334 -16888
rect 31616 -16922 31712 -16888
rect 31838 -15270 31934 -15236
rect 33216 -15270 33312 -15236
rect 31838 -15332 31872 -15270
rect 33278 -15332 33312 -15270
rect 32053 -15404 32069 -15370
rect 32445 -15404 32461 -15370
rect 32689 -15404 32705 -15370
rect 33081 -15404 33097 -15370
rect 31976 -15432 32010 -15416
rect 31976 -15616 32010 -15600
rect 32504 -15432 32538 -15416
rect 32504 -15616 32538 -15600
rect 32612 -15432 32646 -15416
rect 32612 -15616 32646 -15600
rect 33140 -15432 33174 -15416
rect 33140 -15616 33174 -15600
rect 32053 -15662 32069 -15628
rect 32445 -15662 32461 -15628
rect 32689 -15662 32705 -15628
rect 33081 -15662 33097 -15628
rect 31838 -15762 31872 -15700
rect 33278 -15762 33312 -15700
rect 31838 -15796 31934 -15762
rect 33216 -15796 33312 -15762
rect 31838 -15858 31872 -15796
rect 33278 -15858 33312 -15796
rect 32053 -15930 32069 -15896
rect 32445 -15930 32461 -15896
rect 32689 -15930 32705 -15896
rect 33081 -15930 33097 -15896
rect 31976 -15958 32010 -15942
rect 31976 -16742 32010 -16726
rect 32504 -15958 32538 -15942
rect 32504 -16742 32538 -16726
rect 32612 -15958 32646 -15942
rect 32612 -16742 32646 -16726
rect 33140 -15958 33174 -15942
rect 33140 -16742 33174 -16726
rect 32053 -16788 32069 -16754
rect 32445 -16788 32461 -16754
rect 32689 -16788 32705 -16754
rect 33081 -16788 33097 -16754
rect 31838 -16888 31872 -16826
rect 33278 -16888 33312 -16826
rect 31838 -16922 31934 -16888
rect 33216 -16922 33312 -16888
rect 33438 -15270 33534 -15236
rect 34816 -15270 34912 -15236
rect 33438 -15332 33472 -15270
rect 34878 -15332 34912 -15270
rect 33653 -15404 33669 -15370
rect 34045 -15404 34061 -15370
rect 34289 -15404 34305 -15370
rect 34681 -15404 34697 -15370
rect 33576 -15432 33610 -15416
rect 33576 -15616 33610 -15600
rect 34104 -15432 34138 -15416
rect 34104 -15616 34138 -15600
rect 34212 -15432 34246 -15416
rect 34212 -15616 34246 -15600
rect 34740 -15432 34774 -15416
rect 34740 -15616 34774 -15600
rect 33653 -15662 33669 -15628
rect 34045 -15662 34061 -15628
rect 34289 -15662 34305 -15628
rect 34681 -15662 34697 -15628
rect 33438 -15762 33472 -15700
rect 34878 -15762 34912 -15700
rect 33438 -15796 33534 -15762
rect 34816 -15796 34912 -15762
rect 33438 -15858 33472 -15796
rect 34878 -15858 34912 -15796
rect 33653 -15930 33669 -15896
rect 34045 -15930 34061 -15896
rect 34289 -15930 34305 -15896
rect 34681 -15930 34697 -15896
rect 33576 -15958 33610 -15942
rect 33576 -16742 33610 -16726
rect 34104 -15958 34138 -15942
rect 34104 -16742 34138 -16726
rect 34212 -15958 34246 -15942
rect 34212 -16742 34246 -16726
rect 34740 -15958 34774 -15942
rect 34740 -16742 34774 -16726
rect 33653 -16788 33669 -16754
rect 34045 -16788 34061 -16754
rect 34289 -16788 34305 -16754
rect 34681 -16788 34697 -16754
rect 33438 -16888 33472 -16826
rect 34878 -16888 34912 -16826
rect 33438 -16922 33534 -16888
rect 34816 -16922 34912 -16888
rect 35038 -15270 35134 -15236
rect 36416 -15270 36734 -15236
rect 38016 -15270 38112 -15236
rect 35038 -15332 35072 -15270
rect 36478 -15332 38112 -15270
rect 35253 -15404 35269 -15370
rect 35645 -15404 35661 -15370
rect 35889 -15404 35905 -15370
rect 36281 -15404 36297 -15370
rect 35176 -15432 35210 -15416
rect 35176 -15616 35210 -15600
rect 35704 -15432 35738 -15416
rect 35704 -15616 35738 -15600
rect 35812 -15432 35846 -15416
rect 35812 -15616 35846 -15600
rect 36340 -15432 36374 -15416
rect 36340 -15616 36374 -15600
rect 35253 -15662 35269 -15628
rect 35645 -15662 35661 -15628
rect 35889 -15662 35905 -15628
rect 36281 -15662 36297 -15628
rect 35038 -15762 35072 -15700
rect 36512 -15700 36638 -15332
rect 36672 -15370 38078 -15332
rect 36672 -15404 36869 -15370
rect 37245 -15404 37505 -15370
rect 37881 -15404 38078 -15370
rect 36672 -15432 38078 -15404
rect 36672 -15600 36776 -15432
rect 36810 -15600 37304 -15432
rect 37338 -15600 37412 -15432
rect 37446 -15600 37940 -15432
rect 37974 -15600 38078 -15432
rect 36672 -15628 38078 -15600
rect 36672 -15662 36869 -15628
rect 37245 -15662 37505 -15628
rect 37881 -15662 38078 -15628
rect 36672 -15700 38078 -15662
rect 36478 -15762 38112 -15700
rect 35038 -15796 35134 -15762
rect 36416 -15796 36734 -15762
rect 38016 -15796 38112 -15762
rect 35038 -15858 35072 -15796
rect 36478 -15858 38112 -15796
rect 35253 -15930 35269 -15896
rect 35645 -15930 35661 -15896
rect 35889 -15930 35905 -15896
rect 36281 -15930 36297 -15896
rect 35176 -15958 35210 -15942
rect 35176 -16742 35210 -16726
rect 35704 -15958 35738 -15942
rect 35704 -16742 35738 -16726
rect 35812 -15958 35846 -15942
rect 35812 -16742 35846 -16726
rect 36340 -15958 36374 -15942
rect 36340 -16742 36374 -16726
rect 35253 -16788 35269 -16754
rect 35645 -16788 35661 -16754
rect 35889 -16788 35905 -16754
rect 36281 -16788 36297 -16754
rect 35038 -16888 35072 -16826
rect 36512 -16826 36638 -15858
rect 36672 -15896 38078 -15858
rect 36672 -15930 36869 -15896
rect 37245 -15930 37505 -15896
rect 37881 -15930 38078 -15896
rect 36672 -15958 38078 -15930
rect 36672 -16726 36776 -15958
rect 36810 -16726 37304 -15958
rect 37338 -16726 37412 -15958
rect 37446 -16726 37940 -15958
rect 37974 -16726 38078 -15958
rect 36672 -16754 38078 -16726
rect 36672 -16788 36869 -16754
rect 37245 -16788 37505 -16754
rect 37881 -16788 38078 -16754
rect 36672 -16826 38078 -16788
rect 36478 -16888 38112 -16826
rect 35038 -16922 35134 -16888
rect 36416 -16922 36734 -16888
rect 38016 -16922 38112 -16888
rect -140 -17036 1460 -16922
rect 36500 -17036 38100 -16922
rect -162 -17070 -66 -17036
rect 1216 -17070 1534 -17036
rect 2816 -17070 2912 -17036
rect -162 -17132 1472 -17070
rect -128 -17170 1278 -17132
rect -128 -17204 69 -17170
rect 445 -17204 705 -17170
rect 1081 -17204 1278 -17170
rect -128 -17232 1278 -17204
rect -128 -17400 -24 -17232
rect 10 -17400 504 -17232
rect 538 -17400 612 -17232
rect 646 -17400 1140 -17232
rect 1174 -17400 1278 -17232
rect -128 -17428 1278 -17400
rect -128 -17462 69 -17428
rect 445 -17462 705 -17428
rect 1081 -17462 1278 -17428
rect -128 -17500 1278 -17462
rect 1312 -17500 1438 -17132
rect 2878 -17132 2912 -17070
rect 1653 -17204 1669 -17170
rect 2045 -17204 2061 -17170
rect 2289 -17204 2305 -17170
rect 2681 -17204 2697 -17170
rect 1576 -17232 1610 -17216
rect 1576 -17416 1610 -17400
rect 2104 -17232 2138 -17216
rect 2104 -17416 2138 -17400
rect 2212 -17232 2246 -17216
rect 2212 -17416 2246 -17400
rect 2740 -17232 2774 -17216
rect 2740 -17416 2774 -17400
rect 1653 -17462 1669 -17428
rect 2045 -17462 2061 -17428
rect 2289 -17462 2305 -17428
rect 2681 -17462 2697 -17428
rect -162 -17562 1472 -17500
rect 2878 -17562 2912 -17500
rect -162 -17596 -66 -17562
rect 1216 -17596 1534 -17562
rect 2816 -17596 2912 -17562
rect -162 -17658 1472 -17596
rect -128 -17696 1278 -17658
rect -128 -17730 69 -17696
rect 445 -17730 705 -17696
rect 1081 -17730 1278 -17696
rect -128 -17758 1278 -17730
rect -128 -18526 -24 -17758
rect 10 -18526 504 -17758
rect 538 -18526 612 -17758
rect 646 -18526 1140 -17758
rect 1174 -18526 1278 -17758
rect -128 -18554 1278 -18526
rect -128 -18588 69 -18554
rect 445 -18588 705 -18554
rect 1081 -18588 1278 -18554
rect -128 -18626 1278 -18588
rect 1312 -18626 1438 -17658
rect 2878 -17658 2912 -17596
rect 1653 -17730 1669 -17696
rect 2045 -17730 2061 -17696
rect 2289 -17730 2305 -17696
rect 2681 -17730 2697 -17696
rect 1576 -17758 1610 -17742
rect 1576 -18542 1610 -18526
rect 2104 -17758 2138 -17742
rect 2104 -18542 2138 -18526
rect 2212 -17758 2246 -17742
rect 2212 -18542 2246 -18526
rect 2740 -17758 2774 -17742
rect 2740 -18542 2774 -18526
rect 1653 -18588 1669 -18554
rect 2045 -18588 2061 -18554
rect 2289 -18588 2305 -18554
rect 2681 -18588 2697 -18554
rect -162 -18688 1472 -18626
rect 2878 -18688 2912 -18626
rect -162 -18722 -66 -18688
rect 1216 -18722 1534 -18688
rect 2816 -18722 2912 -18688
rect 3038 -17070 3134 -17036
rect 4416 -17070 4512 -17036
rect 3038 -17132 3072 -17070
rect 4478 -17132 4512 -17070
rect 3253 -17204 3269 -17170
rect 3645 -17204 3661 -17170
rect 3889 -17204 3905 -17170
rect 4281 -17204 4297 -17170
rect 3176 -17232 3210 -17216
rect 3176 -17416 3210 -17400
rect 3704 -17232 3738 -17216
rect 3704 -17416 3738 -17400
rect 3812 -17232 3846 -17216
rect 3812 -17416 3846 -17400
rect 4340 -17232 4374 -17216
rect 4340 -17416 4374 -17400
rect 3253 -17462 3269 -17428
rect 3645 -17462 3661 -17428
rect 3889 -17462 3905 -17428
rect 4281 -17462 4297 -17428
rect 3038 -17562 3072 -17500
rect 4478 -17562 4512 -17500
rect 3038 -17596 3134 -17562
rect 4416 -17596 4512 -17562
rect 3038 -17658 3072 -17596
rect 4478 -17658 4512 -17596
rect 3253 -17730 3269 -17696
rect 3645 -17730 3661 -17696
rect 3889 -17730 3905 -17696
rect 4281 -17730 4297 -17696
rect 3176 -17758 3210 -17742
rect 3176 -18542 3210 -18526
rect 3704 -17758 3738 -17742
rect 3704 -18542 3738 -18526
rect 3812 -17758 3846 -17742
rect 3812 -18542 3846 -18526
rect 4340 -17758 4374 -17742
rect 4340 -18542 4374 -18526
rect 3253 -18588 3269 -18554
rect 3645 -18588 3661 -18554
rect 3889 -18588 3905 -18554
rect 4281 -18588 4297 -18554
rect 3038 -18688 3072 -18626
rect 4478 -18688 4512 -18626
rect 3038 -18722 3134 -18688
rect 4416 -18722 4512 -18688
rect 4638 -17070 4734 -17036
rect 6016 -17070 6112 -17036
rect 4638 -17132 4672 -17070
rect 6078 -17132 6112 -17070
rect 4853 -17204 4869 -17170
rect 5245 -17204 5261 -17170
rect 5489 -17204 5505 -17170
rect 5881 -17204 5897 -17170
rect 4776 -17232 4810 -17216
rect 4776 -17416 4810 -17400
rect 5304 -17232 5338 -17216
rect 5304 -17416 5338 -17400
rect 5412 -17232 5446 -17216
rect 5412 -17416 5446 -17400
rect 5940 -17232 5974 -17216
rect 5940 -17416 5974 -17400
rect 4853 -17462 4869 -17428
rect 5245 -17462 5261 -17428
rect 5489 -17462 5505 -17428
rect 5881 -17462 5897 -17428
rect 4638 -17562 4672 -17500
rect 6078 -17562 6112 -17500
rect 4638 -17596 4734 -17562
rect 6016 -17596 6112 -17562
rect 4638 -17658 4672 -17596
rect 6078 -17658 6112 -17596
rect 4853 -17730 4869 -17696
rect 5245 -17730 5261 -17696
rect 5489 -17730 5505 -17696
rect 5881 -17730 5897 -17696
rect 4776 -17758 4810 -17742
rect 4776 -18542 4810 -18526
rect 5304 -17758 5338 -17742
rect 5304 -18542 5338 -18526
rect 5412 -17758 5446 -17742
rect 5412 -18542 5446 -18526
rect 5940 -17758 5974 -17742
rect 5940 -18542 5974 -18526
rect 4853 -18588 4869 -18554
rect 5245 -18588 5261 -18554
rect 5489 -18588 5505 -18554
rect 5881 -18588 5897 -18554
rect 4638 -18688 4672 -18626
rect 6078 -18688 6112 -18626
rect 4638 -18722 4734 -18688
rect 6016 -18722 6112 -18688
rect 6238 -17070 6334 -17036
rect 7616 -17070 7712 -17036
rect 6238 -17132 6272 -17070
rect 7678 -17132 7712 -17070
rect 6453 -17204 6469 -17170
rect 6845 -17204 6861 -17170
rect 7089 -17204 7105 -17170
rect 7481 -17204 7497 -17170
rect 6376 -17232 6410 -17216
rect 6376 -17416 6410 -17400
rect 6904 -17232 6938 -17216
rect 6904 -17416 6938 -17400
rect 7012 -17232 7046 -17216
rect 7012 -17416 7046 -17400
rect 7540 -17232 7574 -17216
rect 7540 -17416 7574 -17400
rect 6453 -17462 6469 -17428
rect 6845 -17462 6861 -17428
rect 7089 -17462 7105 -17428
rect 7481 -17462 7497 -17428
rect 6238 -17562 6272 -17500
rect 7678 -17562 7712 -17500
rect 6238 -17596 6334 -17562
rect 7616 -17596 7712 -17562
rect 6238 -17658 6272 -17596
rect 7678 -17658 7712 -17596
rect 6453 -17730 6469 -17696
rect 6845 -17730 6861 -17696
rect 7089 -17730 7105 -17696
rect 7481 -17730 7497 -17696
rect 6376 -17758 6410 -17742
rect 6376 -18542 6410 -18526
rect 6904 -17758 6938 -17742
rect 6904 -18542 6938 -18526
rect 7012 -17758 7046 -17742
rect 7012 -18542 7046 -18526
rect 7540 -17758 7574 -17742
rect 7540 -18542 7574 -18526
rect 6453 -18588 6469 -18554
rect 6845 -18588 6861 -18554
rect 7089 -18588 7105 -18554
rect 7481 -18588 7497 -18554
rect 6238 -18688 6272 -18626
rect 7678 -18688 7712 -18626
rect 6238 -18722 6334 -18688
rect 7616 -18722 7712 -18688
rect 7838 -17070 7934 -17036
rect 9216 -17070 9312 -17036
rect 7838 -17132 7872 -17070
rect 9278 -17132 9312 -17070
rect 8053 -17204 8069 -17170
rect 8445 -17204 8461 -17170
rect 8689 -17204 8705 -17170
rect 9081 -17204 9097 -17170
rect 7976 -17232 8010 -17216
rect 7976 -17416 8010 -17400
rect 8504 -17232 8538 -17216
rect 8504 -17416 8538 -17400
rect 8612 -17232 8646 -17216
rect 8612 -17416 8646 -17400
rect 9140 -17232 9174 -17216
rect 9140 -17416 9174 -17400
rect 8053 -17462 8069 -17428
rect 8445 -17462 8461 -17428
rect 8689 -17462 8705 -17428
rect 9081 -17462 9097 -17428
rect 7838 -17562 7872 -17500
rect 9278 -17562 9312 -17500
rect 7838 -17596 7934 -17562
rect 9216 -17596 9312 -17562
rect 7838 -17658 7872 -17596
rect 9278 -17658 9312 -17596
rect 8053 -17730 8069 -17696
rect 8445 -17730 8461 -17696
rect 8689 -17730 8705 -17696
rect 9081 -17730 9097 -17696
rect 7976 -17758 8010 -17742
rect 7976 -18542 8010 -18526
rect 8504 -17758 8538 -17742
rect 8504 -18542 8538 -18526
rect 8612 -17758 8646 -17742
rect 8612 -18542 8646 -18526
rect 9140 -17758 9174 -17742
rect 9140 -18542 9174 -18526
rect 8053 -18588 8069 -18554
rect 8445 -18588 8461 -18554
rect 8689 -18588 8705 -18554
rect 9081 -18588 9097 -18554
rect 7838 -18688 7872 -18626
rect 9278 -18688 9312 -18626
rect 7838 -18722 7934 -18688
rect 9216 -18722 9312 -18688
rect 9438 -17070 9534 -17036
rect 10816 -17070 10912 -17036
rect 9438 -17132 9472 -17070
rect 10878 -17132 10912 -17070
rect 9653 -17204 9669 -17170
rect 10045 -17204 10061 -17170
rect 10289 -17204 10305 -17170
rect 10681 -17204 10697 -17170
rect 9576 -17232 9610 -17216
rect 9576 -17416 9610 -17400
rect 10104 -17232 10138 -17216
rect 10104 -17416 10138 -17400
rect 10212 -17232 10246 -17216
rect 10212 -17416 10246 -17400
rect 10740 -17232 10774 -17216
rect 10740 -17416 10774 -17400
rect 9653 -17462 9669 -17428
rect 10045 -17462 10061 -17428
rect 10289 -17462 10305 -17428
rect 10681 -17462 10697 -17428
rect 9438 -17562 9472 -17500
rect 10878 -17562 10912 -17500
rect 9438 -17596 9534 -17562
rect 10816 -17596 10912 -17562
rect 9438 -17658 9472 -17596
rect 10878 -17658 10912 -17596
rect 9653 -17730 9669 -17696
rect 10045 -17730 10061 -17696
rect 10289 -17730 10305 -17696
rect 10681 -17730 10697 -17696
rect 9576 -17758 9610 -17742
rect 9576 -18542 9610 -18526
rect 10104 -17758 10138 -17742
rect 10104 -18542 10138 -18526
rect 10212 -17758 10246 -17742
rect 10212 -18542 10246 -18526
rect 10740 -17758 10774 -17742
rect 10740 -18542 10774 -18526
rect 9653 -18588 9669 -18554
rect 10045 -18588 10061 -18554
rect 10289 -18588 10305 -18554
rect 10681 -18588 10697 -18554
rect 9438 -18688 9472 -18626
rect 10878 -18688 10912 -18626
rect 9438 -18722 9534 -18688
rect 10816 -18722 10912 -18688
rect 11038 -17070 11134 -17036
rect 12416 -17070 12512 -17036
rect 11038 -17132 11072 -17070
rect 12478 -17132 12512 -17070
rect 11253 -17204 11269 -17170
rect 11645 -17204 11661 -17170
rect 11889 -17204 11905 -17170
rect 12281 -17204 12297 -17170
rect 11176 -17232 11210 -17216
rect 11176 -17416 11210 -17400
rect 11704 -17232 11738 -17216
rect 11704 -17416 11738 -17400
rect 11812 -17232 11846 -17216
rect 11812 -17416 11846 -17400
rect 12340 -17232 12374 -17216
rect 12340 -17416 12374 -17400
rect 11253 -17462 11269 -17428
rect 11645 -17462 11661 -17428
rect 11889 -17462 11905 -17428
rect 12281 -17462 12297 -17428
rect 11038 -17562 11072 -17500
rect 12478 -17562 12512 -17500
rect 11038 -17596 11134 -17562
rect 12416 -17596 12512 -17562
rect 11038 -17658 11072 -17596
rect 12478 -17658 12512 -17596
rect 11253 -17730 11269 -17696
rect 11645 -17730 11661 -17696
rect 11889 -17730 11905 -17696
rect 12281 -17730 12297 -17696
rect 11176 -17758 11210 -17742
rect 11176 -18542 11210 -18526
rect 11704 -17758 11738 -17742
rect 11704 -18542 11738 -18526
rect 11812 -17758 11846 -17742
rect 11812 -18542 11846 -18526
rect 12340 -17758 12374 -17742
rect 12340 -18542 12374 -18526
rect 11253 -18588 11269 -18554
rect 11645 -18588 11661 -18554
rect 11889 -18588 11905 -18554
rect 12281 -18588 12297 -18554
rect 11038 -18688 11072 -18626
rect 12478 -18688 12512 -18626
rect 11038 -18722 11134 -18688
rect 12416 -18722 12512 -18688
rect 12638 -17070 12734 -17036
rect 14016 -17070 14112 -17036
rect 12638 -17132 12672 -17070
rect 14078 -17132 14112 -17070
rect 12853 -17204 12869 -17170
rect 13245 -17204 13261 -17170
rect 13489 -17204 13505 -17170
rect 13881 -17204 13897 -17170
rect 12776 -17232 12810 -17216
rect 12776 -17416 12810 -17400
rect 13304 -17232 13338 -17216
rect 13304 -17416 13338 -17400
rect 13412 -17232 13446 -17216
rect 13412 -17416 13446 -17400
rect 13940 -17232 13974 -17216
rect 13940 -17416 13974 -17400
rect 12853 -17462 12869 -17428
rect 13245 -17462 13261 -17428
rect 13489 -17462 13505 -17428
rect 13881 -17462 13897 -17428
rect 12638 -17562 12672 -17500
rect 14078 -17562 14112 -17500
rect 12638 -17596 12734 -17562
rect 14016 -17596 14112 -17562
rect 12638 -17658 12672 -17596
rect 14078 -17658 14112 -17596
rect 12853 -17730 12869 -17696
rect 13245 -17730 13261 -17696
rect 13489 -17730 13505 -17696
rect 13881 -17730 13897 -17696
rect 12776 -17758 12810 -17742
rect 12776 -18542 12810 -18526
rect 13304 -17758 13338 -17742
rect 13304 -18542 13338 -18526
rect 13412 -17758 13446 -17742
rect 13412 -18542 13446 -18526
rect 13940 -17758 13974 -17742
rect 13940 -18542 13974 -18526
rect 12853 -18588 12869 -18554
rect 13245 -18588 13261 -18554
rect 13489 -18588 13505 -18554
rect 13881 -18588 13897 -18554
rect 12638 -18688 12672 -18626
rect 14078 -18688 14112 -18626
rect 12638 -18722 12734 -18688
rect 14016 -18722 14112 -18688
rect 14238 -17070 14334 -17036
rect 15616 -17070 15712 -17036
rect 14238 -17132 14272 -17070
rect 15678 -17132 15712 -17070
rect 14453 -17204 14469 -17170
rect 14845 -17204 14861 -17170
rect 15089 -17204 15105 -17170
rect 15481 -17204 15497 -17170
rect 14376 -17232 14410 -17216
rect 14376 -17416 14410 -17400
rect 14904 -17232 14938 -17216
rect 14904 -17416 14938 -17400
rect 15012 -17232 15046 -17216
rect 15012 -17416 15046 -17400
rect 15540 -17232 15574 -17216
rect 15540 -17416 15574 -17400
rect 14453 -17462 14469 -17428
rect 14845 -17462 14861 -17428
rect 15089 -17462 15105 -17428
rect 15481 -17462 15497 -17428
rect 14238 -17562 14272 -17500
rect 15678 -17562 15712 -17500
rect 14238 -17596 14334 -17562
rect 15616 -17596 15712 -17562
rect 14238 -17658 14272 -17596
rect 15678 -17658 15712 -17596
rect 14453 -17730 14469 -17696
rect 14845 -17730 14861 -17696
rect 15089 -17730 15105 -17696
rect 15481 -17730 15497 -17696
rect 14376 -17758 14410 -17742
rect 14376 -18542 14410 -18526
rect 14904 -17758 14938 -17742
rect 14904 -18542 14938 -18526
rect 15012 -17758 15046 -17742
rect 15012 -18542 15046 -18526
rect 15540 -17758 15574 -17742
rect 15540 -18542 15574 -18526
rect 14453 -18588 14469 -18554
rect 14845 -18588 14861 -18554
rect 15089 -18588 15105 -18554
rect 15481 -18588 15497 -18554
rect 14238 -18688 14272 -18626
rect 15678 -18688 15712 -18626
rect 14238 -18722 14334 -18688
rect 15616 -18722 15712 -18688
rect 15838 -17070 15934 -17036
rect 17216 -17070 17312 -17036
rect 15838 -17132 15872 -17070
rect 17278 -17132 17312 -17070
rect 16053 -17204 16069 -17170
rect 16445 -17204 16461 -17170
rect 16689 -17204 16705 -17170
rect 17081 -17204 17097 -17170
rect 15976 -17232 16010 -17216
rect 15976 -17416 16010 -17400
rect 16504 -17232 16538 -17216
rect 16504 -17416 16538 -17400
rect 16612 -17232 16646 -17216
rect 16612 -17416 16646 -17400
rect 17140 -17232 17174 -17216
rect 17140 -17416 17174 -17400
rect 16053 -17462 16069 -17428
rect 16445 -17462 16461 -17428
rect 16689 -17462 16705 -17428
rect 17081 -17462 17097 -17428
rect 15838 -17562 15872 -17500
rect 17278 -17562 17312 -17500
rect 15838 -17596 15934 -17562
rect 17216 -17596 17312 -17562
rect 15838 -17658 15872 -17596
rect 17278 -17658 17312 -17596
rect 16053 -17730 16069 -17696
rect 16445 -17730 16461 -17696
rect 16689 -17730 16705 -17696
rect 17081 -17730 17097 -17696
rect 15976 -17758 16010 -17742
rect 15976 -18542 16010 -18526
rect 16504 -17758 16538 -17742
rect 16504 -18542 16538 -18526
rect 16612 -17758 16646 -17742
rect 16612 -18542 16646 -18526
rect 17140 -17758 17174 -17742
rect 17140 -18542 17174 -18526
rect 16053 -18588 16069 -18554
rect 16445 -18588 16461 -18554
rect 16689 -18588 16705 -18554
rect 17081 -18588 17097 -18554
rect 15838 -18688 15872 -18626
rect 17278 -18688 17312 -18626
rect 15838 -18722 15934 -18688
rect 17216 -18722 17312 -18688
rect 17438 -17070 17534 -17036
rect 18816 -17070 18912 -17036
rect 17438 -17132 17472 -17070
rect 18878 -17132 18912 -17070
rect 17653 -17204 17669 -17170
rect 18045 -17204 18061 -17170
rect 18289 -17204 18305 -17170
rect 18681 -17204 18697 -17170
rect 17576 -17232 17610 -17216
rect 17576 -17416 17610 -17400
rect 18104 -17232 18138 -17216
rect 18104 -17416 18138 -17400
rect 18212 -17232 18246 -17216
rect 18212 -17416 18246 -17400
rect 18740 -17232 18774 -17216
rect 18740 -17416 18774 -17400
rect 17653 -17462 17669 -17428
rect 18045 -17462 18061 -17428
rect 18289 -17462 18305 -17428
rect 18681 -17462 18697 -17428
rect 17438 -17562 17472 -17500
rect 18878 -17562 18912 -17500
rect 17438 -17596 17534 -17562
rect 18816 -17596 18912 -17562
rect 17438 -17658 17472 -17596
rect 18878 -17658 18912 -17596
rect 17653 -17730 17669 -17696
rect 18045 -17730 18061 -17696
rect 18289 -17730 18305 -17696
rect 18681 -17730 18697 -17696
rect 17576 -17758 17610 -17742
rect 17576 -18542 17610 -18526
rect 18104 -17758 18138 -17742
rect 18104 -18542 18138 -18526
rect 18212 -17758 18246 -17742
rect 18212 -18542 18246 -18526
rect 18740 -17758 18774 -17742
rect 18740 -18542 18774 -18526
rect 17653 -18588 17669 -18554
rect 18045 -18588 18061 -18554
rect 18289 -18588 18305 -18554
rect 18681 -18588 18697 -18554
rect 17438 -18688 17472 -18626
rect 18878 -18688 18912 -18626
rect 17438 -18722 17534 -18688
rect 18816 -18722 18912 -18688
rect 19038 -17070 19134 -17036
rect 20416 -17070 20512 -17036
rect 19038 -17132 19072 -17070
rect 20478 -17132 20512 -17070
rect 19253 -17204 19269 -17170
rect 19645 -17204 19661 -17170
rect 19889 -17204 19905 -17170
rect 20281 -17204 20297 -17170
rect 19176 -17232 19210 -17216
rect 19176 -17416 19210 -17400
rect 19704 -17232 19738 -17216
rect 19704 -17416 19738 -17400
rect 19812 -17232 19846 -17216
rect 19812 -17416 19846 -17400
rect 20340 -17232 20374 -17216
rect 20340 -17416 20374 -17400
rect 19253 -17462 19269 -17428
rect 19645 -17462 19661 -17428
rect 19889 -17462 19905 -17428
rect 20281 -17462 20297 -17428
rect 19038 -17562 19072 -17500
rect 20478 -17562 20512 -17500
rect 19038 -17596 19134 -17562
rect 20416 -17596 20512 -17562
rect 19038 -17658 19072 -17596
rect 20478 -17658 20512 -17596
rect 19253 -17730 19269 -17696
rect 19645 -17730 19661 -17696
rect 19889 -17730 19905 -17696
rect 20281 -17730 20297 -17696
rect 19176 -17758 19210 -17742
rect 19176 -18542 19210 -18526
rect 19704 -17758 19738 -17742
rect 19704 -18542 19738 -18526
rect 19812 -17758 19846 -17742
rect 19812 -18542 19846 -18526
rect 20340 -17758 20374 -17742
rect 20340 -18542 20374 -18526
rect 19253 -18588 19269 -18554
rect 19645 -18588 19661 -18554
rect 19889 -18588 19905 -18554
rect 20281 -18588 20297 -18554
rect 19038 -18688 19072 -18626
rect 20478 -18688 20512 -18626
rect 19038 -18722 19134 -18688
rect 20416 -18722 20512 -18688
rect 20638 -17070 20734 -17036
rect 22016 -17070 22112 -17036
rect 20638 -17132 20672 -17070
rect 22078 -17132 22112 -17070
rect 20853 -17204 20869 -17170
rect 21245 -17204 21261 -17170
rect 21489 -17204 21505 -17170
rect 21881 -17204 21897 -17170
rect 20776 -17232 20810 -17216
rect 20776 -17416 20810 -17400
rect 21304 -17232 21338 -17216
rect 21304 -17416 21338 -17400
rect 21412 -17232 21446 -17216
rect 21412 -17416 21446 -17400
rect 21940 -17232 21974 -17216
rect 21940 -17416 21974 -17400
rect 20853 -17462 20869 -17428
rect 21245 -17462 21261 -17428
rect 21489 -17462 21505 -17428
rect 21881 -17462 21897 -17428
rect 20638 -17562 20672 -17500
rect 22078 -17562 22112 -17500
rect 20638 -17596 20734 -17562
rect 22016 -17596 22112 -17562
rect 20638 -17658 20672 -17596
rect 22078 -17658 22112 -17596
rect 20853 -17730 20869 -17696
rect 21245 -17730 21261 -17696
rect 21489 -17730 21505 -17696
rect 21881 -17730 21897 -17696
rect 20776 -17758 20810 -17742
rect 20776 -18542 20810 -18526
rect 21304 -17758 21338 -17742
rect 21304 -18542 21338 -18526
rect 21412 -17758 21446 -17742
rect 21412 -18542 21446 -18526
rect 21940 -17758 21974 -17742
rect 21940 -18542 21974 -18526
rect 20853 -18588 20869 -18554
rect 21245 -18588 21261 -18554
rect 21489 -18588 21505 -18554
rect 21881 -18588 21897 -18554
rect 20638 -18688 20672 -18626
rect 22078 -18688 22112 -18626
rect 20638 -18722 20734 -18688
rect 22016 -18722 22112 -18688
rect 22238 -17070 22334 -17036
rect 23616 -17070 23712 -17036
rect 22238 -17132 22272 -17070
rect 23678 -17132 23712 -17070
rect 22453 -17204 22469 -17170
rect 22845 -17204 22861 -17170
rect 23089 -17204 23105 -17170
rect 23481 -17204 23497 -17170
rect 22376 -17232 22410 -17216
rect 22376 -17416 22410 -17400
rect 22904 -17232 22938 -17216
rect 22904 -17416 22938 -17400
rect 23012 -17232 23046 -17216
rect 23012 -17416 23046 -17400
rect 23540 -17232 23574 -17216
rect 23540 -17416 23574 -17400
rect 22453 -17462 22469 -17428
rect 22845 -17462 22861 -17428
rect 23089 -17462 23105 -17428
rect 23481 -17462 23497 -17428
rect 22238 -17562 22272 -17500
rect 23678 -17562 23712 -17500
rect 22238 -17596 22334 -17562
rect 23616 -17596 23712 -17562
rect 22238 -17658 22272 -17596
rect 23678 -17658 23712 -17596
rect 22453 -17730 22469 -17696
rect 22845 -17730 22861 -17696
rect 23089 -17730 23105 -17696
rect 23481 -17730 23497 -17696
rect 22376 -17758 22410 -17742
rect 22376 -18542 22410 -18526
rect 22904 -17758 22938 -17742
rect 22904 -18542 22938 -18526
rect 23012 -17758 23046 -17742
rect 23012 -18542 23046 -18526
rect 23540 -17758 23574 -17742
rect 23540 -18542 23574 -18526
rect 22453 -18588 22469 -18554
rect 22845 -18588 22861 -18554
rect 23089 -18588 23105 -18554
rect 23481 -18588 23497 -18554
rect 22238 -18688 22272 -18626
rect 23678 -18688 23712 -18626
rect 22238 -18722 22334 -18688
rect 23616 -18722 23712 -18688
rect 23838 -17070 23934 -17036
rect 25216 -17070 25312 -17036
rect 23838 -17132 23872 -17070
rect 25278 -17132 25312 -17070
rect 24053 -17204 24069 -17170
rect 24445 -17204 24461 -17170
rect 24689 -17204 24705 -17170
rect 25081 -17204 25097 -17170
rect 23976 -17232 24010 -17216
rect 23976 -17416 24010 -17400
rect 24504 -17232 24538 -17216
rect 24504 -17416 24538 -17400
rect 24612 -17232 24646 -17216
rect 24612 -17416 24646 -17400
rect 25140 -17232 25174 -17216
rect 25140 -17416 25174 -17400
rect 24053 -17462 24069 -17428
rect 24445 -17462 24461 -17428
rect 24689 -17462 24705 -17428
rect 25081 -17462 25097 -17428
rect 23838 -17562 23872 -17500
rect 25278 -17562 25312 -17500
rect 23838 -17596 23934 -17562
rect 25216 -17596 25312 -17562
rect 23838 -17658 23872 -17596
rect 25278 -17658 25312 -17596
rect 24053 -17730 24069 -17696
rect 24445 -17730 24461 -17696
rect 24689 -17730 24705 -17696
rect 25081 -17730 25097 -17696
rect 23976 -17758 24010 -17742
rect 23976 -18542 24010 -18526
rect 24504 -17758 24538 -17742
rect 24504 -18542 24538 -18526
rect 24612 -17758 24646 -17742
rect 24612 -18542 24646 -18526
rect 25140 -17758 25174 -17742
rect 25140 -18542 25174 -18526
rect 24053 -18588 24069 -18554
rect 24445 -18588 24461 -18554
rect 24689 -18588 24705 -18554
rect 25081 -18588 25097 -18554
rect 23838 -18688 23872 -18626
rect 25278 -18688 25312 -18626
rect 23838 -18722 23934 -18688
rect 25216 -18722 25312 -18688
rect 25438 -17070 25534 -17036
rect 26816 -17070 26912 -17036
rect 25438 -17132 25472 -17070
rect 26878 -17132 26912 -17070
rect 25653 -17204 25669 -17170
rect 26045 -17204 26061 -17170
rect 26289 -17204 26305 -17170
rect 26681 -17204 26697 -17170
rect 25576 -17232 25610 -17216
rect 25576 -17416 25610 -17400
rect 26104 -17232 26138 -17216
rect 26104 -17416 26138 -17400
rect 26212 -17232 26246 -17216
rect 26212 -17416 26246 -17400
rect 26740 -17232 26774 -17216
rect 26740 -17416 26774 -17400
rect 25653 -17462 25669 -17428
rect 26045 -17462 26061 -17428
rect 26289 -17462 26305 -17428
rect 26681 -17462 26697 -17428
rect 25438 -17562 25472 -17500
rect 26878 -17562 26912 -17500
rect 25438 -17596 25534 -17562
rect 26816 -17596 26912 -17562
rect 25438 -17658 25472 -17596
rect 26878 -17658 26912 -17596
rect 25653 -17730 25669 -17696
rect 26045 -17730 26061 -17696
rect 26289 -17730 26305 -17696
rect 26681 -17730 26697 -17696
rect 25576 -17758 25610 -17742
rect 25576 -18542 25610 -18526
rect 26104 -17758 26138 -17742
rect 26104 -18542 26138 -18526
rect 26212 -17758 26246 -17742
rect 26212 -18542 26246 -18526
rect 26740 -17758 26774 -17742
rect 26740 -18542 26774 -18526
rect 25653 -18588 25669 -18554
rect 26045 -18588 26061 -18554
rect 26289 -18588 26305 -18554
rect 26681 -18588 26697 -18554
rect 25438 -18688 25472 -18626
rect 26878 -18688 26912 -18626
rect 25438 -18722 25534 -18688
rect 26816 -18722 26912 -18688
rect 27038 -17070 27134 -17036
rect 28416 -17070 28512 -17036
rect 27038 -17132 27072 -17070
rect 28478 -17132 28512 -17070
rect 27253 -17204 27269 -17170
rect 27645 -17204 27661 -17170
rect 27889 -17204 27905 -17170
rect 28281 -17204 28297 -17170
rect 27176 -17232 27210 -17216
rect 27176 -17416 27210 -17400
rect 27704 -17232 27738 -17216
rect 27704 -17416 27738 -17400
rect 27812 -17232 27846 -17216
rect 27812 -17416 27846 -17400
rect 28340 -17232 28374 -17216
rect 28340 -17416 28374 -17400
rect 27253 -17462 27269 -17428
rect 27645 -17462 27661 -17428
rect 27889 -17462 27905 -17428
rect 28281 -17462 28297 -17428
rect 27038 -17562 27072 -17500
rect 28478 -17562 28512 -17500
rect 27038 -17596 27134 -17562
rect 28416 -17596 28512 -17562
rect 27038 -17658 27072 -17596
rect 28478 -17658 28512 -17596
rect 27253 -17730 27269 -17696
rect 27645 -17730 27661 -17696
rect 27889 -17730 27905 -17696
rect 28281 -17730 28297 -17696
rect 27176 -17758 27210 -17742
rect 27176 -18542 27210 -18526
rect 27704 -17758 27738 -17742
rect 27704 -18542 27738 -18526
rect 27812 -17758 27846 -17742
rect 27812 -18542 27846 -18526
rect 28340 -17758 28374 -17742
rect 28340 -18542 28374 -18526
rect 27253 -18588 27269 -18554
rect 27645 -18588 27661 -18554
rect 27889 -18588 27905 -18554
rect 28281 -18588 28297 -18554
rect 27038 -18688 27072 -18626
rect 28478 -18688 28512 -18626
rect 27038 -18722 27134 -18688
rect 28416 -18722 28512 -18688
rect 28638 -17070 28734 -17036
rect 30016 -17070 30112 -17036
rect 28638 -17132 28672 -17070
rect 30078 -17132 30112 -17070
rect 28853 -17204 28869 -17170
rect 29245 -17204 29261 -17170
rect 29489 -17204 29505 -17170
rect 29881 -17204 29897 -17170
rect 28776 -17232 28810 -17216
rect 28776 -17416 28810 -17400
rect 29304 -17232 29338 -17216
rect 29304 -17416 29338 -17400
rect 29412 -17232 29446 -17216
rect 29412 -17416 29446 -17400
rect 29940 -17232 29974 -17216
rect 29940 -17416 29974 -17400
rect 28853 -17462 28869 -17428
rect 29245 -17462 29261 -17428
rect 29489 -17462 29505 -17428
rect 29881 -17462 29897 -17428
rect 28638 -17562 28672 -17500
rect 30078 -17562 30112 -17500
rect 28638 -17596 28734 -17562
rect 30016 -17596 30112 -17562
rect 28638 -17658 28672 -17596
rect 30078 -17658 30112 -17596
rect 28853 -17730 28869 -17696
rect 29245 -17730 29261 -17696
rect 29489 -17730 29505 -17696
rect 29881 -17730 29897 -17696
rect 28776 -17758 28810 -17742
rect 28776 -18542 28810 -18526
rect 29304 -17758 29338 -17742
rect 29304 -18542 29338 -18526
rect 29412 -17758 29446 -17742
rect 29412 -18542 29446 -18526
rect 29940 -17758 29974 -17742
rect 29940 -18542 29974 -18526
rect 28853 -18588 28869 -18554
rect 29245 -18588 29261 -18554
rect 29489 -18588 29505 -18554
rect 29881 -18588 29897 -18554
rect 28638 -18688 28672 -18626
rect 30078 -18688 30112 -18626
rect 28638 -18722 28734 -18688
rect 30016 -18722 30112 -18688
rect 30238 -17070 30334 -17036
rect 31616 -17070 31712 -17036
rect 30238 -17132 30272 -17070
rect 31678 -17132 31712 -17070
rect 30453 -17204 30469 -17170
rect 30845 -17204 30861 -17170
rect 31089 -17204 31105 -17170
rect 31481 -17204 31497 -17170
rect 30376 -17232 30410 -17216
rect 30376 -17416 30410 -17400
rect 30904 -17232 30938 -17216
rect 30904 -17416 30938 -17400
rect 31012 -17232 31046 -17216
rect 31012 -17416 31046 -17400
rect 31540 -17232 31574 -17216
rect 31540 -17416 31574 -17400
rect 30453 -17462 30469 -17428
rect 30845 -17462 30861 -17428
rect 31089 -17462 31105 -17428
rect 31481 -17462 31497 -17428
rect 30238 -17562 30272 -17500
rect 31678 -17562 31712 -17500
rect 30238 -17596 30334 -17562
rect 31616 -17596 31712 -17562
rect 30238 -17658 30272 -17596
rect 31678 -17658 31712 -17596
rect 30453 -17730 30469 -17696
rect 30845 -17730 30861 -17696
rect 31089 -17730 31105 -17696
rect 31481 -17730 31497 -17696
rect 30376 -17758 30410 -17742
rect 30376 -18542 30410 -18526
rect 30904 -17758 30938 -17742
rect 30904 -18542 30938 -18526
rect 31012 -17758 31046 -17742
rect 31012 -18542 31046 -18526
rect 31540 -17758 31574 -17742
rect 31540 -18542 31574 -18526
rect 30453 -18588 30469 -18554
rect 30845 -18588 30861 -18554
rect 31089 -18588 31105 -18554
rect 31481 -18588 31497 -18554
rect 30238 -18688 30272 -18626
rect 31678 -18688 31712 -18626
rect 30238 -18722 30334 -18688
rect 31616 -18722 31712 -18688
rect 31838 -17070 31934 -17036
rect 33216 -17070 33312 -17036
rect 31838 -17132 31872 -17070
rect 33278 -17132 33312 -17070
rect 32053 -17204 32069 -17170
rect 32445 -17204 32461 -17170
rect 32689 -17204 32705 -17170
rect 33081 -17204 33097 -17170
rect 31976 -17232 32010 -17216
rect 31976 -17416 32010 -17400
rect 32504 -17232 32538 -17216
rect 32504 -17416 32538 -17400
rect 32612 -17232 32646 -17216
rect 32612 -17416 32646 -17400
rect 33140 -17232 33174 -17216
rect 33140 -17416 33174 -17400
rect 32053 -17462 32069 -17428
rect 32445 -17462 32461 -17428
rect 32689 -17462 32705 -17428
rect 33081 -17462 33097 -17428
rect 31838 -17562 31872 -17500
rect 33278 -17562 33312 -17500
rect 31838 -17596 31934 -17562
rect 33216 -17596 33312 -17562
rect 31838 -17658 31872 -17596
rect 33278 -17658 33312 -17596
rect 32053 -17730 32069 -17696
rect 32445 -17730 32461 -17696
rect 32689 -17730 32705 -17696
rect 33081 -17730 33097 -17696
rect 31976 -17758 32010 -17742
rect 31976 -18542 32010 -18526
rect 32504 -17758 32538 -17742
rect 32504 -18542 32538 -18526
rect 32612 -17758 32646 -17742
rect 32612 -18542 32646 -18526
rect 33140 -17758 33174 -17742
rect 33140 -18542 33174 -18526
rect 32053 -18588 32069 -18554
rect 32445 -18588 32461 -18554
rect 32689 -18588 32705 -18554
rect 33081 -18588 33097 -18554
rect 31838 -18688 31872 -18626
rect 33278 -18688 33312 -18626
rect 31838 -18722 31934 -18688
rect 33216 -18722 33312 -18688
rect 33438 -17070 33534 -17036
rect 34816 -17070 34912 -17036
rect 33438 -17132 33472 -17070
rect 34878 -17132 34912 -17070
rect 33653 -17204 33669 -17170
rect 34045 -17204 34061 -17170
rect 34289 -17204 34305 -17170
rect 34681 -17204 34697 -17170
rect 33576 -17232 33610 -17216
rect 33576 -17416 33610 -17400
rect 34104 -17232 34138 -17216
rect 34104 -17416 34138 -17400
rect 34212 -17232 34246 -17216
rect 34212 -17416 34246 -17400
rect 34740 -17232 34774 -17216
rect 34740 -17416 34774 -17400
rect 33653 -17462 33669 -17428
rect 34045 -17462 34061 -17428
rect 34289 -17462 34305 -17428
rect 34681 -17462 34697 -17428
rect 33438 -17562 33472 -17500
rect 34878 -17562 34912 -17500
rect 33438 -17596 33534 -17562
rect 34816 -17596 34912 -17562
rect 33438 -17658 33472 -17596
rect 34878 -17658 34912 -17596
rect 33653 -17730 33669 -17696
rect 34045 -17730 34061 -17696
rect 34289 -17730 34305 -17696
rect 34681 -17730 34697 -17696
rect 33576 -17758 33610 -17742
rect 33576 -18542 33610 -18526
rect 34104 -17758 34138 -17742
rect 34104 -18542 34138 -18526
rect 34212 -17758 34246 -17742
rect 34212 -18542 34246 -18526
rect 34740 -17758 34774 -17742
rect 34740 -18542 34774 -18526
rect 33653 -18588 33669 -18554
rect 34045 -18588 34061 -18554
rect 34289 -18588 34305 -18554
rect 34681 -18588 34697 -18554
rect 33438 -18688 33472 -18626
rect 34878 -18688 34912 -18626
rect 33438 -18722 33534 -18688
rect 34816 -18722 34912 -18688
rect 35038 -17070 35134 -17036
rect 36416 -17070 36734 -17036
rect 38016 -17070 38112 -17036
rect 35038 -17132 35072 -17070
rect 36478 -17132 38112 -17070
rect 35253 -17204 35269 -17170
rect 35645 -17204 35661 -17170
rect 35889 -17204 35905 -17170
rect 36281 -17204 36297 -17170
rect 35176 -17232 35210 -17216
rect 35176 -17416 35210 -17400
rect 35704 -17232 35738 -17216
rect 35704 -17416 35738 -17400
rect 35812 -17232 35846 -17216
rect 35812 -17416 35846 -17400
rect 36340 -17232 36374 -17216
rect 36340 -17416 36374 -17400
rect 35253 -17462 35269 -17428
rect 35645 -17462 35661 -17428
rect 35889 -17462 35905 -17428
rect 36281 -17462 36297 -17428
rect 35038 -17562 35072 -17500
rect 36512 -17500 36638 -17132
rect 36672 -17170 38078 -17132
rect 36672 -17204 36869 -17170
rect 37245 -17204 37505 -17170
rect 37881 -17204 38078 -17170
rect 36672 -17232 38078 -17204
rect 36672 -17400 36776 -17232
rect 36810 -17400 37304 -17232
rect 37338 -17400 37412 -17232
rect 37446 -17400 37940 -17232
rect 37974 -17400 38078 -17232
rect 36672 -17428 38078 -17400
rect 36672 -17462 36869 -17428
rect 37245 -17462 37505 -17428
rect 37881 -17462 38078 -17428
rect 36672 -17500 38078 -17462
rect 36478 -17562 38112 -17500
rect 35038 -17596 35134 -17562
rect 36416 -17596 36734 -17562
rect 38016 -17596 38112 -17562
rect 35038 -17658 35072 -17596
rect 36478 -17658 38112 -17596
rect 35253 -17730 35269 -17696
rect 35645 -17730 35661 -17696
rect 35889 -17730 35905 -17696
rect 36281 -17730 36297 -17696
rect 35176 -17758 35210 -17742
rect 35176 -18542 35210 -18526
rect 35704 -17758 35738 -17742
rect 35704 -18542 35738 -18526
rect 35812 -17758 35846 -17742
rect 35812 -18542 35846 -18526
rect 36340 -17758 36374 -17742
rect 36340 -18542 36374 -18526
rect 35253 -18588 35269 -18554
rect 35645 -18588 35661 -18554
rect 35889 -18588 35905 -18554
rect 36281 -18588 36297 -18554
rect 35038 -18688 35072 -18626
rect 36512 -18626 36638 -17658
rect 36672 -17696 38078 -17658
rect 36672 -17730 36869 -17696
rect 37245 -17730 37505 -17696
rect 37881 -17730 38078 -17696
rect 36672 -17758 38078 -17730
rect 36672 -18526 36776 -17758
rect 36810 -18526 37304 -17758
rect 37338 -18526 37412 -17758
rect 37446 -18526 37940 -17758
rect 37974 -18526 38078 -17758
rect 36672 -18554 38078 -18526
rect 36672 -18588 36869 -18554
rect 37245 -18588 37505 -18554
rect 37881 -18588 38078 -18554
rect 36672 -18626 38078 -18588
rect 36478 -18688 38112 -18626
rect 35038 -18722 35134 -18688
rect 36416 -18722 36734 -18688
rect 38016 -18722 38112 -18688
rect -140 -18836 1460 -18722
rect 36500 -18836 38100 -18722
rect -162 -18870 -66 -18836
rect 1216 -18870 1534 -18836
rect 2816 -18870 2912 -18836
rect -162 -18932 1472 -18870
rect -128 -18970 1278 -18932
rect -128 -19004 69 -18970
rect 445 -19004 705 -18970
rect 1081 -19004 1278 -18970
rect -128 -19032 1278 -19004
rect -128 -19200 -24 -19032
rect 10 -19200 504 -19032
rect 538 -19200 612 -19032
rect 646 -19200 1140 -19032
rect 1174 -19200 1278 -19032
rect -128 -19228 1278 -19200
rect -128 -19262 69 -19228
rect 445 -19262 705 -19228
rect 1081 -19262 1278 -19228
rect -128 -19300 1278 -19262
rect 1312 -19300 1438 -18932
rect 2878 -18932 2912 -18870
rect 1653 -19004 1669 -18970
rect 2045 -19004 2061 -18970
rect 2289 -19004 2305 -18970
rect 2681 -19004 2697 -18970
rect 1576 -19032 1610 -19016
rect 1576 -19216 1610 -19200
rect 2104 -19032 2138 -19016
rect 2104 -19216 2138 -19200
rect 2212 -19032 2246 -19016
rect 2212 -19216 2246 -19200
rect 2740 -19032 2774 -19016
rect 2740 -19216 2774 -19200
rect 1653 -19262 1669 -19228
rect 2045 -19262 2061 -19228
rect 2289 -19262 2305 -19228
rect 2681 -19262 2697 -19228
rect -162 -19362 1472 -19300
rect 2878 -19362 2912 -19300
rect -162 -19396 -66 -19362
rect 1216 -19396 1534 -19362
rect 2816 -19396 2912 -19362
rect -162 -19458 1472 -19396
rect -128 -19496 1278 -19458
rect -128 -19530 69 -19496
rect 445 -19530 705 -19496
rect 1081 -19530 1278 -19496
rect -128 -19558 1278 -19530
rect -128 -20326 -24 -19558
rect 10 -20326 504 -19558
rect 538 -20326 612 -19558
rect 646 -20326 1140 -19558
rect 1174 -20326 1278 -19558
rect -128 -20354 1278 -20326
rect -128 -20388 69 -20354
rect 445 -20388 705 -20354
rect 1081 -20388 1278 -20354
rect -128 -20426 1278 -20388
rect 1312 -20426 1438 -19458
rect 2878 -19458 2912 -19396
rect 1653 -19530 1669 -19496
rect 2045 -19530 2061 -19496
rect 2289 -19530 2305 -19496
rect 2681 -19530 2697 -19496
rect 1576 -19558 1610 -19542
rect 1576 -20342 1610 -20326
rect 2104 -19558 2138 -19542
rect 2104 -20342 2138 -20326
rect 2212 -19558 2246 -19542
rect 2212 -20342 2246 -20326
rect 2740 -19558 2774 -19542
rect 2740 -20342 2774 -20326
rect 1653 -20388 1669 -20354
rect 2045 -20388 2061 -20354
rect 2289 -20388 2305 -20354
rect 2681 -20388 2697 -20354
rect -162 -20488 1472 -20426
rect 2878 -20488 2912 -20426
rect -162 -20522 -66 -20488
rect 1216 -20522 1534 -20488
rect 2816 -20522 2912 -20488
rect 3038 -18870 3134 -18836
rect 4416 -18870 4512 -18836
rect 3038 -18932 3072 -18870
rect 4478 -18932 4512 -18870
rect 3253 -19004 3269 -18970
rect 3645 -19004 3661 -18970
rect 3889 -19004 3905 -18970
rect 4281 -19004 4297 -18970
rect 3176 -19032 3210 -19016
rect 3176 -19216 3210 -19200
rect 3704 -19032 3738 -19016
rect 3704 -19216 3738 -19200
rect 3812 -19032 3846 -19016
rect 3812 -19216 3846 -19200
rect 4340 -19032 4374 -19016
rect 4340 -19216 4374 -19200
rect 3253 -19262 3269 -19228
rect 3645 -19262 3661 -19228
rect 3889 -19262 3905 -19228
rect 4281 -19262 4297 -19228
rect 3038 -19362 3072 -19300
rect 4478 -19362 4512 -19300
rect 3038 -19396 3134 -19362
rect 4416 -19396 4512 -19362
rect 3038 -19458 3072 -19396
rect 4478 -19458 4512 -19396
rect 3253 -19530 3269 -19496
rect 3645 -19530 3661 -19496
rect 3889 -19530 3905 -19496
rect 4281 -19530 4297 -19496
rect 3176 -19558 3210 -19542
rect 3176 -20342 3210 -20326
rect 3704 -19558 3738 -19542
rect 3704 -20342 3738 -20326
rect 3812 -19558 3846 -19542
rect 3812 -20342 3846 -20326
rect 4340 -19558 4374 -19542
rect 4340 -20342 4374 -20326
rect 3253 -20388 3269 -20354
rect 3645 -20388 3661 -20354
rect 3889 -20388 3905 -20354
rect 4281 -20388 4297 -20354
rect 3038 -20488 3072 -20426
rect 4478 -20488 4512 -20426
rect 3038 -20522 3134 -20488
rect 4416 -20522 4512 -20488
rect 4638 -18870 4734 -18836
rect 6016 -18870 6112 -18836
rect 4638 -18932 4672 -18870
rect 6078 -18932 6112 -18870
rect 4853 -19004 4869 -18970
rect 5245 -19004 5261 -18970
rect 5489 -19004 5505 -18970
rect 5881 -19004 5897 -18970
rect 4776 -19032 4810 -19016
rect 4776 -19216 4810 -19200
rect 5304 -19032 5338 -19016
rect 5304 -19216 5338 -19200
rect 5412 -19032 5446 -19016
rect 5412 -19216 5446 -19200
rect 5940 -19032 5974 -19016
rect 5940 -19216 5974 -19200
rect 4853 -19262 4869 -19228
rect 5245 -19262 5261 -19228
rect 5489 -19262 5505 -19228
rect 5881 -19262 5897 -19228
rect 4638 -19362 4672 -19300
rect 6078 -19362 6112 -19300
rect 4638 -19396 4734 -19362
rect 6016 -19396 6112 -19362
rect 4638 -19458 4672 -19396
rect 6078 -19458 6112 -19396
rect 4853 -19530 4869 -19496
rect 5245 -19530 5261 -19496
rect 5489 -19530 5505 -19496
rect 5881 -19530 5897 -19496
rect 4776 -19558 4810 -19542
rect 4776 -20342 4810 -20326
rect 5304 -19558 5338 -19542
rect 5304 -20342 5338 -20326
rect 5412 -19558 5446 -19542
rect 5412 -20342 5446 -20326
rect 5940 -19558 5974 -19542
rect 5940 -20342 5974 -20326
rect 4853 -20388 4869 -20354
rect 5245 -20388 5261 -20354
rect 5489 -20388 5505 -20354
rect 5881 -20388 5897 -20354
rect 4638 -20488 4672 -20426
rect 6078 -20488 6112 -20426
rect 4638 -20522 4734 -20488
rect 6016 -20522 6112 -20488
rect 6238 -18870 6334 -18836
rect 7616 -18870 7712 -18836
rect 6238 -18932 6272 -18870
rect 7678 -18932 7712 -18870
rect 6453 -19004 6469 -18970
rect 6845 -19004 6861 -18970
rect 7089 -19004 7105 -18970
rect 7481 -19004 7497 -18970
rect 6376 -19032 6410 -19016
rect 6376 -19216 6410 -19200
rect 6904 -19032 6938 -19016
rect 6904 -19216 6938 -19200
rect 7012 -19032 7046 -19016
rect 7012 -19216 7046 -19200
rect 7540 -19032 7574 -19016
rect 7540 -19216 7574 -19200
rect 6453 -19262 6469 -19228
rect 6845 -19262 6861 -19228
rect 7089 -19262 7105 -19228
rect 7481 -19262 7497 -19228
rect 6238 -19362 6272 -19300
rect 7678 -19362 7712 -19300
rect 6238 -19396 6334 -19362
rect 7616 -19396 7712 -19362
rect 6238 -19458 6272 -19396
rect 7678 -19458 7712 -19396
rect 6453 -19530 6469 -19496
rect 6845 -19530 6861 -19496
rect 7089 -19530 7105 -19496
rect 7481 -19530 7497 -19496
rect 6376 -19558 6410 -19542
rect 6376 -20342 6410 -20326
rect 6904 -19558 6938 -19542
rect 6904 -20342 6938 -20326
rect 7012 -19558 7046 -19542
rect 7012 -20342 7046 -20326
rect 7540 -19558 7574 -19542
rect 7540 -20342 7574 -20326
rect 6453 -20388 6469 -20354
rect 6845 -20388 6861 -20354
rect 7089 -20388 7105 -20354
rect 7481 -20388 7497 -20354
rect 6238 -20488 6272 -20426
rect 7678 -20488 7712 -20426
rect 6238 -20522 6334 -20488
rect 7616 -20522 7712 -20488
rect 7838 -18870 7934 -18836
rect 9216 -18870 9312 -18836
rect 7838 -18932 7872 -18870
rect 9278 -18932 9312 -18870
rect 8053 -19004 8069 -18970
rect 8445 -19004 8461 -18970
rect 8689 -19004 8705 -18970
rect 9081 -19004 9097 -18970
rect 7976 -19032 8010 -19016
rect 7976 -19216 8010 -19200
rect 8504 -19032 8538 -19016
rect 8504 -19216 8538 -19200
rect 8612 -19032 8646 -19016
rect 8612 -19216 8646 -19200
rect 9140 -19032 9174 -19016
rect 9140 -19216 9174 -19200
rect 8053 -19262 8069 -19228
rect 8445 -19262 8461 -19228
rect 8689 -19262 8705 -19228
rect 9081 -19262 9097 -19228
rect 7838 -19362 7872 -19300
rect 9278 -19362 9312 -19300
rect 7838 -19396 7934 -19362
rect 9216 -19396 9312 -19362
rect 7838 -19458 7872 -19396
rect 9278 -19458 9312 -19396
rect 8053 -19530 8069 -19496
rect 8445 -19530 8461 -19496
rect 8689 -19530 8705 -19496
rect 9081 -19530 9097 -19496
rect 7976 -19558 8010 -19542
rect 7976 -20342 8010 -20326
rect 8504 -19558 8538 -19542
rect 8504 -20342 8538 -20326
rect 8612 -19558 8646 -19542
rect 8612 -20342 8646 -20326
rect 9140 -19558 9174 -19542
rect 9140 -20342 9174 -20326
rect 8053 -20388 8069 -20354
rect 8445 -20388 8461 -20354
rect 8689 -20388 8705 -20354
rect 9081 -20388 9097 -20354
rect 7838 -20488 7872 -20426
rect 9278 -20488 9312 -20426
rect 7838 -20522 7934 -20488
rect 9216 -20522 9312 -20488
rect 9438 -18870 9534 -18836
rect 10816 -18870 10912 -18836
rect 9438 -18932 9472 -18870
rect 10878 -18932 10912 -18870
rect 9653 -19004 9669 -18970
rect 10045 -19004 10061 -18970
rect 10289 -19004 10305 -18970
rect 10681 -19004 10697 -18970
rect 9576 -19032 9610 -19016
rect 9576 -19216 9610 -19200
rect 10104 -19032 10138 -19016
rect 10104 -19216 10138 -19200
rect 10212 -19032 10246 -19016
rect 10212 -19216 10246 -19200
rect 10740 -19032 10774 -19016
rect 10740 -19216 10774 -19200
rect 9653 -19262 9669 -19228
rect 10045 -19262 10061 -19228
rect 10289 -19262 10305 -19228
rect 10681 -19262 10697 -19228
rect 9438 -19362 9472 -19300
rect 10878 -19362 10912 -19300
rect 9438 -19396 9534 -19362
rect 10816 -19396 10912 -19362
rect 9438 -19458 9472 -19396
rect 10878 -19458 10912 -19396
rect 9653 -19530 9669 -19496
rect 10045 -19530 10061 -19496
rect 10289 -19530 10305 -19496
rect 10681 -19530 10697 -19496
rect 9576 -19558 9610 -19542
rect 9576 -20342 9610 -20326
rect 10104 -19558 10138 -19542
rect 10104 -20342 10138 -20326
rect 10212 -19558 10246 -19542
rect 10212 -20342 10246 -20326
rect 10740 -19558 10774 -19542
rect 10740 -20342 10774 -20326
rect 9653 -20388 9669 -20354
rect 10045 -20388 10061 -20354
rect 10289 -20388 10305 -20354
rect 10681 -20388 10697 -20354
rect 9438 -20488 9472 -20426
rect 10878 -20488 10912 -20426
rect 9438 -20522 9534 -20488
rect 10816 -20522 10912 -20488
rect 11038 -18870 11134 -18836
rect 12416 -18870 12512 -18836
rect 11038 -18932 11072 -18870
rect 12478 -18932 12512 -18870
rect 11253 -19004 11269 -18970
rect 11645 -19004 11661 -18970
rect 11889 -19004 11905 -18970
rect 12281 -19004 12297 -18970
rect 11176 -19032 11210 -19016
rect 11176 -19216 11210 -19200
rect 11704 -19032 11738 -19016
rect 11704 -19216 11738 -19200
rect 11812 -19032 11846 -19016
rect 11812 -19216 11846 -19200
rect 12340 -19032 12374 -19016
rect 12340 -19216 12374 -19200
rect 11253 -19262 11269 -19228
rect 11645 -19262 11661 -19228
rect 11889 -19262 11905 -19228
rect 12281 -19262 12297 -19228
rect 11038 -19362 11072 -19300
rect 12478 -19362 12512 -19300
rect 11038 -19396 11134 -19362
rect 12416 -19396 12512 -19362
rect 11038 -19458 11072 -19396
rect 12478 -19458 12512 -19396
rect 11253 -19530 11269 -19496
rect 11645 -19530 11661 -19496
rect 11889 -19530 11905 -19496
rect 12281 -19530 12297 -19496
rect 11176 -19558 11210 -19542
rect 11176 -20342 11210 -20326
rect 11704 -19558 11738 -19542
rect 11704 -20342 11738 -20326
rect 11812 -19558 11846 -19542
rect 11812 -20342 11846 -20326
rect 12340 -19558 12374 -19542
rect 12340 -20342 12374 -20326
rect 11253 -20388 11269 -20354
rect 11645 -20388 11661 -20354
rect 11889 -20388 11905 -20354
rect 12281 -20388 12297 -20354
rect 11038 -20488 11072 -20426
rect 12478 -20488 12512 -20426
rect 11038 -20522 11134 -20488
rect 12416 -20522 12512 -20488
rect 12638 -18870 12734 -18836
rect 14016 -18870 14112 -18836
rect 12638 -18932 12672 -18870
rect 14078 -18932 14112 -18870
rect 12853 -19004 12869 -18970
rect 13245 -19004 13261 -18970
rect 13489 -19004 13505 -18970
rect 13881 -19004 13897 -18970
rect 12776 -19032 12810 -19016
rect 12776 -19216 12810 -19200
rect 13304 -19032 13338 -19016
rect 13304 -19216 13338 -19200
rect 13412 -19032 13446 -19016
rect 13412 -19216 13446 -19200
rect 13940 -19032 13974 -19016
rect 13940 -19216 13974 -19200
rect 12853 -19262 12869 -19228
rect 13245 -19262 13261 -19228
rect 13489 -19262 13505 -19228
rect 13881 -19262 13897 -19228
rect 12638 -19362 12672 -19300
rect 14078 -19362 14112 -19300
rect 12638 -19396 12734 -19362
rect 14016 -19396 14112 -19362
rect 12638 -19458 12672 -19396
rect 14078 -19458 14112 -19396
rect 12853 -19530 12869 -19496
rect 13245 -19530 13261 -19496
rect 13489 -19530 13505 -19496
rect 13881 -19530 13897 -19496
rect 12776 -19558 12810 -19542
rect 12776 -20342 12810 -20326
rect 13304 -19558 13338 -19542
rect 13304 -20342 13338 -20326
rect 13412 -19558 13446 -19542
rect 13412 -20342 13446 -20326
rect 13940 -19558 13974 -19542
rect 13940 -20342 13974 -20326
rect 12853 -20388 12869 -20354
rect 13245 -20388 13261 -20354
rect 13489 -20388 13505 -20354
rect 13881 -20388 13897 -20354
rect 12638 -20488 12672 -20426
rect 14078 -20488 14112 -20426
rect 12638 -20522 12734 -20488
rect 14016 -20522 14112 -20488
rect 14238 -18870 14334 -18836
rect 15616 -18870 15712 -18836
rect 14238 -18932 14272 -18870
rect 15678 -18932 15712 -18870
rect 14453 -19004 14469 -18970
rect 14845 -19004 14861 -18970
rect 15089 -19004 15105 -18970
rect 15481 -19004 15497 -18970
rect 14376 -19032 14410 -19016
rect 14376 -19216 14410 -19200
rect 14904 -19032 14938 -19016
rect 14904 -19216 14938 -19200
rect 15012 -19032 15046 -19016
rect 15012 -19216 15046 -19200
rect 15540 -19032 15574 -19016
rect 15540 -19216 15574 -19200
rect 14453 -19262 14469 -19228
rect 14845 -19262 14861 -19228
rect 15089 -19262 15105 -19228
rect 15481 -19262 15497 -19228
rect 14238 -19362 14272 -19300
rect 15678 -19362 15712 -19300
rect 14238 -19396 14334 -19362
rect 15616 -19396 15712 -19362
rect 14238 -19458 14272 -19396
rect 15678 -19458 15712 -19396
rect 14453 -19530 14469 -19496
rect 14845 -19530 14861 -19496
rect 15089 -19530 15105 -19496
rect 15481 -19530 15497 -19496
rect 14376 -19558 14410 -19542
rect 14376 -20342 14410 -20326
rect 14904 -19558 14938 -19542
rect 14904 -20342 14938 -20326
rect 15012 -19558 15046 -19542
rect 15012 -20342 15046 -20326
rect 15540 -19558 15574 -19542
rect 15540 -20342 15574 -20326
rect 14453 -20388 14469 -20354
rect 14845 -20388 14861 -20354
rect 15089 -20388 15105 -20354
rect 15481 -20388 15497 -20354
rect 14238 -20488 14272 -20426
rect 15678 -20488 15712 -20426
rect 14238 -20522 14334 -20488
rect 15616 -20522 15712 -20488
rect 15838 -18870 15934 -18836
rect 17216 -18870 17312 -18836
rect 15838 -18932 15872 -18870
rect 17278 -18932 17312 -18870
rect 16053 -19004 16069 -18970
rect 16445 -19004 16461 -18970
rect 16689 -19004 16705 -18970
rect 17081 -19004 17097 -18970
rect 15976 -19032 16010 -19016
rect 15976 -19216 16010 -19200
rect 16504 -19032 16538 -19016
rect 16504 -19216 16538 -19200
rect 16612 -19032 16646 -19016
rect 16612 -19216 16646 -19200
rect 17140 -19032 17174 -19016
rect 17140 -19216 17174 -19200
rect 16053 -19262 16069 -19228
rect 16445 -19262 16461 -19228
rect 16689 -19262 16705 -19228
rect 17081 -19262 17097 -19228
rect 15838 -19362 15872 -19300
rect 17278 -19362 17312 -19300
rect 15838 -19396 15934 -19362
rect 17216 -19396 17312 -19362
rect 15838 -19458 15872 -19396
rect 17278 -19458 17312 -19396
rect 16053 -19530 16069 -19496
rect 16445 -19530 16461 -19496
rect 16689 -19530 16705 -19496
rect 17081 -19530 17097 -19496
rect 15976 -19558 16010 -19542
rect 15976 -20342 16010 -20326
rect 16504 -19558 16538 -19542
rect 16504 -20342 16538 -20326
rect 16612 -19558 16646 -19542
rect 16612 -20342 16646 -20326
rect 17140 -19558 17174 -19542
rect 17140 -20342 17174 -20326
rect 16053 -20388 16069 -20354
rect 16445 -20388 16461 -20354
rect 16689 -20388 16705 -20354
rect 17081 -20388 17097 -20354
rect 15838 -20488 15872 -20426
rect 17278 -20488 17312 -20426
rect 15838 -20522 15934 -20488
rect 17216 -20522 17312 -20488
rect 17438 -18870 17534 -18836
rect 18816 -18870 18912 -18836
rect 17438 -18932 17472 -18870
rect 18878 -18932 18912 -18870
rect 17653 -19004 17669 -18970
rect 18045 -19004 18061 -18970
rect 18289 -19004 18305 -18970
rect 18681 -19004 18697 -18970
rect 17576 -19032 17610 -19016
rect 17576 -19216 17610 -19200
rect 18104 -19032 18138 -19016
rect 18104 -19216 18138 -19200
rect 18212 -19032 18246 -19016
rect 18212 -19216 18246 -19200
rect 18740 -19032 18774 -19016
rect 18740 -19216 18774 -19200
rect 17653 -19262 17669 -19228
rect 18045 -19262 18061 -19228
rect 18289 -19262 18305 -19228
rect 18681 -19262 18697 -19228
rect 17438 -19362 17472 -19300
rect 18878 -19362 18912 -19300
rect 17438 -19396 17534 -19362
rect 18816 -19396 18912 -19362
rect 17438 -19458 17472 -19396
rect 18878 -19458 18912 -19396
rect 17653 -19530 17669 -19496
rect 18045 -19530 18061 -19496
rect 18289 -19530 18305 -19496
rect 18681 -19530 18697 -19496
rect 17576 -19558 17610 -19542
rect 17576 -20342 17610 -20326
rect 18104 -19558 18138 -19542
rect 18104 -20342 18138 -20326
rect 18212 -19558 18246 -19542
rect 18212 -20342 18246 -20326
rect 18740 -19558 18774 -19542
rect 18740 -20342 18774 -20326
rect 17653 -20388 17669 -20354
rect 18045 -20388 18061 -20354
rect 18289 -20388 18305 -20354
rect 18681 -20388 18697 -20354
rect 17438 -20488 17472 -20426
rect 18878 -20488 18912 -20426
rect 17438 -20522 17534 -20488
rect 18816 -20522 18912 -20488
rect 19038 -18870 19134 -18836
rect 20416 -18870 20512 -18836
rect 19038 -18932 19072 -18870
rect 20478 -18932 20512 -18870
rect 19253 -19004 19269 -18970
rect 19645 -19004 19661 -18970
rect 19889 -19004 19905 -18970
rect 20281 -19004 20297 -18970
rect 19176 -19032 19210 -19016
rect 19176 -19216 19210 -19200
rect 19704 -19032 19738 -19016
rect 19704 -19216 19738 -19200
rect 19812 -19032 19846 -19016
rect 19812 -19216 19846 -19200
rect 20340 -19032 20374 -19016
rect 20340 -19216 20374 -19200
rect 19253 -19262 19269 -19228
rect 19645 -19262 19661 -19228
rect 19889 -19262 19905 -19228
rect 20281 -19262 20297 -19228
rect 19038 -19362 19072 -19300
rect 20478 -19362 20512 -19300
rect 19038 -19396 19134 -19362
rect 20416 -19396 20512 -19362
rect 19038 -19458 19072 -19396
rect 20478 -19458 20512 -19396
rect 19253 -19530 19269 -19496
rect 19645 -19530 19661 -19496
rect 19889 -19530 19905 -19496
rect 20281 -19530 20297 -19496
rect 19176 -19558 19210 -19542
rect 19176 -20342 19210 -20326
rect 19704 -19558 19738 -19542
rect 19704 -20342 19738 -20326
rect 19812 -19558 19846 -19542
rect 19812 -20342 19846 -20326
rect 20340 -19558 20374 -19542
rect 20340 -20342 20374 -20326
rect 19253 -20388 19269 -20354
rect 19645 -20388 19661 -20354
rect 19889 -20388 19905 -20354
rect 20281 -20388 20297 -20354
rect 19038 -20488 19072 -20426
rect 20478 -20488 20512 -20426
rect 19038 -20522 19134 -20488
rect 20416 -20522 20512 -20488
rect 20638 -18870 20734 -18836
rect 22016 -18870 22112 -18836
rect 20638 -18932 20672 -18870
rect 22078 -18932 22112 -18870
rect 20853 -19004 20869 -18970
rect 21245 -19004 21261 -18970
rect 21489 -19004 21505 -18970
rect 21881 -19004 21897 -18970
rect 20776 -19032 20810 -19016
rect 20776 -19216 20810 -19200
rect 21304 -19032 21338 -19016
rect 21304 -19216 21338 -19200
rect 21412 -19032 21446 -19016
rect 21412 -19216 21446 -19200
rect 21940 -19032 21974 -19016
rect 21940 -19216 21974 -19200
rect 20853 -19262 20869 -19228
rect 21245 -19262 21261 -19228
rect 21489 -19262 21505 -19228
rect 21881 -19262 21897 -19228
rect 20638 -19362 20672 -19300
rect 22078 -19362 22112 -19300
rect 20638 -19396 20734 -19362
rect 22016 -19396 22112 -19362
rect 20638 -19458 20672 -19396
rect 22078 -19458 22112 -19396
rect 20853 -19530 20869 -19496
rect 21245 -19530 21261 -19496
rect 21489 -19530 21505 -19496
rect 21881 -19530 21897 -19496
rect 20776 -19558 20810 -19542
rect 20776 -20342 20810 -20326
rect 21304 -19558 21338 -19542
rect 21304 -20342 21338 -20326
rect 21412 -19558 21446 -19542
rect 21412 -20342 21446 -20326
rect 21940 -19558 21974 -19542
rect 21940 -20342 21974 -20326
rect 20853 -20388 20869 -20354
rect 21245 -20388 21261 -20354
rect 21489 -20388 21505 -20354
rect 21881 -20388 21897 -20354
rect 20638 -20488 20672 -20426
rect 22078 -20488 22112 -20426
rect 20638 -20522 20734 -20488
rect 22016 -20522 22112 -20488
rect 22238 -18870 22334 -18836
rect 23616 -18870 23712 -18836
rect 22238 -18932 22272 -18870
rect 23678 -18932 23712 -18870
rect 22453 -19004 22469 -18970
rect 22845 -19004 22861 -18970
rect 23089 -19004 23105 -18970
rect 23481 -19004 23497 -18970
rect 22376 -19032 22410 -19016
rect 22376 -19216 22410 -19200
rect 22904 -19032 22938 -19016
rect 22904 -19216 22938 -19200
rect 23012 -19032 23046 -19016
rect 23012 -19216 23046 -19200
rect 23540 -19032 23574 -19016
rect 23540 -19216 23574 -19200
rect 22453 -19262 22469 -19228
rect 22845 -19262 22861 -19228
rect 23089 -19262 23105 -19228
rect 23481 -19262 23497 -19228
rect 22238 -19362 22272 -19300
rect 23678 -19362 23712 -19300
rect 22238 -19396 22334 -19362
rect 23616 -19396 23712 -19362
rect 22238 -19458 22272 -19396
rect 23678 -19458 23712 -19396
rect 22453 -19530 22469 -19496
rect 22845 -19530 22861 -19496
rect 23089 -19530 23105 -19496
rect 23481 -19530 23497 -19496
rect 22376 -19558 22410 -19542
rect 22376 -20342 22410 -20326
rect 22904 -19558 22938 -19542
rect 22904 -20342 22938 -20326
rect 23012 -19558 23046 -19542
rect 23012 -20342 23046 -20326
rect 23540 -19558 23574 -19542
rect 23540 -20342 23574 -20326
rect 22453 -20388 22469 -20354
rect 22845 -20388 22861 -20354
rect 23089 -20388 23105 -20354
rect 23481 -20388 23497 -20354
rect 22238 -20488 22272 -20426
rect 23678 -20488 23712 -20426
rect 22238 -20522 22334 -20488
rect 23616 -20522 23712 -20488
rect 23838 -18870 23934 -18836
rect 25216 -18870 25312 -18836
rect 23838 -18932 23872 -18870
rect 25278 -18932 25312 -18870
rect 24053 -19004 24069 -18970
rect 24445 -19004 24461 -18970
rect 24689 -19004 24705 -18970
rect 25081 -19004 25097 -18970
rect 23976 -19032 24010 -19016
rect 23976 -19216 24010 -19200
rect 24504 -19032 24538 -19016
rect 24504 -19216 24538 -19200
rect 24612 -19032 24646 -19016
rect 24612 -19216 24646 -19200
rect 25140 -19032 25174 -19016
rect 25140 -19216 25174 -19200
rect 24053 -19262 24069 -19228
rect 24445 -19262 24461 -19228
rect 24689 -19262 24705 -19228
rect 25081 -19262 25097 -19228
rect 23838 -19362 23872 -19300
rect 25278 -19362 25312 -19300
rect 23838 -19396 23934 -19362
rect 25216 -19396 25312 -19362
rect 23838 -19458 23872 -19396
rect 25278 -19458 25312 -19396
rect 24053 -19530 24069 -19496
rect 24445 -19530 24461 -19496
rect 24689 -19530 24705 -19496
rect 25081 -19530 25097 -19496
rect 23976 -19558 24010 -19542
rect 23976 -20342 24010 -20326
rect 24504 -19558 24538 -19542
rect 24504 -20342 24538 -20326
rect 24612 -19558 24646 -19542
rect 24612 -20342 24646 -20326
rect 25140 -19558 25174 -19542
rect 25140 -20342 25174 -20326
rect 24053 -20388 24069 -20354
rect 24445 -20388 24461 -20354
rect 24689 -20388 24705 -20354
rect 25081 -20388 25097 -20354
rect 23838 -20488 23872 -20426
rect 25278 -20488 25312 -20426
rect 23838 -20522 23934 -20488
rect 25216 -20522 25312 -20488
rect 25438 -18870 25534 -18836
rect 26816 -18870 26912 -18836
rect 25438 -18932 25472 -18870
rect 26878 -18932 26912 -18870
rect 25653 -19004 25669 -18970
rect 26045 -19004 26061 -18970
rect 26289 -19004 26305 -18970
rect 26681 -19004 26697 -18970
rect 25576 -19032 25610 -19016
rect 25576 -19216 25610 -19200
rect 26104 -19032 26138 -19016
rect 26104 -19216 26138 -19200
rect 26212 -19032 26246 -19016
rect 26212 -19216 26246 -19200
rect 26740 -19032 26774 -19016
rect 26740 -19216 26774 -19200
rect 25653 -19262 25669 -19228
rect 26045 -19262 26061 -19228
rect 26289 -19262 26305 -19228
rect 26681 -19262 26697 -19228
rect 25438 -19362 25472 -19300
rect 26878 -19362 26912 -19300
rect 25438 -19396 25534 -19362
rect 26816 -19396 26912 -19362
rect 25438 -19458 25472 -19396
rect 26878 -19458 26912 -19396
rect 25653 -19530 25669 -19496
rect 26045 -19530 26061 -19496
rect 26289 -19530 26305 -19496
rect 26681 -19530 26697 -19496
rect 25576 -19558 25610 -19542
rect 25576 -20342 25610 -20326
rect 26104 -19558 26138 -19542
rect 26104 -20342 26138 -20326
rect 26212 -19558 26246 -19542
rect 26212 -20342 26246 -20326
rect 26740 -19558 26774 -19542
rect 26740 -20342 26774 -20326
rect 25653 -20388 25669 -20354
rect 26045 -20388 26061 -20354
rect 26289 -20388 26305 -20354
rect 26681 -20388 26697 -20354
rect 25438 -20488 25472 -20426
rect 26878 -20488 26912 -20426
rect 25438 -20522 25534 -20488
rect 26816 -20522 26912 -20488
rect 27038 -18870 27134 -18836
rect 28416 -18870 28512 -18836
rect 27038 -18932 27072 -18870
rect 28478 -18932 28512 -18870
rect 27253 -19004 27269 -18970
rect 27645 -19004 27661 -18970
rect 27889 -19004 27905 -18970
rect 28281 -19004 28297 -18970
rect 27176 -19032 27210 -19016
rect 27176 -19216 27210 -19200
rect 27704 -19032 27738 -19016
rect 27704 -19216 27738 -19200
rect 27812 -19032 27846 -19016
rect 27812 -19216 27846 -19200
rect 28340 -19032 28374 -19016
rect 28340 -19216 28374 -19200
rect 27253 -19262 27269 -19228
rect 27645 -19262 27661 -19228
rect 27889 -19262 27905 -19228
rect 28281 -19262 28297 -19228
rect 27038 -19362 27072 -19300
rect 28478 -19362 28512 -19300
rect 27038 -19396 27134 -19362
rect 28416 -19396 28512 -19362
rect 27038 -19458 27072 -19396
rect 28478 -19458 28512 -19396
rect 27253 -19530 27269 -19496
rect 27645 -19530 27661 -19496
rect 27889 -19530 27905 -19496
rect 28281 -19530 28297 -19496
rect 27176 -19558 27210 -19542
rect 27176 -20342 27210 -20326
rect 27704 -19558 27738 -19542
rect 27704 -20342 27738 -20326
rect 27812 -19558 27846 -19542
rect 27812 -20342 27846 -20326
rect 28340 -19558 28374 -19542
rect 28340 -20342 28374 -20326
rect 27253 -20388 27269 -20354
rect 27645 -20388 27661 -20354
rect 27889 -20388 27905 -20354
rect 28281 -20388 28297 -20354
rect 27038 -20488 27072 -20426
rect 28478 -20488 28512 -20426
rect 27038 -20522 27134 -20488
rect 28416 -20522 28512 -20488
rect 28638 -18870 28734 -18836
rect 30016 -18870 30112 -18836
rect 28638 -18932 28672 -18870
rect 30078 -18932 30112 -18870
rect 28853 -19004 28869 -18970
rect 29245 -19004 29261 -18970
rect 29489 -19004 29505 -18970
rect 29881 -19004 29897 -18970
rect 28776 -19032 28810 -19016
rect 28776 -19216 28810 -19200
rect 29304 -19032 29338 -19016
rect 29304 -19216 29338 -19200
rect 29412 -19032 29446 -19016
rect 29412 -19216 29446 -19200
rect 29940 -19032 29974 -19016
rect 29940 -19216 29974 -19200
rect 28853 -19262 28869 -19228
rect 29245 -19262 29261 -19228
rect 29489 -19262 29505 -19228
rect 29881 -19262 29897 -19228
rect 28638 -19362 28672 -19300
rect 30078 -19362 30112 -19300
rect 28638 -19396 28734 -19362
rect 30016 -19396 30112 -19362
rect 28638 -19458 28672 -19396
rect 30078 -19458 30112 -19396
rect 28853 -19530 28869 -19496
rect 29245 -19530 29261 -19496
rect 29489 -19530 29505 -19496
rect 29881 -19530 29897 -19496
rect 28776 -19558 28810 -19542
rect 28776 -20342 28810 -20326
rect 29304 -19558 29338 -19542
rect 29304 -20342 29338 -20326
rect 29412 -19558 29446 -19542
rect 29412 -20342 29446 -20326
rect 29940 -19558 29974 -19542
rect 29940 -20342 29974 -20326
rect 28853 -20388 28869 -20354
rect 29245 -20388 29261 -20354
rect 29489 -20388 29505 -20354
rect 29881 -20388 29897 -20354
rect 28638 -20488 28672 -20426
rect 30078 -20488 30112 -20426
rect 28638 -20522 28734 -20488
rect 30016 -20522 30112 -20488
rect 30238 -18870 30334 -18836
rect 31616 -18870 31712 -18836
rect 30238 -18932 30272 -18870
rect 31678 -18932 31712 -18870
rect 30453 -19004 30469 -18970
rect 30845 -19004 30861 -18970
rect 31089 -19004 31105 -18970
rect 31481 -19004 31497 -18970
rect 30376 -19032 30410 -19016
rect 30376 -19216 30410 -19200
rect 30904 -19032 30938 -19016
rect 30904 -19216 30938 -19200
rect 31012 -19032 31046 -19016
rect 31012 -19216 31046 -19200
rect 31540 -19032 31574 -19016
rect 31540 -19216 31574 -19200
rect 30453 -19262 30469 -19228
rect 30845 -19262 30861 -19228
rect 31089 -19262 31105 -19228
rect 31481 -19262 31497 -19228
rect 30238 -19362 30272 -19300
rect 31678 -19362 31712 -19300
rect 30238 -19396 30334 -19362
rect 31616 -19396 31712 -19362
rect 30238 -19458 30272 -19396
rect 31678 -19458 31712 -19396
rect 30453 -19530 30469 -19496
rect 30845 -19530 30861 -19496
rect 31089 -19530 31105 -19496
rect 31481 -19530 31497 -19496
rect 30376 -19558 30410 -19542
rect 30376 -20342 30410 -20326
rect 30904 -19558 30938 -19542
rect 30904 -20342 30938 -20326
rect 31012 -19558 31046 -19542
rect 31012 -20342 31046 -20326
rect 31540 -19558 31574 -19542
rect 31540 -20342 31574 -20326
rect 30453 -20388 30469 -20354
rect 30845 -20388 30861 -20354
rect 31089 -20388 31105 -20354
rect 31481 -20388 31497 -20354
rect 30238 -20488 30272 -20426
rect 31678 -20488 31712 -20426
rect 30238 -20522 30334 -20488
rect 31616 -20522 31712 -20488
rect 31838 -18870 31934 -18836
rect 33216 -18870 33312 -18836
rect 31838 -18932 31872 -18870
rect 33278 -18932 33312 -18870
rect 32053 -19004 32069 -18970
rect 32445 -19004 32461 -18970
rect 32689 -19004 32705 -18970
rect 33081 -19004 33097 -18970
rect 31976 -19032 32010 -19016
rect 31976 -19216 32010 -19200
rect 32504 -19032 32538 -19016
rect 32504 -19216 32538 -19200
rect 32612 -19032 32646 -19016
rect 32612 -19216 32646 -19200
rect 33140 -19032 33174 -19016
rect 33140 -19216 33174 -19200
rect 32053 -19262 32069 -19228
rect 32445 -19262 32461 -19228
rect 32689 -19262 32705 -19228
rect 33081 -19262 33097 -19228
rect 31838 -19362 31872 -19300
rect 33278 -19362 33312 -19300
rect 31838 -19396 31934 -19362
rect 33216 -19396 33312 -19362
rect 31838 -19458 31872 -19396
rect 33278 -19458 33312 -19396
rect 32053 -19530 32069 -19496
rect 32445 -19530 32461 -19496
rect 32689 -19530 32705 -19496
rect 33081 -19530 33097 -19496
rect 31976 -19558 32010 -19542
rect 31976 -20342 32010 -20326
rect 32504 -19558 32538 -19542
rect 32504 -20342 32538 -20326
rect 32612 -19558 32646 -19542
rect 32612 -20342 32646 -20326
rect 33140 -19558 33174 -19542
rect 33140 -20342 33174 -20326
rect 32053 -20388 32069 -20354
rect 32445 -20388 32461 -20354
rect 32689 -20388 32705 -20354
rect 33081 -20388 33097 -20354
rect 31838 -20488 31872 -20426
rect 33278 -20488 33312 -20426
rect 31838 -20522 31934 -20488
rect 33216 -20522 33312 -20488
rect 33438 -18870 33534 -18836
rect 34816 -18870 34912 -18836
rect 33438 -18932 33472 -18870
rect 34878 -18932 34912 -18870
rect 33653 -19004 33669 -18970
rect 34045 -19004 34061 -18970
rect 34289 -19004 34305 -18970
rect 34681 -19004 34697 -18970
rect 33576 -19032 33610 -19016
rect 33576 -19216 33610 -19200
rect 34104 -19032 34138 -19016
rect 34104 -19216 34138 -19200
rect 34212 -19032 34246 -19016
rect 34212 -19216 34246 -19200
rect 34740 -19032 34774 -19016
rect 34740 -19216 34774 -19200
rect 33653 -19262 33669 -19228
rect 34045 -19262 34061 -19228
rect 34289 -19262 34305 -19228
rect 34681 -19262 34697 -19228
rect 33438 -19362 33472 -19300
rect 34878 -19362 34912 -19300
rect 33438 -19396 33534 -19362
rect 34816 -19396 34912 -19362
rect 33438 -19458 33472 -19396
rect 34878 -19458 34912 -19396
rect 33653 -19530 33669 -19496
rect 34045 -19530 34061 -19496
rect 34289 -19530 34305 -19496
rect 34681 -19530 34697 -19496
rect 33576 -19558 33610 -19542
rect 33576 -20342 33610 -20326
rect 34104 -19558 34138 -19542
rect 34104 -20342 34138 -20326
rect 34212 -19558 34246 -19542
rect 34212 -20342 34246 -20326
rect 34740 -19558 34774 -19542
rect 34740 -20342 34774 -20326
rect 33653 -20388 33669 -20354
rect 34045 -20388 34061 -20354
rect 34289 -20388 34305 -20354
rect 34681 -20388 34697 -20354
rect 33438 -20488 33472 -20426
rect 34878 -20488 34912 -20426
rect 33438 -20522 33534 -20488
rect 34816 -20522 34912 -20488
rect 35038 -18870 35134 -18836
rect 36416 -18870 36734 -18836
rect 38016 -18870 38112 -18836
rect 35038 -18932 35072 -18870
rect 36478 -18932 38112 -18870
rect 35253 -19004 35269 -18970
rect 35645 -19004 35661 -18970
rect 35889 -19004 35905 -18970
rect 36281 -19004 36297 -18970
rect 35176 -19032 35210 -19016
rect 35176 -19216 35210 -19200
rect 35704 -19032 35738 -19016
rect 35704 -19216 35738 -19200
rect 35812 -19032 35846 -19016
rect 35812 -19216 35846 -19200
rect 36340 -19032 36374 -19016
rect 36340 -19216 36374 -19200
rect 35253 -19262 35269 -19228
rect 35645 -19262 35661 -19228
rect 35889 -19262 35905 -19228
rect 36281 -19262 36297 -19228
rect 35038 -19362 35072 -19300
rect 36512 -19300 36638 -18932
rect 36672 -18970 38078 -18932
rect 36672 -19004 36869 -18970
rect 37245 -19004 37505 -18970
rect 37881 -19004 38078 -18970
rect 36672 -19032 38078 -19004
rect 36672 -19200 36776 -19032
rect 36810 -19200 37304 -19032
rect 37338 -19200 37412 -19032
rect 37446 -19200 37940 -19032
rect 37974 -19200 38078 -19032
rect 36672 -19228 38078 -19200
rect 36672 -19262 36869 -19228
rect 37245 -19262 37505 -19228
rect 37881 -19262 38078 -19228
rect 36672 -19300 38078 -19262
rect 36478 -19362 38112 -19300
rect 35038 -19396 35134 -19362
rect 36416 -19396 36734 -19362
rect 38016 -19396 38112 -19362
rect 35038 -19458 35072 -19396
rect 36478 -19458 38112 -19396
rect 35253 -19530 35269 -19496
rect 35645 -19530 35661 -19496
rect 35889 -19530 35905 -19496
rect 36281 -19530 36297 -19496
rect 35176 -19558 35210 -19542
rect 35176 -20342 35210 -20326
rect 35704 -19558 35738 -19542
rect 35704 -20342 35738 -20326
rect 35812 -19558 35846 -19542
rect 35812 -20342 35846 -20326
rect 36340 -19558 36374 -19542
rect 36340 -20342 36374 -20326
rect 35253 -20388 35269 -20354
rect 35645 -20388 35661 -20354
rect 35889 -20388 35905 -20354
rect 36281 -20388 36297 -20354
rect 35038 -20488 35072 -20426
rect 36512 -20426 36638 -19458
rect 36672 -19496 38078 -19458
rect 36672 -19530 36869 -19496
rect 37245 -19530 37505 -19496
rect 37881 -19530 38078 -19496
rect 36672 -19558 38078 -19530
rect 36672 -20326 36776 -19558
rect 36810 -20326 37304 -19558
rect 37338 -20326 37412 -19558
rect 37446 -20326 37940 -19558
rect 37974 -20326 38078 -19558
rect 36672 -20354 38078 -20326
rect 36672 -20388 36869 -20354
rect 37245 -20388 37505 -20354
rect 37881 -20388 38078 -20354
rect 36672 -20426 38078 -20388
rect 36478 -20488 38112 -20426
rect 35038 -20522 35134 -20488
rect 36416 -20522 36734 -20488
rect 38016 -20522 38112 -20488
rect -140 -20636 1460 -20522
rect 36500 -20636 38100 -20522
rect -162 -20670 -66 -20636
rect 1216 -20670 1534 -20636
rect 2816 -20670 2912 -20636
rect -162 -20732 1472 -20670
rect -128 -20770 1278 -20732
rect -128 -20804 69 -20770
rect 445 -20804 705 -20770
rect 1081 -20804 1278 -20770
rect -128 -20832 1278 -20804
rect -128 -21000 -24 -20832
rect 10 -21000 504 -20832
rect 538 -21000 612 -20832
rect 646 -21000 1140 -20832
rect 1174 -21000 1278 -20832
rect -128 -21028 1278 -21000
rect -128 -21062 69 -21028
rect 445 -21062 705 -21028
rect 1081 -21062 1278 -21028
rect -128 -21100 1278 -21062
rect 1312 -21100 1438 -20732
rect 2878 -20732 2912 -20670
rect 1653 -20804 1669 -20770
rect 2045 -20804 2061 -20770
rect 2289 -20804 2305 -20770
rect 2681 -20804 2697 -20770
rect 1576 -20832 1610 -20816
rect 1576 -21016 1610 -21000
rect 2104 -20832 2138 -20816
rect 2104 -21016 2138 -21000
rect 2212 -20832 2246 -20816
rect 2212 -21016 2246 -21000
rect 2740 -20832 2774 -20816
rect 2740 -21016 2774 -21000
rect 1653 -21062 1669 -21028
rect 2045 -21062 2061 -21028
rect 2289 -21062 2305 -21028
rect 2681 -21062 2697 -21028
rect -162 -21162 1472 -21100
rect 2878 -21162 2912 -21100
rect -162 -21196 -66 -21162
rect 1216 -21196 1534 -21162
rect 2816 -21196 2912 -21162
rect -162 -21258 1472 -21196
rect -128 -21296 1278 -21258
rect -128 -21330 69 -21296
rect 445 -21330 705 -21296
rect 1081 -21330 1278 -21296
rect -128 -21358 1278 -21330
rect -128 -22126 -24 -21358
rect 10 -22126 504 -21358
rect 538 -22126 612 -21358
rect 646 -22126 1140 -21358
rect 1174 -22126 1278 -21358
rect -128 -22154 1278 -22126
rect -128 -22188 69 -22154
rect 445 -22188 705 -22154
rect 1081 -22188 1278 -22154
rect -128 -22226 1278 -22188
rect 1312 -22226 1438 -21258
rect 2878 -21258 2912 -21196
rect 1653 -21330 1669 -21296
rect 2045 -21330 2061 -21296
rect 2289 -21330 2305 -21296
rect 2681 -21330 2697 -21296
rect 1576 -21358 1610 -21342
rect 1576 -22142 1610 -22126
rect 2104 -21358 2138 -21342
rect 2104 -22142 2138 -22126
rect 2212 -21358 2246 -21342
rect 2212 -22142 2246 -22126
rect 2740 -21358 2774 -21342
rect 2740 -22142 2774 -22126
rect 1653 -22188 1669 -22154
rect 2045 -22188 2061 -22154
rect 2289 -22188 2305 -22154
rect 2681 -22188 2697 -22154
rect -162 -22288 1472 -22226
rect 2878 -22288 2912 -22226
rect -162 -22322 -66 -22288
rect 1216 -22322 1534 -22288
rect 2816 -22300 2912 -22288
rect 3038 -20670 3134 -20636
rect 4416 -20670 4512 -20636
rect 3038 -20732 3072 -20670
rect 4478 -20732 4512 -20670
rect 3253 -20804 3269 -20770
rect 3645 -20804 3661 -20770
rect 3889 -20804 3905 -20770
rect 4281 -20804 4297 -20770
rect 3176 -20832 3210 -20816
rect 3176 -21016 3210 -21000
rect 3704 -20832 3738 -20816
rect 3704 -21016 3738 -21000
rect 3812 -20832 3846 -20816
rect 3812 -21016 3846 -21000
rect 4340 -20832 4374 -20816
rect 4340 -21016 4374 -21000
rect 3253 -21062 3269 -21028
rect 3645 -21062 3661 -21028
rect 3889 -21062 3905 -21028
rect 4281 -21062 4297 -21028
rect 3038 -21162 3072 -21100
rect 4478 -21162 4512 -21100
rect 3038 -21196 3134 -21162
rect 4416 -21196 4512 -21162
rect 3038 -21258 3072 -21196
rect 4478 -21258 4512 -21196
rect 3253 -21330 3269 -21296
rect 3645 -21330 3661 -21296
rect 3889 -21330 3905 -21296
rect 4281 -21330 4297 -21296
rect 3176 -21358 3210 -21342
rect 3176 -22142 3210 -22126
rect 3704 -21358 3738 -21342
rect 3704 -22142 3738 -22126
rect 3812 -21358 3846 -21342
rect 3812 -22142 3846 -22126
rect 4340 -21358 4374 -21342
rect 4340 -22142 4374 -22126
rect 3253 -22188 3269 -22154
rect 3645 -22188 3661 -22154
rect 3889 -22188 3905 -22154
rect 4281 -22188 4297 -22154
rect 3038 -22288 3072 -22226
rect 4478 -22280 4512 -22226
rect 4638 -20670 4734 -20636
rect 6016 -20670 6112 -20636
rect 4638 -20732 4672 -20670
rect 6078 -20732 6112 -20670
rect 4853 -20804 4869 -20770
rect 5245 -20804 5261 -20770
rect 5489 -20804 5505 -20770
rect 5881 -20804 5897 -20770
rect 4776 -20832 4810 -20816
rect 4776 -21016 4810 -21000
rect 5304 -20832 5338 -20816
rect 5304 -21016 5338 -21000
rect 5412 -20832 5446 -20816
rect 5412 -21016 5446 -21000
rect 5940 -20832 5974 -20816
rect 5940 -21016 5974 -21000
rect 4853 -21062 4869 -21028
rect 5245 -21062 5261 -21028
rect 5489 -21062 5505 -21028
rect 5881 -21062 5897 -21028
rect 4638 -21162 4672 -21100
rect 6078 -21162 6112 -21100
rect 4638 -21196 4734 -21162
rect 6016 -21196 6112 -21162
rect 4638 -21258 4672 -21196
rect 6078 -21258 6112 -21196
rect 4853 -21330 4869 -21296
rect 5245 -21330 5261 -21296
rect 5489 -21330 5505 -21296
rect 5881 -21330 5897 -21296
rect 4776 -21358 4810 -21342
rect 4776 -22142 4810 -22126
rect 5304 -21358 5338 -21342
rect 5304 -22142 5338 -22126
rect 5412 -21358 5446 -21342
rect 5412 -22142 5446 -22126
rect 5940 -21358 5974 -21342
rect 5940 -22142 5974 -22126
rect 4853 -22188 4869 -22154
rect 5245 -22188 5261 -22154
rect 5489 -22188 5505 -22154
rect 5881 -22188 5897 -22154
rect 4638 -22280 4672 -22226
rect 6078 -22280 6112 -22226
rect 6238 -20670 6334 -20636
rect 7616 -20670 7712 -20636
rect 6238 -20732 6272 -20670
rect 7678 -20732 7712 -20670
rect 6453 -20804 6469 -20770
rect 6845 -20804 6861 -20770
rect 7089 -20804 7105 -20770
rect 7481 -20804 7497 -20770
rect 6376 -20832 6410 -20816
rect 6376 -21016 6410 -21000
rect 6904 -20832 6938 -20816
rect 6904 -21016 6938 -21000
rect 7012 -20832 7046 -20816
rect 7012 -21016 7046 -21000
rect 7540 -20832 7574 -20816
rect 7540 -21016 7574 -21000
rect 6453 -21062 6469 -21028
rect 6845 -21062 6861 -21028
rect 7089 -21062 7105 -21028
rect 7481 -21062 7497 -21028
rect 6238 -21162 6272 -21100
rect 7678 -21162 7712 -21100
rect 6238 -21196 6334 -21162
rect 7616 -21196 7712 -21162
rect 6238 -21258 6272 -21196
rect 7678 -21258 7712 -21196
rect 6453 -21330 6469 -21296
rect 6845 -21330 6861 -21296
rect 7089 -21330 7105 -21296
rect 7481 -21330 7497 -21296
rect 6376 -21358 6410 -21342
rect 6376 -22142 6410 -22126
rect 6904 -21358 6938 -21342
rect 6904 -22142 6938 -22126
rect 7012 -21358 7046 -21342
rect 7012 -22142 7046 -22126
rect 7540 -21358 7574 -21342
rect 7540 -22142 7574 -22126
rect 6453 -22188 6469 -22154
rect 6845 -22188 6861 -22154
rect 7089 -22188 7105 -22154
rect 7481 -22188 7497 -22154
rect 6238 -22280 6272 -22226
rect 7678 -22280 7712 -22226
rect 7838 -20670 7934 -20636
rect 9216 -20670 9312 -20636
rect 7838 -20732 7872 -20670
rect 9278 -20732 9312 -20670
rect 8053 -20804 8069 -20770
rect 8445 -20804 8461 -20770
rect 8689 -20804 8705 -20770
rect 9081 -20804 9097 -20770
rect 7976 -20832 8010 -20816
rect 7976 -21016 8010 -21000
rect 8504 -20832 8538 -20816
rect 8504 -21016 8538 -21000
rect 8612 -20832 8646 -20816
rect 8612 -21016 8646 -21000
rect 9140 -20832 9174 -20816
rect 9140 -21016 9174 -21000
rect 8053 -21062 8069 -21028
rect 8445 -21062 8461 -21028
rect 8689 -21062 8705 -21028
rect 9081 -21062 9097 -21028
rect 7838 -21162 7872 -21100
rect 9278 -21162 9312 -21100
rect 7838 -21196 7934 -21162
rect 9216 -21196 9312 -21162
rect 7838 -21258 7872 -21196
rect 9278 -21258 9312 -21196
rect 8053 -21330 8069 -21296
rect 8445 -21330 8461 -21296
rect 8689 -21330 8705 -21296
rect 9081 -21330 9097 -21296
rect 7976 -21358 8010 -21342
rect 7976 -22142 8010 -22126
rect 8504 -21358 8538 -21342
rect 8504 -22142 8538 -22126
rect 8612 -21358 8646 -21342
rect 8612 -22142 8646 -22126
rect 9140 -21358 9174 -21342
rect 9140 -22142 9174 -22126
rect 8053 -22188 8069 -22154
rect 8445 -22188 8461 -22154
rect 8689 -22188 8705 -22154
rect 9081 -22188 9097 -22154
rect 7838 -22280 7872 -22226
rect 9278 -22280 9312 -22226
rect 9438 -20670 9534 -20636
rect 10816 -20670 10912 -20636
rect 9438 -20732 9472 -20670
rect 10878 -20732 10912 -20670
rect 9653 -20804 9669 -20770
rect 10045 -20804 10061 -20770
rect 10289 -20804 10305 -20770
rect 10681 -20804 10697 -20770
rect 9576 -20832 9610 -20816
rect 9576 -21016 9610 -21000
rect 10104 -20832 10138 -20816
rect 10104 -21016 10138 -21000
rect 10212 -20832 10246 -20816
rect 10212 -21016 10246 -21000
rect 10740 -20832 10774 -20816
rect 10740 -21016 10774 -21000
rect 9653 -21062 9669 -21028
rect 10045 -21062 10061 -21028
rect 10289 -21062 10305 -21028
rect 10681 -21062 10697 -21028
rect 9438 -21162 9472 -21100
rect 10878 -21162 10912 -21100
rect 9438 -21196 9534 -21162
rect 10816 -21196 10912 -21162
rect 9438 -21258 9472 -21196
rect 10878 -21258 10912 -21196
rect 9653 -21330 9669 -21296
rect 10045 -21330 10061 -21296
rect 10289 -21330 10305 -21296
rect 10681 -21330 10697 -21296
rect 9576 -21358 9610 -21342
rect 9576 -22142 9610 -22126
rect 10104 -21358 10138 -21342
rect 10104 -22142 10138 -22126
rect 10212 -21358 10246 -21342
rect 10212 -22142 10246 -22126
rect 10740 -21358 10774 -21342
rect 10740 -22142 10774 -22126
rect 9653 -22188 9669 -22154
rect 10045 -22188 10061 -22154
rect 10289 -22188 10305 -22154
rect 10681 -22188 10697 -22154
rect 9438 -22280 9472 -22226
rect 10878 -22280 10912 -22226
rect 11038 -20670 11134 -20636
rect 12416 -20670 12512 -20636
rect 11038 -20732 11072 -20670
rect 12478 -20732 12512 -20670
rect 11253 -20804 11269 -20770
rect 11645 -20804 11661 -20770
rect 11889 -20804 11905 -20770
rect 12281 -20804 12297 -20770
rect 11176 -20832 11210 -20816
rect 11176 -21016 11210 -21000
rect 11704 -20832 11738 -20816
rect 11704 -21016 11738 -21000
rect 11812 -20832 11846 -20816
rect 11812 -21016 11846 -21000
rect 12340 -20832 12374 -20816
rect 12340 -21016 12374 -21000
rect 11253 -21062 11269 -21028
rect 11645 -21062 11661 -21028
rect 11889 -21062 11905 -21028
rect 12281 -21062 12297 -21028
rect 11038 -21162 11072 -21100
rect 12478 -21162 12512 -21100
rect 11038 -21196 11134 -21162
rect 12416 -21196 12512 -21162
rect 11038 -21258 11072 -21196
rect 12478 -21258 12512 -21196
rect 11253 -21330 11269 -21296
rect 11645 -21330 11661 -21296
rect 11889 -21330 11905 -21296
rect 12281 -21330 12297 -21296
rect 11176 -21358 11210 -21342
rect 11176 -22142 11210 -22126
rect 11704 -21358 11738 -21342
rect 11704 -22142 11738 -22126
rect 11812 -21358 11846 -21342
rect 11812 -22142 11846 -22126
rect 12340 -21358 12374 -21342
rect 12340 -22142 12374 -22126
rect 11253 -22188 11269 -22154
rect 11645 -22188 11661 -22154
rect 11889 -22188 11905 -22154
rect 12281 -22188 12297 -22154
rect 11038 -22280 11072 -22226
rect 12478 -22280 12512 -22226
rect 12638 -20670 12734 -20636
rect 14016 -20670 14112 -20636
rect 12638 -20732 12672 -20670
rect 14078 -20732 14112 -20670
rect 12853 -20804 12869 -20770
rect 13245 -20804 13261 -20770
rect 13489 -20804 13505 -20770
rect 13881 -20804 13897 -20770
rect 12776 -20832 12810 -20816
rect 12776 -21016 12810 -21000
rect 13304 -20832 13338 -20816
rect 13304 -21016 13338 -21000
rect 13412 -20832 13446 -20816
rect 13412 -21016 13446 -21000
rect 13940 -20832 13974 -20816
rect 13940 -21016 13974 -21000
rect 12853 -21062 12869 -21028
rect 13245 -21062 13261 -21028
rect 13489 -21062 13505 -21028
rect 13881 -21062 13897 -21028
rect 12638 -21162 12672 -21100
rect 14078 -21162 14112 -21100
rect 12638 -21196 12734 -21162
rect 14016 -21196 14112 -21162
rect 12638 -21258 12672 -21196
rect 14078 -21258 14112 -21196
rect 12853 -21330 12869 -21296
rect 13245 -21330 13261 -21296
rect 13489 -21330 13505 -21296
rect 13881 -21330 13897 -21296
rect 12776 -21358 12810 -21342
rect 12776 -22142 12810 -22126
rect 13304 -21358 13338 -21342
rect 13304 -22142 13338 -22126
rect 13412 -21358 13446 -21342
rect 13412 -22142 13446 -22126
rect 13940 -21358 13974 -21342
rect 13940 -22142 13974 -22126
rect 12853 -22188 12869 -22154
rect 13245 -22188 13261 -22154
rect 13489 -22188 13505 -22154
rect 13881 -22188 13897 -22154
rect 12638 -22280 12672 -22226
rect 14078 -22280 14112 -22226
rect 14238 -20670 14334 -20636
rect 15616 -20670 15712 -20636
rect 14238 -20732 14272 -20670
rect 15678 -20732 15712 -20670
rect 14453 -20804 14469 -20770
rect 14845 -20804 14861 -20770
rect 15089 -20804 15105 -20770
rect 15481 -20804 15497 -20770
rect 14376 -20832 14410 -20816
rect 14376 -21016 14410 -21000
rect 14904 -20832 14938 -20816
rect 14904 -21016 14938 -21000
rect 15012 -20832 15046 -20816
rect 15012 -21016 15046 -21000
rect 15540 -20832 15574 -20816
rect 15540 -21016 15574 -21000
rect 14453 -21062 14469 -21028
rect 14845 -21062 14861 -21028
rect 15089 -21062 15105 -21028
rect 15481 -21062 15497 -21028
rect 14238 -21162 14272 -21100
rect 15678 -21162 15712 -21100
rect 14238 -21196 14334 -21162
rect 15616 -21196 15712 -21162
rect 14238 -21258 14272 -21196
rect 15678 -21258 15712 -21196
rect 14453 -21330 14469 -21296
rect 14845 -21330 14861 -21296
rect 15089 -21330 15105 -21296
rect 15481 -21330 15497 -21296
rect 14376 -21358 14410 -21342
rect 14376 -22142 14410 -22126
rect 14904 -21358 14938 -21342
rect 14904 -22142 14938 -22126
rect 15012 -21358 15046 -21342
rect 15012 -22142 15046 -22126
rect 15540 -21358 15574 -21342
rect 15540 -22142 15574 -22126
rect 14453 -22188 14469 -22154
rect 14845 -22188 14861 -22154
rect 15089 -22188 15105 -22154
rect 15481 -22188 15497 -22154
rect 14238 -22280 14272 -22226
rect 15678 -22280 15712 -22226
rect 15838 -20670 15934 -20636
rect 17216 -20670 17312 -20636
rect 15838 -20732 15872 -20670
rect 17278 -20732 17312 -20670
rect 16053 -20804 16069 -20770
rect 16445 -20804 16461 -20770
rect 16689 -20804 16705 -20770
rect 17081 -20804 17097 -20770
rect 15976 -20832 16010 -20816
rect 15976 -21016 16010 -21000
rect 16504 -20832 16538 -20816
rect 16504 -21016 16538 -21000
rect 16612 -20832 16646 -20816
rect 16612 -21016 16646 -21000
rect 17140 -20832 17174 -20816
rect 17140 -21016 17174 -21000
rect 16053 -21062 16069 -21028
rect 16445 -21062 16461 -21028
rect 16689 -21062 16705 -21028
rect 17081 -21062 17097 -21028
rect 15838 -21162 15872 -21100
rect 17278 -21162 17312 -21100
rect 15838 -21196 15934 -21162
rect 17216 -21196 17312 -21162
rect 15838 -21258 15872 -21196
rect 17278 -21258 17312 -21196
rect 16053 -21330 16069 -21296
rect 16445 -21330 16461 -21296
rect 16689 -21330 16705 -21296
rect 17081 -21330 17097 -21296
rect 15976 -21358 16010 -21342
rect 15976 -22142 16010 -22126
rect 16504 -21358 16538 -21342
rect 16504 -22142 16538 -22126
rect 16612 -21358 16646 -21342
rect 16612 -22142 16646 -22126
rect 17140 -21358 17174 -21342
rect 17140 -22142 17174 -22126
rect 16053 -22188 16069 -22154
rect 16445 -22188 16461 -22154
rect 16689 -22188 16705 -22154
rect 17081 -22188 17097 -22154
rect 15838 -22280 15872 -22226
rect 17278 -22280 17312 -22226
rect 17438 -20670 17534 -20636
rect 18816 -20670 18912 -20636
rect 17438 -20732 17472 -20670
rect 18878 -20732 18912 -20670
rect 17653 -20804 17669 -20770
rect 18045 -20804 18061 -20770
rect 18289 -20804 18305 -20770
rect 18681 -20804 18697 -20770
rect 17576 -20832 17610 -20816
rect 17576 -21016 17610 -21000
rect 18104 -20832 18138 -20816
rect 18104 -21016 18138 -21000
rect 18212 -20832 18246 -20816
rect 18212 -21016 18246 -21000
rect 18740 -20832 18774 -20816
rect 18740 -21016 18774 -21000
rect 17653 -21062 17669 -21028
rect 18045 -21062 18061 -21028
rect 18289 -21062 18305 -21028
rect 18681 -21062 18697 -21028
rect 17438 -21162 17472 -21100
rect 18878 -21162 18912 -21100
rect 17438 -21196 17534 -21162
rect 18816 -21196 18912 -21162
rect 17438 -21258 17472 -21196
rect 18878 -21258 18912 -21196
rect 17653 -21330 17669 -21296
rect 18045 -21330 18061 -21296
rect 18289 -21330 18305 -21296
rect 18681 -21330 18697 -21296
rect 17576 -21358 17610 -21342
rect 17576 -22142 17610 -22126
rect 18104 -21358 18138 -21342
rect 18104 -22142 18138 -22126
rect 18212 -21358 18246 -21342
rect 18212 -22142 18246 -22126
rect 18740 -21358 18774 -21342
rect 18740 -22142 18774 -22126
rect 17653 -22188 17669 -22154
rect 18045 -22188 18061 -22154
rect 18289 -22188 18305 -22154
rect 18681 -22188 18697 -22154
rect 17438 -22280 17472 -22226
rect 18878 -22280 18912 -22226
rect 19038 -20670 19134 -20636
rect 20416 -20670 20512 -20636
rect 19038 -20732 19072 -20670
rect 20478 -20732 20512 -20670
rect 19253 -20804 19269 -20770
rect 19645 -20804 19661 -20770
rect 19889 -20804 19905 -20770
rect 20281 -20804 20297 -20770
rect 19176 -20832 19210 -20816
rect 19176 -21016 19210 -21000
rect 19704 -20832 19738 -20816
rect 19704 -21016 19738 -21000
rect 19812 -20832 19846 -20816
rect 19812 -21016 19846 -21000
rect 20340 -20832 20374 -20816
rect 20340 -21016 20374 -21000
rect 19253 -21062 19269 -21028
rect 19645 -21062 19661 -21028
rect 19889 -21062 19905 -21028
rect 20281 -21062 20297 -21028
rect 19038 -21162 19072 -21100
rect 20478 -21162 20512 -21100
rect 19038 -21196 19134 -21162
rect 20416 -21196 20512 -21162
rect 19038 -21258 19072 -21196
rect 20478 -21258 20512 -21196
rect 19253 -21330 19269 -21296
rect 19645 -21330 19661 -21296
rect 19889 -21330 19905 -21296
rect 20281 -21330 20297 -21296
rect 19176 -21358 19210 -21342
rect 19176 -22142 19210 -22126
rect 19704 -21358 19738 -21342
rect 19704 -22142 19738 -22126
rect 19812 -21358 19846 -21342
rect 19812 -22142 19846 -22126
rect 20340 -21358 20374 -21342
rect 20340 -22142 20374 -22126
rect 19253 -22188 19269 -22154
rect 19645 -22188 19661 -22154
rect 19889 -22188 19905 -22154
rect 20281 -22188 20297 -22154
rect 19038 -22280 19072 -22226
rect 20478 -22280 20512 -22226
rect 20638 -20670 20734 -20636
rect 22016 -20670 22112 -20636
rect 20638 -20732 20672 -20670
rect 22078 -20732 22112 -20670
rect 20853 -20804 20869 -20770
rect 21245 -20804 21261 -20770
rect 21489 -20804 21505 -20770
rect 21881 -20804 21897 -20770
rect 20776 -20832 20810 -20816
rect 20776 -21016 20810 -21000
rect 21304 -20832 21338 -20816
rect 21304 -21016 21338 -21000
rect 21412 -20832 21446 -20816
rect 21412 -21016 21446 -21000
rect 21940 -20832 21974 -20816
rect 21940 -21016 21974 -21000
rect 20853 -21062 20869 -21028
rect 21245 -21062 21261 -21028
rect 21489 -21062 21505 -21028
rect 21881 -21062 21897 -21028
rect 20638 -21162 20672 -21100
rect 22078 -21162 22112 -21100
rect 20638 -21196 20734 -21162
rect 22016 -21196 22112 -21162
rect 20638 -21258 20672 -21196
rect 22078 -21258 22112 -21196
rect 20853 -21330 20869 -21296
rect 21245 -21330 21261 -21296
rect 21489 -21330 21505 -21296
rect 21881 -21330 21897 -21296
rect 20776 -21358 20810 -21342
rect 20776 -22142 20810 -22126
rect 21304 -21358 21338 -21342
rect 21304 -22142 21338 -22126
rect 21412 -21358 21446 -21342
rect 21412 -22142 21446 -22126
rect 21940 -21358 21974 -21342
rect 21940 -22142 21974 -22126
rect 20853 -22188 20869 -22154
rect 21245 -22188 21261 -22154
rect 21489 -22188 21505 -22154
rect 21881 -22188 21897 -22154
rect 20638 -22280 20672 -22226
rect 22078 -22280 22112 -22226
rect 3300 -22288 22112 -22280
rect 3038 -22300 3134 -22288
rect 2816 -22322 3134 -22300
rect 4416 -22322 4734 -22288
rect 6016 -22322 6334 -22288
rect 7616 -22322 7934 -22288
rect 9216 -22322 9534 -22288
rect 10816 -22322 11134 -22288
rect 12416 -22322 12734 -22288
rect 14016 -22322 14334 -22288
rect 15616 -22322 15934 -22288
rect 17216 -22322 17534 -22288
rect 18816 -22322 19134 -22288
rect 20416 -22322 20734 -22288
rect 22016 -22322 22112 -22288
rect 22238 -20670 22334 -20636
rect 23616 -20670 23712 -20636
rect 22238 -20732 22272 -20670
rect 23678 -20732 23712 -20670
rect 22453 -20804 22469 -20770
rect 22845 -20804 22861 -20770
rect 23089 -20804 23105 -20770
rect 23481 -20804 23497 -20770
rect 22376 -20832 22410 -20816
rect 22376 -21016 22410 -21000
rect 22904 -20832 22938 -20816
rect 22904 -21016 22938 -21000
rect 23012 -20832 23046 -20816
rect 23012 -21016 23046 -21000
rect 23540 -20832 23574 -20816
rect 23540 -21016 23574 -21000
rect 22453 -21062 22469 -21028
rect 22845 -21062 22861 -21028
rect 23089 -21062 23105 -21028
rect 23481 -21062 23497 -21028
rect 22238 -21162 22272 -21100
rect 23678 -21162 23712 -21100
rect 22238 -21196 22334 -21162
rect 23616 -21196 23712 -21162
rect 22238 -21258 22272 -21196
rect 23678 -21258 23712 -21196
rect 22453 -21330 22469 -21296
rect 22845 -21330 22861 -21296
rect 23089 -21330 23105 -21296
rect 23481 -21330 23497 -21296
rect 22376 -21358 22410 -21342
rect 22376 -22142 22410 -22126
rect 22904 -21358 22938 -21342
rect 22904 -22142 22938 -22126
rect 23012 -21358 23046 -21342
rect 23012 -22142 23046 -22126
rect 23540 -21358 23574 -21342
rect 23540 -22142 23574 -22126
rect 22453 -22188 22469 -22154
rect 22845 -22188 22861 -22154
rect 23089 -22188 23105 -22154
rect 23481 -22188 23497 -22154
rect 22238 -22288 22272 -22226
rect 23678 -22288 23712 -22226
rect 22238 -22322 22334 -22288
rect 23616 -22322 23712 -22288
rect 23838 -20670 23934 -20636
rect 25216 -20670 25312 -20636
rect 23838 -20732 23872 -20670
rect 25278 -20732 25312 -20670
rect 24053 -20804 24069 -20770
rect 24445 -20804 24461 -20770
rect 24689 -20804 24705 -20770
rect 25081 -20804 25097 -20770
rect 23976 -20832 24010 -20816
rect 23976 -21016 24010 -21000
rect 24504 -20832 24538 -20816
rect 24504 -21016 24538 -21000
rect 24612 -20832 24646 -20816
rect 24612 -21016 24646 -21000
rect 25140 -20832 25174 -20816
rect 25140 -21016 25174 -21000
rect 24053 -21062 24069 -21028
rect 24445 -21062 24461 -21028
rect 24689 -21062 24705 -21028
rect 25081 -21062 25097 -21028
rect 23838 -21162 23872 -21100
rect 25278 -21162 25312 -21100
rect 23838 -21196 23934 -21162
rect 25216 -21196 25312 -21162
rect 23838 -21258 23872 -21196
rect 25278 -21258 25312 -21196
rect 24053 -21330 24069 -21296
rect 24445 -21330 24461 -21296
rect 24689 -21330 24705 -21296
rect 25081 -21330 25097 -21296
rect 23976 -21358 24010 -21342
rect 23976 -22142 24010 -22126
rect 24504 -21358 24538 -21342
rect 24504 -22142 24538 -22126
rect 24612 -21358 24646 -21342
rect 24612 -22142 24646 -22126
rect 25140 -21358 25174 -21342
rect 25140 -22142 25174 -22126
rect 24053 -22188 24069 -22154
rect 24445 -22188 24461 -22154
rect 24689 -22188 24705 -22154
rect 25081 -22188 25097 -22154
rect 23838 -22288 23872 -22226
rect 25278 -22288 25312 -22226
rect 23838 -22322 23934 -22288
rect 25216 -22322 25312 -22288
rect 25438 -20670 25534 -20636
rect 26816 -20670 26912 -20636
rect 25438 -20732 25472 -20670
rect 26878 -20732 26912 -20670
rect 25653 -20804 25669 -20770
rect 26045 -20804 26061 -20770
rect 26289 -20804 26305 -20770
rect 26681 -20804 26697 -20770
rect 25576 -20832 25610 -20816
rect 25576 -21016 25610 -21000
rect 26104 -20832 26138 -20816
rect 26104 -21016 26138 -21000
rect 26212 -20832 26246 -20816
rect 26212 -21016 26246 -21000
rect 26740 -20832 26774 -20816
rect 26740 -21016 26774 -21000
rect 25653 -21062 25669 -21028
rect 26045 -21062 26061 -21028
rect 26289 -21062 26305 -21028
rect 26681 -21062 26697 -21028
rect 25438 -21162 25472 -21100
rect 26878 -21162 26912 -21100
rect 25438 -21196 25534 -21162
rect 26816 -21196 26912 -21162
rect 25438 -21258 25472 -21196
rect 26878 -21258 26912 -21196
rect 25653 -21330 25669 -21296
rect 26045 -21330 26061 -21296
rect 26289 -21330 26305 -21296
rect 26681 -21330 26697 -21296
rect 25576 -21358 25610 -21342
rect 25576 -22142 25610 -22126
rect 26104 -21358 26138 -21342
rect 26104 -22142 26138 -22126
rect 26212 -21358 26246 -21342
rect 26212 -22142 26246 -22126
rect 26740 -21358 26774 -21342
rect 26740 -22142 26774 -22126
rect 25653 -22188 25669 -22154
rect 26045 -22188 26061 -22154
rect 26289 -22188 26305 -22154
rect 26681 -22188 26697 -22154
rect 25438 -22288 25472 -22226
rect 26878 -22288 26912 -22226
rect 25438 -22322 25534 -22288
rect 26816 -22322 26912 -22288
rect 27038 -20670 27134 -20636
rect 28416 -20670 28512 -20636
rect 27038 -20732 27072 -20670
rect 28478 -20732 28512 -20670
rect 27253 -20804 27269 -20770
rect 27645 -20804 27661 -20770
rect 27889 -20804 27905 -20770
rect 28281 -20804 28297 -20770
rect 27176 -20832 27210 -20816
rect 27176 -21016 27210 -21000
rect 27704 -20832 27738 -20816
rect 27704 -21016 27738 -21000
rect 27812 -20832 27846 -20816
rect 27812 -21016 27846 -21000
rect 28340 -20832 28374 -20816
rect 28340 -21016 28374 -21000
rect 27253 -21062 27269 -21028
rect 27645 -21062 27661 -21028
rect 27889 -21062 27905 -21028
rect 28281 -21062 28297 -21028
rect 27038 -21162 27072 -21100
rect 28478 -21162 28512 -21100
rect 27038 -21196 27134 -21162
rect 28416 -21196 28512 -21162
rect 27038 -21258 27072 -21196
rect 28478 -21258 28512 -21196
rect 27253 -21330 27269 -21296
rect 27645 -21330 27661 -21296
rect 27889 -21330 27905 -21296
rect 28281 -21330 28297 -21296
rect 27176 -21358 27210 -21342
rect 27176 -22142 27210 -22126
rect 27704 -21358 27738 -21342
rect 27704 -22142 27738 -22126
rect 27812 -21358 27846 -21342
rect 27812 -22142 27846 -22126
rect 28340 -21358 28374 -21342
rect 28340 -22142 28374 -22126
rect 27253 -22188 27269 -22154
rect 27645 -22188 27661 -22154
rect 27889 -22188 27905 -22154
rect 28281 -22188 28297 -22154
rect 27038 -22288 27072 -22226
rect 28478 -22288 28512 -22226
rect 27038 -22322 27134 -22288
rect 28416 -22300 28512 -22288
rect 28638 -20670 28734 -20636
rect 30016 -20670 30112 -20636
rect 28638 -20732 28672 -20670
rect 30078 -20732 30112 -20670
rect 28853 -20804 28869 -20770
rect 29245 -20804 29261 -20770
rect 29489 -20804 29505 -20770
rect 29881 -20804 29897 -20770
rect 28776 -20832 28810 -20816
rect 28776 -21016 28810 -21000
rect 29304 -20832 29338 -20816
rect 29304 -21016 29338 -21000
rect 29412 -20832 29446 -20816
rect 29412 -21016 29446 -21000
rect 29940 -20832 29974 -20816
rect 29940 -21016 29974 -21000
rect 28853 -21062 28869 -21028
rect 29245 -21062 29261 -21028
rect 29489 -21062 29505 -21028
rect 29881 -21062 29897 -21028
rect 28638 -21162 28672 -21100
rect 30078 -21162 30112 -21100
rect 28638 -21196 28734 -21162
rect 30016 -21196 30112 -21162
rect 28638 -21258 28672 -21196
rect 30078 -21258 30112 -21196
rect 28853 -21330 28869 -21296
rect 29245 -21330 29261 -21296
rect 29489 -21330 29505 -21296
rect 29881 -21330 29897 -21296
rect 28776 -21358 28810 -21342
rect 28776 -22142 28810 -22126
rect 29304 -21358 29338 -21342
rect 29304 -22142 29338 -22126
rect 29412 -21358 29446 -21342
rect 29412 -22142 29446 -22126
rect 29940 -21358 29974 -21342
rect 29940 -22142 29974 -22126
rect 28853 -22188 28869 -22154
rect 29245 -22188 29261 -22154
rect 29489 -22188 29505 -22154
rect 29881 -22188 29897 -22154
rect 28638 -22288 28672 -22226
rect 30078 -22288 30112 -22226
rect 28638 -22300 28734 -22288
rect 28416 -22322 28734 -22300
rect 30016 -22322 30112 -22288
rect 30238 -20670 30334 -20636
rect 31616 -20670 31712 -20636
rect 30238 -20732 30272 -20670
rect 31678 -20732 31712 -20670
rect 30453 -20804 30469 -20770
rect 30845 -20804 30861 -20770
rect 31089 -20804 31105 -20770
rect 31481 -20804 31497 -20770
rect 30376 -20832 30410 -20816
rect 30376 -21016 30410 -21000
rect 30904 -20832 30938 -20816
rect 30904 -21016 30938 -21000
rect 31012 -20832 31046 -20816
rect 31012 -21016 31046 -21000
rect 31540 -20832 31574 -20816
rect 31540 -21016 31574 -21000
rect 30453 -21062 30469 -21028
rect 30845 -21062 30861 -21028
rect 31089 -21062 31105 -21028
rect 31481 -21062 31497 -21028
rect 30238 -21162 30272 -21100
rect 31678 -21162 31712 -21100
rect 30238 -21196 30334 -21162
rect 31616 -21196 31712 -21162
rect 30238 -21258 30272 -21196
rect 31678 -21258 31712 -21196
rect 30453 -21330 30469 -21296
rect 30845 -21330 30861 -21296
rect 31089 -21330 31105 -21296
rect 31481 -21330 31497 -21296
rect 30376 -21358 30410 -21342
rect 30376 -22142 30410 -22126
rect 30904 -21358 30938 -21342
rect 30904 -22142 30938 -22126
rect 31012 -21358 31046 -21342
rect 31012 -22142 31046 -22126
rect 31540 -21358 31574 -21342
rect 31540 -22142 31574 -22126
rect 30453 -22188 30469 -22154
rect 30845 -22188 30861 -22154
rect 31089 -22188 31105 -22154
rect 31481 -22188 31497 -22154
rect 30238 -22288 30272 -22226
rect 31678 -22288 31712 -22226
rect 30238 -22322 30334 -22288
rect 31616 -22322 31712 -22288
rect 31838 -20670 31934 -20636
rect 33216 -20670 33312 -20636
rect 31838 -20732 31872 -20670
rect 33278 -20732 33312 -20670
rect 32053 -20804 32069 -20770
rect 32445 -20804 32461 -20770
rect 32689 -20804 32705 -20770
rect 33081 -20804 33097 -20770
rect 31976 -20832 32010 -20816
rect 31976 -21016 32010 -21000
rect 32504 -20832 32538 -20816
rect 32504 -21016 32538 -21000
rect 32612 -20832 32646 -20816
rect 32612 -21016 32646 -21000
rect 33140 -20832 33174 -20816
rect 33140 -21016 33174 -21000
rect 32053 -21062 32069 -21028
rect 32445 -21062 32461 -21028
rect 32689 -21062 32705 -21028
rect 33081 -21062 33097 -21028
rect 31838 -21162 31872 -21100
rect 33278 -21162 33312 -21100
rect 31838 -21196 31934 -21162
rect 33216 -21196 33312 -21162
rect 31838 -21258 31872 -21196
rect 33278 -21258 33312 -21196
rect 32053 -21330 32069 -21296
rect 32445 -21330 32461 -21296
rect 32689 -21330 32705 -21296
rect 33081 -21330 33097 -21296
rect 31976 -21358 32010 -21342
rect 31976 -22142 32010 -22126
rect 32504 -21358 32538 -21342
rect 32504 -22142 32538 -22126
rect 32612 -21358 32646 -21342
rect 32612 -22142 32646 -22126
rect 33140 -21358 33174 -21342
rect 33140 -22142 33174 -22126
rect 32053 -22188 32069 -22154
rect 32445 -22188 32461 -22154
rect 32689 -22188 32705 -22154
rect 33081 -22188 33097 -22154
rect 31838 -22288 31872 -22226
rect 33278 -22288 33312 -22226
rect 31838 -22322 31934 -22288
rect 33216 -22300 33312 -22288
rect 33438 -20670 33534 -20636
rect 34816 -20670 34912 -20636
rect 33438 -20732 33472 -20670
rect 34878 -20732 34912 -20670
rect 33653 -20804 33669 -20770
rect 34045 -20804 34061 -20770
rect 34289 -20804 34305 -20770
rect 34681 -20804 34697 -20770
rect 33576 -20832 33610 -20816
rect 33576 -21016 33610 -21000
rect 34104 -20832 34138 -20816
rect 34104 -21016 34138 -21000
rect 34212 -20832 34246 -20816
rect 34212 -21016 34246 -21000
rect 34740 -20832 34774 -20816
rect 34740 -21016 34774 -21000
rect 33653 -21062 33669 -21028
rect 34045 -21062 34061 -21028
rect 34289 -21062 34305 -21028
rect 34681 -21062 34697 -21028
rect 33438 -21162 33472 -21100
rect 34878 -21162 34912 -21100
rect 33438 -21196 33534 -21162
rect 34816 -21196 34912 -21162
rect 33438 -21258 33472 -21196
rect 34878 -21258 34912 -21196
rect 33653 -21330 33669 -21296
rect 34045 -21330 34061 -21296
rect 34289 -21330 34305 -21296
rect 34681 -21330 34697 -21296
rect 33576 -21358 33610 -21342
rect 33576 -22142 33610 -22126
rect 34104 -21358 34138 -21342
rect 34104 -22142 34138 -22126
rect 34212 -21358 34246 -21342
rect 34212 -22142 34246 -22126
rect 34740 -21358 34774 -21342
rect 34740 -22142 34774 -22126
rect 33653 -22188 33669 -22154
rect 34045 -22188 34061 -22154
rect 34289 -22188 34305 -22154
rect 34681 -22188 34697 -22154
rect 33438 -22288 33472 -22226
rect 34878 -22288 34912 -22226
rect 33438 -22300 33534 -22288
rect 33216 -22322 33534 -22300
rect 34816 -22322 34912 -22288
rect 35038 -20670 35134 -20636
rect 36416 -20670 36734 -20636
rect 38016 -20670 38112 -20636
rect 35038 -20732 35072 -20670
rect 36478 -20732 38112 -20670
rect 35253 -20804 35269 -20770
rect 35645 -20804 35661 -20770
rect 35889 -20804 35905 -20770
rect 36281 -20804 36297 -20770
rect 35176 -20832 35210 -20816
rect 35176 -21016 35210 -21000
rect 35704 -20832 35738 -20816
rect 35704 -21016 35738 -21000
rect 35812 -20832 35846 -20816
rect 35812 -21016 35846 -21000
rect 36340 -20832 36374 -20816
rect 36340 -21016 36374 -21000
rect 35253 -21062 35269 -21028
rect 35645 -21062 35661 -21028
rect 35889 -21062 35905 -21028
rect 36281 -21062 36297 -21028
rect 35038 -21162 35072 -21100
rect 36512 -21100 36638 -20732
rect 36672 -20770 38078 -20732
rect 36672 -20804 36869 -20770
rect 37245 -20804 37505 -20770
rect 37881 -20804 38078 -20770
rect 36672 -20832 38078 -20804
rect 36672 -21000 36776 -20832
rect 36810 -21000 37304 -20832
rect 37338 -21000 37412 -20832
rect 37446 -21000 37940 -20832
rect 37974 -21000 38078 -20832
rect 36672 -21028 38078 -21000
rect 36672 -21062 36869 -21028
rect 37245 -21062 37505 -21028
rect 37881 -21062 38078 -21028
rect 36672 -21100 38078 -21062
rect 36478 -21162 38112 -21100
rect 35038 -21196 35134 -21162
rect 36416 -21196 36734 -21162
rect 38016 -21196 38112 -21162
rect 35038 -21258 35072 -21196
rect 36478 -21258 38112 -21196
rect 35253 -21330 35269 -21296
rect 35645 -21330 35661 -21296
rect 35889 -21330 35905 -21296
rect 36281 -21330 36297 -21296
rect 35176 -21358 35210 -21342
rect 35176 -22142 35210 -22126
rect 35704 -21358 35738 -21342
rect 35704 -22142 35738 -22126
rect 35812 -21358 35846 -21342
rect 35812 -22142 35846 -22126
rect 36340 -21358 36374 -21342
rect 36340 -22142 36374 -22126
rect 35253 -22188 35269 -22154
rect 35645 -22188 35661 -22154
rect 35889 -22188 35905 -22154
rect 36281 -22188 36297 -22154
rect 35038 -22288 35072 -22226
rect 36512 -22226 36638 -21258
rect 36672 -21296 38078 -21258
rect 36672 -21330 36869 -21296
rect 37245 -21330 37505 -21296
rect 37881 -21330 38078 -21296
rect 36672 -21358 38078 -21330
rect 36672 -22126 36776 -21358
rect 36810 -22126 37304 -21358
rect 37338 -22126 37412 -21358
rect 37446 -22126 37940 -21358
rect 37974 -22126 38078 -21358
rect 36672 -22154 38078 -22126
rect 36672 -22188 36869 -22154
rect 37245 -22188 37505 -22154
rect 37881 -22188 38078 -22154
rect 36672 -22226 38078 -22188
rect 36478 -22288 38112 -22226
rect 35038 -22322 35134 -22288
rect 36416 -22300 36734 -22288
rect 36416 -22322 36512 -22300
rect 36638 -22322 36734 -22300
rect 38016 -22322 38112 -22288
rect 60 -23920 22110 -22322
rect 28260 -22524 29140 -22322
rect 32240 -22404 34110 -22322
rect 32240 -22430 32594 -22404
rect 32330 -22438 32594 -22430
rect 33336 -22424 34110 -22404
rect 33336 -22438 33964 -22424
rect 32330 -22500 32532 -22438
rect 28218 -22558 28314 -22524
rect 29056 -22558 29152 -22524
rect 28218 -22620 28252 -22558
rect 29118 -22620 29152 -22558
rect 28352 -22684 28386 -22668
rect 28352 -23476 28386 -23460
rect 28510 -22684 28544 -22668
rect 28510 -23476 28544 -23460
rect 28668 -22684 28702 -22668
rect 28668 -23476 28702 -23460
rect 28826 -22684 28860 -22668
rect 28826 -23476 28860 -23460
rect 28984 -22684 29018 -22668
rect 28984 -23476 29018 -23460
rect 28398 -23553 28414 -23519
rect 28482 -23553 28498 -23519
rect 28556 -23553 28572 -23519
rect 28640 -23553 28656 -23519
rect 28714 -23553 28730 -23519
rect 28798 -23553 28814 -23519
rect 28872 -23553 28888 -23519
rect 28956 -23553 28972 -23519
rect 28218 -23658 28252 -23596
rect 32330 -23146 32498 -22500
rect 33398 -22458 33964 -22438
rect 34390 -22458 34486 -22424
rect 33398 -22500 33902 -22458
rect 32678 -22576 32694 -22542
rect 32762 -22576 32778 -22542
rect 32836 -22576 32852 -22542
rect 32920 -22576 32936 -22542
rect 32994 -22576 33010 -22542
rect 33078 -22576 33094 -22542
rect 33152 -22576 33168 -22542
rect 33236 -22576 33252 -22542
rect 32632 -22635 32666 -22619
rect 32632 -23027 32666 -23011
rect 32790 -22635 32824 -22619
rect 32790 -23027 32824 -23011
rect 32948 -22635 32982 -22619
rect 32948 -23027 32982 -23011
rect 33106 -22635 33140 -22619
rect 33106 -23027 33140 -23011
rect 33264 -22635 33298 -22619
rect 33264 -23027 33298 -23011
rect 32678 -23104 32694 -23070
rect 32762 -23104 32778 -23070
rect 32836 -23104 32852 -23070
rect 32920 -23104 32936 -23070
rect 32994 -23104 33010 -23070
rect 33078 -23104 33094 -23070
rect 33152 -23104 33168 -23070
rect 33236 -23104 33252 -23070
rect 32330 -23208 32532 -23146
rect 33432 -22520 33902 -22500
rect 33432 -23146 33868 -22520
rect 33398 -23166 33868 -23146
rect 34452 -22520 34486 -22458
rect 34048 -22596 34064 -22562
rect 34132 -22596 34148 -22562
rect 34206 -22596 34222 -22562
rect 34290 -22596 34306 -22562
rect 34002 -22655 34036 -22639
rect 34002 -23047 34036 -23031
rect 34160 -22655 34194 -22639
rect 34160 -23047 34194 -23031
rect 34318 -22655 34352 -22639
rect 34318 -23047 34352 -23031
rect 34048 -23124 34064 -23090
rect 34132 -23124 34148 -23090
rect 34206 -23124 34222 -23090
rect 34290 -23124 34306 -23090
rect 33398 -23208 33902 -23166
rect 32330 -23242 32594 -23208
rect 33336 -23228 33902 -23208
rect 34452 -23228 34486 -23166
rect 33336 -23242 33957 -23228
rect 32330 -23300 32520 -23242
rect 33410 -23262 33957 -23242
rect 34397 -23262 34486 -23228
rect 33410 -23330 33880 -23262
rect 29118 -23658 29152 -23596
rect 28218 -23692 28314 -23658
rect 29056 -23692 29152 -23658
rect 33036 -23580 33132 -23546
rect 34190 -23580 34286 -23546
rect 33036 -23642 33070 -23580
rect 60 -24172 22220 -23920
rect 48 -24206 144 -24172
rect 1990 -24206 2344 -24172
rect 4190 -24206 4544 -24172
rect 6390 -24206 6744 -24172
rect 8590 -24206 8944 -24172
rect 10790 -24206 11144 -24172
rect 12990 -24206 13344 -24172
rect 15190 -24206 15544 -24172
rect 17390 -24206 17744 -24172
rect 19590 -24206 19944 -24172
rect 21790 -24206 22220 -24172
rect 48 -24268 22220 -24206
rect 82 -24306 2052 -24268
rect 82 -24340 279 -24306
rect 1855 -24340 2052 -24306
rect 82 -24368 2052 -24340
rect 82 -24636 186 -24368
rect 220 -24636 1914 -24368
rect 1948 -24636 2052 -24368
rect 82 -24664 2052 -24636
rect 82 -24698 279 -24664
rect 1855 -24698 2052 -24664
rect 82 -24736 2052 -24698
rect 2086 -24736 2248 -24268
rect 2282 -24306 4252 -24268
rect 2282 -24340 2479 -24306
rect 4055 -24340 4252 -24306
rect 2282 -24368 4252 -24340
rect 2282 -24636 2386 -24368
rect 2420 -24636 4114 -24368
rect 4148 -24636 4252 -24368
rect 2282 -24664 4252 -24636
rect 2282 -24698 2479 -24664
rect 4055 -24698 4252 -24664
rect 2282 -24736 4252 -24698
rect 4286 -24736 4448 -24268
rect 4482 -24306 6452 -24268
rect 4482 -24340 4679 -24306
rect 6255 -24340 6452 -24306
rect 4482 -24368 6452 -24340
rect 4482 -24636 4586 -24368
rect 4620 -24636 6314 -24368
rect 6348 -24636 6452 -24368
rect 4482 -24664 6452 -24636
rect 4482 -24698 4679 -24664
rect 6255 -24698 6452 -24664
rect 4482 -24736 6452 -24698
rect 6486 -24736 6648 -24268
rect 6682 -24306 8652 -24268
rect 6682 -24340 6879 -24306
rect 8455 -24340 8652 -24306
rect 6682 -24368 8652 -24340
rect 6682 -24636 6786 -24368
rect 6820 -24636 8514 -24368
rect 8548 -24636 8652 -24368
rect 6682 -24664 8652 -24636
rect 6682 -24698 6879 -24664
rect 8455 -24698 8652 -24664
rect 6682 -24736 8652 -24698
rect 8686 -24736 8848 -24268
rect 8882 -24306 10852 -24268
rect 8882 -24340 9079 -24306
rect 10655 -24340 10852 -24306
rect 8882 -24368 10852 -24340
rect 8882 -24636 8986 -24368
rect 9020 -24636 10714 -24368
rect 10748 -24636 10852 -24368
rect 8882 -24664 10852 -24636
rect 8882 -24698 9079 -24664
rect 10655 -24698 10852 -24664
rect 8882 -24736 10852 -24698
rect 10886 -24736 11048 -24268
rect 11082 -24306 13052 -24268
rect 11082 -24340 11279 -24306
rect 12855 -24340 13052 -24306
rect 11082 -24368 13052 -24340
rect 11082 -24636 11186 -24368
rect 11220 -24636 12914 -24368
rect 12948 -24636 13052 -24368
rect 11082 -24664 13052 -24636
rect 11082 -24698 11279 -24664
rect 12855 -24698 13052 -24664
rect 11082 -24736 13052 -24698
rect 13086 -24736 13248 -24268
rect 13282 -24306 15252 -24268
rect 13282 -24340 13479 -24306
rect 15055 -24340 15252 -24306
rect 13282 -24368 15252 -24340
rect 13282 -24636 13386 -24368
rect 13420 -24636 15114 -24368
rect 15148 -24636 15252 -24368
rect 13282 -24664 15252 -24636
rect 13282 -24698 13479 -24664
rect 15055 -24698 15252 -24664
rect 13282 -24736 15252 -24698
rect 15286 -24736 15448 -24268
rect 15482 -24306 17452 -24268
rect 15482 -24340 15679 -24306
rect 17255 -24340 17452 -24306
rect 15482 -24368 17452 -24340
rect 15482 -24636 15586 -24368
rect 15620 -24636 17314 -24368
rect 17348 -24636 17452 -24368
rect 15482 -24664 17452 -24636
rect 15482 -24698 15679 -24664
rect 17255 -24698 17452 -24664
rect 15482 -24736 17452 -24698
rect 17486 -24736 17648 -24268
rect 17682 -24306 19652 -24268
rect 17682 -24340 17879 -24306
rect 19455 -24340 19652 -24306
rect 17682 -24368 19652 -24340
rect 17682 -24636 17786 -24368
rect 17820 -24636 19514 -24368
rect 19548 -24636 19652 -24368
rect 17682 -24664 19652 -24636
rect 17682 -24698 17879 -24664
rect 19455 -24698 19652 -24664
rect 17682 -24736 19652 -24698
rect 19686 -24736 19848 -24268
rect 19882 -24306 21852 -24268
rect 19882 -24340 20079 -24306
rect 21655 -24340 21852 -24306
rect 19882 -24368 21852 -24340
rect 19882 -24636 19986 -24368
rect 20020 -24636 21714 -24368
rect 21748 -24636 21852 -24368
rect 19882 -24664 21852 -24636
rect 19882 -24698 20079 -24664
rect 21655 -24698 21852 -24664
rect 19882 -24736 21852 -24698
rect 21886 -24500 22220 -24268
rect 34252 -23642 34286 -23580
rect 33216 -23718 33232 -23684
rect 33300 -23718 33316 -23684
rect 33374 -23718 33390 -23684
rect 33458 -23718 33474 -23684
rect 33532 -23718 33548 -23684
rect 33616 -23718 33632 -23684
rect 33690 -23718 33706 -23684
rect 33774 -23718 33790 -23684
rect 33848 -23718 33864 -23684
rect 33932 -23718 33948 -23684
rect 34006 -23718 34022 -23684
rect 34090 -23718 34106 -23684
rect 33170 -23777 33204 -23761
rect 33170 -24169 33204 -24153
rect 33328 -23777 33362 -23761
rect 33328 -24169 33362 -24153
rect 33486 -23777 33520 -23761
rect 33486 -24169 33520 -24153
rect 33644 -23777 33678 -23761
rect 33644 -24169 33678 -24153
rect 33802 -23777 33836 -23761
rect 33802 -24169 33836 -24153
rect 33960 -23777 33994 -23761
rect 33960 -24169 33994 -24153
rect 34118 -23777 34152 -23761
rect 34118 -24169 34152 -24153
rect 33216 -24246 33232 -24212
rect 33300 -24246 33316 -24212
rect 33374 -24246 33390 -24212
rect 33458 -24246 33474 -24212
rect 33532 -24246 33548 -24212
rect 33616 -24246 33632 -24212
rect 33690 -24246 33706 -24212
rect 33774 -24246 33790 -24212
rect 33848 -24246 33864 -24212
rect 33932 -24246 33948 -24212
rect 34006 -24246 34022 -24212
rect 34090 -24246 34106 -24212
rect 27580 -24320 29820 -24300
rect 21886 -24514 22900 -24500
rect 27020 -24514 27130 -24320
rect 21886 -24548 22292 -24514
rect 26968 -24548 27130 -24514
rect 21886 -24610 22900 -24548
rect 21886 -24736 22196 -24610
rect 48 -24798 22196 -24736
rect 48 -24832 144 -24798
rect 1990 -24820 2344 -24798
rect 1990 -24832 2086 -24820
rect 2248 -24832 2344 -24820
rect 4190 -24820 4544 -24798
rect 4190 -24832 4286 -24820
rect 4448 -24832 4544 -24820
rect 6390 -24820 6744 -24798
rect 6390 -24832 6486 -24820
rect 6648 -24832 6744 -24820
rect 8590 -24820 8944 -24798
rect 8590 -24832 8686 -24820
rect 8848 -24832 8944 -24820
rect 10790 -24820 11144 -24798
rect 10790 -24832 10886 -24820
rect 11048 -24832 11144 -24820
rect 12990 -24820 13344 -24798
rect 12990 -24832 13086 -24820
rect 13248 -24832 13344 -24820
rect 15190 -24820 15544 -24798
rect 15190 -24832 15286 -24820
rect 15448 -24832 15544 -24820
rect 17390 -24820 17744 -24798
rect 17390 -24832 17486 -24820
rect 17648 -24832 17744 -24820
rect 19590 -24820 19944 -24798
rect 19590 -24832 19686 -24820
rect 19848 -24832 19944 -24820
rect 21790 -24832 22196 -24798
rect 60 -24972 2060 -24832
rect 19860 -24972 22196 -24832
rect 22230 -24665 22900 -24610
rect 26360 -24665 26900 -24548
rect 27020 -24610 27130 -24548
rect 48 -25006 144 -24972
rect 1990 -25006 2086 -24972
rect 48 -25068 2086 -25006
rect 82 -25106 2052 -25068
rect 82 -25140 279 -25106
rect 1855 -25140 2052 -25106
rect 82 -25168 2052 -25140
rect 82 -25436 186 -25168
rect 220 -25436 1914 -25168
rect 1948 -25436 2052 -25168
rect 82 -25464 2052 -25436
rect 82 -25498 279 -25464
rect 1855 -25498 2052 -25464
rect 82 -25536 2052 -25498
rect 48 -25598 2086 -25536
rect 48 -25632 144 -25598
rect 1990 -25632 2086 -25598
rect 2248 -25006 2344 -24972
rect 4190 -25006 4286 -24972
rect 2248 -25068 2282 -25006
rect 4252 -25068 4286 -25006
rect 2463 -25140 2479 -25106
rect 4055 -25140 4071 -25106
rect 2386 -25168 2420 -25152
rect 2386 -25452 2420 -25436
rect 4114 -25168 4148 -25152
rect 4114 -25452 4148 -25436
rect 2463 -25498 2479 -25464
rect 4055 -25498 4071 -25464
rect 2248 -25598 2282 -25536
rect 4252 -25598 4286 -25536
rect 2248 -25632 2344 -25598
rect 4190 -25632 4286 -25598
rect 4448 -25006 4544 -24972
rect 6390 -25006 6486 -24972
rect 4448 -25068 4482 -25006
rect 6452 -25068 6486 -25006
rect 4663 -25140 4679 -25106
rect 6255 -25140 6271 -25106
rect 4586 -25168 4620 -25152
rect 4586 -25452 4620 -25436
rect 6314 -25168 6348 -25152
rect 6314 -25452 6348 -25436
rect 4663 -25498 4679 -25464
rect 6255 -25498 6271 -25464
rect 4448 -25598 4482 -25536
rect 6452 -25598 6486 -25536
rect 4448 -25632 4544 -25598
rect 6390 -25632 6486 -25598
rect 6648 -25006 6744 -24972
rect 8590 -25006 8686 -24972
rect 6648 -25068 6682 -25006
rect 8652 -25068 8686 -25006
rect 6863 -25140 6879 -25106
rect 8455 -25140 8471 -25106
rect 6786 -25168 6820 -25152
rect 6786 -25452 6820 -25436
rect 8514 -25168 8548 -25152
rect 8514 -25452 8548 -25436
rect 6863 -25498 6879 -25464
rect 8455 -25498 8471 -25464
rect 6648 -25598 6682 -25536
rect 8652 -25598 8686 -25536
rect 6648 -25632 6744 -25598
rect 8590 -25632 8686 -25598
rect 8848 -25006 8944 -24972
rect 10790 -25006 10886 -24972
rect 8848 -25068 8882 -25006
rect 10852 -25068 10886 -25006
rect 9063 -25140 9079 -25106
rect 10655 -25140 10671 -25106
rect 8986 -25168 9020 -25152
rect 8986 -25452 9020 -25436
rect 10714 -25168 10748 -25152
rect 10714 -25452 10748 -25436
rect 9063 -25498 9079 -25464
rect 10655 -25498 10671 -25464
rect 8848 -25598 8882 -25536
rect 10852 -25598 10886 -25536
rect 8848 -25632 8944 -25598
rect 10790 -25632 10886 -25598
rect 11048 -25006 11144 -24972
rect 12990 -25006 13086 -24972
rect 11048 -25068 11082 -25006
rect 13052 -25068 13086 -25006
rect 11263 -25140 11279 -25106
rect 12855 -25140 12871 -25106
rect 11186 -25168 11220 -25152
rect 11186 -25452 11220 -25436
rect 12914 -25168 12948 -25152
rect 12914 -25452 12948 -25436
rect 11263 -25498 11279 -25464
rect 12855 -25498 12871 -25464
rect 11048 -25598 11082 -25536
rect 13052 -25598 13086 -25536
rect 11048 -25632 11144 -25598
rect 12990 -25632 13086 -25598
rect 13248 -25006 13344 -24972
rect 15190 -25006 15286 -24972
rect 13248 -25068 13282 -25006
rect 15252 -25068 15286 -25006
rect 13463 -25140 13479 -25106
rect 15055 -25140 15071 -25106
rect 13386 -25168 13420 -25152
rect 13386 -25452 13420 -25436
rect 15114 -25168 15148 -25152
rect 15114 -25452 15148 -25436
rect 13463 -25498 13479 -25464
rect 15055 -25498 15071 -25464
rect 13248 -25598 13282 -25536
rect 15252 -25598 15286 -25536
rect 13248 -25632 13344 -25598
rect 15190 -25632 15286 -25598
rect 15448 -25006 15544 -24972
rect 17390 -25006 17486 -24972
rect 15448 -25068 15482 -25006
rect 17452 -25068 17486 -25006
rect 15663 -25140 15679 -25106
rect 17255 -25140 17271 -25106
rect 15586 -25168 15620 -25152
rect 15586 -25452 15620 -25436
rect 17314 -25168 17348 -25152
rect 17314 -25452 17348 -25436
rect 15663 -25498 15679 -25464
rect 17255 -25498 17271 -25464
rect 15448 -25598 15482 -25536
rect 17452 -25598 17486 -25536
rect 15448 -25632 15544 -25598
rect 17390 -25632 17486 -25598
rect 17648 -25006 17744 -24972
rect 19590 -25006 19686 -24972
rect 17648 -25068 17682 -25006
rect 19652 -25068 19686 -25006
rect 17863 -25140 17879 -25106
rect 19455 -25140 19471 -25106
rect 17786 -25168 17820 -25152
rect 17786 -25452 17820 -25436
rect 19514 -25168 19548 -25152
rect 19514 -25452 19548 -25436
rect 17863 -25498 17879 -25464
rect 19455 -25498 19471 -25464
rect 17648 -25598 17682 -25536
rect 19652 -25598 19686 -25536
rect 17648 -25632 17744 -25598
rect 19590 -25632 19686 -25598
rect 19848 -25006 19944 -24972
rect 21790 -25006 22196 -24972
rect 19848 -25068 22196 -25006
rect 19882 -25106 21852 -25068
rect 19882 -25140 20079 -25106
rect 21655 -25140 21852 -25106
rect 19882 -25168 21852 -25140
rect 19882 -25436 19986 -25168
rect 20020 -25436 21714 -25168
rect 21748 -25436 21852 -25168
rect 19882 -25464 21852 -25436
rect 19882 -25498 20079 -25464
rect 21655 -25498 21852 -25464
rect 19882 -25536 21852 -25498
rect 21886 -25536 22196 -25068
rect 19848 -25598 22196 -25536
rect 19848 -25632 19944 -25598
rect 21790 -25632 22196 -25598
rect 60 -25772 2060 -25632
rect 19860 -25772 22196 -25632
rect 48 -25806 144 -25772
rect 1990 -25806 2086 -25772
rect 48 -25868 2086 -25806
rect 82 -25906 2052 -25868
rect 82 -25940 279 -25906
rect 1855 -25940 2052 -25906
rect 82 -25968 2052 -25940
rect 82 -26236 186 -25968
rect 220 -26236 1914 -25968
rect 1948 -26236 2052 -25968
rect 82 -26264 2052 -26236
rect 82 -26298 279 -26264
rect 1855 -26298 2052 -26264
rect 82 -26336 2052 -26298
rect 48 -26398 2086 -26336
rect 48 -26432 144 -26398
rect 1990 -26432 2086 -26398
rect 2248 -25806 2344 -25772
rect 4190 -25806 4286 -25772
rect 2248 -25868 2282 -25806
rect 4252 -25868 4286 -25806
rect 2463 -25940 2479 -25906
rect 4055 -25940 4071 -25906
rect 2386 -25968 2420 -25952
rect 2386 -26252 2420 -26236
rect 4114 -25968 4148 -25952
rect 4114 -26252 4148 -26236
rect 2463 -26298 2479 -26264
rect 4055 -26298 4071 -26264
rect 2248 -26398 2282 -26336
rect 4252 -26398 4286 -26336
rect 2248 -26432 2344 -26398
rect 4190 -26432 4286 -26398
rect 4448 -25806 4544 -25772
rect 6390 -25806 6486 -25772
rect 4448 -25868 4482 -25806
rect 6452 -25868 6486 -25806
rect 4663 -25940 4679 -25906
rect 6255 -25940 6271 -25906
rect 4586 -25968 4620 -25952
rect 4586 -26252 4620 -26236
rect 6314 -25968 6348 -25952
rect 6314 -26252 6348 -26236
rect 4663 -26298 4679 -26264
rect 6255 -26298 6271 -26264
rect 4448 -26398 4482 -26336
rect 6452 -26398 6486 -26336
rect 4448 -26432 4544 -26398
rect 6390 -26432 6486 -26398
rect 6648 -25806 6744 -25772
rect 8590 -25806 8686 -25772
rect 6648 -25868 6682 -25806
rect 8652 -25868 8686 -25806
rect 6863 -25940 6879 -25906
rect 8455 -25940 8471 -25906
rect 6786 -25968 6820 -25952
rect 6786 -26252 6820 -26236
rect 8514 -25968 8548 -25952
rect 8514 -26252 8548 -26236
rect 6863 -26298 6879 -26264
rect 8455 -26298 8471 -26264
rect 6648 -26398 6682 -26336
rect 8652 -26398 8686 -26336
rect 6648 -26432 6744 -26398
rect 8590 -26432 8686 -26398
rect 8848 -25806 8944 -25772
rect 10790 -25806 10886 -25772
rect 8848 -25868 8882 -25806
rect 10852 -25868 10886 -25806
rect 9063 -25940 9079 -25906
rect 10655 -25940 10671 -25906
rect 8986 -25968 9020 -25952
rect 8986 -26252 9020 -26236
rect 10714 -25968 10748 -25952
rect 10714 -26252 10748 -26236
rect 9063 -26298 9079 -26264
rect 10655 -26298 10671 -26264
rect 8848 -26398 8882 -26336
rect 10852 -26398 10886 -26336
rect 8848 -26432 8944 -26398
rect 10790 -26432 10886 -26398
rect 11048 -25806 11144 -25772
rect 12990 -25806 13086 -25772
rect 11048 -25868 11082 -25806
rect 13052 -25868 13086 -25806
rect 11263 -25940 11279 -25906
rect 12855 -25940 12871 -25906
rect 11186 -25968 11220 -25952
rect 11186 -26252 11220 -26236
rect 12914 -25968 12948 -25952
rect 12914 -26252 12948 -26236
rect 11263 -26298 11279 -26264
rect 12855 -26298 12871 -26264
rect 11048 -26398 11082 -26336
rect 13052 -26398 13086 -26336
rect 11048 -26432 11144 -26398
rect 12990 -26432 13086 -26398
rect 13248 -25806 13344 -25772
rect 15190 -25806 15286 -25772
rect 13248 -25868 13282 -25806
rect 15252 -25868 15286 -25806
rect 13463 -25940 13479 -25906
rect 15055 -25940 15071 -25906
rect 13386 -25968 13420 -25952
rect 13386 -26252 13420 -26236
rect 15114 -25968 15148 -25952
rect 15114 -26252 15148 -26236
rect 13463 -26298 13479 -26264
rect 15055 -26298 15071 -26264
rect 13248 -26398 13282 -26336
rect 15252 -26398 15286 -26336
rect 13248 -26432 13344 -26398
rect 15190 -26432 15286 -26398
rect 15448 -25806 15544 -25772
rect 17390 -25806 17486 -25772
rect 15448 -25868 15482 -25806
rect 17452 -25868 17486 -25806
rect 15663 -25940 15679 -25906
rect 17255 -25940 17271 -25906
rect 15586 -25968 15620 -25952
rect 15586 -26252 15620 -26236
rect 17314 -25968 17348 -25952
rect 17314 -26252 17348 -26236
rect 15663 -26298 15679 -26264
rect 17255 -26298 17271 -26264
rect 15448 -26398 15482 -26336
rect 17452 -26398 17486 -26336
rect 15448 -26432 15544 -26398
rect 17390 -26432 17486 -26398
rect 17648 -25806 17744 -25772
rect 19590 -25806 19686 -25772
rect 17648 -25868 17682 -25806
rect 19652 -25868 19686 -25806
rect 17863 -25940 17879 -25906
rect 19455 -25940 19471 -25906
rect 17786 -25968 17820 -25952
rect 17786 -26252 17820 -26236
rect 19514 -25968 19548 -25952
rect 19514 -26252 19548 -26236
rect 17863 -26298 17879 -26264
rect 19455 -26298 19471 -26264
rect 17648 -26398 17682 -26336
rect 19652 -26398 19686 -26336
rect 17648 -26432 17744 -26398
rect 19590 -26432 19686 -26398
rect 19848 -25806 19944 -25772
rect 21790 -25806 22196 -25772
rect 19848 -25868 22196 -25806
rect 19882 -25906 21852 -25868
rect 19882 -25940 20079 -25906
rect 21655 -25940 21852 -25906
rect 19882 -25968 21852 -25940
rect 19882 -26236 19986 -25968
rect 20020 -26236 21714 -25968
rect 21748 -26236 21852 -25968
rect 19882 -26264 21852 -26236
rect 19882 -26298 20079 -26264
rect 21655 -26298 21852 -26264
rect 19882 -26336 21852 -26298
rect 21886 -26336 22196 -25868
rect 19848 -26398 22196 -26336
rect 19848 -26432 19944 -26398
rect 21790 -26432 22196 -26398
rect 60 -26572 2060 -26432
rect 19860 -26572 22196 -26432
rect 48 -26606 144 -26572
rect 1990 -26606 2086 -26572
rect 48 -26668 2086 -26606
rect 82 -26706 2052 -26668
rect 82 -26740 279 -26706
rect 1855 -26740 2052 -26706
rect 82 -26768 2052 -26740
rect 82 -27036 186 -26768
rect 220 -27036 1914 -26768
rect 1948 -27036 2052 -26768
rect 82 -27064 2052 -27036
rect 82 -27098 279 -27064
rect 1855 -27098 2052 -27064
rect 82 -27136 2052 -27098
rect 48 -27198 2086 -27136
rect 48 -27232 144 -27198
rect 1990 -27232 2086 -27198
rect 2248 -26606 2344 -26572
rect 4190 -26606 4286 -26572
rect 2248 -26668 2282 -26606
rect 4252 -26668 4286 -26606
rect 2463 -26740 2479 -26706
rect 4055 -26740 4071 -26706
rect 2386 -26768 2420 -26752
rect 2386 -27052 2420 -27036
rect 4114 -26768 4148 -26752
rect 4114 -27052 4148 -27036
rect 2463 -27098 2479 -27064
rect 4055 -27098 4071 -27064
rect 2248 -27198 2282 -27136
rect 4252 -27198 4286 -27136
rect 2248 -27232 2344 -27198
rect 4190 -27232 4286 -27198
rect 4448 -26606 4544 -26572
rect 6390 -26606 6486 -26572
rect 4448 -26668 4482 -26606
rect 6452 -26668 6486 -26606
rect 4663 -26740 4679 -26706
rect 6255 -26740 6271 -26706
rect 4586 -26768 4620 -26752
rect 4586 -27052 4620 -27036
rect 6314 -26768 6348 -26752
rect 6314 -27052 6348 -27036
rect 4663 -27098 4679 -27064
rect 6255 -27098 6271 -27064
rect 4448 -27198 4482 -27136
rect 6452 -27198 6486 -27136
rect 4448 -27232 4544 -27198
rect 6390 -27232 6486 -27198
rect 6648 -26606 6744 -26572
rect 8590 -26606 8686 -26572
rect 6648 -26668 6682 -26606
rect 8652 -26668 8686 -26606
rect 6863 -26740 6879 -26706
rect 8455 -26740 8471 -26706
rect 6786 -26768 6820 -26752
rect 6786 -27052 6820 -27036
rect 8514 -26768 8548 -26752
rect 8514 -27052 8548 -27036
rect 6863 -27098 6879 -27064
rect 8455 -27098 8471 -27064
rect 6648 -27198 6682 -27136
rect 8652 -27198 8686 -27136
rect 6648 -27232 6744 -27198
rect 8590 -27232 8686 -27198
rect 8848 -26606 8944 -26572
rect 10790 -26606 10886 -26572
rect 8848 -26668 8882 -26606
rect 10852 -26668 10886 -26606
rect 9063 -26740 9079 -26706
rect 10655 -26740 10671 -26706
rect 8986 -26768 9020 -26752
rect 8986 -27052 9020 -27036
rect 10714 -26768 10748 -26752
rect 10714 -27052 10748 -27036
rect 9063 -27098 9079 -27064
rect 10655 -27098 10671 -27064
rect 8848 -27198 8882 -27136
rect 10852 -27198 10886 -27136
rect 8848 -27232 8944 -27198
rect 10790 -27232 10886 -27198
rect 11048 -26606 11144 -26572
rect 12990 -26606 13086 -26572
rect 11048 -26668 11082 -26606
rect 13052 -26668 13086 -26606
rect 11263 -26740 11279 -26706
rect 12855 -26740 12871 -26706
rect 11186 -26768 11220 -26752
rect 11186 -27052 11220 -27036
rect 12914 -26768 12948 -26752
rect 12914 -27052 12948 -27036
rect 11263 -27098 11279 -27064
rect 12855 -27098 12871 -27064
rect 11048 -27198 11082 -27136
rect 13052 -27198 13086 -27136
rect 11048 -27232 11144 -27198
rect 12990 -27232 13086 -27198
rect 13248 -26606 13344 -26572
rect 15190 -26606 15286 -26572
rect 13248 -26668 13282 -26606
rect 15252 -26668 15286 -26606
rect 13463 -26740 13479 -26706
rect 15055 -26740 15071 -26706
rect 13386 -26768 13420 -26752
rect 13386 -27052 13420 -27036
rect 15114 -26768 15148 -26752
rect 15114 -27052 15148 -27036
rect 13463 -27098 13479 -27064
rect 15055 -27098 15071 -27064
rect 13248 -27198 13282 -27136
rect 15252 -27198 15286 -27136
rect 13248 -27232 13344 -27198
rect 15190 -27232 15286 -27198
rect 15448 -26606 15544 -26572
rect 17390 -26606 17486 -26572
rect 15448 -26668 15482 -26606
rect 17452 -26668 17486 -26606
rect 15663 -26740 15679 -26706
rect 17255 -26740 17271 -26706
rect 15586 -26768 15620 -26752
rect 15586 -27052 15620 -27036
rect 17314 -26768 17348 -26752
rect 17314 -27052 17348 -27036
rect 15663 -27098 15679 -27064
rect 17255 -27098 17271 -27064
rect 15448 -27198 15482 -27136
rect 17452 -27198 17486 -27136
rect 15448 -27232 15544 -27198
rect 17390 -27232 17486 -27198
rect 17648 -26606 17744 -26572
rect 19590 -26606 19686 -26572
rect 17648 -26668 17682 -26606
rect 19652 -26668 19686 -26606
rect 17863 -26740 17879 -26706
rect 19455 -26740 19471 -26706
rect 17786 -26768 17820 -26752
rect 17786 -27052 17820 -27036
rect 19514 -26768 19548 -26752
rect 19514 -27052 19548 -27036
rect 17863 -27098 17879 -27064
rect 19455 -27098 19471 -27064
rect 17648 -27198 17682 -27136
rect 19652 -27198 19686 -27136
rect 17648 -27232 17744 -27198
rect 19590 -27232 19686 -27198
rect 19848 -26606 19944 -26572
rect 21790 -26606 22196 -26572
rect 19848 -26668 22196 -26606
rect 19882 -26706 21852 -26668
rect 19882 -26740 20079 -26706
rect 21655 -26740 21852 -26706
rect 19882 -26768 21852 -26740
rect 19882 -27036 19986 -26768
rect 20020 -27036 21714 -26768
rect 21748 -27036 21852 -26768
rect 19882 -27064 21852 -27036
rect 19882 -27098 20079 -27064
rect 21655 -27098 21852 -27064
rect 19882 -27136 21852 -27098
rect 21886 -27136 22196 -26668
rect 19848 -27198 22196 -27136
rect 19848 -27232 19944 -27198
rect 21790 -27232 22196 -27198
rect 60 -27372 2060 -27232
rect 19860 -27372 22196 -27232
rect 48 -27406 144 -27372
rect 1990 -27406 2086 -27372
rect 48 -27468 2086 -27406
rect 82 -27506 2052 -27468
rect 82 -27540 279 -27506
rect 1855 -27540 2052 -27506
rect 82 -27568 2052 -27540
rect 82 -27836 186 -27568
rect 220 -27836 1914 -27568
rect 1948 -27836 2052 -27568
rect 82 -27864 2052 -27836
rect 82 -27898 279 -27864
rect 1855 -27898 2052 -27864
rect 82 -27936 2052 -27898
rect 48 -27998 2086 -27936
rect 48 -28032 144 -27998
rect 1990 -28032 2086 -27998
rect 2248 -27406 2344 -27372
rect 4190 -27406 4286 -27372
rect 2248 -27468 2282 -27406
rect 4252 -27468 4286 -27406
rect 2463 -27540 2479 -27506
rect 4055 -27540 4071 -27506
rect 2386 -27568 2420 -27552
rect 2386 -27852 2420 -27836
rect 4114 -27568 4148 -27552
rect 4114 -27852 4148 -27836
rect 2463 -27898 2479 -27864
rect 4055 -27898 4071 -27864
rect 2248 -27998 2282 -27936
rect 4252 -27998 4286 -27936
rect 2248 -28032 2344 -27998
rect 4190 -28032 4286 -27998
rect 4448 -27406 4544 -27372
rect 6390 -27406 6486 -27372
rect 4448 -27468 4482 -27406
rect 6452 -27468 6486 -27406
rect 4663 -27540 4679 -27506
rect 6255 -27540 6271 -27506
rect 4586 -27568 4620 -27552
rect 4586 -27852 4620 -27836
rect 6314 -27568 6348 -27552
rect 6314 -27852 6348 -27836
rect 4663 -27898 4679 -27864
rect 6255 -27898 6271 -27864
rect 4448 -27998 4482 -27936
rect 6452 -27998 6486 -27936
rect 4448 -28032 4544 -27998
rect 6390 -28032 6486 -27998
rect 6648 -27406 6744 -27372
rect 8590 -27406 8686 -27372
rect 6648 -27468 6682 -27406
rect 8652 -27468 8686 -27406
rect 6863 -27540 6879 -27506
rect 8455 -27540 8471 -27506
rect 6786 -27568 6820 -27552
rect 6786 -27852 6820 -27836
rect 8514 -27568 8548 -27552
rect 8514 -27852 8548 -27836
rect 6863 -27898 6879 -27864
rect 8455 -27898 8471 -27864
rect 6648 -27998 6682 -27936
rect 8652 -27998 8686 -27936
rect 6648 -28032 6744 -27998
rect 8590 -28032 8686 -27998
rect 8848 -27406 8944 -27372
rect 10790 -27406 10886 -27372
rect 8848 -27468 8882 -27406
rect 10852 -27468 10886 -27406
rect 9063 -27540 9079 -27506
rect 10655 -27540 10671 -27506
rect 8986 -27568 9020 -27552
rect 8986 -27852 9020 -27836
rect 10714 -27568 10748 -27552
rect 10714 -27852 10748 -27836
rect 9063 -27898 9079 -27864
rect 10655 -27898 10671 -27864
rect 8848 -27998 8882 -27936
rect 10852 -27998 10886 -27936
rect 8848 -28032 8944 -27998
rect 10790 -28032 10886 -27998
rect 11048 -27406 11144 -27372
rect 12990 -27406 13086 -27372
rect 11048 -27468 11082 -27406
rect 13052 -27468 13086 -27406
rect 11263 -27540 11279 -27506
rect 12855 -27540 12871 -27506
rect 11186 -27568 11220 -27552
rect 11186 -27852 11220 -27836
rect 12914 -27568 12948 -27552
rect 12914 -27852 12948 -27836
rect 11263 -27898 11279 -27864
rect 12855 -27898 12871 -27864
rect 11048 -27998 11082 -27936
rect 13052 -27998 13086 -27936
rect 11048 -28032 11144 -27998
rect 12990 -28032 13086 -27998
rect 13248 -27406 13344 -27372
rect 15190 -27406 15286 -27372
rect 13248 -27468 13282 -27406
rect 15252 -27468 15286 -27406
rect 13463 -27540 13479 -27506
rect 15055 -27540 15071 -27506
rect 13386 -27568 13420 -27552
rect 13386 -27852 13420 -27836
rect 15114 -27568 15148 -27552
rect 15114 -27852 15148 -27836
rect 13463 -27898 13479 -27864
rect 15055 -27898 15071 -27864
rect 13248 -27998 13282 -27936
rect 15252 -27998 15286 -27936
rect 13248 -28032 13344 -27998
rect 15190 -28032 15286 -27998
rect 15448 -27406 15544 -27372
rect 17390 -27406 17486 -27372
rect 15448 -27468 15482 -27406
rect 17452 -27468 17486 -27406
rect 15663 -27540 15679 -27506
rect 17255 -27540 17271 -27506
rect 15586 -27568 15620 -27552
rect 15586 -27852 15620 -27836
rect 17314 -27568 17348 -27552
rect 17314 -27852 17348 -27836
rect 15663 -27898 15679 -27864
rect 17255 -27898 17271 -27864
rect 15448 -27998 15482 -27936
rect 17452 -27998 17486 -27936
rect 15448 -28032 15544 -27998
rect 17390 -28032 17486 -27998
rect 17648 -27406 17744 -27372
rect 19590 -27406 19686 -27372
rect 17648 -27468 17682 -27406
rect 19652 -27468 19686 -27406
rect 17863 -27540 17879 -27506
rect 19455 -27540 19471 -27506
rect 17786 -27568 17820 -27552
rect 17786 -27852 17820 -27836
rect 19514 -27568 19548 -27552
rect 19514 -27852 19548 -27836
rect 17863 -27898 17879 -27864
rect 19455 -27898 19471 -27864
rect 17648 -27998 17682 -27936
rect 19652 -27998 19686 -27936
rect 17648 -28032 17744 -27998
rect 19590 -28032 19686 -27998
rect 19848 -27406 19944 -27372
rect 21790 -27406 22196 -27372
rect 19848 -27468 22196 -27406
rect 19882 -27506 21852 -27468
rect 19882 -27540 20079 -27506
rect 21655 -27540 21852 -27506
rect 19882 -27568 21852 -27540
rect 19882 -27836 19986 -27568
rect 20020 -27836 21714 -27568
rect 21748 -27836 21852 -27568
rect 19882 -27864 21852 -27836
rect 19882 -27898 20079 -27864
rect 21655 -27898 21852 -27864
rect 19882 -27936 21852 -27898
rect 21886 -27936 22196 -27468
rect 19848 -27998 22196 -27936
rect 19848 -28032 19944 -27998
rect 21790 -28032 22196 -27998
rect 60 -28172 2060 -28032
rect 19860 -28172 22196 -28032
rect 48 -28206 144 -28172
rect 1990 -28206 2086 -28172
rect 48 -28268 2086 -28206
rect 82 -28306 2052 -28268
rect 82 -28340 279 -28306
rect 1855 -28340 2052 -28306
rect 82 -28368 2052 -28340
rect 82 -28636 186 -28368
rect 220 -28636 1914 -28368
rect 1948 -28636 2052 -28368
rect 82 -28664 2052 -28636
rect 82 -28698 279 -28664
rect 1855 -28698 2052 -28664
rect 82 -28736 2052 -28698
rect 48 -28798 2086 -28736
rect 48 -28832 144 -28798
rect 1990 -28832 2086 -28798
rect 2248 -28206 2344 -28172
rect 4190 -28206 4286 -28172
rect 2248 -28268 2282 -28206
rect 4252 -28268 4286 -28206
rect 2463 -28340 2479 -28306
rect 4055 -28340 4071 -28306
rect 2386 -28368 2420 -28352
rect 2386 -28652 2420 -28636
rect 4114 -28368 4148 -28352
rect 4114 -28652 4148 -28636
rect 2463 -28698 2479 -28664
rect 4055 -28698 4071 -28664
rect 2248 -28798 2282 -28736
rect 4252 -28798 4286 -28736
rect 2248 -28832 2344 -28798
rect 4190 -28832 4286 -28798
rect 4448 -28206 4544 -28172
rect 6390 -28206 6486 -28172
rect 4448 -28268 4482 -28206
rect 6452 -28268 6486 -28206
rect 4663 -28340 4679 -28306
rect 6255 -28340 6271 -28306
rect 4586 -28368 4620 -28352
rect 4586 -28652 4620 -28636
rect 6314 -28368 6348 -28352
rect 6314 -28652 6348 -28636
rect 4663 -28698 4679 -28664
rect 6255 -28698 6271 -28664
rect 4448 -28798 4482 -28736
rect 6452 -28798 6486 -28736
rect 4448 -28832 4544 -28798
rect 6390 -28832 6486 -28798
rect 6648 -28206 6744 -28172
rect 8590 -28206 8686 -28172
rect 6648 -28268 6682 -28206
rect 8652 -28268 8686 -28206
rect 6863 -28340 6879 -28306
rect 8455 -28340 8471 -28306
rect 6786 -28368 6820 -28352
rect 6786 -28652 6820 -28636
rect 8514 -28368 8548 -28352
rect 8514 -28652 8548 -28636
rect 6863 -28698 6879 -28664
rect 8455 -28698 8471 -28664
rect 6648 -28798 6682 -28736
rect 8652 -28798 8686 -28736
rect 6648 -28832 6744 -28798
rect 8590 -28832 8686 -28798
rect 8848 -28206 8944 -28172
rect 10790 -28206 10886 -28172
rect 8848 -28268 8882 -28206
rect 10852 -28268 10886 -28206
rect 9063 -28340 9079 -28306
rect 10655 -28340 10671 -28306
rect 8986 -28368 9020 -28352
rect 8986 -28652 9020 -28636
rect 10714 -28368 10748 -28352
rect 10714 -28652 10748 -28636
rect 9063 -28698 9079 -28664
rect 10655 -28698 10671 -28664
rect 8848 -28798 8882 -28736
rect 10852 -28798 10886 -28736
rect 8848 -28832 8944 -28798
rect 10790 -28832 10886 -28798
rect 11048 -28206 11144 -28172
rect 12990 -28206 13086 -28172
rect 11048 -28268 11082 -28206
rect 13052 -28268 13086 -28206
rect 11263 -28340 11279 -28306
rect 12855 -28340 12871 -28306
rect 11186 -28368 11220 -28352
rect 11186 -28652 11220 -28636
rect 12914 -28368 12948 -28352
rect 12914 -28652 12948 -28636
rect 11263 -28698 11279 -28664
rect 12855 -28698 12871 -28664
rect 11048 -28798 11082 -28736
rect 13052 -28798 13086 -28736
rect 11048 -28832 11144 -28798
rect 12990 -28832 13086 -28798
rect 13248 -28206 13344 -28172
rect 15190 -28206 15286 -28172
rect 13248 -28268 13282 -28206
rect 15252 -28268 15286 -28206
rect 13463 -28340 13479 -28306
rect 15055 -28340 15071 -28306
rect 13386 -28368 13420 -28352
rect 13386 -28652 13420 -28636
rect 15114 -28368 15148 -28352
rect 15114 -28652 15148 -28636
rect 13463 -28698 13479 -28664
rect 15055 -28698 15071 -28664
rect 13248 -28798 13282 -28736
rect 15252 -28798 15286 -28736
rect 13248 -28832 13344 -28798
rect 15190 -28832 15286 -28798
rect 15448 -28206 15544 -28172
rect 17390 -28206 17486 -28172
rect 15448 -28268 15482 -28206
rect 17452 -28268 17486 -28206
rect 15663 -28340 15679 -28306
rect 17255 -28340 17271 -28306
rect 15586 -28368 15620 -28352
rect 15586 -28652 15620 -28636
rect 17314 -28368 17348 -28352
rect 17314 -28652 17348 -28636
rect 15663 -28698 15679 -28664
rect 17255 -28698 17271 -28664
rect 15448 -28798 15482 -28736
rect 17452 -28798 17486 -28736
rect 15448 -28832 15544 -28798
rect 17390 -28832 17486 -28798
rect 17648 -28206 17744 -28172
rect 19590 -28206 19686 -28172
rect 17648 -28268 17682 -28206
rect 19652 -28268 19686 -28206
rect 17863 -28340 17879 -28306
rect 19455 -28340 19471 -28306
rect 17786 -28368 17820 -28352
rect 17786 -28652 17820 -28636
rect 19514 -28368 19548 -28352
rect 19514 -28652 19548 -28636
rect 17863 -28698 17879 -28664
rect 19455 -28698 19471 -28664
rect 17648 -28798 17682 -28736
rect 19652 -28798 19686 -28736
rect 17648 -28832 17744 -28798
rect 19590 -28832 19686 -28798
rect 19848 -28206 19944 -28172
rect 21790 -28206 22196 -28172
rect 19848 -28268 22196 -28206
rect 19882 -28306 21852 -28268
rect 19882 -28340 20079 -28306
rect 21655 -28340 21852 -28306
rect 19882 -28368 21852 -28340
rect 19882 -28636 19986 -28368
rect 20020 -28636 21714 -28368
rect 21748 -28636 21852 -28368
rect 19882 -28664 21852 -28636
rect 19882 -28698 20079 -28664
rect 21655 -28698 21852 -28664
rect 19882 -28736 21852 -28698
rect 21886 -28736 22196 -28268
rect 19848 -28798 22196 -28736
rect 19848 -28832 19944 -28798
rect 21790 -28832 22196 -28798
rect 60 -28972 2060 -28832
rect 19860 -28972 22196 -28832
rect 48 -29006 144 -28972
rect 1990 -29006 2086 -28972
rect 48 -29068 2086 -29006
rect 82 -29106 2052 -29068
rect 82 -29140 279 -29106
rect 1855 -29140 2052 -29106
rect 82 -29168 2052 -29140
rect 82 -29436 186 -29168
rect 220 -29436 1914 -29168
rect 1948 -29436 2052 -29168
rect 82 -29464 2052 -29436
rect 82 -29498 279 -29464
rect 1855 -29498 2052 -29464
rect 82 -29536 2052 -29498
rect 48 -29598 2086 -29536
rect 48 -29632 144 -29598
rect 1990 -29632 2086 -29598
rect 2248 -29006 2344 -28972
rect 4190 -29006 4286 -28972
rect 2248 -29068 2282 -29006
rect 4252 -29068 4286 -29006
rect 2463 -29140 2479 -29106
rect 4055 -29140 4071 -29106
rect 2386 -29168 2420 -29152
rect 2386 -29452 2420 -29436
rect 4114 -29168 4148 -29152
rect 4114 -29452 4148 -29436
rect 2463 -29498 2479 -29464
rect 4055 -29498 4071 -29464
rect 2248 -29598 2282 -29536
rect 4252 -29598 4286 -29536
rect 2248 -29632 2344 -29598
rect 4190 -29632 4286 -29598
rect 4448 -29006 4544 -28972
rect 6390 -29006 6486 -28972
rect 4448 -29068 4482 -29006
rect 6452 -29068 6486 -29006
rect 4663 -29140 4679 -29106
rect 6255 -29140 6271 -29106
rect 4586 -29168 4620 -29152
rect 4586 -29452 4620 -29436
rect 6314 -29168 6348 -29152
rect 6314 -29452 6348 -29436
rect 4663 -29498 4679 -29464
rect 6255 -29498 6271 -29464
rect 4448 -29598 4482 -29536
rect 6452 -29598 6486 -29536
rect 4448 -29632 4544 -29598
rect 6390 -29632 6486 -29598
rect 6648 -29006 6744 -28972
rect 8590 -29006 8686 -28972
rect 6648 -29068 6682 -29006
rect 8652 -29068 8686 -29006
rect 6863 -29140 6879 -29106
rect 8455 -29140 8471 -29106
rect 6786 -29168 6820 -29152
rect 6786 -29452 6820 -29436
rect 8514 -29168 8548 -29152
rect 8514 -29452 8548 -29436
rect 6863 -29498 6879 -29464
rect 8455 -29498 8471 -29464
rect 6648 -29598 6682 -29536
rect 8652 -29598 8686 -29536
rect 6648 -29632 6744 -29598
rect 8590 -29632 8686 -29598
rect 8848 -29006 8944 -28972
rect 10790 -29006 10886 -28972
rect 8848 -29068 8882 -29006
rect 10852 -29068 10886 -29006
rect 9063 -29140 9079 -29106
rect 10655 -29140 10671 -29106
rect 8986 -29168 9020 -29152
rect 8986 -29452 9020 -29436
rect 10714 -29168 10748 -29152
rect 10714 -29452 10748 -29436
rect 9063 -29498 9079 -29464
rect 10655 -29498 10671 -29464
rect 8848 -29598 8882 -29536
rect 10852 -29598 10886 -29536
rect 8848 -29632 8944 -29598
rect 10790 -29632 10886 -29598
rect 11048 -29006 11144 -28972
rect 12990 -29006 13086 -28972
rect 11048 -29068 11082 -29006
rect 13052 -29068 13086 -29006
rect 11263 -29140 11279 -29106
rect 12855 -29140 12871 -29106
rect 11186 -29168 11220 -29152
rect 11186 -29452 11220 -29436
rect 12914 -29168 12948 -29152
rect 12914 -29452 12948 -29436
rect 11263 -29498 11279 -29464
rect 12855 -29498 12871 -29464
rect 11048 -29598 11082 -29536
rect 13052 -29598 13086 -29536
rect 11048 -29632 11144 -29598
rect 12990 -29632 13086 -29598
rect 13248 -29006 13344 -28972
rect 15190 -29006 15286 -28972
rect 13248 -29068 13282 -29006
rect 15252 -29068 15286 -29006
rect 13463 -29140 13479 -29106
rect 15055 -29140 15071 -29106
rect 13386 -29168 13420 -29152
rect 13386 -29452 13420 -29436
rect 15114 -29168 15148 -29152
rect 15114 -29452 15148 -29436
rect 13463 -29498 13479 -29464
rect 15055 -29498 15071 -29464
rect 13248 -29598 13282 -29536
rect 15252 -29598 15286 -29536
rect 13248 -29632 13344 -29598
rect 15190 -29632 15286 -29598
rect 15448 -29006 15544 -28972
rect 17390 -29006 17486 -28972
rect 15448 -29068 15482 -29006
rect 17452 -29068 17486 -29006
rect 15663 -29140 15679 -29106
rect 17255 -29140 17271 -29106
rect 15586 -29168 15620 -29152
rect 15586 -29452 15620 -29436
rect 17314 -29168 17348 -29152
rect 17314 -29452 17348 -29436
rect 15663 -29498 15679 -29464
rect 17255 -29498 17271 -29464
rect 15448 -29598 15482 -29536
rect 17452 -29598 17486 -29536
rect 15448 -29632 15544 -29598
rect 17390 -29632 17486 -29598
rect 17648 -29006 17744 -28972
rect 19590 -29006 19686 -28972
rect 17648 -29068 17682 -29006
rect 19652 -29068 19686 -29006
rect 17863 -29140 17879 -29106
rect 19455 -29140 19471 -29106
rect 17786 -29168 17820 -29152
rect 17786 -29452 17820 -29436
rect 19514 -29168 19548 -29152
rect 19514 -29452 19548 -29436
rect 17863 -29498 17879 -29464
rect 19455 -29498 19471 -29464
rect 17648 -29598 17682 -29536
rect 19652 -29598 19686 -29536
rect 17648 -29632 17744 -29598
rect 19590 -29632 19686 -29598
rect 19848 -29006 19944 -28972
rect 21790 -29006 22196 -28972
rect 19848 -29068 22196 -29006
rect 19882 -29106 21852 -29068
rect 19882 -29140 20079 -29106
rect 21655 -29140 21852 -29106
rect 19882 -29168 21852 -29140
rect 19882 -29436 19986 -29168
rect 20020 -29436 21714 -29168
rect 21748 -29436 21852 -29168
rect 19882 -29464 21852 -29436
rect 19882 -29498 20079 -29464
rect 21655 -29498 21852 -29464
rect 19882 -29536 21852 -29498
rect 21886 -29536 22196 -29068
rect 19848 -29598 22196 -29536
rect 19848 -29632 19944 -29598
rect 21790 -29632 22196 -29598
rect 60 -29772 2060 -29632
rect 19860 -29772 22196 -29632
rect 48 -29806 144 -29772
rect 1990 -29806 2086 -29772
rect 48 -29868 2086 -29806
rect 82 -29906 2052 -29868
rect 82 -29940 279 -29906
rect 1855 -29940 2052 -29906
rect 82 -29968 2052 -29940
rect 82 -30236 186 -29968
rect 220 -30236 1914 -29968
rect 1948 -30236 2052 -29968
rect 82 -30264 2052 -30236
rect 82 -30298 279 -30264
rect 1855 -30298 2052 -30264
rect 82 -30336 2052 -30298
rect 48 -30398 2086 -30336
rect 48 -30432 144 -30398
rect 1990 -30432 2086 -30398
rect 2248 -29806 2344 -29772
rect 4190 -29806 4286 -29772
rect 2248 -29868 2282 -29806
rect 4252 -29868 4286 -29806
rect 2463 -29940 2479 -29906
rect 4055 -29940 4071 -29906
rect 2386 -29968 2420 -29952
rect 2386 -30252 2420 -30236
rect 4114 -29968 4148 -29952
rect 4114 -30252 4148 -30236
rect 2463 -30298 2479 -30264
rect 4055 -30298 4071 -30264
rect 2248 -30398 2282 -30336
rect 4252 -30398 4286 -30336
rect 2248 -30432 2344 -30398
rect 4190 -30432 4286 -30398
rect 4448 -29806 4544 -29772
rect 6390 -29806 6486 -29772
rect 4448 -29868 4482 -29806
rect 6452 -29868 6486 -29806
rect 4663 -29940 4679 -29906
rect 6255 -29940 6271 -29906
rect 4586 -29968 4620 -29952
rect 4586 -30252 4620 -30236
rect 6314 -29968 6348 -29952
rect 6314 -30252 6348 -30236
rect 4663 -30298 4679 -30264
rect 6255 -30298 6271 -30264
rect 4448 -30398 4482 -30336
rect 6452 -30398 6486 -30336
rect 4448 -30432 4544 -30398
rect 6390 -30432 6486 -30398
rect 6648 -29806 6744 -29772
rect 8590 -29806 8686 -29772
rect 6648 -29868 6682 -29806
rect 8652 -29868 8686 -29806
rect 6863 -29940 6879 -29906
rect 8455 -29940 8471 -29906
rect 6786 -29968 6820 -29952
rect 6786 -30252 6820 -30236
rect 8514 -29968 8548 -29952
rect 8514 -30252 8548 -30236
rect 6863 -30298 6879 -30264
rect 8455 -30298 8471 -30264
rect 6648 -30398 6682 -30336
rect 8652 -30398 8686 -30336
rect 6648 -30432 6744 -30398
rect 8590 -30432 8686 -30398
rect 8848 -29806 8944 -29772
rect 10790 -29806 10886 -29772
rect 8848 -29868 8882 -29806
rect 10852 -29868 10886 -29806
rect 9063 -29940 9079 -29906
rect 10655 -29940 10671 -29906
rect 8986 -29968 9020 -29952
rect 8986 -30252 9020 -30236
rect 10714 -29968 10748 -29952
rect 10714 -30252 10748 -30236
rect 9063 -30298 9079 -30264
rect 10655 -30298 10671 -30264
rect 8848 -30398 8882 -30336
rect 10852 -30398 10886 -30336
rect 8848 -30432 8944 -30398
rect 10790 -30432 10886 -30398
rect 11048 -29806 11144 -29772
rect 12990 -29806 13086 -29772
rect 11048 -29868 11082 -29806
rect 13052 -29868 13086 -29806
rect 11263 -29940 11279 -29906
rect 12855 -29940 12871 -29906
rect 11186 -29968 11220 -29952
rect 11186 -30252 11220 -30236
rect 12914 -29968 12948 -29952
rect 12914 -30252 12948 -30236
rect 11263 -30298 11279 -30264
rect 12855 -30298 12871 -30264
rect 11048 -30398 11082 -30336
rect 13052 -30398 13086 -30336
rect 11048 -30432 11144 -30398
rect 12990 -30432 13086 -30398
rect 13248 -29806 13344 -29772
rect 15190 -29806 15286 -29772
rect 13248 -29868 13282 -29806
rect 15252 -29868 15286 -29806
rect 13463 -29940 13479 -29906
rect 15055 -29940 15071 -29906
rect 13386 -29968 13420 -29952
rect 13386 -30252 13420 -30236
rect 15114 -29968 15148 -29952
rect 15114 -30252 15148 -30236
rect 13463 -30298 13479 -30264
rect 15055 -30298 15071 -30264
rect 13248 -30398 13282 -30336
rect 15252 -30398 15286 -30336
rect 13248 -30432 13344 -30398
rect 15190 -30432 15286 -30398
rect 15448 -29806 15544 -29772
rect 17390 -29806 17486 -29772
rect 15448 -29868 15482 -29806
rect 17452 -29868 17486 -29806
rect 15663 -29940 15679 -29906
rect 17255 -29940 17271 -29906
rect 15586 -29968 15620 -29952
rect 15586 -30252 15620 -30236
rect 17314 -29968 17348 -29952
rect 17314 -30252 17348 -30236
rect 15663 -30298 15679 -30264
rect 17255 -30298 17271 -30264
rect 15448 -30398 15482 -30336
rect 17452 -30398 17486 -30336
rect 15448 -30432 15544 -30398
rect 17390 -30432 17486 -30398
rect 17648 -29806 17744 -29772
rect 19590 -29806 19686 -29772
rect 17648 -29868 17682 -29806
rect 19652 -29868 19686 -29806
rect 17863 -29940 17879 -29906
rect 19455 -29940 19471 -29906
rect 17786 -29968 17820 -29952
rect 17786 -30252 17820 -30236
rect 19514 -29968 19548 -29952
rect 19514 -30252 19548 -30236
rect 17863 -30298 17879 -30264
rect 19455 -30298 19471 -30264
rect 17648 -30398 17682 -30336
rect 19652 -30398 19686 -30336
rect 17648 -30432 17744 -30398
rect 19590 -30432 19686 -30398
rect 19848 -29806 19944 -29772
rect 21790 -29806 22196 -29772
rect 19848 -29868 22196 -29806
rect 19882 -29906 21852 -29868
rect 19882 -29940 20079 -29906
rect 21655 -29940 21852 -29906
rect 19882 -29968 21852 -29940
rect 19882 -30236 19986 -29968
rect 20020 -30236 21714 -29968
rect 21748 -30236 21852 -29968
rect 19882 -30264 21852 -30236
rect 19882 -30298 20079 -30264
rect 21655 -30298 21852 -30264
rect 19882 -30336 21852 -30298
rect 21886 -30336 22196 -29868
rect 19848 -30398 22196 -30336
rect 19848 -30432 19944 -30398
rect 21790 -30432 22196 -30398
rect 60 -30572 2060 -30432
rect 19860 -30572 22196 -30432
rect 48 -30606 144 -30572
rect 1990 -30606 2086 -30572
rect 48 -30668 2086 -30606
rect 82 -30706 2052 -30668
rect 82 -30740 279 -30706
rect 1855 -30740 2052 -30706
rect 82 -30768 2052 -30740
rect 82 -31036 186 -30768
rect 220 -31036 1914 -30768
rect 1948 -31036 2052 -30768
rect 82 -31064 2052 -31036
rect 82 -31098 279 -31064
rect 1855 -31098 2052 -31064
rect 82 -31136 2052 -31098
rect 48 -31198 2086 -31136
rect 48 -31232 144 -31198
rect 1990 -31232 2086 -31198
rect 2248 -30606 2344 -30572
rect 4190 -30606 4286 -30572
rect 2248 -30668 2282 -30606
rect 4252 -30668 4286 -30606
rect 2463 -30740 2479 -30706
rect 4055 -30740 4071 -30706
rect 2386 -30768 2420 -30752
rect 2386 -31052 2420 -31036
rect 4114 -30768 4148 -30752
rect 4114 -31052 4148 -31036
rect 2463 -31098 2479 -31064
rect 4055 -31098 4071 -31064
rect 2248 -31198 2282 -31136
rect 4252 -31198 4286 -31136
rect 2248 -31232 2344 -31198
rect 4190 -31232 4286 -31198
rect 4448 -30606 4544 -30572
rect 6390 -30606 6486 -30572
rect 4448 -30668 4482 -30606
rect 6452 -30668 6486 -30606
rect 4663 -30740 4679 -30706
rect 6255 -30740 6271 -30706
rect 4586 -30768 4620 -30752
rect 4586 -31052 4620 -31036
rect 6314 -30768 6348 -30752
rect 6314 -31052 6348 -31036
rect 4663 -31098 4679 -31064
rect 6255 -31098 6271 -31064
rect 4448 -31198 4482 -31136
rect 6452 -31198 6486 -31136
rect 4448 -31232 4544 -31198
rect 6390 -31232 6486 -31198
rect 6648 -30606 6744 -30572
rect 8590 -30606 8686 -30572
rect 6648 -30668 6682 -30606
rect 8652 -30668 8686 -30606
rect 6863 -30740 6879 -30706
rect 8455 -30740 8471 -30706
rect 6786 -30768 6820 -30752
rect 6786 -31052 6820 -31036
rect 8514 -30768 8548 -30752
rect 8514 -31052 8548 -31036
rect 6863 -31098 6879 -31064
rect 8455 -31098 8471 -31064
rect 6648 -31198 6682 -31136
rect 8652 -31198 8686 -31136
rect 6648 -31232 6744 -31198
rect 8590 -31232 8686 -31198
rect 8848 -30606 8944 -30572
rect 10790 -30606 10886 -30572
rect 8848 -30668 8882 -30606
rect 10852 -30668 10886 -30606
rect 9063 -30740 9079 -30706
rect 10655 -30740 10671 -30706
rect 8986 -30768 9020 -30752
rect 8986 -31052 9020 -31036
rect 10714 -30768 10748 -30752
rect 10714 -31052 10748 -31036
rect 9063 -31098 9079 -31064
rect 10655 -31098 10671 -31064
rect 8848 -31198 8882 -31136
rect 10852 -31198 10886 -31136
rect 8848 -31232 8944 -31198
rect 10790 -31232 10886 -31198
rect 11048 -30606 11144 -30572
rect 12990 -30606 13086 -30572
rect 11048 -30668 11082 -30606
rect 13052 -30668 13086 -30606
rect 11263 -30740 11279 -30706
rect 12855 -30740 12871 -30706
rect 11186 -30768 11220 -30752
rect 11186 -31052 11220 -31036
rect 12914 -30768 12948 -30752
rect 12914 -31052 12948 -31036
rect 11263 -31098 11279 -31064
rect 12855 -31098 12871 -31064
rect 11048 -31198 11082 -31136
rect 13052 -31198 13086 -31136
rect 11048 -31232 11144 -31198
rect 12990 -31232 13086 -31198
rect 13248 -30606 13344 -30572
rect 15190 -30606 15286 -30572
rect 13248 -30668 13282 -30606
rect 15252 -30668 15286 -30606
rect 13463 -30740 13479 -30706
rect 15055 -30740 15071 -30706
rect 13386 -30768 13420 -30752
rect 13386 -31052 13420 -31036
rect 15114 -30768 15148 -30752
rect 15114 -31052 15148 -31036
rect 13463 -31098 13479 -31064
rect 15055 -31098 15071 -31064
rect 13248 -31198 13282 -31136
rect 15252 -31198 15286 -31136
rect 13248 -31232 13344 -31198
rect 15190 -31232 15286 -31198
rect 15448 -30606 15544 -30572
rect 17390 -30606 17486 -30572
rect 15448 -30668 15482 -30606
rect 17452 -30668 17486 -30606
rect 15663 -30740 15679 -30706
rect 17255 -30740 17271 -30706
rect 15586 -30768 15620 -30752
rect 15586 -31052 15620 -31036
rect 17314 -30768 17348 -30752
rect 17314 -31052 17348 -31036
rect 15663 -31098 15679 -31064
rect 17255 -31098 17271 -31064
rect 15448 -31198 15482 -31136
rect 17452 -31198 17486 -31136
rect 15448 -31232 15544 -31198
rect 17390 -31232 17486 -31198
rect 17648 -30606 17744 -30572
rect 19590 -30606 19686 -30572
rect 17648 -30668 17682 -30606
rect 19652 -30668 19686 -30606
rect 17863 -30740 17879 -30706
rect 19455 -30740 19471 -30706
rect 17786 -30768 17820 -30752
rect 17786 -31052 17820 -31036
rect 19514 -30768 19548 -30752
rect 19514 -31052 19548 -31036
rect 17863 -31098 17879 -31064
rect 19455 -31098 19471 -31064
rect 17648 -31198 17682 -31136
rect 19652 -31198 19686 -31136
rect 17648 -31232 17744 -31198
rect 19590 -31232 19686 -31198
rect 19848 -30606 19944 -30572
rect 21790 -30606 22196 -30572
rect 19848 -30668 22196 -30606
rect 19882 -30706 21852 -30668
rect 19882 -30740 20079 -30706
rect 21655 -30740 21852 -30706
rect 19882 -30768 21852 -30740
rect 19882 -31036 19986 -30768
rect 20020 -31036 21714 -30768
rect 21748 -31036 21852 -30768
rect 19882 -31064 21852 -31036
rect 19882 -31098 20079 -31064
rect 21655 -31098 21852 -31064
rect 19882 -31136 21852 -31098
rect 21886 -31136 22196 -30668
rect 19848 -31198 22196 -31136
rect 19848 -31232 19944 -31198
rect 21790 -31232 22196 -31198
rect 60 -31372 2060 -31232
rect 19860 -31372 22196 -31232
rect 48 -31406 144 -31372
rect 1990 -31380 2086 -31372
rect 2248 -31380 2344 -31372
rect 1990 -31406 2344 -31380
rect 4190 -31380 4286 -31372
rect 4448 -31380 4544 -31372
rect 4190 -31406 4544 -31380
rect 6390 -31380 6486 -31372
rect 6648 -31380 6744 -31372
rect 6390 -31406 6744 -31380
rect 8590 -31380 8686 -31372
rect 8848 -31380 8944 -31372
rect 8590 -31406 8944 -31380
rect 10790 -31380 10886 -31372
rect 11048 -31380 11144 -31372
rect 10790 -31406 11144 -31380
rect 12990 -31380 13086 -31372
rect 13248 -31380 13344 -31372
rect 12990 -31406 13344 -31380
rect 15190 -31380 15286 -31372
rect 15448 -31380 15544 -31372
rect 15190 -31406 15544 -31380
rect 17390 -31380 17486 -31372
rect 17648 -31380 17744 -31372
rect 17390 -31406 17744 -31380
rect 19590 -31380 19686 -31372
rect 19848 -31380 19944 -31372
rect 19590 -31406 19944 -31380
rect 21790 -31406 22196 -31372
rect 48 -31468 22196 -31406
rect 82 -31506 2052 -31468
rect 82 -31540 279 -31506
rect 1855 -31540 2052 -31506
rect 82 -31568 2052 -31540
rect 82 -31836 186 -31568
rect 220 -31836 1914 -31568
rect 1948 -31836 2052 -31568
rect 82 -31864 2052 -31836
rect 82 -31898 279 -31864
rect 1855 -31898 2052 -31864
rect 82 -31936 2052 -31898
rect 2086 -31936 2248 -31468
rect 2282 -31506 4252 -31468
rect 2282 -31540 2479 -31506
rect 4055 -31540 4252 -31506
rect 2282 -31568 4252 -31540
rect 2282 -31836 2386 -31568
rect 2420 -31836 4114 -31568
rect 4148 -31836 4252 -31568
rect 2282 -31864 4252 -31836
rect 2282 -31898 2479 -31864
rect 4055 -31898 4252 -31864
rect 2282 -31936 4252 -31898
rect 4286 -31936 4448 -31468
rect 4482 -31506 6452 -31468
rect 4482 -31540 4679 -31506
rect 6255 -31540 6452 -31506
rect 4482 -31568 6452 -31540
rect 4482 -31836 4586 -31568
rect 4620 -31836 6314 -31568
rect 6348 -31836 6452 -31568
rect 4482 -31864 6452 -31836
rect 4482 -31898 4679 -31864
rect 6255 -31898 6452 -31864
rect 4482 -31936 6452 -31898
rect 6486 -31936 6648 -31468
rect 6682 -31506 8652 -31468
rect 6682 -31540 6879 -31506
rect 8455 -31540 8652 -31506
rect 6682 -31568 8652 -31540
rect 6682 -31836 6786 -31568
rect 6820 -31836 8514 -31568
rect 8548 -31836 8652 -31568
rect 6682 -31864 8652 -31836
rect 6682 -31898 6879 -31864
rect 8455 -31898 8652 -31864
rect 6682 -31936 8652 -31898
rect 8686 -31936 8848 -31468
rect 8882 -31506 10852 -31468
rect 8882 -31540 9079 -31506
rect 10655 -31540 10852 -31506
rect 8882 -31568 10852 -31540
rect 8882 -31836 8986 -31568
rect 9020 -31836 10714 -31568
rect 10748 -31836 10852 -31568
rect 8882 -31864 10852 -31836
rect 8882 -31898 9079 -31864
rect 10655 -31898 10852 -31864
rect 8882 -31936 10852 -31898
rect 10886 -31936 11048 -31468
rect 11082 -31506 13052 -31468
rect 11082 -31540 11279 -31506
rect 12855 -31540 13052 -31506
rect 11082 -31568 13052 -31540
rect 11082 -31836 11186 -31568
rect 11220 -31836 12914 -31568
rect 12948 -31836 13052 -31568
rect 11082 -31864 13052 -31836
rect 11082 -31898 11279 -31864
rect 12855 -31898 13052 -31864
rect 11082 -31936 13052 -31898
rect 13086 -31936 13248 -31468
rect 13282 -31506 15252 -31468
rect 13282 -31540 13479 -31506
rect 15055 -31540 15252 -31506
rect 13282 -31568 15252 -31540
rect 13282 -31836 13386 -31568
rect 13420 -31836 15114 -31568
rect 15148 -31836 15252 -31568
rect 13282 -31864 15252 -31836
rect 13282 -31898 13479 -31864
rect 15055 -31898 15252 -31864
rect 13282 -31936 15252 -31898
rect 15286 -31936 15448 -31468
rect 15482 -31506 17452 -31468
rect 15482 -31540 15679 -31506
rect 17255 -31540 17452 -31506
rect 15482 -31568 17452 -31540
rect 15482 -31836 15586 -31568
rect 15620 -31836 17314 -31568
rect 17348 -31836 17452 -31568
rect 15482 -31864 17452 -31836
rect 15482 -31898 15679 -31864
rect 17255 -31898 17452 -31864
rect 15482 -31936 17452 -31898
rect 17486 -31936 17648 -31468
rect 17682 -31506 19652 -31468
rect 17682 -31540 17879 -31506
rect 19455 -31540 19652 -31506
rect 17682 -31568 19652 -31540
rect 17682 -31836 17786 -31568
rect 17820 -31836 19514 -31568
rect 19548 -31836 19652 -31568
rect 17682 -31864 19652 -31836
rect 17682 -31898 17879 -31864
rect 19455 -31898 19652 -31864
rect 17682 -31936 19652 -31898
rect 19686 -31936 19848 -31468
rect 19882 -31506 21852 -31468
rect 19882 -31540 20079 -31506
rect 21655 -31540 21852 -31506
rect 19882 -31568 21852 -31540
rect 19882 -31836 19986 -31568
rect 20020 -31836 21714 -31568
rect 21748 -31836 21852 -31568
rect 19882 -31864 21852 -31836
rect 19882 -31898 20079 -31864
rect 21655 -31898 21852 -31864
rect 19882 -31936 21852 -31898
rect 21886 -31936 22196 -31468
rect 22230 -25060 22347 -24665
rect 27020 -24680 27030 -24610
rect 26913 -25080 27030 -24680
rect 48 -31968 22196 -31936
rect 22230 -31900 22347 -31500
rect 27020 -31500 27030 -25080
rect 26913 -31880 27030 -31500
rect 48 -31998 22230 -31968
rect 48 -32032 144 -31998
rect 1990 -32020 2344 -31998
rect 1990 -32032 2086 -32020
rect 2248 -32032 2344 -32020
rect 4190 -32020 4544 -31998
rect 4190 -32032 4286 -32020
rect 4448 -32032 4544 -32020
rect 6390 -32020 6744 -31998
rect 6390 -32032 6486 -32020
rect 6648 -32032 6744 -32020
rect 8590 -32020 8944 -31998
rect 8590 -32032 8686 -32020
rect 8848 -32032 8944 -32020
rect 10790 -32020 11144 -31998
rect 10790 -32032 10886 -32020
rect 11048 -32032 11144 -32020
rect 12990 -32020 13344 -31998
rect 12990 -32032 13086 -32020
rect 13248 -32032 13344 -32020
rect 15190 -32020 15544 -31998
rect 15190 -32032 15286 -32020
rect 15448 -32032 15544 -32020
rect 17390 -32020 17744 -31998
rect 17390 -32032 17486 -32020
rect 17648 -32032 17744 -32020
rect 19590 -32020 19944 -31998
rect 19590 -32032 19686 -32020
rect 19848 -32032 19944 -32020
rect 21790 -32010 22230 -31998
rect 21790 -32020 22040 -32010
rect 22140 -32020 22230 -32010
rect 21790 -32032 21886 -32020
rect 22196 -32030 22230 -32020
rect 22360 -32030 22900 -31913
rect 26360 -32030 26900 -31913
rect 27020 -31968 27030 -31880
rect 27064 -31968 27130 -24610
rect 27020 -32030 27130 -31968
rect 22196 -32064 22292 -32030
rect 26968 -32060 27130 -32030
rect 27430 -24502 29820 -24320
rect 33036 -24350 33070 -24288
rect 34252 -24350 34286 -24288
rect 33036 -24384 33132 -24350
rect 34190 -24384 34286 -24350
rect 34408 -23578 34504 -23544
rect 37142 -23578 37238 -23544
rect 34408 -23640 34442 -23578
rect 37204 -23640 37238 -23578
rect 34588 -23716 34604 -23682
rect 34672 -23716 34688 -23682
rect 34746 -23716 34762 -23682
rect 34830 -23716 34846 -23682
rect 34904 -23716 34920 -23682
rect 34988 -23716 35004 -23682
rect 35062 -23716 35078 -23682
rect 35146 -23716 35162 -23682
rect 35220 -23716 35236 -23682
rect 35304 -23716 35320 -23682
rect 35378 -23716 35394 -23682
rect 35462 -23716 35478 -23682
rect 35536 -23716 35552 -23682
rect 35620 -23716 35636 -23682
rect 35694 -23716 35710 -23682
rect 35778 -23716 35794 -23682
rect 35852 -23716 35868 -23682
rect 35936 -23716 35952 -23682
rect 36010 -23716 36026 -23682
rect 36094 -23716 36110 -23682
rect 36168 -23716 36184 -23682
rect 36252 -23716 36268 -23682
rect 36326 -23716 36342 -23682
rect 36410 -23716 36426 -23682
rect 36484 -23716 36500 -23682
rect 36568 -23716 36584 -23682
rect 36642 -23716 36658 -23682
rect 36726 -23716 36742 -23682
rect 36800 -23716 36816 -23682
rect 36884 -23716 36900 -23682
rect 36958 -23716 36974 -23682
rect 37042 -23716 37058 -23682
rect 34542 -23775 34576 -23759
rect 34542 -24167 34576 -24151
rect 34700 -23775 34734 -23759
rect 34700 -24167 34734 -24151
rect 34858 -23775 34892 -23759
rect 34858 -24167 34892 -24151
rect 35016 -23775 35050 -23759
rect 35016 -24167 35050 -24151
rect 35174 -23775 35208 -23759
rect 35174 -24167 35208 -24151
rect 35332 -23775 35366 -23759
rect 35332 -24167 35366 -24151
rect 35490 -23775 35524 -23759
rect 35490 -24167 35524 -24151
rect 35648 -23775 35682 -23759
rect 35648 -24167 35682 -24151
rect 35806 -23775 35840 -23759
rect 35806 -24167 35840 -24151
rect 35964 -23775 35998 -23759
rect 35964 -24167 35998 -24151
rect 36122 -23775 36156 -23759
rect 36122 -24167 36156 -24151
rect 36280 -23775 36314 -23759
rect 36280 -24167 36314 -24151
rect 36438 -23775 36472 -23759
rect 36438 -24167 36472 -24151
rect 36596 -23775 36630 -23759
rect 36596 -24167 36630 -24151
rect 36754 -23775 36788 -23759
rect 36754 -24167 36788 -24151
rect 36912 -23775 36946 -23759
rect 36912 -24167 36946 -24151
rect 37070 -23775 37104 -23759
rect 37070 -24167 37104 -24151
rect 34588 -24244 34604 -24210
rect 34672 -24244 34688 -24210
rect 34746 -24244 34762 -24210
rect 34830 -24244 34846 -24210
rect 34904 -24244 34920 -24210
rect 34988 -24244 35004 -24210
rect 35062 -24244 35078 -24210
rect 35146 -24244 35162 -24210
rect 35220 -24244 35236 -24210
rect 35304 -24244 35320 -24210
rect 35378 -24244 35394 -24210
rect 35462 -24244 35478 -24210
rect 35536 -24244 35552 -24210
rect 35620 -24244 35636 -24210
rect 35694 -24244 35710 -24210
rect 35778 -24244 35794 -24210
rect 35852 -24244 35868 -24210
rect 35936 -24244 35952 -24210
rect 36010 -24244 36026 -24210
rect 36094 -24244 36110 -24210
rect 36168 -24244 36184 -24210
rect 36252 -24244 36268 -24210
rect 36326 -24244 36342 -24210
rect 36410 -24244 36426 -24210
rect 36484 -24244 36500 -24210
rect 36568 -24244 36584 -24210
rect 36642 -24244 36658 -24210
rect 36726 -24244 36742 -24210
rect 36800 -24244 36816 -24210
rect 36884 -24244 36900 -24210
rect 36958 -24244 36974 -24210
rect 37042 -24244 37058 -24210
rect 34408 -24348 34442 -24286
rect 37204 -24348 37238 -24286
rect 34408 -24382 34504 -24348
rect 37142 -24382 37238 -24348
rect 27430 -24536 27884 -24502
rect 28852 -24536 29820 -24502
rect 27430 -24598 27822 -24536
rect 27430 -25226 27788 -24598
rect 28914 -24598 29820 -24536
rect 27968 -24674 27984 -24640
rect 28752 -24674 28768 -24640
rect 27922 -24724 27956 -24708
rect 27922 -25116 27956 -25100
rect 28780 -24724 28814 -24708
rect 28780 -25116 28814 -25100
rect 27968 -25184 27984 -25150
rect 28752 -25184 28768 -25150
rect 27430 -25288 27822 -25226
rect 28948 -25226 29820 -24598
rect 28914 -25288 29820 -25226
rect 27430 -25322 27884 -25288
rect 28852 -25322 29820 -25288
rect 27430 -25408 29820 -25322
rect 27430 -25442 27884 -25408
rect 28850 -25442 29820 -25408
rect 27430 -25504 27822 -25442
rect 27430 -26246 27788 -25504
rect 28912 -25504 29820 -25442
rect 27932 -25576 27948 -25542
rect 28724 -25576 28740 -25542
rect 28774 -25604 28808 -25588
rect 28774 -25688 28808 -25672
rect 27932 -25734 27948 -25700
rect 28724 -25734 28740 -25700
rect 28774 -25762 28808 -25746
rect 28774 -25846 28808 -25830
rect 27932 -25892 27948 -25858
rect 28724 -25892 28740 -25858
rect 28774 -25920 28808 -25904
rect 28774 -26004 28808 -25988
rect 27932 -26050 27948 -26016
rect 28724 -26050 28740 -26016
rect 28774 -26078 28808 -26062
rect 28774 -26162 28808 -26146
rect 27932 -26208 27948 -26174
rect 28724 -26208 28740 -26174
rect 27430 -26308 27822 -26246
rect 28946 -26246 29820 -25504
rect 28912 -26308 29820 -26246
rect 27430 -26342 27884 -26308
rect 28850 -26342 29820 -26308
rect 27430 -26448 29820 -26342
rect 27430 -26482 27884 -26448
rect 28850 -26482 29820 -26448
rect 27430 -26544 27822 -26482
rect 27430 -27286 27788 -26544
rect 28912 -26544 29820 -26482
rect 27932 -26616 27948 -26582
rect 28724 -26616 28740 -26582
rect 28774 -26644 28808 -26628
rect 28774 -26728 28808 -26712
rect 27932 -26774 27948 -26740
rect 28724 -26774 28740 -26740
rect 28774 -26802 28808 -26786
rect 28774 -26886 28808 -26870
rect 27932 -26932 27948 -26898
rect 28724 -26932 28740 -26898
rect 28774 -26960 28808 -26944
rect 28774 -27044 28808 -27028
rect 27932 -27090 27948 -27056
rect 28724 -27090 28740 -27056
rect 28774 -27118 28808 -27102
rect 28774 -27202 28808 -27186
rect 27932 -27248 27948 -27214
rect 28724 -27248 28740 -27214
rect 27430 -27348 27822 -27286
rect 28946 -27286 29820 -26544
rect 34758 -24730 34854 -24696
rect 35900 -24730 35996 -24696
rect 34758 -24792 34792 -24730
rect 35962 -24792 35996 -24730
rect 34973 -24864 34989 -24830
rect 35765 -24864 35781 -24830
rect 34896 -24892 34930 -24876
rect 34896 -25076 34930 -25060
rect 35824 -24892 35858 -24876
rect 35824 -25076 35858 -25060
rect 34973 -25122 34989 -25088
rect 35765 -25122 35781 -25088
rect 34896 -25150 34930 -25134
rect 34896 -25334 34930 -25318
rect 35824 -25150 35858 -25134
rect 35824 -25334 35858 -25318
rect 34973 -25380 34989 -25346
rect 35765 -25380 35781 -25346
rect 34896 -25408 34930 -25392
rect 34896 -25592 34930 -25576
rect 35824 -25408 35858 -25392
rect 35824 -25592 35858 -25576
rect 34973 -25638 34989 -25604
rect 35765 -25638 35781 -25604
rect 34896 -25666 34930 -25650
rect 34896 -25850 34930 -25834
rect 35824 -25666 35858 -25650
rect 35824 -25850 35858 -25834
rect 34973 -25896 34989 -25862
rect 35765 -25896 35781 -25862
rect 34896 -25924 34930 -25908
rect 34896 -26108 34930 -26092
rect 35824 -25924 35858 -25908
rect 35824 -26108 35858 -26092
rect 34973 -26154 34989 -26120
rect 35765 -26154 35781 -26120
rect 34896 -26182 34930 -26166
rect 34896 -26366 34930 -26350
rect 35824 -26182 35858 -26166
rect 35824 -26366 35858 -26350
rect 34973 -26412 34989 -26378
rect 35765 -26412 35781 -26378
rect 34896 -26440 34930 -26424
rect 34896 -26624 34930 -26608
rect 35824 -26440 35858 -26424
rect 35824 -26624 35858 -26608
rect 34973 -26670 34989 -26636
rect 35765 -26670 35781 -26636
rect 34896 -26698 34930 -26682
rect 34896 -26882 34930 -26866
rect 35824 -26698 35858 -26682
rect 35824 -26882 35858 -26866
rect 34973 -26928 34989 -26894
rect 35765 -26928 35781 -26894
rect 34758 -27028 34792 -26966
rect 35962 -27028 35996 -26966
rect 34758 -27062 34854 -27028
rect 35900 -27062 35996 -27028
rect 36098 -24730 36194 -24696
rect 37240 -24730 37336 -24696
rect 36098 -24792 36132 -24730
rect 37302 -24792 37336 -24730
rect 36313 -24864 36329 -24830
rect 37105 -24864 37121 -24830
rect 36236 -24892 36270 -24876
rect 36236 -25076 36270 -25060
rect 37164 -24892 37198 -24876
rect 37164 -25076 37198 -25060
rect 36313 -25122 36329 -25088
rect 37105 -25122 37121 -25088
rect 36236 -25150 36270 -25134
rect 36236 -25334 36270 -25318
rect 37164 -25150 37198 -25134
rect 37164 -25334 37198 -25318
rect 36313 -25380 36329 -25346
rect 37105 -25380 37121 -25346
rect 36236 -25408 36270 -25392
rect 36236 -25592 36270 -25576
rect 37164 -25408 37198 -25392
rect 37164 -25592 37198 -25576
rect 36313 -25638 36329 -25604
rect 37105 -25638 37121 -25604
rect 36236 -25666 36270 -25650
rect 36236 -25850 36270 -25834
rect 37164 -25666 37198 -25650
rect 37164 -25850 37198 -25834
rect 36313 -25896 36329 -25862
rect 37105 -25896 37121 -25862
rect 36236 -25924 36270 -25908
rect 36236 -26108 36270 -26092
rect 37164 -25924 37198 -25908
rect 37164 -26108 37198 -26092
rect 36313 -26154 36329 -26120
rect 37105 -26154 37121 -26120
rect 36236 -26182 36270 -26166
rect 36236 -26366 36270 -26350
rect 37164 -26182 37198 -26166
rect 37164 -26366 37198 -26350
rect 36313 -26412 36329 -26378
rect 37105 -26412 37121 -26378
rect 36236 -26440 36270 -26424
rect 36236 -26624 36270 -26608
rect 37164 -26440 37198 -26424
rect 37164 -26624 37198 -26608
rect 36313 -26670 36329 -26636
rect 37105 -26670 37121 -26636
rect 36236 -26698 36270 -26682
rect 36236 -26882 36270 -26866
rect 37164 -26698 37198 -26682
rect 37164 -26882 37198 -26866
rect 36313 -26928 36329 -26894
rect 37105 -26928 37121 -26894
rect 36098 -27028 36132 -26966
rect 37302 -27028 37336 -26966
rect 36098 -27062 36194 -27028
rect 37240 -27062 37336 -27028
rect 28912 -27348 29820 -27286
rect 27430 -27382 27884 -27348
rect 28850 -27382 29820 -27348
rect 27430 -27488 29820 -27382
rect 27430 -27522 27884 -27488
rect 28850 -27522 29820 -27488
rect 27430 -27584 27822 -27522
rect 27430 -28326 27788 -27584
rect 28912 -27584 29820 -27522
rect 27932 -27656 27948 -27622
rect 28724 -27656 28740 -27622
rect 28774 -27684 28808 -27668
rect 28774 -27768 28808 -27752
rect 27932 -27814 27948 -27780
rect 28724 -27814 28740 -27780
rect 28774 -27842 28808 -27826
rect 28774 -27926 28808 -27910
rect 27932 -27972 27948 -27938
rect 28724 -27972 28740 -27938
rect 28774 -28000 28808 -27984
rect 28774 -28084 28808 -28068
rect 27932 -28130 27948 -28096
rect 28724 -28130 28740 -28096
rect 28774 -28158 28808 -28142
rect 28774 -28242 28808 -28226
rect 27932 -28288 27948 -28254
rect 28724 -28288 28740 -28254
rect 27430 -28388 27822 -28326
rect 28946 -28326 29820 -27584
rect 28912 -28388 29820 -28326
rect 27430 -28422 27884 -28388
rect 28850 -28422 29820 -28388
rect 27430 -28528 29820 -28422
rect 27430 -28562 27884 -28528
rect 28850 -28562 29820 -28528
rect 27430 -28624 27822 -28562
rect 27430 -29366 27788 -28624
rect 28912 -28624 29820 -28562
rect 27932 -28696 27948 -28662
rect 28724 -28696 28740 -28662
rect 28774 -28724 28808 -28708
rect 28774 -28808 28808 -28792
rect 27932 -28854 27948 -28820
rect 28724 -28854 28740 -28820
rect 28774 -28882 28808 -28866
rect 28774 -28966 28808 -28950
rect 27932 -29012 27948 -28978
rect 28724 -29012 28740 -28978
rect 28774 -29040 28808 -29024
rect 28774 -29124 28808 -29108
rect 27932 -29170 27948 -29136
rect 28724 -29170 28740 -29136
rect 28774 -29198 28808 -29182
rect 28774 -29282 28808 -29266
rect 27932 -29328 27948 -29294
rect 28724 -29328 28740 -29294
rect 27430 -29428 27822 -29366
rect 28946 -29366 29820 -28624
rect 31678 -28398 31712 -28302
rect 32104 -28398 32152 -28302
rect 31858 -28474 31874 -28440
rect 31942 -28474 31958 -28440
rect 31812 -28533 31846 -28517
rect 31812 -28925 31846 -28909
rect 31970 -28533 32004 -28517
rect 31970 -28925 32004 -28909
rect 31858 -29002 31874 -28968
rect 31942 -29002 31958 -28968
rect 31678 -29106 31712 -29044
rect 32138 -29044 32152 -28398
rect 32298 -28474 32314 -28440
rect 32382 -28474 32398 -28440
rect 32252 -28533 32286 -28517
rect 32252 -28925 32286 -28909
rect 32410 -28533 32444 -28517
rect 32410 -28925 32444 -28909
rect 32298 -29002 32314 -28968
rect 32382 -29002 32398 -28968
rect 32104 -29106 32152 -29044
rect 32544 -29106 32592 -28302
rect 32738 -28474 32754 -28440
rect 32822 -28474 32838 -28440
rect 32692 -28533 32726 -28517
rect 32692 -28925 32726 -28909
rect 32850 -28533 32884 -28517
rect 32984 -28602 33018 -28302
rect 33878 -28398 33912 -28302
rect 32850 -28925 32884 -28909
rect 32972 -28636 33068 -28602
rect 33636 -28636 33732 -28602
rect 32972 -28683 33018 -28636
rect 32738 -29002 32754 -28968
rect 32822 -29002 32838 -28968
rect 33006 -29059 33018 -28683
rect 33698 -28698 33732 -28636
rect 33152 -28774 33168 -28740
rect 33536 -28774 33552 -28740
rect 33106 -28833 33140 -28817
rect 33106 -28925 33140 -28909
rect 33564 -28833 33598 -28817
rect 33564 -28925 33598 -28909
rect 33152 -29002 33168 -28968
rect 33536 -29002 33552 -28968
rect 32972 -29106 33018 -29059
rect 33698 -29106 33732 -29044
rect 31678 -29140 31774 -29106
rect 32042 -29140 32214 -29106
rect 32482 -29140 32654 -29106
rect 32922 -29140 33068 -29106
rect 33636 -29140 33732 -29106
rect 34304 -28398 34352 -28302
rect 34058 -28474 34074 -28440
rect 34142 -28474 34158 -28440
rect 34012 -28533 34046 -28517
rect 34012 -28925 34046 -28909
rect 34170 -28533 34204 -28517
rect 34170 -28925 34204 -28909
rect 34058 -29002 34074 -28968
rect 34142 -29002 34158 -28968
rect 33878 -29106 33912 -29044
rect 34338 -29044 34352 -28398
rect 34498 -28474 34514 -28440
rect 34582 -28474 34598 -28440
rect 34452 -28533 34486 -28517
rect 34452 -28925 34486 -28909
rect 34610 -28533 34644 -28517
rect 34610 -28925 34644 -28909
rect 34498 -29002 34514 -28968
rect 34582 -29002 34598 -28968
rect 34304 -29106 34352 -29044
rect 34744 -29106 34792 -28302
rect 34938 -28474 34954 -28440
rect 35022 -28474 35038 -28440
rect 34892 -28533 34926 -28517
rect 34892 -28925 34926 -28909
rect 35050 -28533 35084 -28517
rect 35184 -28602 35218 -28302
rect 36078 -28398 36112 -28302
rect 35050 -28925 35084 -28909
rect 35172 -28636 35268 -28602
rect 35836 -28636 35932 -28602
rect 35172 -28683 35218 -28636
rect 34938 -29002 34954 -28968
rect 35022 -29002 35038 -28968
rect 35206 -29059 35218 -28683
rect 35898 -28698 35932 -28636
rect 35352 -28774 35368 -28740
rect 35736 -28774 35752 -28740
rect 35306 -28833 35340 -28817
rect 35306 -28925 35340 -28909
rect 35764 -28833 35798 -28817
rect 35764 -28925 35798 -28909
rect 35352 -29002 35368 -28968
rect 35736 -29002 35752 -28968
rect 35172 -29106 35218 -29059
rect 35898 -29106 35932 -29044
rect 33878 -29140 33974 -29106
rect 34242 -29140 34414 -29106
rect 34682 -29140 34854 -29106
rect 35122 -29140 35268 -29106
rect 35836 -29140 35932 -29106
rect 36504 -28398 36552 -28302
rect 36258 -28474 36274 -28440
rect 36342 -28474 36358 -28440
rect 36212 -28533 36246 -28517
rect 36212 -28925 36246 -28909
rect 36370 -28533 36404 -28517
rect 36370 -28925 36404 -28909
rect 36258 -29002 36274 -28968
rect 36342 -29002 36358 -28968
rect 36078 -29106 36112 -29044
rect 36538 -29044 36552 -28398
rect 36698 -28474 36714 -28440
rect 36782 -28474 36798 -28440
rect 36652 -28533 36686 -28517
rect 36652 -28925 36686 -28909
rect 36810 -28533 36844 -28517
rect 36810 -28925 36844 -28909
rect 36698 -29002 36714 -28968
rect 36782 -29002 36798 -28968
rect 36504 -29106 36552 -29044
rect 36944 -29106 36992 -28302
rect 37138 -28474 37154 -28440
rect 37222 -28474 37238 -28440
rect 37092 -28533 37126 -28517
rect 37092 -28925 37126 -28909
rect 37250 -28533 37284 -28517
rect 37384 -28602 37418 -28302
rect 37250 -28925 37284 -28909
rect 37372 -28636 37468 -28602
rect 38036 -28636 38132 -28602
rect 37372 -28683 37418 -28636
rect 37138 -29002 37154 -28968
rect 37222 -29002 37238 -28968
rect 37406 -29059 37418 -28683
rect 38098 -28698 38132 -28636
rect 37552 -28774 37568 -28740
rect 37936 -28774 37952 -28740
rect 37506 -28833 37540 -28817
rect 37506 -28925 37540 -28909
rect 37964 -28833 37998 -28817
rect 37964 -28925 37998 -28909
rect 37552 -29002 37568 -28968
rect 37936 -29002 37952 -28968
rect 37372 -29106 37418 -29059
rect 38098 -29106 38132 -29044
rect 36078 -29140 36174 -29106
rect 36442 -29140 36614 -29106
rect 36882 -29140 37054 -29106
rect 37322 -29140 37468 -29106
rect 38036 -29140 38132 -29106
rect 28912 -29428 29820 -29366
rect 27430 -29462 27884 -29428
rect 28850 -29462 29820 -29428
rect 27430 -29568 29820 -29462
rect 27430 -29602 27884 -29568
rect 28850 -29602 29820 -29568
rect 27430 -29664 27822 -29602
rect 27430 -30406 27788 -29664
rect 28912 -29664 29820 -29602
rect 27932 -29736 27948 -29702
rect 28724 -29736 28740 -29702
rect 28774 -29764 28808 -29748
rect 28774 -29848 28808 -29832
rect 27932 -29894 27948 -29860
rect 28724 -29894 28740 -29860
rect 28774 -29922 28808 -29906
rect 28774 -30006 28808 -29990
rect 27932 -30052 27948 -30018
rect 28724 -30052 28740 -30018
rect 28774 -30080 28808 -30064
rect 28774 -30164 28808 -30148
rect 27932 -30210 27948 -30176
rect 28724 -30210 28740 -30176
rect 28774 -30238 28808 -30222
rect 28774 -30322 28808 -30306
rect 27932 -30368 27948 -30334
rect 28724 -30368 28740 -30334
rect 27430 -30468 27822 -30406
rect 28946 -30406 29820 -29664
rect 28912 -30468 29820 -30406
rect 27430 -30502 27884 -30468
rect 28850 -30502 29820 -30468
rect 27430 -30608 29820 -30502
rect 27430 -30642 27884 -30608
rect 28850 -30642 29820 -30608
rect 27430 -30704 27822 -30642
rect 27430 -31446 27788 -30704
rect 28912 -30704 29820 -30642
rect 27932 -30776 27948 -30742
rect 28724 -30776 28740 -30742
rect 28774 -30804 28808 -30788
rect 28774 -30888 28808 -30872
rect 27932 -30934 27948 -30900
rect 28724 -30934 28740 -30900
rect 28774 -30962 28808 -30946
rect 28774 -31046 28808 -31030
rect 27932 -31092 27948 -31058
rect 28724 -31092 28740 -31058
rect 28774 -31120 28808 -31104
rect 28774 -31204 28808 -31188
rect 27932 -31250 27948 -31216
rect 28724 -31250 28740 -31216
rect 28774 -31278 28808 -31262
rect 28774 -31362 28808 -31346
rect 27932 -31408 27948 -31374
rect 28724 -31408 28740 -31374
rect 27430 -31508 27822 -31446
rect 28946 -31446 29820 -30704
rect 30840 -29331 38300 -29300
rect 30840 -29365 31775 -29331
rect 32043 -29365 32215 -29331
rect 32483 -29365 32655 -29331
rect 32923 -29365 33094 -29331
rect 33678 -29365 33975 -29331
rect 34243 -29365 34415 -29331
rect 34683 -29365 34855 -29331
rect 35123 -29365 35294 -29331
rect 35878 -29365 36175 -29331
rect 36443 -29365 36615 -29331
rect 36883 -29365 37055 -29331
rect 37323 -29365 37494 -29331
rect 38078 -29365 38300 -29331
rect 30840 -29427 31713 -29365
rect 30840 -29855 31679 -29427
rect 32105 -29420 32153 -29365
rect 32105 -29427 32119 -29420
rect 31859 -29503 31875 -29469
rect 31943 -29503 31959 -29469
rect 31813 -29553 31847 -29537
rect 31813 -29745 31847 -29729
rect 31971 -29553 32005 -29537
rect 31971 -29745 32005 -29729
rect 31859 -29813 31875 -29779
rect 31943 -29813 31959 -29779
rect 30840 -29951 31713 -29855
rect 32299 -29503 32315 -29469
rect 32383 -29503 32399 -29469
rect 32253 -29553 32287 -29537
rect 32253 -29745 32287 -29729
rect 32411 -29553 32445 -29537
rect 32411 -29745 32445 -29729
rect 32299 -29813 32315 -29779
rect 32383 -29813 32399 -29779
rect 32105 -29862 32119 -29855
rect 32105 -29917 32153 -29862
rect 32545 -29917 32593 -29365
rect 32985 -29420 33032 -29365
rect 32739 -29503 32755 -29469
rect 32823 -29503 32839 -29469
rect 32693 -29553 32727 -29537
rect 32693 -29745 32727 -29729
rect 32851 -29553 32885 -29537
rect 32851 -29745 32885 -29729
rect 32739 -29813 32755 -29779
rect 32823 -29813 32839 -29779
rect 32985 -29862 32998 -29420
rect 33740 -29427 33913 -29365
rect 33178 -29503 33194 -29469
rect 33262 -29503 33278 -29469
rect 33336 -29503 33352 -29469
rect 33420 -29503 33436 -29469
rect 33494 -29503 33510 -29469
rect 33578 -29503 33594 -29469
rect 33132 -29553 33166 -29537
rect 33132 -29745 33166 -29729
rect 33290 -29553 33324 -29537
rect 33290 -29745 33324 -29729
rect 33448 -29553 33482 -29537
rect 33448 -29745 33482 -29729
rect 33606 -29553 33640 -29537
rect 33606 -29745 33640 -29729
rect 33178 -29813 33194 -29779
rect 33262 -29813 33278 -29779
rect 33336 -29813 33352 -29779
rect 33420 -29813 33436 -29779
rect 33494 -29813 33510 -29779
rect 33578 -29813 33594 -29779
rect 32985 -29917 33032 -29862
rect 33774 -29855 33879 -29427
rect 34305 -29420 34353 -29365
rect 34305 -29427 34319 -29420
rect 34059 -29503 34075 -29469
rect 34143 -29503 34159 -29469
rect 34013 -29553 34047 -29537
rect 34013 -29745 34047 -29729
rect 34171 -29553 34205 -29537
rect 34171 -29745 34205 -29729
rect 34059 -29813 34075 -29779
rect 34143 -29813 34159 -29779
rect 33740 -29917 33913 -29855
rect 34499 -29503 34515 -29469
rect 34583 -29503 34599 -29469
rect 34453 -29553 34487 -29537
rect 34453 -29745 34487 -29729
rect 34611 -29553 34645 -29537
rect 34611 -29745 34645 -29729
rect 34499 -29813 34515 -29779
rect 34583 -29813 34599 -29779
rect 34305 -29862 34319 -29855
rect 34305 -29917 34353 -29862
rect 34745 -29917 34793 -29365
rect 35185 -29420 35232 -29365
rect 34939 -29503 34955 -29469
rect 35023 -29503 35039 -29469
rect 34893 -29553 34927 -29537
rect 34893 -29745 34927 -29729
rect 35051 -29553 35085 -29537
rect 35051 -29745 35085 -29729
rect 34939 -29813 34955 -29779
rect 35023 -29813 35039 -29779
rect 35185 -29862 35198 -29420
rect 35940 -29427 36113 -29365
rect 35378 -29503 35394 -29469
rect 35462 -29503 35478 -29469
rect 35536 -29503 35552 -29469
rect 35620 -29503 35636 -29469
rect 35694 -29503 35710 -29469
rect 35778 -29503 35794 -29469
rect 35332 -29553 35366 -29537
rect 35332 -29745 35366 -29729
rect 35490 -29553 35524 -29537
rect 35490 -29745 35524 -29729
rect 35648 -29553 35682 -29537
rect 35648 -29745 35682 -29729
rect 35806 -29553 35840 -29537
rect 35806 -29745 35840 -29729
rect 35378 -29813 35394 -29779
rect 35462 -29813 35478 -29779
rect 35536 -29813 35552 -29779
rect 35620 -29813 35636 -29779
rect 35694 -29813 35710 -29779
rect 35778 -29813 35794 -29779
rect 35185 -29917 35232 -29862
rect 35974 -29855 36079 -29427
rect 36505 -29420 36553 -29365
rect 36505 -29427 36519 -29420
rect 36259 -29503 36275 -29469
rect 36343 -29503 36359 -29469
rect 36213 -29553 36247 -29537
rect 36213 -29745 36247 -29729
rect 36371 -29553 36405 -29537
rect 36371 -29745 36405 -29729
rect 36259 -29813 36275 -29779
rect 36343 -29813 36359 -29779
rect 35940 -29917 36113 -29855
rect 36699 -29503 36715 -29469
rect 36783 -29503 36799 -29469
rect 36653 -29553 36687 -29537
rect 36653 -29745 36687 -29729
rect 36811 -29553 36845 -29537
rect 36811 -29745 36845 -29729
rect 36699 -29813 36715 -29779
rect 36783 -29813 36799 -29779
rect 36505 -29862 36519 -29855
rect 36505 -29917 36553 -29862
rect 36945 -29917 36993 -29365
rect 37385 -29420 37432 -29365
rect 37139 -29503 37155 -29469
rect 37223 -29503 37239 -29469
rect 37093 -29553 37127 -29537
rect 37093 -29745 37127 -29729
rect 37251 -29553 37285 -29537
rect 37251 -29745 37285 -29729
rect 37139 -29813 37155 -29779
rect 37223 -29813 37239 -29779
rect 37385 -29862 37398 -29420
rect 38140 -29427 38300 -29365
rect 37578 -29503 37594 -29469
rect 37662 -29503 37678 -29469
rect 37736 -29503 37752 -29469
rect 37820 -29503 37836 -29469
rect 37894 -29503 37910 -29469
rect 37978 -29503 37994 -29469
rect 37532 -29553 37566 -29537
rect 37532 -29745 37566 -29729
rect 37690 -29553 37724 -29537
rect 37690 -29745 37724 -29729
rect 37848 -29553 37882 -29537
rect 37848 -29745 37882 -29729
rect 38006 -29553 38040 -29537
rect 38006 -29745 38040 -29729
rect 37578 -29813 37594 -29779
rect 37662 -29813 37678 -29779
rect 37736 -29813 37752 -29779
rect 37820 -29813 37836 -29779
rect 37894 -29813 37910 -29779
rect 37978 -29813 37994 -29779
rect 37385 -29917 37432 -29862
rect 38174 -29855 38300 -29427
rect 38140 -29917 38300 -29855
rect 32105 -29951 32192 -29917
rect 32506 -29951 32593 -29917
rect 32985 -29951 33094 -29917
rect 33678 -29951 33913 -29917
rect 34305 -29951 34392 -29917
rect 34706 -29951 34793 -29917
rect 35185 -29951 35294 -29917
rect 35878 -29951 36113 -29917
rect 36505 -29951 36592 -29917
rect 36906 -29951 36993 -29917
rect 37385 -29951 37494 -29917
rect 38078 -29951 38300 -29917
rect 30840 -30073 38300 -29951
rect 30840 -30107 31744 -30073
rect 32328 -30107 32437 -30073
rect 32829 -30107 32916 -30073
rect 33230 -30107 33317 -30073
rect 33709 -30107 33944 -30073
rect 34528 -30107 34637 -30073
rect 35029 -30107 35116 -30073
rect 35430 -30107 35517 -30073
rect 35909 -30107 36144 -30073
rect 36728 -30107 36837 -30073
rect 37229 -30107 37316 -30073
rect 37630 -30107 37717 -30073
rect 30840 -30169 31682 -30107
rect 30840 -30597 31648 -30169
rect 32390 -30162 32437 -30107
rect 31828 -30245 31844 -30211
rect 31912 -30245 31928 -30211
rect 31986 -30245 32002 -30211
rect 32070 -30245 32086 -30211
rect 32144 -30245 32160 -30211
rect 32228 -30245 32244 -30211
rect 31782 -30295 31816 -30279
rect 31782 -30487 31816 -30471
rect 31940 -30295 31974 -30279
rect 31940 -30487 31974 -30471
rect 32098 -30295 32132 -30279
rect 32098 -30487 32132 -30471
rect 32256 -30295 32290 -30279
rect 32256 -30487 32290 -30471
rect 31828 -30555 31844 -30521
rect 31912 -30555 31928 -30521
rect 31986 -30555 32002 -30521
rect 32070 -30555 32086 -30521
rect 32144 -30555 32160 -30521
rect 32228 -30555 32244 -30521
rect 30840 -30659 31682 -30597
rect 32424 -30604 32437 -30162
rect 32583 -30245 32599 -30211
rect 32667 -30245 32683 -30211
rect 32537 -30295 32571 -30279
rect 32537 -30487 32571 -30471
rect 32695 -30295 32729 -30279
rect 32695 -30487 32729 -30471
rect 32583 -30555 32599 -30521
rect 32667 -30555 32683 -30521
rect 32390 -30659 32437 -30604
rect 32829 -30659 32877 -30107
rect 33269 -30162 33317 -30107
rect 33303 -30169 33317 -30162
rect 33023 -30245 33039 -30211
rect 33107 -30245 33123 -30211
rect 32977 -30295 33011 -30279
rect 32977 -30487 33011 -30471
rect 33135 -30295 33169 -30279
rect 33135 -30487 33169 -30471
rect 33023 -30555 33039 -30521
rect 33107 -30555 33123 -30521
rect 33709 -30169 33882 -30107
rect 33463 -30245 33479 -30211
rect 33547 -30245 33563 -30211
rect 33417 -30295 33451 -30279
rect 33417 -30487 33451 -30471
rect 33575 -30295 33609 -30279
rect 33575 -30487 33609 -30471
rect 33463 -30555 33479 -30521
rect 33547 -30555 33563 -30521
rect 33303 -30604 33317 -30597
rect 33269 -30659 33317 -30604
rect 33743 -30597 33848 -30169
rect 34590 -30162 34637 -30107
rect 34028 -30245 34044 -30211
rect 34112 -30245 34128 -30211
rect 34186 -30245 34202 -30211
rect 34270 -30245 34286 -30211
rect 34344 -30245 34360 -30211
rect 34428 -30245 34444 -30211
rect 33982 -30295 34016 -30279
rect 33982 -30487 34016 -30471
rect 34140 -30295 34174 -30279
rect 34140 -30487 34174 -30471
rect 34298 -30295 34332 -30279
rect 34298 -30487 34332 -30471
rect 34456 -30295 34490 -30279
rect 34456 -30487 34490 -30471
rect 34028 -30555 34044 -30521
rect 34112 -30555 34128 -30521
rect 34186 -30555 34202 -30521
rect 34270 -30555 34286 -30521
rect 34344 -30555 34360 -30521
rect 34428 -30555 34444 -30521
rect 33709 -30659 33882 -30597
rect 34624 -30604 34637 -30162
rect 34783 -30245 34799 -30211
rect 34867 -30245 34883 -30211
rect 34737 -30295 34771 -30279
rect 34737 -30487 34771 -30471
rect 34895 -30295 34929 -30279
rect 34895 -30487 34929 -30471
rect 34783 -30555 34799 -30521
rect 34867 -30555 34883 -30521
rect 34590 -30659 34637 -30604
rect 35029 -30659 35077 -30107
rect 35469 -30162 35517 -30107
rect 35503 -30169 35517 -30162
rect 35223 -30245 35239 -30211
rect 35307 -30245 35323 -30211
rect 35177 -30295 35211 -30279
rect 35177 -30487 35211 -30471
rect 35335 -30295 35369 -30279
rect 35335 -30487 35369 -30471
rect 35223 -30555 35239 -30521
rect 35307 -30555 35323 -30521
rect 35909 -30169 36082 -30107
rect 35663 -30245 35679 -30211
rect 35747 -30245 35763 -30211
rect 35617 -30295 35651 -30279
rect 35617 -30487 35651 -30471
rect 35775 -30295 35809 -30279
rect 35775 -30487 35809 -30471
rect 35663 -30555 35679 -30521
rect 35747 -30555 35763 -30521
rect 35503 -30604 35517 -30597
rect 35469 -30659 35517 -30604
rect 35943 -30597 36048 -30169
rect 36790 -30162 36837 -30107
rect 36228 -30245 36244 -30211
rect 36312 -30245 36328 -30211
rect 36386 -30245 36402 -30211
rect 36470 -30245 36486 -30211
rect 36544 -30245 36560 -30211
rect 36628 -30245 36644 -30211
rect 36182 -30295 36216 -30279
rect 36182 -30487 36216 -30471
rect 36340 -30295 36374 -30279
rect 36340 -30487 36374 -30471
rect 36498 -30295 36532 -30279
rect 36498 -30487 36532 -30471
rect 36656 -30295 36690 -30279
rect 36656 -30487 36690 -30471
rect 36228 -30555 36244 -30521
rect 36312 -30555 36328 -30521
rect 36386 -30555 36402 -30521
rect 36470 -30555 36486 -30521
rect 36544 -30555 36560 -30521
rect 36628 -30555 36644 -30521
rect 35909 -30659 36082 -30597
rect 36824 -30604 36837 -30162
rect 36983 -30245 36999 -30211
rect 37067 -30245 37083 -30211
rect 36937 -30295 36971 -30279
rect 36937 -30487 36971 -30471
rect 37095 -30295 37129 -30279
rect 37095 -30487 37129 -30471
rect 36983 -30555 36999 -30521
rect 37067 -30555 37083 -30521
rect 36790 -30659 36837 -30604
rect 37229 -30659 37277 -30107
rect 37669 -30162 37717 -30107
rect 37703 -30169 37717 -30162
rect 37423 -30245 37439 -30211
rect 37507 -30245 37523 -30211
rect 37377 -30295 37411 -30279
rect 37377 -30487 37411 -30471
rect 37535 -30295 37569 -30279
rect 37535 -30487 37569 -30471
rect 37423 -30555 37439 -30521
rect 37507 -30555 37523 -30521
rect 38109 -30169 38300 -30073
rect 37863 -30245 37879 -30211
rect 37947 -30245 37963 -30211
rect 37817 -30295 37851 -30279
rect 37817 -30487 37851 -30471
rect 37975 -30295 38009 -30279
rect 37975 -30487 38009 -30471
rect 37863 -30555 37879 -30521
rect 37947 -30555 37963 -30521
rect 37703 -30604 37717 -30597
rect 37669 -30659 37717 -30604
rect 38143 -30597 38300 -30169
rect 38109 -30659 38300 -30597
rect 30840 -30693 31744 -30659
rect 32328 -30693 32499 -30659
rect 32767 -30693 32939 -30659
rect 33207 -30693 33379 -30659
rect 33647 -30693 33944 -30659
rect 34528 -30693 34699 -30659
rect 34967 -30693 35139 -30659
rect 35407 -30693 35579 -30659
rect 35847 -30693 36144 -30659
rect 36728 -30693 36899 -30659
rect 37167 -30693 37339 -30659
rect 37607 -30693 37779 -30659
rect 38047 -30693 38300 -30659
rect 30840 -30740 38300 -30693
rect 31690 -30918 31786 -30884
rect 32354 -30918 32500 -30884
rect 32768 -30918 32940 -30884
rect 33208 -30918 33380 -30884
rect 33648 -30918 33744 -30884
rect 31690 -30980 31724 -30918
rect 32404 -30965 32450 -30918
rect 31870 -31056 31886 -31022
rect 32254 -31056 32270 -31022
rect 31824 -31115 31858 -31099
rect 31824 -31207 31858 -31191
rect 32282 -31115 32316 -31099
rect 32282 -31207 32316 -31191
rect 31870 -31284 31886 -31250
rect 32254 -31284 32270 -31250
rect 31690 -31388 31724 -31326
rect 32404 -31341 32416 -30965
rect 32584 -31056 32600 -31022
rect 32668 -31056 32684 -31022
rect 32404 -31388 32450 -31341
rect 31690 -31422 31786 -31388
rect 32354 -31422 32450 -31388
rect 32538 -31115 32572 -31099
rect 28912 -31508 29820 -31446
rect 27430 -31542 27884 -31508
rect 28850 -31542 29820 -31508
rect 27430 -31660 29820 -31542
rect 27430 -32060 27700 -31660
rect 32404 -31722 32438 -31422
rect 32538 -31507 32572 -31491
rect 32696 -31115 32730 -31099
rect 32696 -31507 32730 -31491
rect 32584 -31584 32600 -31550
rect 32668 -31584 32684 -31550
rect 32830 -31722 32878 -30918
rect 33270 -30980 33318 -30918
rect 33024 -31056 33040 -31022
rect 33108 -31056 33124 -31022
rect 32978 -31115 33012 -31099
rect 32978 -31507 33012 -31491
rect 33136 -31115 33170 -31099
rect 33136 -31507 33170 -31491
rect 33024 -31584 33040 -31550
rect 33108 -31584 33124 -31550
rect 33270 -31626 33284 -30980
rect 33710 -30980 33744 -30918
rect 33464 -31056 33480 -31022
rect 33548 -31056 33564 -31022
rect 33418 -31115 33452 -31099
rect 33418 -31507 33452 -31491
rect 33576 -31115 33610 -31099
rect 33576 -31507 33610 -31491
rect 33464 -31584 33480 -31550
rect 33548 -31584 33564 -31550
rect 33270 -31722 33318 -31626
rect 33890 -30918 33986 -30884
rect 34554 -30918 34700 -30884
rect 34968 -30918 35140 -30884
rect 35408 -30918 35580 -30884
rect 35848 -30918 35944 -30884
rect 33890 -30980 33924 -30918
rect 34604 -30965 34650 -30918
rect 34070 -31056 34086 -31022
rect 34454 -31056 34470 -31022
rect 34024 -31115 34058 -31099
rect 34024 -31207 34058 -31191
rect 34482 -31115 34516 -31099
rect 34482 -31207 34516 -31191
rect 34070 -31284 34086 -31250
rect 34454 -31284 34470 -31250
rect 33890 -31388 33924 -31326
rect 34604 -31341 34616 -30965
rect 34784 -31056 34800 -31022
rect 34868 -31056 34884 -31022
rect 34604 -31388 34650 -31341
rect 33890 -31422 33986 -31388
rect 34554 -31422 34650 -31388
rect 34738 -31115 34772 -31099
rect 33710 -31722 33744 -31626
rect 34604 -31722 34638 -31422
rect 34738 -31507 34772 -31491
rect 34896 -31115 34930 -31099
rect 34896 -31507 34930 -31491
rect 34784 -31584 34800 -31550
rect 34868 -31584 34884 -31550
rect 35030 -31722 35078 -30918
rect 35470 -30980 35518 -30918
rect 35224 -31056 35240 -31022
rect 35308 -31056 35324 -31022
rect 35178 -31115 35212 -31099
rect 35178 -31507 35212 -31491
rect 35336 -31115 35370 -31099
rect 35336 -31507 35370 -31491
rect 35224 -31584 35240 -31550
rect 35308 -31584 35324 -31550
rect 35470 -31626 35484 -30980
rect 35910 -30980 35944 -30918
rect 35664 -31056 35680 -31022
rect 35748 -31056 35764 -31022
rect 35618 -31115 35652 -31099
rect 35618 -31507 35652 -31491
rect 35776 -31115 35810 -31099
rect 35776 -31507 35810 -31491
rect 35664 -31584 35680 -31550
rect 35748 -31584 35764 -31550
rect 35470 -31722 35518 -31626
rect 36090 -30918 36186 -30884
rect 36754 -30918 36900 -30884
rect 37168 -30918 37340 -30884
rect 37608 -30918 37780 -30884
rect 38048 -30918 38144 -30884
rect 36090 -30980 36124 -30918
rect 36804 -30965 36850 -30918
rect 36270 -31056 36286 -31022
rect 36654 -31056 36670 -31022
rect 36224 -31115 36258 -31099
rect 36224 -31207 36258 -31191
rect 36682 -31115 36716 -31099
rect 36682 -31207 36716 -31191
rect 36270 -31284 36286 -31250
rect 36654 -31284 36670 -31250
rect 36090 -31388 36124 -31326
rect 36804 -31341 36816 -30965
rect 36984 -31056 37000 -31022
rect 37068 -31056 37084 -31022
rect 36804 -31388 36850 -31341
rect 36090 -31422 36186 -31388
rect 36754 -31422 36850 -31388
rect 36938 -31115 36972 -31099
rect 35910 -31722 35944 -31626
rect 36804 -31722 36838 -31422
rect 36938 -31507 36972 -31491
rect 37096 -31115 37130 -31099
rect 37096 -31507 37130 -31491
rect 36984 -31584 37000 -31550
rect 37068 -31584 37084 -31550
rect 37230 -31722 37278 -30918
rect 37670 -30980 37718 -30918
rect 37424 -31056 37440 -31022
rect 37508 -31056 37524 -31022
rect 37378 -31115 37412 -31099
rect 37378 -31507 37412 -31491
rect 37536 -31115 37570 -31099
rect 37536 -31507 37570 -31491
rect 37424 -31584 37440 -31550
rect 37508 -31584 37524 -31550
rect 37670 -31626 37684 -30980
rect 38110 -30980 38144 -30918
rect 37864 -31056 37880 -31022
rect 37948 -31056 37964 -31022
rect 37818 -31115 37852 -31099
rect 37818 -31507 37852 -31491
rect 37976 -31115 38010 -31099
rect 37976 -31507 38010 -31491
rect 37864 -31584 37880 -31550
rect 37948 -31584 37964 -31550
rect 37670 -31722 37718 -31626
rect 38110 -31722 38144 -31626
rect 26968 -32064 27064 -32060
<< viali >>
rect 22508 11910 26790 11944
rect -70 10870 -10 10930
rect 2130 10870 2190 10930
rect 2470 10940 4046 10974
rect 2386 10644 2420 10912
rect 4096 10644 4130 10912
rect 2470 10582 4046 10616
rect 4330 10870 4390 10930
rect 4670 10940 6246 10974
rect 4586 10644 4620 10912
rect 6296 10644 6330 10912
rect 4670 10582 6246 10616
rect 6530 10870 6590 10930
rect 6870 10940 8446 10974
rect 6786 10644 6820 10912
rect 8496 10644 8530 10912
rect 6870 10582 8446 10616
rect 8730 10870 8790 10930
rect 9070 10940 10646 10974
rect 8986 10644 9020 10912
rect 10696 10644 10730 10912
rect 9070 10582 10646 10616
rect 10930 10870 10990 10930
rect 11270 10940 12846 10974
rect 11186 10644 11220 10912
rect 12896 10644 12930 10912
rect 11270 10582 12846 10616
rect 13130 10870 13190 10930
rect 13470 10940 15046 10974
rect 13386 10644 13420 10912
rect 15096 10644 15130 10912
rect 13470 10582 15046 10616
rect 15330 10870 15390 10930
rect 15670 10940 17246 10974
rect 15586 10644 15620 10912
rect 17296 10644 17330 10912
rect 15670 10582 17246 10616
rect 17530 10870 17590 10930
rect 17870 10940 19446 10974
rect 17786 10644 17820 10912
rect 19496 10644 19530 10912
rect 17870 10582 19446 10616
rect 19730 10870 19790 10930
rect 21930 10870 21990 10930
rect -70 10070 -10 10130
rect 2130 10070 2190 10130
rect 2470 10140 4046 10174
rect 2386 9844 2420 10112
rect 4096 9844 4130 10112
rect 2470 9782 4046 9816
rect 4330 10070 4390 10130
rect 4670 10140 6246 10174
rect 4586 9844 4620 10112
rect 6296 9844 6330 10112
rect 4670 9782 6246 9816
rect 6530 10070 6590 10130
rect 6870 10140 8446 10174
rect 6786 9844 6820 10112
rect 8496 9844 8530 10112
rect 6870 9782 8446 9816
rect 8730 10070 8790 10130
rect 9070 10140 10646 10174
rect 8986 9844 9020 10112
rect 10696 9844 10730 10112
rect 9070 9782 10646 9816
rect 10930 10070 10990 10130
rect 11270 10140 12846 10174
rect 11186 9844 11220 10112
rect 12896 9844 12930 10112
rect 11270 9782 12846 9816
rect 13130 10070 13190 10130
rect 13470 10140 15046 10174
rect 13386 9844 13420 10112
rect 15096 9844 15130 10112
rect 13470 9782 15046 9816
rect 15330 10070 15390 10130
rect 15670 10140 17246 10174
rect 15586 9844 15620 10112
rect 17296 9844 17330 10112
rect 15670 9782 17246 9816
rect 17530 10070 17590 10130
rect 17870 10140 19446 10174
rect 17786 9844 17820 10112
rect 19496 9844 19530 10112
rect 17870 9782 19446 9816
rect 19730 10070 19790 10130
rect 21930 10070 21990 10130
rect -70 9270 -10 9330
rect 2130 9270 2190 9330
rect 2470 9340 4046 9374
rect 2386 9044 2420 9312
rect 4096 9044 4130 9312
rect 2470 8982 4046 9016
rect 4330 9270 4390 9330
rect 4670 9340 6246 9374
rect 4586 9044 4620 9312
rect 6296 9044 6330 9312
rect 4670 8982 6246 9016
rect 6530 9270 6590 9330
rect 6870 9340 8446 9374
rect 6786 9044 6820 9312
rect 8496 9044 8530 9312
rect 6870 8982 8446 9016
rect 8730 9270 8790 9330
rect 9070 9340 10646 9374
rect 8986 9044 9020 9312
rect 10696 9044 10730 9312
rect 9070 8982 10646 9016
rect 10930 9270 10990 9330
rect 11270 9340 12846 9374
rect 11186 9044 11220 9312
rect 12896 9044 12930 9312
rect 11270 8982 12846 9016
rect 13130 9270 13190 9330
rect 13470 9340 15046 9374
rect 13386 9044 13420 9312
rect 15096 9044 15130 9312
rect 13470 8982 15046 9016
rect 15330 9270 15390 9330
rect 15670 9340 17246 9374
rect 15586 9044 15620 9312
rect 17296 9044 17330 9312
rect 15670 8982 17246 9016
rect 17530 9270 17590 9330
rect 17870 9340 19446 9374
rect 17786 9044 17820 9312
rect 19496 9044 19530 9312
rect 17870 8982 19446 9016
rect 19730 9270 19790 9330
rect 21930 9270 21990 9330
rect -70 8470 -10 8530
rect 2130 8470 2190 8530
rect 2470 8540 4046 8574
rect 2386 8244 2420 8512
rect 4096 8244 4130 8512
rect 2470 8182 4046 8216
rect 4330 8470 4390 8530
rect 4670 8540 6246 8574
rect 4586 8244 4620 8512
rect 6296 8244 6330 8512
rect 4670 8182 6246 8216
rect 6530 8470 6590 8530
rect 6870 8540 8446 8574
rect 6786 8244 6820 8512
rect 8496 8244 8530 8512
rect 6870 8182 8446 8216
rect 8730 8470 8790 8530
rect 9070 8540 10646 8574
rect 8986 8244 9020 8512
rect 10696 8244 10730 8512
rect 9070 8182 10646 8216
rect 10930 8470 10990 8530
rect 11270 8540 12846 8574
rect 11186 8244 11220 8512
rect 12896 8244 12930 8512
rect 11270 8182 12846 8216
rect 13130 8470 13190 8530
rect 13470 8540 15046 8574
rect 13386 8244 13420 8512
rect 15096 8244 15130 8512
rect 13470 8182 15046 8216
rect 15330 8470 15390 8530
rect 15670 8540 17246 8574
rect 15586 8244 15620 8512
rect 17296 8244 17330 8512
rect 15670 8182 17246 8216
rect 17530 8470 17590 8530
rect 17870 8540 19446 8574
rect 17786 8244 17820 8512
rect 19496 8244 19530 8512
rect 17870 8182 19446 8216
rect 19730 8470 19790 8530
rect 21930 8470 21990 8530
rect -70 7670 -10 7730
rect 2130 7670 2190 7730
rect 2470 7740 4046 7774
rect 2386 7444 2420 7712
rect 4096 7444 4130 7712
rect 2470 7382 4046 7416
rect 4330 7670 4390 7730
rect 4670 7740 6246 7774
rect 4586 7444 4620 7712
rect 6296 7444 6330 7712
rect 4670 7382 6246 7416
rect 6530 7670 6590 7730
rect 6870 7740 8446 7774
rect 6786 7444 6820 7712
rect 8496 7444 8530 7712
rect 6870 7382 8446 7416
rect 8730 7670 8790 7730
rect 9070 7740 10646 7774
rect 8986 7444 9020 7712
rect 10696 7444 10730 7712
rect 9070 7382 10646 7416
rect 10930 7670 10990 7730
rect 11270 7740 12846 7774
rect 11186 7444 11220 7712
rect 12896 7444 12930 7712
rect 11270 7382 12846 7416
rect 13130 7670 13190 7730
rect 13470 7740 15046 7774
rect 13386 7444 13420 7712
rect 15096 7444 15130 7712
rect 13470 7382 15046 7416
rect 15330 7670 15390 7730
rect 15670 7740 17246 7774
rect 15586 7444 15620 7712
rect 17296 7444 17330 7712
rect 15670 7382 17246 7416
rect 17530 7670 17590 7730
rect 17870 7740 19446 7774
rect 17786 7444 17820 7712
rect 19496 7444 19530 7712
rect 17870 7382 19446 7416
rect 19730 7670 19790 7730
rect 21930 7670 21990 7730
rect -70 6870 -10 6930
rect 2130 6870 2190 6930
rect 2470 6940 4046 6974
rect 2386 6644 2420 6912
rect 4096 6644 4130 6912
rect 2470 6582 4046 6616
rect 4330 6870 4390 6930
rect 4670 6940 6246 6974
rect 4586 6644 4620 6912
rect 6296 6644 6330 6912
rect 4670 6582 6246 6616
rect 6530 6870 6590 6930
rect 6870 6940 8446 6974
rect 6786 6644 6820 6912
rect 8496 6644 8530 6912
rect 6870 6582 8446 6616
rect 8730 6870 8790 6930
rect 9070 6940 10646 6974
rect 8986 6644 9020 6912
rect 10696 6644 10730 6912
rect 9070 6582 10646 6616
rect 10930 6870 10990 6930
rect 11270 6940 12846 6974
rect 11186 6644 11220 6912
rect 12896 6644 12930 6912
rect 11270 6582 12846 6616
rect 13130 6870 13190 6930
rect 13470 6940 15046 6974
rect 13386 6644 13420 6912
rect 15096 6644 15130 6912
rect 13470 6582 15046 6616
rect 15330 6870 15390 6930
rect 15670 6940 17246 6974
rect 15586 6644 15620 6912
rect 17296 6644 17330 6912
rect 15670 6582 17246 6616
rect 17530 6870 17590 6930
rect 17870 6940 19446 6974
rect 17786 6644 17820 6912
rect 19496 6644 19530 6912
rect 17870 6582 19446 6616
rect 19730 6870 19790 6930
rect 21930 6870 21990 6930
rect -70 6070 -10 6130
rect 2130 6070 2190 6130
rect 2470 6140 4046 6174
rect 2386 5844 2420 6112
rect 4096 5844 4130 6112
rect 2470 5782 4046 5816
rect 4330 6070 4390 6130
rect 4670 6140 6246 6174
rect 4586 5844 4620 6112
rect 6296 5844 6330 6112
rect 4670 5782 6246 5816
rect 6530 6070 6590 6130
rect 6870 6140 8446 6174
rect 6786 5844 6820 6112
rect 8496 5844 8530 6112
rect 6870 5782 8446 5816
rect 8730 6070 8790 6130
rect 9070 6140 10646 6174
rect 8986 5844 9020 6112
rect 10696 5844 10730 6112
rect 9070 5782 10646 5816
rect 10930 6070 10990 6130
rect 11270 6140 12846 6174
rect 11186 5844 11220 6112
rect 12896 5844 12930 6112
rect 11270 5782 12846 5816
rect 13130 6070 13190 6130
rect 13470 6140 15046 6174
rect 13386 5844 13420 6112
rect 15096 5844 15130 6112
rect 13470 5782 15046 5816
rect 15330 6070 15390 6130
rect 15670 6140 17246 6174
rect 15586 5844 15620 6112
rect 17296 5844 17330 6112
rect 15670 5782 17246 5816
rect 17530 6070 17590 6130
rect 17870 6140 19446 6174
rect 17786 5844 17820 6112
rect 19496 5844 19530 6112
rect 17870 5782 19446 5816
rect 19730 6070 19790 6130
rect 21930 6070 21990 6130
rect -70 5270 -10 5330
rect 2130 5270 2190 5330
rect 2470 5340 4046 5374
rect 2386 5044 2420 5312
rect 4096 5044 4130 5312
rect 2470 4982 4046 5016
rect 4330 5270 4390 5330
rect 4670 5340 6246 5374
rect 4586 5044 4620 5312
rect 6296 5044 6330 5312
rect 4670 4982 6246 5016
rect 6530 5270 6590 5330
rect 6870 5340 8446 5374
rect 6786 5044 6820 5312
rect 8496 5044 8530 5312
rect 6870 4982 8446 5016
rect 8730 5270 8790 5330
rect 9070 5340 10646 5374
rect 8986 5044 9020 5312
rect 10696 5044 10730 5312
rect 9070 4982 10646 5016
rect 10930 5270 10990 5330
rect 11270 5340 12846 5374
rect 11186 5044 11220 5312
rect 12896 5044 12930 5312
rect 11270 4982 12846 5016
rect 13130 5270 13190 5330
rect 13470 5340 15046 5374
rect 13386 5044 13420 5312
rect 15096 5044 15130 5312
rect 13470 4982 15046 5016
rect 15330 5270 15390 5330
rect 15670 5340 17246 5374
rect 15586 5044 15620 5312
rect 17296 5044 17330 5312
rect 15670 4982 17246 5016
rect 17530 5270 17590 5330
rect 17870 5340 19446 5374
rect 17786 5044 17820 5312
rect 19496 5044 19530 5312
rect 17870 4982 19446 5016
rect 19730 5270 19790 5330
rect 21930 5270 21990 5330
rect 22236 4842 22270 11538
rect 22382 11399 22920 11796
rect 23048 11399 23586 11796
rect 23714 11399 24252 11796
rect 24380 11399 24918 11796
rect 25046 11399 25584 11796
rect 25712 11399 26250 11796
rect 26378 11399 26916 11796
rect 9072 4542 10648 4576
rect 8988 4273 9022 4487
rect 10698 4273 10732 4487
rect 9072 4184 10648 4218
rect 11272 4542 12848 4576
rect 11188 4273 11222 4487
rect 12898 4273 12932 4487
rect 11272 4184 12848 4218
rect 22382 4584 22920 4981
rect 23048 4584 23586 4981
rect 23714 4584 24252 4981
rect 24380 4584 24918 4981
rect 25046 4584 25584 4981
rect 25712 4584 26250 4981
rect 26378 4584 26916 4981
rect 27028 4842 27062 11538
rect 30073 11903 30639 11937
rect 30757 11903 30819 11937
rect 30819 11903 31087 11937
rect 31087 11903 31149 11937
rect 31236 11903 31259 11937
rect 31259 11903 31527 11937
rect 31527 11903 31550 11937
rect 31637 11903 31699 11937
rect 31699 11903 31967 11937
rect 31967 11903 32029 11937
rect 27922 11558 28802 11592
rect 27938 11424 28714 11458
rect 28773 11335 28807 11389
rect 27938 11266 28714 11300
rect 28773 11177 28807 11231
rect 27938 11108 28714 11142
rect 28773 11019 28807 11073
rect 27938 10950 28714 10984
rect 28773 10861 28807 10915
rect 27938 10792 28714 10826
rect 30710 11841 30744 11848
rect 30178 11765 30218 11799
rect 30336 11765 30376 11799
rect 30494 11765 30534 11799
rect 30102 11539 30136 11715
rect 30260 11539 30294 11715
rect 30418 11539 30452 11715
rect 30576 11539 30610 11715
rect 30178 11455 30218 11489
rect 30336 11455 30376 11489
rect 30494 11455 30534 11489
rect 30710 11413 30744 11841
rect 30710 11406 30744 11413
rect 30933 11765 30973 11799
rect 30857 11539 30891 11715
rect 31015 11539 31049 11715
rect 30933 11455 30973 11489
rect 31589 11841 31623 11848
rect 31359 11765 31427 11799
rect 31297 11539 31331 11715
rect 31455 11539 31489 11715
rect 31359 11455 31427 11489
rect 31589 11413 31603 11841
rect 31603 11413 31623 11841
rect 31799 11765 31867 11799
rect 31737 11539 31771 11715
rect 31895 11539 31929 11715
rect 31799 11455 31867 11489
rect 31589 11406 31623 11413
rect 32273 11903 32839 11937
rect 32957 11903 33019 11937
rect 33019 11903 33287 11937
rect 33287 11903 33349 11937
rect 33436 11903 33459 11937
rect 33459 11903 33727 11937
rect 33727 11903 33750 11937
rect 33837 11903 33899 11937
rect 33899 11903 34167 11937
rect 34167 11903 34229 11937
rect 32910 11841 32944 11848
rect 32378 11765 32418 11799
rect 32536 11765 32576 11799
rect 32694 11765 32734 11799
rect 32302 11539 32336 11715
rect 32460 11539 32494 11715
rect 32618 11539 32652 11715
rect 32776 11539 32810 11715
rect 32378 11455 32418 11489
rect 32536 11455 32576 11489
rect 32694 11455 32734 11489
rect 32910 11413 32944 11841
rect 32910 11406 32944 11413
rect 33133 11765 33173 11799
rect 33057 11539 33091 11715
rect 33215 11539 33249 11715
rect 33133 11455 33173 11489
rect 33789 11841 33823 11848
rect 33559 11765 33627 11799
rect 33497 11539 33531 11715
rect 33655 11539 33689 11715
rect 33559 11455 33627 11489
rect 33789 11413 33803 11841
rect 33803 11413 33823 11841
rect 33999 11765 34067 11799
rect 33937 11539 33971 11715
rect 34095 11539 34129 11715
rect 33999 11455 34067 11489
rect 33789 11406 33823 11413
rect 34473 11903 35039 11937
rect 35157 11903 35219 11937
rect 35219 11903 35487 11937
rect 35487 11903 35549 11937
rect 35636 11903 35659 11937
rect 35659 11903 35927 11937
rect 35927 11903 35950 11937
rect 36037 11903 36099 11937
rect 36099 11903 36367 11937
rect 36367 11903 36429 11937
rect 35110 11841 35144 11848
rect 34578 11765 34618 11799
rect 34736 11765 34776 11799
rect 34894 11765 34934 11799
rect 34502 11539 34536 11715
rect 34660 11539 34694 11715
rect 34818 11539 34852 11715
rect 34976 11539 35010 11715
rect 34578 11455 34618 11489
rect 34736 11455 34776 11489
rect 34894 11455 34934 11489
rect 35110 11413 35144 11841
rect 35110 11406 35144 11413
rect 35333 11765 35373 11799
rect 35257 11539 35291 11715
rect 35415 11539 35449 11715
rect 35333 11455 35373 11489
rect 35989 11841 36023 11848
rect 35759 11765 35827 11799
rect 35697 11539 35731 11715
rect 35855 11539 35889 11715
rect 35759 11455 35827 11489
rect 35989 11413 36003 11841
rect 36003 11413 36023 11841
rect 36199 11765 36267 11799
rect 36137 11539 36171 11715
rect 36295 11539 36329 11715
rect 36199 11455 36267 11489
rect 35989 11406 36023 11413
rect 27922 10658 28802 10692
rect 30280 10954 30500 10988
rect 30144 10819 30178 10895
rect 30602 10819 30636 10895
rect 30280 10726 30500 10760
rect 30736 11030 30770 11045
rect 30736 10684 30770 11030
rect 30934 10954 30974 10988
rect 30736 10669 30770 10684
rect 30113 10588 30667 10622
rect 27922 10518 28802 10552
rect 27938 10384 28714 10418
rect 28773 10295 28807 10349
rect 27938 10226 28714 10260
rect 28773 10137 28807 10191
rect 27938 10068 28714 10102
rect 28773 9979 28807 10033
rect 27938 9910 28714 9944
rect 28773 9821 28807 9875
rect 27938 9752 28714 9786
rect 30858 10519 30892 10895
rect 31016 10519 31050 10895
rect 30934 10426 30974 10460
rect 30758 10288 30820 10322
rect 30820 10288 31088 10322
rect 31088 10288 31150 10322
rect 31374 10954 31414 10988
rect 31298 10519 31332 10895
rect 31456 10519 31490 10895
rect 31374 10426 31414 10460
rect 31814 10954 31854 10988
rect 31738 10519 31772 10895
rect 31896 10519 31930 10895
rect 31814 10426 31854 10460
rect 31198 10288 31260 10322
rect 31260 10288 31528 10322
rect 31528 10288 31590 10322
rect 32480 10954 32700 10988
rect 32344 10819 32378 10895
rect 32802 10819 32836 10895
rect 32480 10726 32700 10760
rect 32936 11030 32970 11045
rect 32936 10684 32970 11030
rect 33134 10954 33174 10988
rect 32936 10669 32970 10684
rect 32313 10588 32867 10622
rect 31638 10288 31700 10322
rect 31700 10288 31968 10322
rect 31968 10288 32030 10322
rect 33058 10519 33092 10895
rect 33216 10519 33250 10895
rect 33134 10426 33174 10460
rect 32958 10288 33020 10322
rect 33020 10288 33288 10322
rect 33288 10288 33350 10322
rect 33574 10954 33614 10988
rect 33498 10519 33532 10895
rect 33656 10519 33690 10895
rect 33574 10426 33614 10460
rect 34014 10954 34054 10988
rect 33938 10519 33972 10895
rect 34096 10519 34130 10895
rect 34014 10426 34054 10460
rect 33398 10288 33460 10322
rect 33460 10288 33728 10322
rect 33728 10288 33790 10322
rect 34680 10954 34900 10988
rect 34544 10819 34578 10895
rect 35002 10819 35036 10895
rect 34680 10726 34900 10760
rect 35136 11030 35170 11045
rect 35136 10684 35170 11030
rect 35334 10954 35374 10988
rect 35136 10669 35170 10684
rect 34513 10588 35067 10622
rect 33838 10288 33900 10322
rect 33900 10288 34168 10322
rect 34168 10288 34230 10322
rect 35258 10519 35292 10895
rect 35416 10519 35450 10895
rect 35334 10426 35374 10460
rect 35158 10288 35220 10322
rect 35220 10288 35488 10322
rect 35488 10288 35550 10322
rect 35774 10954 35814 10988
rect 35698 10519 35732 10895
rect 35856 10519 35890 10895
rect 35774 10426 35814 10460
rect 36214 10954 36254 10988
rect 36138 10519 36172 10895
rect 36296 10519 36330 10895
rect 36214 10426 36254 10460
rect 35598 10288 35660 10322
rect 35660 10288 35928 10322
rect 35928 10288 35990 10322
rect 36038 10288 36100 10322
rect 36100 10288 36368 10322
rect 36368 10288 36430 10322
rect 29827 9782 31387 9816
rect 27922 9618 28802 9652
rect 29794 9644 30562 9678
rect 30652 9644 31420 9678
rect 27922 9478 28802 9512
rect 27938 9344 28714 9378
rect 28773 9255 28807 9309
rect 27938 9186 28714 9220
rect 28773 9097 28807 9151
rect 27938 9028 28714 9062
rect 28773 8939 28807 8993
rect 27938 8870 28714 8904
rect 28773 8781 28807 8835
rect 27938 8712 28714 8746
rect 29598 9243 29632 9551
rect 29732 9209 29766 9585
rect 30590 9209 30624 9585
rect 31448 9209 31482 9585
rect 31582 9243 31616 9551
rect 29794 9116 30562 9150
rect 30652 9116 31420 9150
rect 29827 8978 31387 9012
rect 32830 9008 32892 9042
rect 32892 9008 33478 9042
rect 33478 9008 33540 9042
rect 29827 8778 31387 8812
rect 29794 8640 30562 8674
rect 30652 8640 31420 8674
rect 27922 8578 28802 8612
rect 27922 8438 28802 8472
rect 27938 8304 28714 8338
rect 28773 8215 28807 8269
rect 27938 8146 28714 8180
rect 28773 8057 28807 8111
rect 27938 7988 28714 8022
rect 28773 7899 28807 7953
rect 27938 7830 28714 7864
rect 28773 7741 28807 7795
rect 27938 7672 28714 7706
rect 27922 7538 28802 7572
rect 29598 7513 29632 8637
rect 29732 8205 29766 8581
rect 30590 8205 30624 8581
rect 31448 8205 31482 8581
rect 29794 8112 30562 8146
rect 30652 8112 31420 8146
rect 29794 8004 30562 8038
rect 30652 8004 31420 8038
rect 29732 7569 29766 7945
rect 30590 7569 30624 7945
rect 31448 7569 31482 7945
rect 31582 7513 31616 8637
rect 33006 8906 33106 8940
rect 33264 8906 33364 8940
rect 32910 8071 32944 8847
rect 33168 8071 33202 8847
rect 33426 8071 33460 8847
rect 33006 7978 33106 8012
rect 33264 7978 33364 8012
rect 33670 9008 33732 9042
rect 33732 9008 34318 9042
rect 34318 9008 34380 9042
rect 33846 8906 33946 8940
rect 34104 8906 34204 8940
rect 33750 8071 33784 8847
rect 34008 8071 34042 8847
rect 34266 8071 34300 8847
rect 33846 7978 33946 8012
rect 34104 7978 34204 8012
rect 34510 8788 34572 8822
rect 34572 8788 34730 8822
rect 34730 8788 34792 8822
rect 34634 8686 34668 8720
rect 34590 8251 34624 8627
rect 34678 8251 34712 8627
rect 34634 8158 34668 8192
rect 34930 8788 34992 8822
rect 34992 8788 35150 8822
rect 35150 8788 35212 8822
rect 35054 8686 35088 8720
rect 35010 8251 35044 8627
rect 35098 8251 35132 8627
rect 35054 8158 35088 8192
rect 35350 8788 35412 8822
rect 35412 8788 35570 8822
rect 35570 8788 35632 8822
rect 35474 8686 35508 8720
rect 35430 8251 35464 8627
rect 35518 8251 35552 8627
rect 35474 8158 35508 8192
rect 29794 7476 30562 7510
rect 30652 7476 31420 7510
rect 27922 7398 28802 7432
rect 27938 7264 28714 7298
rect 28773 7175 28807 7229
rect 27938 7106 28714 7140
rect 28773 7017 28807 7071
rect 27938 6948 28714 6982
rect 28773 6859 28807 6913
rect 27938 6790 28714 6824
rect 28773 6701 28807 6755
rect 27938 6632 28714 6666
rect 29538 7102 29572 7115
rect 29538 6734 29572 7102
rect 29769 7030 30545 7064
rect 29676 6868 29710 6968
rect 30604 6868 30638 6968
rect 29769 6772 30545 6806
rect 29538 6721 29572 6734
rect 31109 7030 31885 7064
rect 31016 6868 31050 6968
rect 31944 6868 31978 6968
rect 31109 6772 31885 6806
rect 33548 7476 33588 7510
rect 33706 7476 33746 7510
rect 33864 7476 33904 7510
rect 34022 7476 34062 7510
rect 33472 7050 33506 7426
rect 33630 7050 33664 7426
rect 33788 7050 33822 7426
rect 33946 7050 33980 7426
rect 34104 7050 34138 7426
rect 33548 6966 33588 7000
rect 33706 6966 33746 7000
rect 33864 6966 33904 7000
rect 34022 6966 34062 7000
rect 34634 7368 34668 7402
rect 34590 7142 34624 7318
rect 34678 7142 34712 7318
rect 34634 7058 34668 7092
rect 34510 6956 34572 6990
rect 34572 6956 34730 6990
rect 34730 6956 34792 6990
rect 35054 7368 35088 7402
rect 35010 7142 35044 7318
rect 35098 7142 35132 7318
rect 35054 7058 35088 7092
rect 34930 6956 34992 6990
rect 34992 6956 35150 6990
rect 35150 6956 35212 6990
rect 35474 7368 35508 7402
rect 35430 7142 35464 7318
rect 35518 7142 35552 7318
rect 35474 7058 35508 7092
rect 35350 6956 35412 6990
rect 35412 6956 35570 6990
rect 35570 6956 35632 6990
rect 33372 6828 33434 6862
rect 33434 6828 34176 6862
rect 34176 6828 34238 6862
rect 27922 6498 28802 6532
rect 27922 6358 28802 6392
rect 27938 6224 28714 6258
rect 28773 6135 28807 6189
rect 27938 6066 28714 6100
rect 28773 5977 28807 6031
rect 27938 5908 28714 5942
rect 28773 5819 28807 5873
rect 27938 5750 28714 5784
rect 28773 5661 28807 5715
rect 27938 5592 28714 5626
rect 27922 5458 28802 5492
rect 22508 4436 26790 4470
rect 27921 5342 28795 5376
rect 27974 5204 28742 5238
rect 27912 4369 27946 5145
rect 28770 4369 28804 5145
rect 27974 4276 28742 4310
rect 28904 4289 28938 5225
rect 29770 6200 30546 6234
rect 29686 6021 29720 6155
rect 30596 6021 30630 6155
rect 29770 5942 30546 5976
rect 31110 6200 31886 6234
rect 31026 6021 31060 6155
rect 31936 6021 31970 6155
rect 31110 5942 31886 5976
rect 29984 5546 30352 5580
rect 29922 5420 29956 5496
rect 30380 5420 30414 5496
rect 29984 5336 30352 5370
rect 31294 5546 31662 5580
rect 31232 5420 31266 5496
rect 31690 5420 31724 5496
rect 31294 5336 31662 5370
rect 29770 4940 30546 4974
rect 29686 4761 29720 4895
rect 30596 4761 30630 4895
rect 29770 4682 30546 4716
rect 31110 4940 31886 4974
rect 31026 4761 31060 4895
rect 31936 4761 31970 4895
rect 31110 4682 31886 4716
rect 27921 4138 28795 4172
rect 32772 4134 33970 4168
rect 34883 4134 35449 4168
rect 32588 3457 32622 4059
rect 32801 3996 32835 4030
rect 32959 3996 32993 4030
rect 33117 3996 33151 4030
rect 33275 3996 33309 4030
rect 33433 3996 33467 4030
rect 33591 3996 33625 4030
rect 33749 3996 33783 4030
rect 33907 3996 33941 4030
rect 32722 3570 32756 3946
rect 32880 3570 32914 3946
rect 33038 3570 33072 3946
rect 33196 3570 33230 3946
rect 33354 3570 33388 3946
rect 33512 3570 33546 3946
rect 33670 3570 33704 3946
rect 33828 3570 33862 3946
rect 33986 3570 34020 3946
rect 32801 3486 32835 3520
rect 32959 3486 32993 3520
rect 33117 3486 33151 3520
rect 33275 3486 33309 3520
rect 33433 3486 33467 3520
rect 33591 3486 33625 3520
rect 33749 3486 33783 3520
rect 33907 3486 33941 3520
rect 17164 3354 17232 3388
rect 17322 3354 17390 3388
rect 17480 3354 17548 3388
rect 17638 3354 17706 3388
rect 17102 2528 17136 3304
rect 17260 2528 17294 3304
rect 17418 2528 17452 3304
rect 17576 2528 17610 3304
rect 17734 2528 17768 3304
rect 34120 3457 34154 4059
rect 34778 3457 34812 4059
rect 34991 3996 35025 4030
rect 35149 3996 35183 4030
rect 35307 3996 35341 4030
rect 34912 3570 34946 3946
rect 35070 3570 35104 3946
rect 35228 3570 35262 3946
rect 35386 3570 35420 3946
rect 34991 3486 35025 3520
rect 35149 3486 35183 3520
rect 35307 3486 35341 3520
rect 35520 3457 35554 4059
rect 36460 5966 36836 6000
rect 36376 5787 36410 5921
rect 36886 5787 36920 5921
rect 36460 5708 36836 5742
rect 36376 5529 36410 5663
rect 36886 5529 36920 5663
rect 36460 5450 36836 5484
rect 36376 5271 36410 5405
rect 36886 5271 36920 5405
rect 36460 5192 36836 5226
rect 36376 5013 36410 5147
rect 36886 5013 36920 5147
rect 36460 4934 36836 4968
rect 36376 4755 36410 4889
rect 36886 4755 36920 4889
rect 36460 4676 36836 4710
rect 36376 4497 36410 4631
rect 36886 4497 36920 4631
rect 36460 4418 36836 4452
rect 36376 4239 36410 4373
rect 36886 4239 36920 4373
rect 36460 4160 36836 4194
rect 36376 3981 36410 4115
rect 36886 3981 36920 4115
rect 36460 3902 36836 3936
rect 37246 5966 37622 6000
rect 37162 5787 37196 5921
rect 37672 5787 37706 5921
rect 37246 5708 37622 5742
rect 37162 5529 37196 5663
rect 37672 5529 37706 5663
rect 37246 5450 37622 5484
rect 37162 5271 37196 5405
rect 37672 5271 37706 5405
rect 37246 5192 37622 5226
rect 37162 5013 37196 5147
rect 37672 5013 37706 5147
rect 37246 4934 37622 4968
rect 37162 4755 37196 4889
rect 37672 4755 37706 4889
rect 37246 4676 37622 4710
rect 37162 4497 37196 4631
rect 37672 4497 37706 4631
rect 37246 4418 37622 4452
rect 37162 4239 37196 4373
rect 37672 4239 37706 4373
rect 37246 4160 37622 4194
rect 37162 3981 37196 4115
rect 37672 3981 37706 4115
rect 37246 3902 37622 3936
rect 32347 3204 32354 3238
rect 32354 3204 32780 3238
rect 32780 3204 32787 3238
rect 33947 3204 33954 3238
rect 33954 3204 34380 3238
rect 34380 3204 34387 3238
rect 35547 3204 35554 3238
rect 35554 3204 35980 3238
rect 35980 3204 35987 3238
rect 32258 2527 32292 3129
rect 32471 3066 32505 3100
rect 32629 3066 32663 3100
rect 32392 2640 32426 3016
rect 32550 2640 32584 3016
rect 32708 2640 32742 3016
rect 32471 2556 32505 2590
rect 32629 2556 32663 2590
rect 32842 2527 32876 3129
rect 33858 2527 33892 3129
rect 34071 3066 34105 3100
rect 34229 3066 34263 3100
rect 33992 2640 34026 3016
rect 34150 2640 34184 3016
rect 34308 2640 34342 3016
rect 34071 2556 34105 2590
rect 34229 2556 34263 2590
rect 34442 2527 34476 3129
rect 35458 2527 35492 3129
rect 35671 3066 35705 3100
rect 35829 3066 35863 3100
rect 35592 2640 35626 3016
rect 35750 2640 35784 3016
rect 35908 2640 35942 3016
rect 35671 2556 35705 2590
rect 35829 2556 35863 2590
rect 36042 2527 36076 3129
rect -117 2195 -55 2229
rect -55 2195 1191 2229
rect 1191 2195 1253 2229
rect 1483 2195 1545 2229
rect 1545 2195 2791 2229
rect 2791 2195 2853 2229
rect 71 2061 447 2095
rect 689 2061 1065 2095
rect -13 1303 21 1995
rect 497 1303 531 1995
rect 605 1303 639 1995
rect 1115 1303 1149 1995
rect 71 1203 447 1237
rect 689 1203 1065 1237
rect 3083 2195 3145 2229
rect 3145 2195 4391 2229
rect 4391 2195 4453 2229
rect 1671 2061 2047 2095
rect 2289 2061 2665 2095
rect 1587 1303 1621 1995
rect 2097 1303 2131 1995
rect 2205 1303 2239 1995
rect 2715 1303 2749 1995
rect 1671 1203 2047 1237
rect 2289 1203 2665 1237
rect 4683 2195 4745 2229
rect 4745 2195 5991 2229
rect 5991 2195 6053 2229
rect 3271 2061 3647 2095
rect 3889 2061 4265 2095
rect 3187 1303 3221 1995
rect 3697 1303 3731 1995
rect 3805 1303 3839 1995
rect 4315 1303 4349 1995
rect 3271 1203 3647 1237
rect 3889 1203 4265 1237
rect 6283 2195 6345 2229
rect 6345 2195 7591 2229
rect 7591 2195 7653 2229
rect 4871 2061 5247 2095
rect 5489 2061 5865 2095
rect 4787 1303 4821 1995
rect 5297 1303 5331 1995
rect 5405 1303 5439 1995
rect 5915 1303 5949 1995
rect 4871 1203 5247 1237
rect 5489 1203 5865 1237
rect 7883 2195 7945 2229
rect 7945 2195 9191 2229
rect 9191 2195 9253 2229
rect 6471 2061 6847 2095
rect 7089 2061 7465 2095
rect 6387 1303 6421 1995
rect 6897 1303 6931 1995
rect 7005 1303 7039 1995
rect 7515 1303 7549 1995
rect 6471 1203 6847 1237
rect 7089 1203 7465 1237
rect 9483 2195 9545 2229
rect 9545 2195 10791 2229
rect 10791 2195 10853 2229
rect 8071 2061 8447 2095
rect 8689 2061 9065 2095
rect 7987 1303 8021 1995
rect 8497 1303 8531 1995
rect 8605 1303 8639 1995
rect 9115 1303 9149 1995
rect 8071 1203 8447 1237
rect 8689 1203 9065 1237
rect 11083 2195 11145 2229
rect 11145 2195 12391 2229
rect 12391 2195 12453 2229
rect 9671 2061 10047 2095
rect 10289 2061 10665 2095
rect 9587 1303 9621 1995
rect 10097 1303 10131 1995
rect 10205 1303 10239 1995
rect 10715 1303 10749 1995
rect 9671 1203 10047 1237
rect 10289 1203 10665 1237
rect 12683 2195 12745 2229
rect 12745 2195 13991 2229
rect 13991 2195 14053 2229
rect 11271 2061 11647 2095
rect 11889 2061 12265 2095
rect 11187 1303 11221 1995
rect 11697 1303 11731 1995
rect 11805 1303 11839 1995
rect 12315 1303 12349 1995
rect 11271 1203 11647 1237
rect 11889 1203 12265 1237
rect 14283 2195 14345 2229
rect 14345 2195 15591 2229
rect 15591 2195 15653 2229
rect 12871 2061 13247 2095
rect 13489 2061 13865 2095
rect 12787 1303 12821 1995
rect 13297 1303 13331 1995
rect 13405 1303 13439 1995
rect 13915 1303 13949 1995
rect 12871 1203 13247 1237
rect 13489 1203 13865 1237
rect 15883 2195 15945 2229
rect 15945 2195 17191 2229
rect 17191 2195 17253 2229
rect 14471 2061 14847 2095
rect 15089 2061 15465 2095
rect 14387 1303 14421 1995
rect 14897 1303 14931 1995
rect 15005 1303 15039 1995
rect 15515 1303 15549 1995
rect 14471 1203 14847 1237
rect 15089 1203 15465 1237
rect 17483 2195 17545 2229
rect 17545 2195 18791 2229
rect 18791 2195 18853 2229
rect 16071 2061 16447 2095
rect 16689 2061 17065 2095
rect 15987 1303 16021 1995
rect 16497 1303 16531 1995
rect 16605 1303 16639 1995
rect 17115 1303 17149 1995
rect 16071 1203 16447 1237
rect 16689 1203 17065 1237
rect 19083 2195 19145 2229
rect 19145 2195 20391 2229
rect 20391 2195 20453 2229
rect 17671 2061 18047 2095
rect 18289 2061 18665 2095
rect 17587 1303 17621 1995
rect 18097 1303 18131 1995
rect 18205 1303 18239 1995
rect 18715 1303 18749 1995
rect 17671 1203 18047 1237
rect 18289 1203 18665 1237
rect 20683 2195 20745 2229
rect 20745 2195 21991 2229
rect 21991 2195 22053 2229
rect 19271 2061 19647 2095
rect 19889 2061 20265 2095
rect 19187 1303 19221 1995
rect 19697 1303 19731 1995
rect 19805 1303 19839 1995
rect 20315 1303 20349 1995
rect 19271 1203 19647 1237
rect 19889 1203 20265 1237
rect 22283 2195 22345 2229
rect 22345 2195 23591 2229
rect 23591 2195 23653 2229
rect 20871 2061 21247 2095
rect 21489 2061 21865 2095
rect 20787 1303 20821 1995
rect 21297 1303 21331 1995
rect 21405 1303 21439 1995
rect 21915 1303 21949 1995
rect 20871 1203 21247 1237
rect 21489 1203 21865 1237
rect 23883 2195 23945 2229
rect 23945 2195 25191 2229
rect 25191 2195 25253 2229
rect 22471 2061 22847 2095
rect 23089 2061 23465 2095
rect 22387 1303 22421 1995
rect 22897 1303 22931 1995
rect 23005 1303 23039 1995
rect 23515 1303 23549 1995
rect 22471 1203 22847 1237
rect 23089 1203 23465 1237
rect 25483 2195 25545 2229
rect 25545 2195 26791 2229
rect 26791 2195 26853 2229
rect 24071 2061 24447 2095
rect 24689 2061 25065 2095
rect 23987 1303 24021 1995
rect 24497 1303 24531 1995
rect 24605 1303 24639 1995
rect 25115 1303 25149 1995
rect 24071 1203 24447 1237
rect 24689 1203 25065 1237
rect 27083 2195 27145 2229
rect 27145 2195 28391 2229
rect 28391 2195 28453 2229
rect 25671 2061 26047 2095
rect 26289 2061 26665 2095
rect 25587 1303 25621 1995
rect 26097 1303 26131 1995
rect 26205 1303 26239 1995
rect 26715 1303 26749 1995
rect 25671 1203 26047 1237
rect 26289 1203 26665 1237
rect 28683 2195 28745 2229
rect 28745 2195 29991 2229
rect 29991 2195 30053 2229
rect 27271 2061 27647 2095
rect 27889 2061 28265 2095
rect 27187 1303 27221 1995
rect 27697 1303 27731 1995
rect 27805 1303 27839 1995
rect 28315 1303 28349 1995
rect 27271 1203 27647 1237
rect 27889 1203 28265 1237
rect 30283 2195 30345 2229
rect 30345 2195 31591 2229
rect 31591 2195 31653 2229
rect 28871 2061 29247 2095
rect 29489 2061 29865 2095
rect 28787 1303 28821 1995
rect 29297 1303 29331 1995
rect 29405 1303 29439 1995
rect 29915 1303 29949 1995
rect 28871 1203 29247 1237
rect 29489 1203 29865 1237
rect 31883 2195 31945 2229
rect 31945 2195 33191 2229
rect 33191 2195 33253 2229
rect 30471 2061 30847 2095
rect 31089 2061 31465 2095
rect 30387 1303 30421 1995
rect 30897 1303 30931 1995
rect 31005 1303 31039 1995
rect 31515 1303 31549 1995
rect 30471 1203 30847 1237
rect 31089 1203 31465 1237
rect 33483 2195 33545 2229
rect 33545 2195 34791 2229
rect 34791 2195 34853 2229
rect 32071 2061 32447 2095
rect 32689 2061 33065 2095
rect 31987 1303 32021 1995
rect 32497 1303 32531 1995
rect 32605 1303 32639 1995
rect 33115 1303 33149 1995
rect 32071 1203 32447 1237
rect 32689 1203 33065 1237
rect 35083 2195 35145 2229
rect 35145 2195 36391 2229
rect 36391 2195 36453 2229
rect 33671 2061 34047 2095
rect 34289 2061 34665 2095
rect 33587 1303 33621 1995
rect 34097 1303 34131 1995
rect 34205 1303 34239 1995
rect 34715 1303 34749 1995
rect 33671 1203 34047 1237
rect 34289 1203 34665 1237
rect 36683 2195 36745 2229
rect 36745 2195 37991 2229
rect 37991 2195 38053 2229
rect 35271 2061 35647 2095
rect 35889 2061 36265 2095
rect 35187 1303 35221 1995
rect 35697 1303 35731 1995
rect 35805 1303 35839 1995
rect 36315 1303 36349 1995
rect 35271 1203 35647 1237
rect 35889 1203 36265 1237
rect 36871 2061 37247 2095
rect 37489 2061 37865 2095
rect 36787 1303 36821 1995
rect 37297 1303 37331 1995
rect 37405 1303 37439 1995
rect 37915 1303 37949 1995
rect 36871 1203 37247 1237
rect 37489 1203 37865 1237
rect 71 915 447 949
rect 689 915 1065 949
rect -13 736 21 870
rect 497 736 531 870
rect 605 736 639 870
rect 1115 736 1149 870
rect 71 657 447 691
rect 689 657 1065 691
rect 1671 915 2047 949
rect 2289 915 2665 949
rect 1587 736 1621 870
rect 2097 736 2131 870
rect 2205 736 2239 870
rect 2715 736 2749 870
rect 1671 657 2047 691
rect 2289 657 2665 691
rect 3271 915 3647 949
rect 3889 915 4265 949
rect 3187 736 3221 870
rect 3697 736 3731 870
rect 3805 736 3839 870
rect 4315 736 4349 870
rect 3271 657 3647 691
rect 3889 657 4265 691
rect 4871 915 5247 949
rect 5489 915 5865 949
rect 4787 736 4821 870
rect 5297 736 5331 870
rect 5405 736 5439 870
rect 5915 736 5949 870
rect 4871 657 5247 691
rect 5489 657 5865 691
rect 6471 915 6847 949
rect 7089 915 7465 949
rect 6387 736 6421 870
rect 6897 736 6931 870
rect 7005 736 7039 870
rect 7515 736 7549 870
rect 6471 657 6847 691
rect 7089 657 7465 691
rect 8071 915 8447 949
rect 8689 915 9065 949
rect 7987 736 8021 870
rect 8497 736 8531 870
rect 8605 736 8639 870
rect 9115 736 9149 870
rect 8071 657 8447 691
rect 8689 657 9065 691
rect 9671 915 10047 949
rect 10289 915 10665 949
rect 9587 736 9621 870
rect 10097 736 10131 870
rect 10205 736 10239 870
rect 10715 736 10749 870
rect 9671 657 10047 691
rect 10289 657 10665 691
rect 11271 915 11647 949
rect 11889 915 12265 949
rect 11187 736 11221 870
rect 11697 736 11731 870
rect 11805 736 11839 870
rect 12315 736 12349 870
rect 11271 657 11647 691
rect 11889 657 12265 691
rect 12871 915 13247 949
rect 13489 915 13865 949
rect 12787 736 12821 870
rect 13297 736 13331 870
rect 13405 736 13439 870
rect 13915 736 13949 870
rect 12871 657 13247 691
rect 13489 657 13865 691
rect 14471 915 14847 949
rect 15089 915 15465 949
rect 14387 736 14421 870
rect 14897 736 14931 870
rect 15005 736 15039 870
rect 15515 736 15549 870
rect 14471 657 14847 691
rect 15089 657 15465 691
rect 16071 915 16447 949
rect 16689 915 17065 949
rect 15987 736 16021 870
rect 16497 736 16531 870
rect 16605 736 16639 870
rect 17115 736 17149 870
rect 16071 657 16447 691
rect 16689 657 17065 691
rect 17671 915 18047 949
rect 18289 915 18665 949
rect 17587 736 17621 870
rect 18097 736 18131 870
rect 18205 736 18239 870
rect 18715 736 18749 870
rect 17671 657 18047 691
rect 18289 657 18665 691
rect 19271 915 19647 949
rect 19889 915 20265 949
rect 19187 736 19221 870
rect 19697 736 19731 870
rect 19805 736 19839 870
rect 20315 736 20349 870
rect 19271 657 19647 691
rect 19889 657 20265 691
rect 20871 915 21247 949
rect 21489 915 21865 949
rect 20787 736 20821 870
rect 21297 736 21331 870
rect 21405 736 21439 870
rect 21915 736 21949 870
rect 20871 657 21247 691
rect 21489 657 21865 691
rect 22471 915 22847 949
rect 23089 915 23465 949
rect 22387 736 22421 870
rect 22897 736 22931 870
rect 23005 736 23039 870
rect 23515 736 23549 870
rect 22471 657 22847 691
rect 23089 657 23465 691
rect 24071 915 24447 949
rect 24689 915 25065 949
rect 23987 736 24021 870
rect 24497 736 24531 870
rect 24605 736 24639 870
rect 25115 736 25149 870
rect 24071 657 24447 691
rect 24689 657 25065 691
rect 25671 915 26047 949
rect 26289 915 26665 949
rect 25587 736 25621 870
rect 26097 736 26131 870
rect 26205 736 26239 870
rect 26715 736 26749 870
rect 25671 657 26047 691
rect 26289 657 26665 691
rect 27271 915 27647 949
rect 27889 915 28265 949
rect 27187 736 27221 870
rect 27697 736 27731 870
rect 27805 736 27839 870
rect 28315 736 28349 870
rect 27271 657 27647 691
rect 27889 657 28265 691
rect 28871 915 29247 949
rect 29489 915 29865 949
rect 28787 736 28821 870
rect 29297 736 29331 870
rect 29405 736 29439 870
rect 29915 736 29949 870
rect 28871 657 29247 691
rect 29489 657 29865 691
rect 30471 915 30847 949
rect 31089 915 31465 949
rect 30387 736 30421 870
rect 30897 736 30931 870
rect 31005 736 31039 870
rect 31515 736 31549 870
rect 30471 657 30847 691
rect 31089 657 31465 691
rect 32071 915 32447 949
rect 32689 915 33065 949
rect 31987 736 32021 870
rect 32497 736 32531 870
rect 32605 736 32639 870
rect 33115 736 33149 870
rect 32071 657 32447 691
rect 32689 657 33065 691
rect 33671 915 34047 949
rect 34289 915 34665 949
rect 33587 736 33621 870
rect 34097 736 34131 870
rect 34205 736 34239 870
rect 34715 736 34749 870
rect 33671 657 34047 691
rect 34289 657 34665 691
rect 35271 915 35647 949
rect 35889 915 36265 949
rect 35187 736 35221 870
rect 35697 736 35731 870
rect 35805 736 35839 870
rect 36315 736 36349 870
rect 35271 657 35647 691
rect 35889 657 36265 691
rect 36871 915 37247 949
rect 37489 915 37865 949
rect 36787 736 36821 870
rect 37297 736 37331 870
rect 37405 736 37439 870
rect 37915 736 37949 870
rect 36871 657 37247 691
rect 37489 657 37865 691
rect -117 395 -55 429
rect -55 395 1191 429
rect 1191 395 1253 429
rect 1483 395 1545 429
rect 1545 395 2791 429
rect 2791 395 2853 429
rect 71 261 447 295
rect 689 261 1065 295
rect -13 -497 21 195
rect 497 -497 531 195
rect 605 -497 639 195
rect 1115 -497 1149 195
rect 71 -597 447 -563
rect 689 -597 1065 -563
rect 3083 395 3145 429
rect 3145 395 4391 429
rect 4391 395 4453 429
rect 1671 261 2047 295
rect 2289 261 2665 295
rect 1587 -497 1621 195
rect 2097 -497 2131 195
rect 2205 -497 2239 195
rect 2715 -497 2749 195
rect 1671 -597 2047 -563
rect 2289 -597 2665 -563
rect 4683 395 4745 429
rect 4745 395 5991 429
rect 5991 395 6053 429
rect 3271 261 3647 295
rect 3889 261 4265 295
rect 3187 -497 3221 195
rect 3697 -497 3731 195
rect 3805 -497 3839 195
rect 4315 -497 4349 195
rect 3271 -597 3647 -563
rect 3889 -597 4265 -563
rect 6283 395 6345 429
rect 6345 395 7591 429
rect 7591 395 7653 429
rect 4871 261 5247 295
rect 5489 261 5865 295
rect 4787 -497 4821 195
rect 5297 -497 5331 195
rect 5405 -497 5439 195
rect 5915 -497 5949 195
rect 4871 -597 5247 -563
rect 5489 -597 5865 -563
rect 7883 395 7945 429
rect 7945 395 9191 429
rect 9191 395 9253 429
rect 6471 261 6847 295
rect 7089 261 7465 295
rect 6387 -497 6421 195
rect 6897 -497 6931 195
rect 7005 -497 7039 195
rect 7515 -497 7549 195
rect 6471 -597 6847 -563
rect 7089 -597 7465 -563
rect 9483 395 9545 429
rect 9545 395 10791 429
rect 10791 395 10853 429
rect 8071 261 8447 295
rect 8689 261 9065 295
rect 7987 -497 8021 195
rect 8497 -497 8531 195
rect 8605 -497 8639 195
rect 9115 -497 9149 195
rect 8071 -597 8447 -563
rect 8689 -597 9065 -563
rect 11083 395 11145 429
rect 11145 395 12391 429
rect 12391 395 12453 429
rect 9671 261 10047 295
rect 10289 261 10665 295
rect 9587 -497 9621 195
rect 10097 -497 10131 195
rect 10205 -497 10239 195
rect 10715 -497 10749 195
rect 9671 -597 10047 -563
rect 10289 -597 10665 -563
rect 12683 395 12745 429
rect 12745 395 13991 429
rect 13991 395 14053 429
rect 11271 261 11647 295
rect 11889 261 12265 295
rect 11187 -497 11221 195
rect 11697 -497 11731 195
rect 11805 -497 11839 195
rect 12315 -497 12349 195
rect 11271 -597 11647 -563
rect 11889 -597 12265 -563
rect 14283 395 14345 429
rect 14345 395 15591 429
rect 15591 395 15653 429
rect 12871 261 13247 295
rect 13489 261 13865 295
rect 12787 -497 12821 195
rect 13297 -497 13331 195
rect 13405 -497 13439 195
rect 13915 -497 13949 195
rect 12871 -597 13247 -563
rect 13489 -597 13865 -563
rect 15883 395 15945 429
rect 15945 395 17191 429
rect 17191 395 17253 429
rect 14471 261 14847 295
rect 15089 261 15465 295
rect 14387 -497 14421 195
rect 14897 -497 14931 195
rect 15005 -497 15039 195
rect 15515 -497 15549 195
rect 14471 -597 14847 -563
rect 15089 -597 15465 -563
rect 17483 395 17545 429
rect 17545 395 18791 429
rect 18791 395 18853 429
rect 16071 261 16447 295
rect 16689 261 17065 295
rect 15987 -497 16021 195
rect 16497 -497 16531 195
rect 16605 -497 16639 195
rect 17115 -497 17149 195
rect 16071 -597 16447 -563
rect 16689 -597 17065 -563
rect 19083 395 19145 429
rect 19145 395 20391 429
rect 20391 395 20453 429
rect 17671 261 18047 295
rect 18289 261 18665 295
rect 17587 -497 17621 195
rect 18097 -497 18131 195
rect 18205 -497 18239 195
rect 18715 -497 18749 195
rect 17671 -597 18047 -563
rect 18289 -597 18665 -563
rect 20683 395 20745 429
rect 20745 395 21991 429
rect 21991 395 22053 429
rect 19271 261 19647 295
rect 19889 261 20265 295
rect 19187 -497 19221 195
rect 19697 -497 19731 195
rect 19805 -497 19839 195
rect 20315 -497 20349 195
rect 19271 -597 19647 -563
rect 19889 -597 20265 -563
rect 22283 395 22345 429
rect 22345 395 23591 429
rect 23591 395 23653 429
rect 20871 261 21247 295
rect 21489 261 21865 295
rect 20787 -497 20821 195
rect 21297 -497 21331 195
rect 21405 -497 21439 195
rect 21915 -497 21949 195
rect 20871 -597 21247 -563
rect 21489 -597 21865 -563
rect 23883 395 23945 429
rect 23945 395 25191 429
rect 25191 395 25253 429
rect 22471 261 22847 295
rect 23089 261 23465 295
rect 22387 -497 22421 195
rect 22897 -497 22931 195
rect 23005 -497 23039 195
rect 23515 -497 23549 195
rect 22471 -597 22847 -563
rect 23089 -597 23465 -563
rect 25483 395 25545 429
rect 25545 395 26791 429
rect 26791 395 26853 429
rect 24071 261 24447 295
rect 24689 261 25065 295
rect 23987 -497 24021 195
rect 24497 -497 24531 195
rect 24605 -497 24639 195
rect 25115 -497 25149 195
rect 24071 -597 24447 -563
rect 24689 -597 25065 -563
rect 27083 395 27145 429
rect 27145 395 28391 429
rect 28391 395 28453 429
rect 25671 261 26047 295
rect 26289 261 26665 295
rect 25587 -497 25621 195
rect 26097 -497 26131 195
rect 26205 -497 26239 195
rect 26715 -497 26749 195
rect 25671 -597 26047 -563
rect 26289 -597 26665 -563
rect 28683 395 28745 429
rect 28745 395 29991 429
rect 29991 395 30053 429
rect 27271 261 27647 295
rect 27889 261 28265 295
rect 27187 -497 27221 195
rect 27697 -497 27731 195
rect 27805 -497 27839 195
rect 28315 -497 28349 195
rect 27271 -597 27647 -563
rect 27889 -597 28265 -563
rect 30283 395 30345 429
rect 30345 395 31591 429
rect 31591 395 31653 429
rect 28871 261 29247 295
rect 29489 261 29865 295
rect 28787 -497 28821 195
rect 29297 -497 29331 195
rect 29405 -497 29439 195
rect 29915 -497 29949 195
rect 28871 -597 29247 -563
rect 29489 -597 29865 -563
rect 31883 395 31945 429
rect 31945 395 33191 429
rect 33191 395 33253 429
rect 30471 261 30847 295
rect 31089 261 31465 295
rect 30387 -497 30421 195
rect 30897 -497 30931 195
rect 31005 -497 31039 195
rect 31515 -497 31549 195
rect 30471 -597 30847 -563
rect 31089 -597 31465 -563
rect 33483 395 33545 429
rect 33545 395 34791 429
rect 34791 395 34853 429
rect 32071 261 32447 295
rect 32689 261 33065 295
rect 31987 -497 32021 195
rect 32497 -497 32531 195
rect 32605 -497 32639 195
rect 33115 -497 33149 195
rect 32071 -597 32447 -563
rect 32689 -597 33065 -563
rect 35083 395 35145 429
rect 35145 395 36391 429
rect 36391 395 36453 429
rect 36683 395 36745 429
rect 36745 395 37991 429
rect 37991 395 38053 429
rect 33671 261 34047 295
rect 34289 261 34665 295
rect 33587 -497 33621 195
rect 34097 -497 34131 195
rect 34205 -497 34239 195
rect 34715 -497 34749 195
rect 33671 -597 34047 -563
rect 34289 -597 34665 -563
rect 35271 261 35647 295
rect 35889 261 36265 295
rect 35187 -497 35221 195
rect 35697 -497 35731 195
rect 35805 -497 35839 195
rect 36315 -497 36349 195
rect 35271 -597 35647 -563
rect 35889 -597 36265 -563
rect 36871 261 37247 295
rect 37489 261 37865 295
rect 36787 -497 36821 195
rect 37297 -497 37331 195
rect 37405 -497 37439 195
rect 37915 -497 37949 195
rect 36871 -597 37247 -563
rect 37489 -597 37865 -563
rect 71 -885 447 -851
rect 689 -885 1065 -851
rect -13 -1064 21 -930
rect 497 -1064 531 -930
rect 605 -1064 639 -930
rect 1115 -1064 1149 -930
rect 71 -1143 447 -1109
rect 689 -1143 1065 -1109
rect 1671 -885 2047 -851
rect 2289 -885 2665 -851
rect 1587 -1064 1621 -930
rect 2097 -1064 2131 -930
rect 2205 -1064 2239 -930
rect 2715 -1064 2749 -930
rect 1671 -1143 2047 -1109
rect 2289 -1143 2665 -1109
rect 3271 -885 3647 -851
rect 3889 -885 4265 -851
rect 3187 -1064 3221 -930
rect 3697 -1064 3731 -930
rect 3805 -1064 3839 -930
rect 4315 -1064 4349 -930
rect 3271 -1143 3647 -1109
rect 3889 -1143 4265 -1109
rect 4871 -885 5247 -851
rect 5489 -885 5865 -851
rect 4787 -1064 4821 -930
rect 5297 -1064 5331 -930
rect 5405 -1064 5439 -930
rect 5915 -1064 5949 -930
rect 4871 -1143 5247 -1109
rect 5489 -1143 5865 -1109
rect 6471 -885 6847 -851
rect 7089 -885 7465 -851
rect 6387 -1064 6421 -930
rect 6897 -1064 6931 -930
rect 7005 -1064 7039 -930
rect 7515 -1064 7549 -930
rect 6471 -1143 6847 -1109
rect 7089 -1143 7465 -1109
rect 8071 -885 8447 -851
rect 8689 -885 9065 -851
rect 7987 -1064 8021 -930
rect 8497 -1064 8531 -930
rect 8605 -1064 8639 -930
rect 9115 -1064 9149 -930
rect 8071 -1143 8447 -1109
rect 8689 -1143 9065 -1109
rect 9671 -885 10047 -851
rect 10289 -885 10665 -851
rect 9587 -1064 9621 -930
rect 10097 -1064 10131 -930
rect 10205 -1064 10239 -930
rect 10715 -1064 10749 -930
rect 9671 -1143 10047 -1109
rect 10289 -1143 10665 -1109
rect 11271 -885 11647 -851
rect 11889 -885 12265 -851
rect 11187 -1064 11221 -930
rect 11697 -1064 11731 -930
rect 11805 -1064 11839 -930
rect 12315 -1064 12349 -930
rect 11271 -1143 11647 -1109
rect 11889 -1143 12265 -1109
rect 12871 -885 13247 -851
rect 13489 -885 13865 -851
rect 12787 -1064 12821 -930
rect 13297 -1064 13331 -930
rect 13405 -1064 13439 -930
rect 13915 -1064 13949 -930
rect 12871 -1143 13247 -1109
rect 13489 -1143 13865 -1109
rect 14471 -885 14847 -851
rect 15089 -885 15465 -851
rect 14387 -1064 14421 -930
rect 14897 -1064 14931 -930
rect 15005 -1064 15039 -930
rect 15515 -1064 15549 -930
rect 14471 -1143 14847 -1109
rect 15089 -1143 15465 -1109
rect 16071 -885 16447 -851
rect 16689 -885 17065 -851
rect 15987 -1064 16021 -930
rect 16497 -1064 16531 -930
rect 16605 -1064 16639 -930
rect 17115 -1064 17149 -930
rect 16071 -1143 16447 -1109
rect 16689 -1143 17065 -1109
rect 17671 -885 18047 -851
rect 18289 -885 18665 -851
rect 17587 -1064 17621 -930
rect 18097 -1064 18131 -930
rect 18205 -1064 18239 -930
rect 18715 -1064 18749 -930
rect 17671 -1143 18047 -1109
rect 18289 -1143 18665 -1109
rect 19271 -885 19647 -851
rect 19889 -885 20265 -851
rect 19187 -1064 19221 -930
rect 19697 -1064 19731 -930
rect 19805 -1064 19839 -930
rect 20315 -1064 20349 -930
rect 19271 -1143 19647 -1109
rect 19889 -1143 20265 -1109
rect 20871 -885 21247 -851
rect 21489 -885 21865 -851
rect 20787 -1064 20821 -930
rect 21297 -1064 21331 -930
rect 21405 -1064 21439 -930
rect 21915 -1064 21949 -930
rect 20871 -1143 21247 -1109
rect 21489 -1143 21865 -1109
rect 22471 -885 22847 -851
rect 23089 -885 23465 -851
rect 22387 -1064 22421 -930
rect 22897 -1064 22931 -930
rect 23005 -1064 23039 -930
rect 23515 -1064 23549 -930
rect 22471 -1143 22847 -1109
rect 23089 -1143 23465 -1109
rect 24071 -885 24447 -851
rect 24689 -885 25065 -851
rect 23987 -1064 24021 -930
rect 24497 -1064 24531 -930
rect 24605 -1064 24639 -930
rect 25115 -1064 25149 -930
rect 24071 -1143 24447 -1109
rect 24689 -1143 25065 -1109
rect 25671 -885 26047 -851
rect 26289 -885 26665 -851
rect 25587 -1064 25621 -930
rect 26097 -1064 26131 -930
rect 26205 -1064 26239 -930
rect 26715 -1064 26749 -930
rect 25671 -1143 26047 -1109
rect 26289 -1143 26665 -1109
rect 27271 -885 27647 -851
rect 27889 -885 28265 -851
rect 27187 -1064 27221 -930
rect 27697 -1064 27731 -930
rect 27805 -1064 27839 -930
rect 28315 -1064 28349 -930
rect 27271 -1143 27647 -1109
rect 27889 -1143 28265 -1109
rect 28871 -885 29247 -851
rect 29489 -885 29865 -851
rect 28787 -1064 28821 -930
rect 29297 -1064 29331 -930
rect 29405 -1064 29439 -930
rect 29915 -1064 29949 -930
rect 28871 -1143 29247 -1109
rect 29489 -1143 29865 -1109
rect 30471 -885 30847 -851
rect 31089 -885 31465 -851
rect 30387 -1064 30421 -930
rect 30897 -1064 30931 -930
rect 31005 -1064 31039 -930
rect 31515 -1064 31549 -930
rect 30471 -1143 30847 -1109
rect 31089 -1143 31465 -1109
rect 32071 -885 32447 -851
rect 32689 -885 33065 -851
rect 31987 -1064 32021 -930
rect 32497 -1064 32531 -930
rect 32605 -1064 32639 -930
rect 33115 -1064 33149 -930
rect 32071 -1143 32447 -1109
rect 32689 -1143 33065 -1109
rect 33671 -885 34047 -851
rect 34289 -885 34665 -851
rect 33587 -1064 33621 -930
rect 34097 -1064 34131 -930
rect 34205 -1064 34239 -930
rect 34715 -1064 34749 -930
rect 33671 -1143 34047 -1109
rect 34289 -1143 34665 -1109
rect 35271 -885 35647 -851
rect 35889 -885 36265 -851
rect 35187 -1064 35221 -930
rect 35697 -1064 35731 -930
rect 35805 -1064 35839 -930
rect 36315 -1064 36349 -930
rect 35271 -1143 35647 -1109
rect 35889 -1143 36265 -1109
rect 36871 -885 37247 -851
rect 37489 -885 37865 -851
rect 36787 -1064 36821 -930
rect 37297 -1064 37331 -930
rect 37405 -1064 37439 -930
rect 37915 -1064 37949 -930
rect 36871 -1143 37247 -1109
rect 37489 -1143 37865 -1109
rect -117 -1405 -55 -1371
rect -55 -1405 1191 -1371
rect 1191 -1405 1253 -1371
rect 1483 -1405 1545 -1371
rect 1545 -1405 2791 -1371
rect 2791 -1405 2853 -1371
rect 71 -1539 447 -1505
rect 689 -1539 1065 -1505
rect -13 -2297 21 -1605
rect 497 -2297 531 -1605
rect 605 -2297 639 -1605
rect 1115 -2297 1149 -1605
rect 71 -2397 447 -2363
rect 689 -2397 1065 -2363
rect 3083 -1405 3145 -1371
rect 3145 -1405 4391 -1371
rect 4391 -1405 4453 -1371
rect 1671 -1539 2047 -1505
rect 2289 -1539 2665 -1505
rect 1587 -2297 1621 -1605
rect 2097 -2297 2131 -1605
rect 2205 -2297 2239 -1605
rect 2715 -2297 2749 -1605
rect 1671 -2397 2047 -2363
rect 2289 -2397 2665 -2363
rect 4683 -1405 4745 -1371
rect 4745 -1405 5991 -1371
rect 5991 -1405 6053 -1371
rect 3271 -1539 3647 -1505
rect 3889 -1539 4265 -1505
rect 3187 -2297 3221 -1605
rect 3697 -2297 3731 -1605
rect 3805 -2297 3839 -1605
rect 4315 -2297 4349 -1605
rect 3271 -2397 3647 -2363
rect 3889 -2397 4265 -2363
rect 6283 -1405 6345 -1371
rect 6345 -1405 7591 -1371
rect 7591 -1405 7653 -1371
rect 4871 -1539 5247 -1505
rect 5489 -1539 5865 -1505
rect 4787 -2297 4821 -1605
rect 5297 -2297 5331 -1605
rect 5405 -2297 5439 -1605
rect 5915 -2297 5949 -1605
rect 4871 -2397 5247 -2363
rect 5489 -2397 5865 -2363
rect 7883 -1405 7945 -1371
rect 7945 -1405 9191 -1371
rect 9191 -1405 9253 -1371
rect 6471 -1539 6847 -1505
rect 7089 -1539 7465 -1505
rect 6387 -2297 6421 -1605
rect 6897 -2297 6931 -1605
rect 7005 -2297 7039 -1605
rect 7515 -2297 7549 -1605
rect 6471 -2397 6847 -2363
rect 7089 -2397 7465 -2363
rect 9483 -1405 9545 -1371
rect 9545 -1405 10791 -1371
rect 10791 -1405 10853 -1371
rect 8071 -1539 8447 -1505
rect 8689 -1539 9065 -1505
rect 7987 -2297 8021 -1605
rect 8497 -2297 8531 -1605
rect 8605 -2297 8639 -1605
rect 9115 -2297 9149 -1605
rect 8071 -2397 8447 -2363
rect 8689 -2397 9065 -2363
rect 11083 -1405 11145 -1371
rect 11145 -1405 12391 -1371
rect 12391 -1405 12453 -1371
rect 9671 -1539 10047 -1505
rect 10289 -1539 10665 -1505
rect 9587 -2297 9621 -1605
rect 10097 -2297 10131 -1605
rect 10205 -2297 10239 -1605
rect 10715 -2297 10749 -1605
rect 9671 -2397 10047 -2363
rect 10289 -2397 10665 -2363
rect 12683 -1405 12745 -1371
rect 12745 -1405 13991 -1371
rect 13991 -1405 14053 -1371
rect 11271 -1539 11647 -1505
rect 11889 -1539 12265 -1505
rect 11187 -2297 11221 -1605
rect 11697 -2297 11731 -1605
rect 11805 -2297 11839 -1605
rect 12315 -2297 12349 -1605
rect 11271 -2397 11647 -2363
rect 11889 -2397 12265 -2363
rect 14283 -1405 14345 -1371
rect 14345 -1405 15591 -1371
rect 15591 -1405 15653 -1371
rect 12871 -1539 13247 -1505
rect 13489 -1539 13865 -1505
rect 12787 -2297 12821 -1605
rect 13297 -2297 13331 -1605
rect 13405 -2297 13439 -1605
rect 13915 -2297 13949 -1605
rect 12871 -2397 13247 -2363
rect 13489 -2397 13865 -2363
rect 15883 -1405 15945 -1371
rect 15945 -1405 17191 -1371
rect 17191 -1405 17253 -1371
rect 14471 -1539 14847 -1505
rect 15089 -1539 15465 -1505
rect 14387 -2297 14421 -1605
rect 14897 -2297 14931 -1605
rect 15005 -2297 15039 -1605
rect 15515 -2297 15549 -1605
rect 14471 -2397 14847 -2363
rect 15089 -2397 15465 -2363
rect 17483 -1405 17545 -1371
rect 17545 -1405 18791 -1371
rect 18791 -1405 18853 -1371
rect 16071 -1539 16447 -1505
rect 16689 -1539 17065 -1505
rect 15987 -2297 16021 -1605
rect 16497 -2297 16531 -1605
rect 16605 -2297 16639 -1605
rect 17115 -2297 17149 -1605
rect 16071 -2397 16447 -2363
rect 16689 -2397 17065 -2363
rect 19083 -1405 19145 -1371
rect 19145 -1405 20391 -1371
rect 20391 -1405 20453 -1371
rect 17671 -1539 18047 -1505
rect 18289 -1539 18665 -1505
rect 17587 -2297 17621 -1605
rect 18097 -2297 18131 -1605
rect 18205 -2297 18239 -1605
rect 18715 -2297 18749 -1605
rect 17671 -2397 18047 -2363
rect 18289 -2397 18665 -2363
rect 20683 -1405 20745 -1371
rect 20745 -1405 21991 -1371
rect 21991 -1405 22053 -1371
rect 19271 -1539 19647 -1505
rect 19889 -1539 20265 -1505
rect 19187 -2297 19221 -1605
rect 19697 -2297 19731 -1605
rect 19805 -2297 19839 -1605
rect 20315 -2297 20349 -1605
rect 19271 -2397 19647 -2363
rect 19889 -2397 20265 -2363
rect 22283 -1405 22345 -1371
rect 22345 -1405 23591 -1371
rect 23591 -1405 23653 -1371
rect 20871 -1539 21247 -1505
rect 21489 -1539 21865 -1505
rect 20787 -2297 20821 -1605
rect 21297 -2297 21331 -1605
rect 21405 -2297 21439 -1605
rect 21915 -2297 21949 -1605
rect 20871 -2397 21247 -2363
rect 21489 -2397 21865 -2363
rect 23883 -1405 23945 -1371
rect 23945 -1405 25191 -1371
rect 25191 -1405 25253 -1371
rect 22471 -1539 22847 -1505
rect 23089 -1539 23465 -1505
rect 22387 -2297 22421 -1605
rect 22897 -2297 22931 -1605
rect 23005 -2297 23039 -1605
rect 23515 -2297 23549 -1605
rect 22471 -2397 22847 -2363
rect 23089 -2397 23465 -2363
rect 25483 -1405 25545 -1371
rect 25545 -1405 26791 -1371
rect 26791 -1405 26853 -1371
rect 24071 -1539 24447 -1505
rect 24689 -1539 25065 -1505
rect 23987 -2297 24021 -1605
rect 24497 -2297 24531 -1605
rect 24605 -2297 24639 -1605
rect 25115 -2297 25149 -1605
rect 24071 -2397 24447 -2363
rect 24689 -2397 25065 -2363
rect 27083 -1405 27145 -1371
rect 27145 -1405 28391 -1371
rect 28391 -1405 28453 -1371
rect 25671 -1539 26047 -1505
rect 26289 -1539 26665 -1505
rect 25587 -2297 25621 -1605
rect 26097 -2297 26131 -1605
rect 26205 -2297 26239 -1605
rect 26715 -2297 26749 -1605
rect 25671 -2397 26047 -2363
rect 26289 -2397 26665 -2363
rect 28683 -1405 28745 -1371
rect 28745 -1405 29991 -1371
rect 29991 -1405 30053 -1371
rect 27271 -1539 27647 -1505
rect 27889 -1539 28265 -1505
rect 27187 -2297 27221 -1605
rect 27697 -2297 27731 -1605
rect 27805 -2297 27839 -1605
rect 28315 -2297 28349 -1605
rect 27271 -2397 27647 -2363
rect 27889 -2397 28265 -2363
rect 30283 -1405 30345 -1371
rect 30345 -1405 31591 -1371
rect 31591 -1405 31653 -1371
rect 28871 -1539 29247 -1505
rect 29489 -1539 29865 -1505
rect 28787 -2297 28821 -1605
rect 29297 -2297 29331 -1605
rect 29405 -2297 29439 -1605
rect 29915 -2297 29949 -1605
rect 28871 -2397 29247 -2363
rect 29489 -2397 29865 -2363
rect 31883 -1405 31945 -1371
rect 31945 -1405 33191 -1371
rect 33191 -1405 33253 -1371
rect 30471 -1539 30847 -1505
rect 31089 -1539 31465 -1505
rect 30387 -2297 30421 -1605
rect 30897 -2297 30931 -1605
rect 31005 -2297 31039 -1605
rect 31515 -2297 31549 -1605
rect 30471 -2397 30847 -2363
rect 31089 -2397 31465 -2363
rect 33483 -1405 33545 -1371
rect 33545 -1405 34791 -1371
rect 34791 -1405 34853 -1371
rect 32071 -1539 32447 -1505
rect 32689 -1539 33065 -1505
rect 31987 -2297 32021 -1605
rect 32497 -2297 32531 -1605
rect 32605 -2297 32639 -1605
rect 33115 -2297 33149 -1605
rect 32071 -2397 32447 -2363
rect 32689 -2397 33065 -2363
rect 35083 -1405 35145 -1371
rect 35145 -1405 36391 -1371
rect 36391 -1405 36453 -1371
rect 36683 -1405 36745 -1371
rect 36745 -1405 37991 -1371
rect 37991 -1405 38053 -1371
rect 33671 -1539 34047 -1505
rect 34289 -1539 34665 -1505
rect 33587 -2297 33621 -1605
rect 34097 -2297 34131 -1605
rect 34205 -2297 34239 -1605
rect 34715 -2297 34749 -1605
rect 33671 -2397 34047 -2363
rect 34289 -2397 34665 -2363
rect 35271 -1539 35647 -1505
rect 35889 -1539 36265 -1505
rect 35187 -2297 35221 -1605
rect 35697 -2297 35731 -1605
rect 35805 -2297 35839 -1605
rect 36315 -2297 36349 -1605
rect 35271 -2397 35647 -2363
rect 35889 -2397 36265 -2363
rect 36871 -1539 37247 -1505
rect 37489 -1539 37865 -1505
rect 36787 -2297 36821 -1605
rect 37297 -2297 37331 -1605
rect 37405 -2297 37439 -1605
rect 37915 -2297 37949 -1605
rect 36871 -2397 37247 -2363
rect 37489 -2397 37865 -2363
rect 71 -2685 447 -2651
rect 689 -2685 1065 -2651
rect -13 -2864 21 -2730
rect 497 -2864 531 -2730
rect 605 -2864 639 -2730
rect 1115 -2864 1149 -2730
rect 71 -2943 447 -2909
rect 689 -2943 1065 -2909
rect 1671 -2685 2047 -2651
rect 2289 -2685 2665 -2651
rect 1587 -2864 1621 -2730
rect 2097 -2864 2131 -2730
rect 2205 -2864 2239 -2730
rect 2715 -2864 2749 -2730
rect 1671 -2943 2047 -2909
rect 2289 -2943 2665 -2909
rect 3271 -2685 3647 -2651
rect 3889 -2685 4265 -2651
rect 3187 -2864 3221 -2730
rect 3697 -2864 3731 -2730
rect 3805 -2864 3839 -2730
rect 4315 -2864 4349 -2730
rect 3271 -2943 3647 -2909
rect 3889 -2943 4265 -2909
rect 4871 -2685 5247 -2651
rect 5489 -2685 5865 -2651
rect 4787 -2864 4821 -2730
rect 5297 -2864 5331 -2730
rect 5405 -2864 5439 -2730
rect 5915 -2864 5949 -2730
rect 4871 -2943 5247 -2909
rect 5489 -2943 5865 -2909
rect 6471 -2685 6847 -2651
rect 7089 -2685 7465 -2651
rect 6387 -2864 6421 -2730
rect 6897 -2864 6931 -2730
rect 7005 -2864 7039 -2730
rect 7515 -2864 7549 -2730
rect 6471 -2943 6847 -2909
rect 7089 -2943 7465 -2909
rect 8071 -2685 8447 -2651
rect 8689 -2685 9065 -2651
rect 7987 -2864 8021 -2730
rect 8497 -2864 8531 -2730
rect 8605 -2864 8639 -2730
rect 9115 -2864 9149 -2730
rect 8071 -2943 8447 -2909
rect 8689 -2943 9065 -2909
rect 9671 -2685 10047 -2651
rect 10289 -2685 10665 -2651
rect 9587 -2864 9621 -2730
rect 10097 -2864 10131 -2730
rect 10205 -2864 10239 -2730
rect 10715 -2864 10749 -2730
rect 9671 -2943 10047 -2909
rect 10289 -2943 10665 -2909
rect 11271 -2685 11647 -2651
rect 11889 -2685 12265 -2651
rect 11187 -2864 11221 -2730
rect 11697 -2864 11731 -2730
rect 11805 -2864 11839 -2730
rect 12315 -2864 12349 -2730
rect 11271 -2943 11647 -2909
rect 11889 -2943 12265 -2909
rect 12871 -2685 13247 -2651
rect 13489 -2685 13865 -2651
rect 12787 -2864 12821 -2730
rect 13297 -2864 13331 -2730
rect 13405 -2864 13439 -2730
rect 13915 -2864 13949 -2730
rect 12871 -2943 13247 -2909
rect 13489 -2943 13865 -2909
rect 14471 -2685 14847 -2651
rect 15089 -2685 15465 -2651
rect 14387 -2864 14421 -2730
rect 14897 -2864 14931 -2730
rect 15005 -2864 15039 -2730
rect 15515 -2864 15549 -2730
rect 14471 -2943 14847 -2909
rect 15089 -2943 15465 -2909
rect 16071 -2685 16447 -2651
rect 16689 -2685 17065 -2651
rect 15987 -2864 16021 -2730
rect 16497 -2864 16531 -2730
rect 16605 -2864 16639 -2730
rect 17115 -2864 17149 -2730
rect 16071 -2943 16447 -2909
rect 16689 -2943 17065 -2909
rect 17671 -2685 18047 -2651
rect 18289 -2685 18665 -2651
rect 17587 -2864 17621 -2730
rect 18097 -2864 18131 -2730
rect 18205 -2864 18239 -2730
rect 18715 -2864 18749 -2730
rect 17671 -2943 18047 -2909
rect 18289 -2943 18665 -2909
rect 19271 -2685 19647 -2651
rect 19889 -2685 20265 -2651
rect 19187 -2864 19221 -2730
rect 19697 -2864 19731 -2730
rect 19805 -2864 19839 -2730
rect 20315 -2864 20349 -2730
rect 19271 -2943 19647 -2909
rect 19889 -2943 20265 -2909
rect 20871 -2685 21247 -2651
rect 21489 -2685 21865 -2651
rect 20787 -2864 20821 -2730
rect 21297 -2864 21331 -2730
rect 21405 -2864 21439 -2730
rect 21915 -2864 21949 -2730
rect 20871 -2943 21247 -2909
rect 21489 -2943 21865 -2909
rect 22471 -2685 22847 -2651
rect 23089 -2685 23465 -2651
rect 22387 -2864 22421 -2730
rect 22897 -2864 22931 -2730
rect 23005 -2864 23039 -2730
rect 23515 -2864 23549 -2730
rect 22471 -2943 22847 -2909
rect 23089 -2943 23465 -2909
rect 24071 -2685 24447 -2651
rect 24689 -2685 25065 -2651
rect 23987 -2864 24021 -2730
rect 24497 -2864 24531 -2730
rect 24605 -2864 24639 -2730
rect 25115 -2864 25149 -2730
rect 24071 -2943 24447 -2909
rect 24689 -2943 25065 -2909
rect 25671 -2685 26047 -2651
rect 26289 -2685 26665 -2651
rect 25587 -2864 25621 -2730
rect 26097 -2864 26131 -2730
rect 26205 -2864 26239 -2730
rect 26715 -2864 26749 -2730
rect 25671 -2943 26047 -2909
rect 26289 -2943 26665 -2909
rect 27271 -2685 27647 -2651
rect 27889 -2685 28265 -2651
rect 27187 -2864 27221 -2730
rect 27697 -2864 27731 -2730
rect 27805 -2864 27839 -2730
rect 28315 -2864 28349 -2730
rect 27271 -2943 27647 -2909
rect 27889 -2943 28265 -2909
rect 28871 -2685 29247 -2651
rect 29489 -2685 29865 -2651
rect 28787 -2864 28821 -2730
rect 29297 -2864 29331 -2730
rect 29405 -2864 29439 -2730
rect 29915 -2864 29949 -2730
rect 28871 -2943 29247 -2909
rect 29489 -2943 29865 -2909
rect 30471 -2685 30847 -2651
rect 31089 -2685 31465 -2651
rect 30387 -2864 30421 -2730
rect 30897 -2864 30931 -2730
rect 31005 -2864 31039 -2730
rect 31515 -2864 31549 -2730
rect 30471 -2943 30847 -2909
rect 31089 -2943 31465 -2909
rect 32071 -2685 32447 -2651
rect 32689 -2685 33065 -2651
rect 31987 -2864 32021 -2730
rect 32497 -2864 32531 -2730
rect 32605 -2864 32639 -2730
rect 33115 -2864 33149 -2730
rect 32071 -2943 32447 -2909
rect 32689 -2943 33065 -2909
rect 33671 -2685 34047 -2651
rect 34289 -2685 34665 -2651
rect 33587 -2864 33621 -2730
rect 34097 -2864 34131 -2730
rect 34205 -2864 34239 -2730
rect 34715 -2864 34749 -2730
rect 33671 -2943 34047 -2909
rect 34289 -2943 34665 -2909
rect 35271 -2685 35647 -2651
rect 35889 -2685 36265 -2651
rect 35187 -2864 35221 -2730
rect 35697 -2864 35731 -2730
rect 35805 -2864 35839 -2730
rect 36315 -2864 36349 -2730
rect 35271 -2943 35647 -2909
rect 35889 -2943 36265 -2909
rect 36871 -2685 37247 -2651
rect 37489 -2685 37865 -2651
rect 36787 -2864 36821 -2730
rect 37297 -2864 37331 -2730
rect 37405 -2864 37439 -2730
rect 37915 -2864 37949 -2730
rect 36871 -2943 37247 -2909
rect 37489 -2943 37865 -2909
rect -117 -3205 -55 -3171
rect -55 -3205 1191 -3171
rect 1191 -3205 1253 -3171
rect 1483 -3205 1545 -3171
rect 1545 -3205 2791 -3171
rect 2791 -3205 2853 -3171
rect 71 -3339 447 -3305
rect 689 -3339 1065 -3305
rect -13 -4097 21 -3405
rect 497 -4097 531 -3405
rect 605 -4097 639 -3405
rect 1115 -4097 1149 -3405
rect 71 -4197 447 -4163
rect 689 -4197 1065 -4163
rect 3083 -3205 3145 -3171
rect 3145 -3205 4391 -3171
rect 4391 -3205 4453 -3171
rect 1671 -3339 2047 -3305
rect 2289 -3339 2665 -3305
rect 1587 -4097 1621 -3405
rect 2097 -4097 2131 -3405
rect 2205 -4097 2239 -3405
rect 2715 -4097 2749 -3405
rect 1671 -4197 2047 -4163
rect 2289 -4197 2665 -4163
rect 4683 -3205 4745 -3171
rect 4745 -3205 5991 -3171
rect 5991 -3205 6053 -3171
rect 3271 -3339 3647 -3305
rect 3889 -3339 4265 -3305
rect 3187 -4097 3221 -3405
rect 3697 -4097 3731 -3405
rect 3805 -4097 3839 -3405
rect 4315 -4097 4349 -3405
rect 3271 -4197 3647 -4163
rect 3889 -4197 4265 -4163
rect 6283 -3205 6345 -3171
rect 6345 -3205 7591 -3171
rect 7591 -3205 7653 -3171
rect 4871 -3339 5247 -3305
rect 5489 -3339 5865 -3305
rect 4787 -4097 4821 -3405
rect 5297 -4097 5331 -3405
rect 5405 -4097 5439 -3405
rect 5915 -4097 5949 -3405
rect 4871 -4197 5247 -4163
rect 5489 -4197 5865 -4163
rect 7883 -3205 7945 -3171
rect 7945 -3205 9191 -3171
rect 9191 -3205 9253 -3171
rect 6471 -3339 6847 -3305
rect 7089 -3339 7465 -3305
rect 6387 -4097 6421 -3405
rect 6897 -4097 6931 -3405
rect 7005 -4097 7039 -3405
rect 7515 -4097 7549 -3405
rect 6471 -4197 6847 -4163
rect 7089 -4197 7465 -4163
rect 9483 -3205 9545 -3171
rect 9545 -3205 10791 -3171
rect 10791 -3205 10853 -3171
rect 8071 -3339 8447 -3305
rect 8689 -3339 9065 -3305
rect 7987 -4097 8021 -3405
rect 8497 -4097 8531 -3405
rect 8605 -4097 8639 -3405
rect 9115 -4097 9149 -3405
rect 8071 -4197 8447 -4163
rect 8689 -4197 9065 -4163
rect 11083 -3205 11145 -3171
rect 11145 -3205 12391 -3171
rect 12391 -3205 12453 -3171
rect 9671 -3339 10047 -3305
rect 10289 -3339 10665 -3305
rect 9587 -4097 9621 -3405
rect 10097 -4097 10131 -3405
rect 10205 -4097 10239 -3405
rect 10715 -4097 10749 -3405
rect 9671 -4197 10047 -4163
rect 10289 -4197 10665 -4163
rect 12683 -3205 12745 -3171
rect 12745 -3205 13991 -3171
rect 13991 -3205 14053 -3171
rect 11271 -3339 11647 -3305
rect 11889 -3339 12265 -3305
rect 11187 -4097 11221 -3405
rect 11697 -4097 11731 -3405
rect 11805 -4097 11839 -3405
rect 12315 -4097 12349 -3405
rect 11271 -4197 11647 -4163
rect 11889 -4197 12265 -4163
rect 14283 -3205 14345 -3171
rect 14345 -3205 15591 -3171
rect 15591 -3205 15653 -3171
rect 12871 -3339 13247 -3305
rect 13489 -3339 13865 -3305
rect 12787 -4097 12821 -3405
rect 13297 -4097 13331 -3405
rect 13405 -4097 13439 -3405
rect 13915 -4097 13949 -3405
rect 12871 -4197 13247 -4163
rect 13489 -4197 13865 -4163
rect 15883 -3205 15945 -3171
rect 15945 -3205 17191 -3171
rect 17191 -3205 17253 -3171
rect 14471 -3339 14847 -3305
rect 15089 -3339 15465 -3305
rect 14387 -4097 14421 -3405
rect 14897 -4097 14931 -3405
rect 15005 -4097 15039 -3405
rect 15515 -4097 15549 -3405
rect 14471 -4197 14847 -4163
rect 15089 -4197 15465 -4163
rect 17483 -3205 17545 -3171
rect 17545 -3205 18791 -3171
rect 18791 -3205 18853 -3171
rect 16071 -3339 16447 -3305
rect 16689 -3339 17065 -3305
rect 15987 -4097 16021 -3405
rect 16497 -4097 16531 -3405
rect 16605 -4097 16639 -3405
rect 17115 -4097 17149 -3405
rect 16071 -4197 16447 -4163
rect 16689 -4197 17065 -4163
rect 19083 -3205 19145 -3171
rect 19145 -3205 20391 -3171
rect 20391 -3205 20453 -3171
rect 17671 -3339 18047 -3305
rect 18289 -3339 18665 -3305
rect 17587 -4097 17621 -3405
rect 18097 -4097 18131 -3405
rect 18205 -4097 18239 -3405
rect 18715 -4097 18749 -3405
rect 17671 -4197 18047 -4163
rect 18289 -4197 18665 -4163
rect 20683 -3205 20745 -3171
rect 20745 -3205 21991 -3171
rect 21991 -3205 22053 -3171
rect 19271 -3339 19647 -3305
rect 19889 -3339 20265 -3305
rect 19187 -4097 19221 -3405
rect 19697 -4097 19731 -3405
rect 19805 -4097 19839 -3405
rect 20315 -4097 20349 -3405
rect 19271 -4197 19647 -4163
rect 19889 -4197 20265 -4163
rect 22283 -3205 22345 -3171
rect 22345 -3205 23591 -3171
rect 23591 -3205 23653 -3171
rect 20871 -3339 21247 -3305
rect 21489 -3339 21865 -3305
rect 20787 -4097 20821 -3405
rect 21297 -4097 21331 -3405
rect 21405 -4097 21439 -3405
rect 21915 -4097 21949 -3405
rect 20871 -4197 21247 -4163
rect 21489 -4197 21865 -4163
rect 23883 -3205 23945 -3171
rect 23945 -3205 25191 -3171
rect 25191 -3205 25253 -3171
rect 22471 -3339 22847 -3305
rect 23089 -3339 23465 -3305
rect 22387 -4097 22421 -3405
rect 22897 -4097 22931 -3405
rect 23005 -4097 23039 -3405
rect 23515 -4097 23549 -3405
rect 22471 -4197 22847 -4163
rect 23089 -4197 23465 -4163
rect 25483 -3205 25545 -3171
rect 25545 -3205 26791 -3171
rect 26791 -3205 26853 -3171
rect 24071 -3339 24447 -3305
rect 24689 -3339 25065 -3305
rect 23987 -4097 24021 -3405
rect 24497 -4097 24531 -3405
rect 24605 -4097 24639 -3405
rect 25115 -4097 25149 -3405
rect 24071 -4197 24447 -4163
rect 24689 -4197 25065 -4163
rect 27083 -3205 27145 -3171
rect 27145 -3205 28391 -3171
rect 28391 -3205 28453 -3171
rect 25671 -3339 26047 -3305
rect 26289 -3339 26665 -3305
rect 25587 -4097 25621 -3405
rect 26097 -4097 26131 -3405
rect 26205 -4097 26239 -3405
rect 26715 -4097 26749 -3405
rect 25671 -4197 26047 -4163
rect 26289 -4197 26665 -4163
rect 28683 -3205 28745 -3171
rect 28745 -3205 29991 -3171
rect 29991 -3205 30053 -3171
rect 27271 -3339 27647 -3305
rect 27889 -3339 28265 -3305
rect 27187 -4097 27221 -3405
rect 27697 -4097 27731 -3405
rect 27805 -4097 27839 -3405
rect 28315 -4097 28349 -3405
rect 27271 -4197 27647 -4163
rect 27889 -4197 28265 -4163
rect 30283 -3205 30345 -3171
rect 30345 -3205 31591 -3171
rect 31591 -3205 31653 -3171
rect 28871 -3339 29247 -3305
rect 29489 -3339 29865 -3305
rect 28787 -4097 28821 -3405
rect 29297 -4097 29331 -3405
rect 29405 -4097 29439 -3405
rect 29915 -4097 29949 -3405
rect 28871 -4197 29247 -4163
rect 29489 -4197 29865 -4163
rect 31883 -3205 31945 -3171
rect 31945 -3205 33191 -3171
rect 33191 -3205 33253 -3171
rect 30471 -3339 30847 -3305
rect 31089 -3339 31465 -3305
rect 30387 -4097 30421 -3405
rect 30897 -4097 30931 -3405
rect 31005 -4097 31039 -3405
rect 31515 -4097 31549 -3405
rect 30471 -4197 30847 -4163
rect 31089 -4197 31465 -4163
rect 33483 -3205 33545 -3171
rect 33545 -3205 34791 -3171
rect 34791 -3205 34853 -3171
rect 32071 -3339 32447 -3305
rect 32689 -3339 33065 -3305
rect 31987 -4097 32021 -3405
rect 32497 -4097 32531 -3405
rect 32605 -4097 32639 -3405
rect 33115 -4097 33149 -3405
rect 32071 -4197 32447 -4163
rect 32689 -4197 33065 -4163
rect 35083 -3205 35145 -3171
rect 35145 -3205 36391 -3171
rect 36391 -3205 36453 -3171
rect 36683 -3205 36745 -3171
rect 36745 -3205 37991 -3171
rect 37991 -3205 38053 -3171
rect 33671 -3339 34047 -3305
rect 34289 -3339 34665 -3305
rect 33587 -4097 33621 -3405
rect 34097 -4097 34131 -3405
rect 34205 -4097 34239 -3405
rect 34715 -4097 34749 -3405
rect 33671 -4197 34047 -4163
rect 34289 -4197 34665 -4163
rect 35271 -3339 35647 -3305
rect 35889 -3339 36265 -3305
rect 35187 -4097 35221 -3405
rect 35697 -4097 35731 -3405
rect 35805 -4097 35839 -3405
rect 36315 -4097 36349 -3405
rect 35271 -4197 35647 -4163
rect 35889 -4197 36265 -4163
rect 36871 -3339 37247 -3305
rect 37489 -3339 37865 -3305
rect 36787 -4097 36821 -3405
rect 37297 -4097 37331 -3405
rect 37405 -4097 37439 -3405
rect 37915 -4097 37949 -3405
rect 36871 -4197 37247 -4163
rect 37489 -4197 37865 -4163
rect 71 -4485 447 -4451
rect 689 -4485 1065 -4451
rect -13 -4664 21 -4530
rect 497 -4664 531 -4530
rect 605 -4664 639 -4530
rect 1115 -4664 1149 -4530
rect 71 -4743 447 -4709
rect 689 -4743 1065 -4709
rect 1671 -4485 2047 -4451
rect 2289 -4485 2665 -4451
rect 1587 -4664 1621 -4530
rect 2097 -4664 2131 -4530
rect 2205 -4664 2239 -4530
rect 2715 -4664 2749 -4530
rect 1671 -4743 2047 -4709
rect 2289 -4743 2665 -4709
rect 3271 -4485 3647 -4451
rect 3889 -4485 4265 -4451
rect 3187 -4664 3221 -4530
rect 3697 -4664 3731 -4530
rect 3805 -4664 3839 -4530
rect 4315 -4664 4349 -4530
rect 3271 -4743 3647 -4709
rect 3889 -4743 4265 -4709
rect 4871 -4485 5247 -4451
rect 5489 -4485 5865 -4451
rect 4787 -4664 4821 -4530
rect 5297 -4664 5331 -4530
rect 5405 -4664 5439 -4530
rect 5915 -4664 5949 -4530
rect 4871 -4743 5247 -4709
rect 5489 -4743 5865 -4709
rect 6471 -4485 6847 -4451
rect 7089 -4485 7465 -4451
rect 6387 -4664 6421 -4530
rect 6897 -4664 6931 -4530
rect 7005 -4664 7039 -4530
rect 7515 -4664 7549 -4530
rect 6471 -4743 6847 -4709
rect 7089 -4743 7465 -4709
rect 8071 -4485 8447 -4451
rect 8689 -4485 9065 -4451
rect 7987 -4664 8021 -4530
rect 8497 -4664 8531 -4530
rect 8605 -4664 8639 -4530
rect 9115 -4664 9149 -4530
rect 8071 -4743 8447 -4709
rect 8689 -4743 9065 -4709
rect 9671 -4485 10047 -4451
rect 10289 -4485 10665 -4451
rect 9587 -4664 9621 -4530
rect 10097 -4664 10131 -4530
rect 10205 -4664 10239 -4530
rect 10715 -4664 10749 -4530
rect 9671 -4743 10047 -4709
rect 10289 -4743 10665 -4709
rect 11271 -4485 11647 -4451
rect 11889 -4485 12265 -4451
rect 11187 -4664 11221 -4530
rect 11697 -4664 11731 -4530
rect 11805 -4664 11839 -4530
rect 12315 -4664 12349 -4530
rect 11271 -4743 11647 -4709
rect 11889 -4743 12265 -4709
rect 12871 -4485 13247 -4451
rect 13489 -4485 13865 -4451
rect 12787 -4664 12821 -4530
rect 13297 -4664 13331 -4530
rect 13405 -4664 13439 -4530
rect 13915 -4664 13949 -4530
rect 12871 -4743 13247 -4709
rect 13489 -4743 13865 -4709
rect 14471 -4485 14847 -4451
rect 15089 -4485 15465 -4451
rect 14387 -4664 14421 -4530
rect 14897 -4664 14931 -4530
rect 15005 -4664 15039 -4530
rect 15515 -4664 15549 -4530
rect 14471 -4743 14847 -4709
rect 15089 -4743 15465 -4709
rect 16071 -4485 16447 -4451
rect 16689 -4485 17065 -4451
rect 15987 -4664 16021 -4530
rect 16497 -4664 16531 -4530
rect 16605 -4664 16639 -4530
rect 17115 -4664 17149 -4530
rect 16071 -4743 16447 -4709
rect 16689 -4743 17065 -4709
rect 17671 -4485 18047 -4451
rect 18289 -4485 18665 -4451
rect 17587 -4664 17621 -4530
rect 18097 -4664 18131 -4530
rect 18205 -4664 18239 -4530
rect 18715 -4664 18749 -4530
rect 17671 -4743 18047 -4709
rect 18289 -4743 18665 -4709
rect 19271 -4485 19647 -4451
rect 19889 -4485 20265 -4451
rect 19187 -4664 19221 -4530
rect 19697 -4664 19731 -4530
rect 19805 -4664 19839 -4530
rect 20315 -4664 20349 -4530
rect 19271 -4743 19647 -4709
rect 19889 -4743 20265 -4709
rect 20871 -4485 21247 -4451
rect 21489 -4485 21865 -4451
rect 20787 -4664 20821 -4530
rect 21297 -4664 21331 -4530
rect 21405 -4664 21439 -4530
rect 21915 -4664 21949 -4530
rect 20871 -4743 21247 -4709
rect 21489 -4743 21865 -4709
rect 22471 -4485 22847 -4451
rect 23089 -4485 23465 -4451
rect 22387 -4664 22421 -4530
rect 22897 -4664 22931 -4530
rect 23005 -4664 23039 -4530
rect 23515 -4664 23549 -4530
rect 22471 -4743 22847 -4709
rect 23089 -4743 23465 -4709
rect 24071 -4485 24447 -4451
rect 24689 -4485 25065 -4451
rect 23987 -4664 24021 -4530
rect 24497 -4664 24531 -4530
rect 24605 -4664 24639 -4530
rect 25115 -4664 25149 -4530
rect 24071 -4743 24447 -4709
rect 24689 -4743 25065 -4709
rect 25671 -4485 26047 -4451
rect 26289 -4485 26665 -4451
rect 25587 -4664 25621 -4530
rect 26097 -4664 26131 -4530
rect 26205 -4664 26239 -4530
rect 26715 -4664 26749 -4530
rect 25671 -4743 26047 -4709
rect 26289 -4743 26665 -4709
rect 27271 -4485 27647 -4451
rect 27889 -4485 28265 -4451
rect 27187 -4664 27221 -4530
rect 27697 -4664 27731 -4530
rect 27805 -4664 27839 -4530
rect 28315 -4664 28349 -4530
rect 27271 -4743 27647 -4709
rect 27889 -4743 28265 -4709
rect 28871 -4485 29247 -4451
rect 29489 -4485 29865 -4451
rect 28787 -4664 28821 -4530
rect 29297 -4664 29331 -4530
rect 29405 -4664 29439 -4530
rect 29915 -4664 29949 -4530
rect 28871 -4743 29247 -4709
rect 29489 -4743 29865 -4709
rect 30471 -4485 30847 -4451
rect 31089 -4485 31465 -4451
rect 30387 -4664 30421 -4530
rect 30897 -4664 30931 -4530
rect 31005 -4664 31039 -4530
rect 31515 -4664 31549 -4530
rect 30471 -4743 30847 -4709
rect 31089 -4743 31465 -4709
rect 32071 -4485 32447 -4451
rect 32689 -4485 33065 -4451
rect 31987 -4664 32021 -4530
rect 32497 -4664 32531 -4530
rect 32605 -4664 32639 -4530
rect 33115 -4664 33149 -4530
rect 32071 -4743 32447 -4709
rect 32689 -4743 33065 -4709
rect 33671 -4485 34047 -4451
rect 34289 -4485 34665 -4451
rect 33587 -4664 33621 -4530
rect 34097 -4664 34131 -4530
rect 34205 -4664 34239 -4530
rect 34715 -4664 34749 -4530
rect 33671 -4743 34047 -4709
rect 34289 -4743 34665 -4709
rect 35271 -4485 35647 -4451
rect 35889 -4485 36265 -4451
rect 35187 -4664 35221 -4530
rect 35697 -4664 35731 -4530
rect 35805 -4664 35839 -4530
rect 36315 -4664 36349 -4530
rect 35271 -4743 35647 -4709
rect 35889 -4743 36265 -4709
rect 36871 -4485 37247 -4451
rect 37489 -4485 37865 -4451
rect 36787 -4664 36821 -4530
rect 37297 -4664 37331 -4530
rect 37405 -4664 37439 -4530
rect 37915 -4664 37949 -4530
rect 36871 -4743 37247 -4709
rect 37489 -4743 37865 -4709
rect 69 -8204 445 -8170
rect 705 -8204 1081 -8170
rect -24 -8375 10 -8257
rect 504 -8375 538 -8257
rect 612 -8375 646 -8257
rect 1140 -8375 1174 -8257
rect 69 -8462 445 -8428
rect 705 -8462 1081 -8428
rect 1669 -8204 2045 -8170
rect 2305 -8204 2681 -8170
rect 1576 -8375 1610 -8257
rect 2104 -8375 2138 -8257
rect 2212 -8375 2246 -8257
rect 2740 -8375 2774 -8257
rect 1669 -8462 2045 -8428
rect 2305 -8462 2681 -8428
rect 69 -8730 445 -8696
rect 705 -8730 1081 -8696
rect -24 -9488 10 -8796
rect 504 -9488 538 -8796
rect 612 -9488 646 -8796
rect 1140 -9488 1174 -8796
rect 69 -9588 445 -9554
rect 705 -9588 1081 -9554
rect 1669 -8730 2045 -8696
rect 2305 -8730 2681 -8696
rect 1576 -9488 1610 -8796
rect 2104 -9488 2138 -8796
rect 2212 -9488 2246 -8796
rect 2740 -9488 2774 -8796
rect 1669 -9588 2045 -9554
rect 2305 -9588 2681 -9554
rect 13 -9722 1137 -9688
rect 1613 -9722 2737 -9688
rect 3269 -8204 3645 -8170
rect 3905 -8204 4281 -8170
rect 3176 -8375 3210 -8257
rect 3704 -8375 3738 -8257
rect 3812 -8375 3846 -8257
rect 4340 -8375 4374 -8257
rect 3269 -8462 3645 -8428
rect 3905 -8462 4281 -8428
rect 3269 -8730 3645 -8696
rect 3905 -8730 4281 -8696
rect 3176 -9488 3210 -8796
rect 3704 -9488 3738 -8796
rect 3812 -9488 3846 -8796
rect 4340 -9488 4374 -8796
rect 3269 -9588 3645 -9554
rect 3905 -9588 4281 -9554
rect 3213 -9722 4337 -9688
rect 4869 -8204 5245 -8170
rect 5505 -8204 5881 -8170
rect 4776 -8375 4810 -8257
rect 5304 -8375 5338 -8257
rect 5412 -8375 5446 -8257
rect 5940 -8375 5974 -8257
rect 4869 -8462 5245 -8428
rect 5505 -8462 5881 -8428
rect 4869 -8730 5245 -8696
rect 5505 -8730 5881 -8696
rect 4776 -9488 4810 -8796
rect 5304 -9488 5338 -8796
rect 5412 -9488 5446 -8796
rect 5940 -9488 5974 -8796
rect 4869 -9588 5245 -9554
rect 5505 -9588 5881 -9554
rect 4813 -9722 5937 -9688
rect 6469 -8204 6845 -8170
rect 7105 -8204 7481 -8170
rect 6376 -8375 6410 -8257
rect 6904 -8375 6938 -8257
rect 7012 -8375 7046 -8257
rect 7540 -8375 7574 -8257
rect 6469 -8462 6845 -8428
rect 7105 -8462 7481 -8428
rect 6469 -8730 6845 -8696
rect 7105 -8730 7481 -8696
rect 6376 -9488 6410 -8796
rect 6904 -9488 6938 -8796
rect 7012 -9488 7046 -8796
rect 7540 -9488 7574 -8796
rect 6469 -9588 6845 -9554
rect 7105 -9588 7481 -9554
rect 6413 -9722 7537 -9688
rect 8069 -8204 8445 -8170
rect 8705 -8204 9081 -8170
rect 7976 -8375 8010 -8257
rect 8504 -8375 8538 -8257
rect 8612 -8375 8646 -8257
rect 9140 -8375 9174 -8257
rect 8069 -8462 8445 -8428
rect 8705 -8462 9081 -8428
rect 8069 -8730 8445 -8696
rect 8705 -8730 9081 -8696
rect 7976 -9488 8010 -8796
rect 8504 -9488 8538 -8796
rect 8612 -9488 8646 -8796
rect 9140 -9488 9174 -8796
rect 8069 -9588 8445 -9554
rect 8705 -9588 9081 -9554
rect 8013 -9722 9137 -9688
rect 9669 -8204 10045 -8170
rect 10305 -8204 10681 -8170
rect 9576 -8375 9610 -8257
rect 10104 -8375 10138 -8257
rect 10212 -8375 10246 -8257
rect 10740 -8375 10774 -8257
rect 9669 -8462 10045 -8428
rect 10305 -8462 10681 -8428
rect 9669 -8730 10045 -8696
rect 10305 -8730 10681 -8696
rect 9576 -9488 9610 -8796
rect 10104 -9488 10138 -8796
rect 10212 -9488 10246 -8796
rect 10740 -9488 10774 -8796
rect 9669 -9588 10045 -9554
rect 10305 -9588 10681 -9554
rect 9613 -9722 10737 -9688
rect 11269 -8204 11645 -8170
rect 11905 -8204 12281 -8170
rect 11176 -8375 11210 -8257
rect 11704 -8375 11738 -8257
rect 11812 -8375 11846 -8257
rect 12340 -8375 12374 -8257
rect 11269 -8462 11645 -8428
rect 11905 -8462 12281 -8428
rect 11269 -8730 11645 -8696
rect 11905 -8730 12281 -8696
rect 11176 -9488 11210 -8796
rect 11704 -9488 11738 -8796
rect 11812 -9488 11846 -8796
rect 12340 -9488 12374 -8796
rect 11269 -9588 11645 -9554
rect 11905 -9588 12281 -9554
rect 11213 -9722 12337 -9688
rect 12869 -8204 13245 -8170
rect 13505 -8204 13881 -8170
rect 12776 -8375 12810 -8257
rect 13304 -8375 13338 -8257
rect 13412 -8375 13446 -8257
rect 13940 -8375 13974 -8257
rect 12869 -8462 13245 -8428
rect 13505 -8462 13881 -8428
rect 12869 -8730 13245 -8696
rect 13505 -8730 13881 -8696
rect 12776 -9488 12810 -8796
rect 13304 -9488 13338 -8796
rect 13412 -9488 13446 -8796
rect 13940 -9488 13974 -8796
rect 12869 -9588 13245 -9554
rect 13505 -9588 13881 -9554
rect 12813 -9722 13937 -9688
rect 14469 -8204 14845 -8170
rect 15105 -8204 15481 -8170
rect 14376 -8375 14410 -8257
rect 14904 -8375 14938 -8257
rect 15012 -8375 15046 -8257
rect 15540 -8375 15574 -8257
rect 14469 -8462 14845 -8428
rect 15105 -8462 15481 -8428
rect 14469 -8730 14845 -8696
rect 15105 -8730 15481 -8696
rect 14376 -9488 14410 -8796
rect 14904 -9488 14938 -8796
rect 15012 -9488 15046 -8796
rect 15540 -9488 15574 -8796
rect 14469 -9588 14845 -9554
rect 15105 -9588 15481 -9554
rect 14413 -9722 15537 -9688
rect 16069 -8204 16445 -8170
rect 16705 -8204 17081 -8170
rect 15976 -8375 16010 -8257
rect 16504 -8375 16538 -8257
rect 16612 -8375 16646 -8257
rect 17140 -8375 17174 -8257
rect 16069 -8462 16445 -8428
rect 16705 -8462 17081 -8428
rect 16069 -8730 16445 -8696
rect 16705 -8730 17081 -8696
rect 15976 -9488 16010 -8796
rect 16504 -9488 16538 -8796
rect 16612 -9488 16646 -8796
rect 17140 -9488 17174 -8796
rect 16069 -9588 16445 -9554
rect 16705 -9588 17081 -9554
rect 16013 -9722 17137 -9688
rect 17669 -8204 18045 -8170
rect 18305 -8204 18681 -8170
rect 17576 -8375 17610 -8257
rect 18104 -8375 18138 -8257
rect 18212 -8375 18246 -8257
rect 18740 -8375 18774 -8257
rect 17669 -8462 18045 -8428
rect 18305 -8462 18681 -8428
rect 17669 -8730 18045 -8696
rect 18305 -8730 18681 -8696
rect 17576 -9488 17610 -8796
rect 18104 -9488 18138 -8796
rect 18212 -9488 18246 -8796
rect 18740 -9488 18774 -8796
rect 17669 -9588 18045 -9554
rect 18305 -9588 18681 -9554
rect 17613 -9722 18737 -9688
rect 19269 -8204 19645 -8170
rect 19905 -8204 20281 -8170
rect 19176 -8375 19210 -8257
rect 19704 -8375 19738 -8257
rect 19812 -8375 19846 -8257
rect 20340 -8375 20374 -8257
rect 19269 -8462 19645 -8428
rect 19905 -8462 20281 -8428
rect 19269 -8730 19645 -8696
rect 19905 -8730 20281 -8696
rect 19176 -9488 19210 -8796
rect 19704 -9488 19738 -8796
rect 19812 -9488 19846 -8796
rect 20340 -9488 20374 -8796
rect 19269 -9588 19645 -9554
rect 19905 -9588 20281 -9554
rect 19213 -9722 20337 -9688
rect 20869 -8204 21245 -8170
rect 21505 -8204 21881 -8170
rect 20776 -8375 20810 -8257
rect 21304 -8375 21338 -8257
rect 21412 -8375 21446 -8257
rect 21940 -8375 21974 -8257
rect 20869 -8462 21245 -8428
rect 21505 -8462 21881 -8428
rect 20869 -8730 21245 -8696
rect 21505 -8730 21881 -8696
rect 20776 -9488 20810 -8796
rect 21304 -9488 21338 -8796
rect 21412 -9488 21446 -8796
rect 21940 -9488 21974 -8796
rect 20869 -9588 21245 -9554
rect 21505 -9588 21881 -9554
rect 20813 -9722 21937 -9688
rect 22469 -8204 22845 -8170
rect 23105 -8204 23481 -8170
rect 22376 -8375 22410 -8257
rect 22904 -8375 22938 -8257
rect 23012 -8375 23046 -8257
rect 23540 -8375 23574 -8257
rect 22469 -8462 22845 -8428
rect 23105 -8462 23481 -8428
rect 22469 -8730 22845 -8696
rect 23105 -8730 23481 -8696
rect 22376 -9488 22410 -8796
rect 22904 -9488 22938 -8796
rect 23012 -9488 23046 -8796
rect 23540 -9488 23574 -8796
rect 22469 -9588 22845 -9554
rect 23105 -9588 23481 -9554
rect 22413 -9722 23537 -9688
rect 24069 -8204 24445 -8170
rect 24705 -8204 25081 -8170
rect 23976 -8375 24010 -8257
rect 24504 -8375 24538 -8257
rect 24612 -8375 24646 -8257
rect 25140 -8375 25174 -8257
rect 24069 -8462 24445 -8428
rect 24705 -8462 25081 -8428
rect 24069 -8730 24445 -8696
rect 24705 -8730 25081 -8696
rect 23976 -9488 24010 -8796
rect 24504 -9488 24538 -8796
rect 24612 -9488 24646 -8796
rect 25140 -9488 25174 -8796
rect 24069 -9588 24445 -9554
rect 24705 -9588 25081 -9554
rect 24013 -9722 25137 -9688
rect 25669 -8204 26045 -8170
rect 26305 -8204 26681 -8170
rect 25576 -8375 25610 -8257
rect 26104 -8375 26138 -8257
rect 26212 -8375 26246 -8257
rect 26740 -8375 26774 -8257
rect 25669 -8462 26045 -8428
rect 26305 -8462 26681 -8428
rect 25669 -8730 26045 -8696
rect 26305 -8730 26681 -8696
rect 25576 -9488 25610 -8796
rect 26104 -9488 26138 -8796
rect 26212 -9488 26246 -8796
rect 26740 -9488 26774 -8796
rect 25669 -9588 26045 -9554
rect 26305 -9588 26681 -9554
rect 25613 -9722 26737 -9688
rect 27269 -8204 27645 -8170
rect 27905 -8204 28281 -8170
rect 27176 -8375 27210 -8257
rect 27704 -8375 27738 -8257
rect 27812 -8375 27846 -8257
rect 28340 -8375 28374 -8257
rect 27269 -8462 27645 -8428
rect 27905 -8462 28281 -8428
rect 27269 -8730 27645 -8696
rect 27905 -8730 28281 -8696
rect 27176 -9488 27210 -8796
rect 27704 -9488 27738 -8796
rect 27812 -9488 27846 -8796
rect 28340 -9488 28374 -8796
rect 27269 -9588 27645 -9554
rect 27905 -9588 28281 -9554
rect 27213 -9722 28337 -9688
rect 28869 -8204 29245 -8170
rect 29505 -8204 29881 -8170
rect 28776 -8375 28810 -8257
rect 29304 -8375 29338 -8257
rect 29412 -8375 29446 -8257
rect 29940 -8375 29974 -8257
rect 28869 -8462 29245 -8428
rect 29505 -8462 29881 -8428
rect 28869 -8730 29245 -8696
rect 29505 -8730 29881 -8696
rect 28776 -9488 28810 -8796
rect 29304 -9488 29338 -8796
rect 29412 -9488 29446 -8796
rect 29940 -9488 29974 -8796
rect 28869 -9588 29245 -9554
rect 29505 -9588 29881 -9554
rect 28813 -9722 29937 -9688
rect 30469 -8204 30845 -8170
rect 31105 -8204 31481 -8170
rect 30376 -8375 30410 -8257
rect 30904 -8375 30938 -8257
rect 31012 -8375 31046 -8257
rect 31540 -8375 31574 -8257
rect 30469 -8462 30845 -8428
rect 31105 -8462 31481 -8428
rect 30469 -8730 30845 -8696
rect 31105 -8730 31481 -8696
rect 30376 -9488 30410 -8796
rect 30904 -9488 30938 -8796
rect 31012 -9488 31046 -8796
rect 31540 -9488 31574 -8796
rect 30469 -9588 30845 -9554
rect 31105 -9588 31481 -9554
rect 30413 -9722 31537 -9688
rect 32069 -8204 32445 -8170
rect 32705 -8204 33081 -8170
rect 31976 -8375 32010 -8257
rect 32504 -8375 32538 -8257
rect 32612 -8375 32646 -8257
rect 33140 -8375 33174 -8257
rect 32069 -8462 32445 -8428
rect 32705 -8462 33081 -8428
rect 32069 -8730 32445 -8696
rect 32705 -8730 33081 -8696
rect 31976 -9488 32010 -8796
rect 32504 -9488 32538 -8796
rect 32612 -9488 32646 -8796
rect 33140 -9488 33174 -8796
rect 32069 -9588 32445 -9554
rect 32705 -9588 33081 -9554
rect 32013 -9722 33137 -9688
rect 33669 -8204 34045 -8170
rect 34305 -8204 34681 -8170
rect 33576 -8375 33610 -8257
rect 34104 -8375 34138 -8257
rect 34212 -8375 34246 -8257
rect 34740 -8375 34774 -8257
rect 33669 -8462 34045 -8428
rect 34305 -8462 34681 -8428
rect 33669 -8730 34045 -8696
rect 34305 -8730 34681 -8696
rect 33576 -9488 33610 -8796
rect 34104 -9488 34138 -8796
rect 34212 -9488 34246 -8796
rect 34740 -9488 34774 -8796
rect 33669 -9588 34045 -9554
rect 34305 -9588 34681 -9554
rect 33613 -9722 34737 -9688
rect 35269 -8204 35645 -8170
rect 35905 -8204 36281 -8170
rect 35176 -8375 35210 -8257
rect 35704 -8375 35738 -8257
rect 35812 -8375 35846 -8257
rect 36340 -8375 36374 -8257
rect 35269 -8462 35645 -8428
rect 35905 -8462 36281 -8428
rect 36869 -8204 37245 -8170
rect 37505 -8204 37881 -8170
rect 36776 -8375 36810 -8257
rect 37304 -8375 37338 -8257
rect 37412 -8375 37446 -8257
rect 37940 -8375 37974 -8257
rect 36869 -8462 37245 -8428
rect 37505 -8462 37881 -8428
rect 35269 -8730 35645 -8696
rect 35905 -8730 36281 -8696
rect 35176 -9488 35210 -8796
rect 35704 -9488 35738 -8796
rect 35812 -9488 35846 -8796
rect 36340 -9488 36374 -8796
rect 35269 -9588 35645 -9554
rect 35905 -9588 36281 -9554
rect 36869 -8730 37245 -8696
rect 37505 -8730 37881 -8696
rect 36776 -9488 36810 -8796
rect 37304 -9488 37338 -8796
rect 37412 -9488 37446 -8796
rect 37940 -9488 37974 -8796
rect 36869 -9588 37245 -9554
rect 37505 -9588 37881 -9554
rect 35213 -9722 36337 -9688
rect 36813 -9722 37937 -9688
rect 69 -10004 445 -9970
rect 705 -10004 1081 -9970
rect -24 -10175 10 -10057
rect 504 -10175 538 -10057
rect 612 -10175 646 -10057
rect 1140 -10175 1174 -10057
rect 69 -10262 445 -10228
rect 705 -10262 1081 -10228
rect 1669 -10004 2045 -9970
rect 2305 -10004 2681 -9970
rect 1576 -10175 1610 -10057
rect 2104 -10175 2138 -10057
rect 2212 -10175 2246 -10057
rect 2740 -10175 2774 -10057
rect 1669 -10262 2045 -10228
rect 2305 -10262 2681 -10228
rect 69 -10530 445 -10496
rect 705 -10530 1081 -10496
rect -24 -11288 10 -10596
rect 504 -11288 538 -10596
rect 612 -11288 646 -10596
rect 1140 -11288 1174 -10596
rect 69 -11388 445 -11354
rect 705 -11388 1081 -11354
rect 1669 -10530 2045 -10496
rect 2305 -10530 2681 -10496
rect 1576 -11288 1610 -10596
rect 2104 -11288 2138 -10596
rect 2212 -11288 2246 -10596
rect 2740 -11288 2774 -10596
rect 1669 -11388 2045 -11354
rect 2305 -11388 2681 -11354
rect 13 -11522 1137 -11488
rect 1613 -11522 2737 -11488
rect 3269 -10004 3645 -9970
rect 3905 -10004 4281 -9970
rect 3176 -10175 3210 -10057
rect 3704 -10175 3738 -10057
rect 3812 -10175 3846 -10057
rect 4340 -10175 4374 -10057
rect 3269 -10262 3645 -10228
rect 3905 -10262 4281 -10228
rect 3269 -10530 3645 -10496
rect 3905 -10530 4281 -10496
rect 3176 -11288 3210 -10596
rect 3704 -11288 3738 -10596
rect 3812 -11288 3846 -10596
rect 4340 -11288 4374 -10596
rect 3269 -11388 3645 -11354
rect 3905 -11388 4281 -11354
rect 3213 -11522 4337 -11488
rect 4869 -10004 5245 -9970
rect 5505 -10004 5881 -9970
rect 4776 -10175 4810 -10057
rect 5304 -10175 5338 -10057
rect 5412 -10175 5446 -10057
rect 5940 -10175 5974 -10057
rect 4869 -10262 5245 -10228
rect 5505 -10262 5881 -10228
rect 4869 -10530 5245 -10496
rect 5505 -10530 5881 -10496
rect 4776 -11288 4810 -10596
rect 5304 -11288 5338 -10596
rect 5412 -11288 5446 -10596
rect 5940 -11288 5974 -10596
rect 4869 -11388 5245 -11354
rect 5505 -11388 5881 -11354
rect 4813 -11522 5937 -11488
rect 6469 -10004 6845 -9970
rect 7105 -10004 7481 -9970
rect 6376 -10175 6410 -10057
rect 6904 -10175 6938 -10057
rect 7012 -10175 7046 -10057
rect 7540 -10175 7574 -10057
rect 6469 -10262 6845 -10228
rect 7105 -10262 7481 -10228
rect 6469 -10530 6845 -10496
rect 7105 -10530 7481 -10496
rect 6376 -11288 6410 -10596
rect 6904 -11288 6938 -10596
rect 7012 -11288 7046 -10596
rect 7540 -11288 7574 -10596
rect 6469 -11388 6845 -11354
rect 7105 -11388 7481 -11354
rect 6413 -11522 7537 -11488
rect 8069 -10004 8445 -9970
rect 8705 -10004 9081 -9970
rect 7976 -10175 8010 -10057
rect 8504 -10175 8538 -10057
rect 8612 -10175 8646 -10057
rect 9140 -10175 9174 -10057
rect 8069 -10262 8445 -10228
rect 8705 -10262 9081 -10228
rect 8069 -10530 8445 -10496
rect 8705 -10530 9081 -10496
rect 7976 -11288 8010 -10596
rect 8504 -11288 8538 -10596
rect 8612 -11288 8646 -10596
rect 9140 -11288 9174 -10596
rect 8069 -11388 8445 -11354
rect 8705 -11388 9081 -11354
rect 8013 -11522 9137 -11488
rect 9669 -10004 10045 -9970
rect 10305 -10004 10681 -9970
rect 9576 -10175 9610 -10057
rect 10104 -10175 10138 -10057
rect 10212 -10175 10246 -10057
rect 10740 -10175 10774 -10057
rect 9669 -10262 10045 -10228
rect 10305 -10262 10681 -10228
rect 9669 -10530 10045 -10496
rect 10305 -10530 10681 -10496
rect 9576 -11288 9610 -10596
rect 10104 -11288 10138 -10596
rect 10212 -11288 10246 -10596
rect 10740 -11288 10774 -10596
rect 9669 -11388 10045 -11354
rect 10305 -11388 10681 -11354
rect 9613 -11522 10737 -11488
rect 11269 -10004 11645 -9970
rect 11905 -10004 12281 -9970
rect 11176 -10175 11210 -10057
rect 11704 -10175 11738 -10057
rect 11812 -10175 11846 -10057
rect 12340 -10175 12374 -10057
rect 11269 -10262 11645 -10228
rect 11905 -10262 12281 -10228
rect 11269 -10530 11645 -10496
rect 11905 -10530 12281 -10496
rect 11176 -11288 11210 -10596
rect 11704 -11288 11738 -10596
rect 11812 -11288 11846 -10596
rect 12340 -11288 12374 -10596
rect 11269 -11388 11645 -11354
rect 11905 -11388 12281 -11354
rect 11213 -11522 12337 -11488
rect 12869 -10004 13245 -9970
rect 13505 -10004 13881 -9970
rect 12776 -10175 12810 -10057
rect 13304 -10175 13338 -10057
rect 13412 -10175 13446 -10057
rect 13940 -10175 13974 -10057
rect 12869 -10262 13245 -10228
rect 13505 -10262 13881 -10228
rect 12869 -10530 13245 -10496
rect 13505 -10530 13881 -10496
rect 12776 -11288 12810 -10596
rect 13304 -11288 13338 -10596
rect 13412 -11288 13446 -10596
rect 13940 -11288 13974 -10596
rect 12869 -11388 13245 -11354
rect 13505 -11388 13881 -11354
rect 12813 -11522 13937 -11488
rect 14469 -10004 14845 -9970
rect 15105 -10004 15481 -9970
rect 14376 -10175 14410 -10057
rect 14904 -10175 14938 -10057
rect 15012 -10175 15046 -10057
rect 15540 -10175 15574 -10057
rect 14469 -10262 14845 -10228
rect 15105 -10262 15481 -10228
rect 14469 -10530 14845 -10496
rect 15105 -10530 15481 -10496
rect 14376 -11288 14410 -10596
rect 14904 -11288 14938 -10596
rect 15012 -11288 15046 -10596
rect 15540 -11288 15574 -10596
rect 14469 -11388 14845 -11354
rect 15105 -11388 15481 -11354
rect 14413 -11522 15537 -11488
rect 16069 -10004 16445 -9970
rect 16705 -10004 17081 -9970
rect 15976 -10175 16010 -10057
rect 16504 -10175 16538 -10057
rect 16612 -10175 16646 -10057
rect 17140 -10175 17174 -10057
rect 16069 -10262 16445 -10228
rect 16705 -10262 17081 -10228
rect 16069 -10530 16445 -10496
rect 16705 -10530 17081 -10496
rect 15976 -11288 16010 -10596
rect 16504 -11288 16538 -10596
rect 16612 -11288 16646 -10596
rect 17140 -11288 17174 -10596
rect 16069 -11388 16445 -11354
rect 16705 -11388 17081 -11354
rect 16013 -11522 17137 -11488
rect 17669 -10004 18045 -9970
rect 18305 -10004 18681 -9970
rect 17576 -10175 17610 -10057
rect 18104 -10175 18138 -10057
rect 18212 -10175 18246 -10057
rect 18740 -10175 18774 -10057
rect 17669 -10262 18045 -10228
rect 18305 -10262 18681 -10228
rect 17669 -10530 18045 -10496
rect 18305 -10530 18681 -10496
rect 17576 -11288 17610 -10596
rect 18104 -11288 18138 -10596
rect 18212 -11288 18246 -10596
rect 18740 -11288 18774 -10596
rect 17669 -11388 18045 -11354
rect 18305 -11388 18681 -11354
rect 17613 -11522 18737 -11488
rect 19269 -10004 19645 -9970
rect 19905 -10004 20281 -9970
rect 19176 -10175 19210 -10057
rect 19704 -10175 19738 -10057
rect 19812 -10175 19846 -10057
rect 20340 -10175 20374 -10057
rect 19269 -10262 19645 -10228
rect 19905 -10262 20281 -10228
rect 19269 -10530 19645 -10496
rect 19905 -10530 20281 -10496
rect 19176 -11288 19210 -10596
rect 19704 -11288 19738 -10596
rect 19812 -11288 19846 -10596
rect 20340 -11288 20374 -10596
rect 19269 -11388 19645 -11354
rect 19905 -11388 20281 -11354
rect 19213 -11522 20337 -11488
rect 20869 -10004 21245 -9970
rect 21505 -10004 21881 -9970
rect 20776 -10175 20810 -10057
rect 21304 -10175 21338 -10057
rect 21412 -10175 21446 -10057
rect 21940 -10175 21974 -10057
rect 20869 -10262 21245 -10228
rect 21505 -10262 21881 -10228
rect 20869 -10530 21245 -10496
rect 21505 -10530 21881 -10496
rect 20776 -11288 20810 -10596
rect 21304 -11288 21338 -10596
rect 21412 -11288 21446 -10596
rect 21940 -11288 21974 -10596
rect 20869 -11388 21245 -11354
rect 21505 -11388 21881 -11354
rect 20813 -11522 21937 -11488
rect 22469 -10004 22845 -9970
rect 23105 -10004 23481 -9970
rect 22376 -10175 22410 -10057
rect 22904 -10175 22938 -10057
rect 23012 -10175 23046 -10057
rect 23540 -10175 23574 -10057
rect 22469 -10262 22845 -10228
rect 23105 -10262 23481 -10228
rect 22469 -10530 22845 -10496
rect 23105 -10530 23481 -10496
rect 22376 -11288 22410 -10596
rect 22904 -11288 22938 -10596
rect 23012 -11288 23046 -10596
rect 23540 -11288 23574 -10596
rect 22469 -11388 22845 -11354
rect 23105 -11388 23481 -11354
rect 22413 -11522 23537 -11488
rect 24069 -10004 24445 -9970
rect 24705 -10004 25081 -9970
rect 23976 -10175 24010 -10057
rect 24504 -10175 24538 -10057
rect 24612 -10175 24646 -10057
rect 25140 -10175 25174 -10057
rect 24069 -10262 24445 -10228
rect 24705 -10262 25081 -10228
rect 24069 -10530 24445 -10496
rect 24705 -10530 25081 -10496
rect 23976 -11288 24010 -10596
rect 24504 -11288 24538 -10596
rect 24612 -11288 24646 -10596
rect 25140 -11288 25174 -10596
rect 24069 -11388 24445 -11354
rect 24705 -11388 25081 -11354
rect 24013 -11522 25137 -11488
rect 25669 -10004 26045 -9970
rect 26305 -10004 26681 -9970
rect 25576 -10175 25610 -10057
rect 26104 -10175 26138 -10057
rect 26212 -10175 26246 -10057
rect 26740 -10175 26774 -10057
rect 25669 -10262 26045 -10228
rect 26305 -10262 26681 -10228
rect 25669 -10530 26045 -10496
rect 26305 -10530 26681 -10496
rect 25576 -11288 25610 -10596
rect 26104 -11288 26138 -10596
rect 26212 -11288 26246 -10596
rect 26740 -11288 26774 -10596
rect 25669 -11388 26045 -11354
rect 26305 -11388 26681 -11354
rect 25613 -11522 26737 -11488
rect 27269 -10004 27645 -9970
rect 27905 -10004 28281 -9970
rect 27176 -10175 27210 -10057
rect 27704 -10175 27738 -10057
rect 27812 -10175 27846 -10057
rect 28340 -10175 28374 -10057
rect 27269 -10262 27645 -10228
rect 27905 -10262 28281 -10228
rect 27269 -10530 27645 -10496
rect 27905 -10530 28281 -10496
rect 27176 -11288 27210 -10596
rect 27704 -11288 27738 -10596
rect 27812 -11288 27846 -10596
rect 28340 -11288 28374 -10596
rect 27269 -11388 27645 -11354
rect 27905 -11388 28281 -11354
rect 27213 -11522 28337 -11488
rect 28869 -10004 29245 -9970
rect 29505 -10004 29881 -9970
rect 28776 -10175 28810 -10057
rect 29304 -10175 29338 -10057
rect 29412 -10175 29446 -10057
rect 29940 -10175 29974 -10057
rect 28869 -10262 29245 -10228
rect 29505 -10262 29881 -10228
rect 28869 -10530 29245 -10496
rect 29505 -10530 29881 -10496
rect 28776 -11288 28810 -10596
rect 29304 -11288 29338 -10596
rect 29412 -11288 29446 -10596
rect 29940 -11288 29974 -10596
rect 28869 -11388 29245 -11354
rect 29505 -11388 29881 -11354
rect 28813 -11522 29937 -11488
rect 30469 -10004 30845 -9970
rect 31105 -10004 31481 -9970
rect 30376 -10175 30410 -10057
rect 30904 -10175 30938 -10057
rect 31012 -10175 31046 -10057
rect 31540 -10175 31574 -10057
rect 30469 -10262 30845 -10228
rect 31105 -10262 31481 -10228
rect 30469 -10530 30845 -10496
rect 31105 -10530 31481 -10496
rect 30376 -11288 30410 -10596
rect 30904 -11288 30938 -10596
rect 31012 -11288 31046 -10596
rect 31540 -11288 31574 -10596
rect 30469 -11388 30845 -11354
rect 31105 -11388 31481 -11354
rect 30413 -11522 31537 -11488
rect 32069 -10004 32445 -9970
rect 32705 -10004 33081 -9970
rect 31976 -10175 32010 -10057
rect 32504 -10175 32538 -10057
rect 32612 -10175 32646 -10057
rect 33140 -10175 33174 -10057
rect 32069 -10262 32445 -10228
rect 32705 -10262 33081 -10228
rect 32069 -10530 32445 -10496
rect 32705 -10530 33081 -10496
rect 31976 -11288 32010 -10596
rect 32504 -11288 32538 -10596
rect 32612 -11288 32646 -10596
rect 33140 -11288 33174 -10596
rect 32069 -11388 32445 -11354
rect 32705 -11388 33081 -11354
rect 32013 -11522 33137 -11488
rect 33669 -10004 34045 -9970
rect 34305 -10004 34681 -9970
rect 33576 -10175 33610 -10057
rect 34104 -10175 34138 -10057
rect 34212 -10175 34246 -10057
rect 34740 -10175 34774 -10057
rect 33669 -10262 34045 -10228
rect 34305 -10262 34681 -10228
rect 33669 -10530 34045 -10496
rect 34305 -10530 34681 -10496
rect 33576 -11288 33610 -10596
rect 34104 -11288 34138 -10596
rect 34212 -11288 34246 -10596
rect 34740 -11288 34774 -10596
rect 33669 -11388 34045 -11354
rect 34305 -11388 34681 -11354
rect 33613 -11522 34737 -11488
rect 35269 -10004 35645 -9970
rect 35905 -10004 36281 -9970
rect 35176 -10175 35210 -10057
rect 35704 -10175 35738 -10057
rect 35812 -10175 35846 -10057
rect 36340 -10175 36374 -10057
rect 35269 -10262 35645 -10228
rect 35905 -10262 36281 -10228
rect 36869 -10004 37245 -9970
rect 37505 -10004 37881 -9970
rect 36776 -10175 36810 -10057
rect 37304 -10175 37338 -10057
rect 37412 -10175 37446 -10057
rect 37940 -10175 37974 -10057
rect 36869 -10262 37245 -10228
rect 37505 -10262 37881 -10228
rect 35269 -10530 35645 -10496
rect 35905 -10530 36281 -10496
rect 35176 -11288 35210 -10596
rect 35704 -11288 35738 -10596
rect 35812 -11288 35846 -10596
rect 36340 -11288 36374 -10596
rect 35269 -11388 35645 -11354
rect 35905 -11388 36281 -11354
rect 36869 -10530 37245 -10496
rect 37505 -10530 37881 -10496
rect 36776 -11288 36810 -10596
rect 37304 -11288 37338 -10596
rect 37412 -11288 37446 -10596
rect 37940 -11288 37974 -10596
rect 36869 -11388 37245 -11354
rect 37505 -11388 37881 -11354
rect 35213 -11522 36337 -11488
rect 36813 -11522 37937 -11488
rect 69 -11804 445 -11770
rect 705 -11804 1081 -11770
rect -24 -11975 10 -11857
rect 504 -11975 538 -11857
rect 612 -11975 646 -11857
rect 1140 -11975 1174 -11857
rect 69 -12062 445 -12028
rect 705 -12062 1081 -12028
rect 1669 -11804 2045 -11770
rect 2305 -11804 2681 -11770
rect 1576 -11975 1610 -11857
rect 2104 -11975 2138 -11857
rect 2212 -11975 2246 -11857
rect 2740 -11975 2774 -11857
rect 1669 -12062 2045 -12028
rect 2305 -12062 2681 -12028
rect 69 -12330 445 -12296
rect 705 -12330 1081 -12296
rect -24 -13088 10 -12396
rect 504 -13088 538 -12396
rect 612 -13088 646 -12396
rect 1140 -13088 1174 -12396
rect 69 -13188 445 -13154
rect 705 -13188 1081 -13154
rect 1669 -12330 2045 -12296
rect 2305 -12330 2681 -12296
rect 1576 -13088 1610 -12396
rect 2104 -13088 2138 -12396
rect 2212 -13088 2246 -12396
rect 2740 -13088 2774 -12396
rect 1669 -13188 2045 -13154
rect 2305 -13188 2681 -13154
rect 13 -13322 1137 -13288
rect 1613 -13322 2737 -13288
rect 3269 -11804 3645 -11770
rect 3905 -11804 4281 -11770
rect 3176 -11975 3210 -11857
rect 3704 -11975 3738 -11857
rect 3812 -11975 3846 -11857
rect 4340 -11975 4374 -11857
rect 3269 -12062 3645 -12028
rect 3905 -12062 4281 -12028
rect 3269 -12330 3645 -12296
rect 3905 -12330 4281 -12296
rect 3176 -13088 3210 -12396
rect 3704 -13088 3738 -12396
rect 3812 -13088 3846 -12396
rect 4340 -13088 4374 -12396
rect 3269 -13188 3645 -13154
rect 3905 -13188 4281 -13154
rect 3213 -13322 4337 -13288
rect 4869 -11804 5245 -11770
rect 5505 -11804 5881 -11770
rect 4776 -11975 4810 -11857
rect 5304 -11975 5338 -11857
rect 5412 -11975 5446 -11857
rect 5940 -11975 5974 -11857
rect 4869 -12062 5245 -12028
rect 5505 -12062 5881 -12028
rect 4869 -12330 5245 -12296
rect 5505 -12330 5881 -12296
rect 4776 -13088 4810 -12396
rect 5304 -13088 5338 -12396
rect 5412 -13088 5446 -12396
rect 5940 -13088 5974 -12396
rect 4869 -13188 5245 -13154
rect 5505 -13188 5881 -13154
rect 4813 -13322 5937 -13288
rect 6469 -11804 6845 -11770
rect 7105 -11804 7481 -11770
rect 6376 -11975 6410 -11857
rect 6904 -11975 6938 -11857
rect 7012 -11975 7046 -11857
rect 7540 -11975 7574 -11857
rect 6469 -12062 6845 -12028
rect 7105 -12062 7481 -12028
rect 6469 -12330 6845 -12296
rect 7105 -12330 7481 -12296
rect 6376 -13088 6410 -12396
rect 6904 -13088 6938 -12396
rect 7012 -13088 7046 -12396
rect 7540 -13088 7574 -12396
rect 6469 -13188 6845 -13154
rect 7105 -13188 7481 -13154
rect 6413 -13322 7537 -13288
rect 8069 -11804 8445 -11770
rect 8705 -11804 9081 -11770
rect 7976 -11975 8010 -11857
rect 8504 -11975 8538 -11857
rect 8612 -11975 8646 -11857
rect 9140 -11975 9174 -11857
rect 8069 -12062 8445 -12028
rect 8705 -12062 9081 -12028
rect 8069 -12330 8445 -12296
rect 8705 -12330 9081 -12296
rect 7976 -13088 8010 -12396
rect 8504 -13088 8538 -12396
rect 8612 -13088 8646 -12396
rect 9140 -13088 9174 -12396
rect 8069 -13188 8445 -13154
rect 8705 -13188 9081 -13154
rect 8013 -13322 9137 -13288
rect 9669 -11804 10045 -11770
rect 10305 -11804 10681 -11770
rect 9576 -11975 9610 -11857
rect 10104 -11975 10138 -11857
rect 10212 -11975 10246 -11857
rect 10740 -11975 10774 -11857
rect 9669 -12062 10045 -12028
rect 10305 -12062 10681 -12028
rect 9669 -12330 10045 -12296
rect 10305 -12330 10681 -12296
rect 9576 -13088 9610 -12396
rect 10104 -13088 10138 -12396
rect 10212 -13088 10246 -12396
rect 10740 -13088 10774 -12396
rect 9669 -13188 10045 -13154
rect 10305 -13188 10681 -13154
rect 9613 -13322 10737 -13288
rect 11269 -11804 11645 -11770
rect 11905 -11804 12281 -11770
rect 11176 -11975 11210 -11857
rect 11704 -11975 11738 -11857
rect 11812 -11975 11846 -11857
rect 12340 -11975 12374 -11857
rect 11269 -12062 11645 -12028
rect 11905 -12062 12281 -12028
rect 11269 -12330 11645 -12296
rect 11905 -12330 12281 -12296
rect 11176 -13088 11210 -12396
rect 11704 -13088 11738 -12396
rect 11812 -13088 11846 -12396
rect 12340 -13088 12374 -12396
rect 11269 -13188 11645 -13154
rect 11905 -13188 12281 -13154
rect 11213 -13322 12337 -13288
rect 12869 -11804 13245 -11770
rect 13505 -11804 13881 -11770
rect 12776 -11975 12810 -11857
rect 13304 -11975 13338 -11857
rect 13412 -11975 13446 -11857
rect 13940 -11975 13974 -11857
rect 12869 -12062 13245 -12028
rect 13505 -12062 13881 -12028
rect 12869 -12330 13245 -12296
rect 13505 -12330 13881 -12296
rect 12776 -13088 12810 -12396
rect 13304 -13088 13338 -12396
rect 13412 -13088 13446 -12396
rect 13940 -13088 13974 -12396
rect 12869 -13188 13245 -13154
rect 13505 -13188 13881 -13154
rect 12813 -13322 13937 -13288
rect 14469 -11804 14845 -11770
rect 15105 -11804 15481 -11770
rect 14376 -11975 14410 -11857
rect 14904 -11975 14938 -11857
rect 15012 -11975 15046 -11857
rect 15540 -11975 15574 -11857
rect 14469 -12062 14845 -12028
rect 15105 -12062 15481 -12028
rect 14469 -12330 14845 -12296
rect 15105 -12330 15481 -12296
rect 14376 -13088 14410 -12396
rect 14904 -13088 14938 -12396
rect 15012 -13088 15046 -12396
rect 15540 -13088 15574 -12396
rect 14469 -13188 14845 -13154
rect 15105 -13188 15481 -13154
rect 14413 -13322 15537 -13288
rect 16069 -11804 16445 -11770
rect 16705 -11804 17081 -11770
rect 15976 -11975 16010 -11857
rect 16504 -11975 16538 -11857
rect 16612 -11975 16646 -11857
rect 17140 -11975 17174 -11857
rect 16069 -12062 16445 -12028
rect 16705 -12062 17081 -12028
rect 16069 -12330 16445 -12296
rect 16705 -12330 17081 -12296
rect 15976 -13088 16010 -12396
rect 16504 -13088 16538 -12396
rect 16612 -13088 16646 -12396
rect 17140 -13088 17174 -12396
rect 16069 -13188 16445 -13154
rect 16705 -13188 17081 -13154
rect 16013 -13322 17137 -13288
rect 17669 -11804 18045 -11770
rect 18305 -11804 18681 -11770
rect 17576 -11975 17610 -11857
rect 18104 -11975 18138 -11857
rect 18212 -11975 18246 -11857
rect 18740 -11975 18774 -11857
rect 17669 -12062 18045 -12028
rect 18305 -12062 18681 -12028
rect 17669 -12330 18045 -12296
rect 18305 -12330 18681 -12296
rect 17576 -13088 17610 -12396
rect 18104 -13088 18138 -12396
rect 18212 -13088 18246 -12396
rect 18740 -13088 18774 -12396
rect 17669 -13188 18045 -13154
rect 18305 -13188 18681 -13154
rect 17613 -13322 18737 -13288
rect 19269 -11804 19645 -11770
rect 19905 -11804 20281 -11770
rect 19176 -11975 19210 -11857
rect 19704 -11975 19738 -11857
rect 19812 -11975 19846 -11857
rect 20340 -11975 20374 -11857
rect 19269 -12062 19645 -12028
rect 19905 -12062 20281 -12028
rect 19269 -12330 19645 -12296
rect 19905 -12330 20281 -12296
rect 19176 -13088 19210 -12396
rect 19704 -13088 19738 -12396
rect 19812 -13088 19846 -12396
rect 20340 -13088 20374 -12396
rect 19269 -13188 19645 -13154
rect 19905 -13188 20281 -13154
rect 19213 -13322 20337 -13288
rect 20869 -11804 21245 -11770
rect 21505 -11804 21881 -11770
rect 20776 -11975 20810 -11857
rect 21304 -11975 21338 -11857
rect 21412 -11975 21446 -11857
rect 21940 -11975 21974 -11857
rect 20869 -12062 21245 -12028
rect 21505 -12062 21881 -12028
rect 20869 -12330 21245 -12296
rect 21505 -12330 21881 -12296
rect 20776 -13088 20810 -12396
rect 21304 -13088 21338 -12396
rect 21412 -13088 21446 -12396
rect 21940 -13088 21974 -12396
rect 20869 -13188 21245 -13154
rect 21505 -13188 21881 -13154
rect 20813 -13322 21937 -13288
rect 22469 -11804 22845 -11770
rect 23105 -11804 23481 -11770
rect 22376 -11975 22410 -11857
rect 22904 -11975 22938 -11857
rect 23012 -11975 23046 -11857
rect 23540 -11975 23574 -11857
rect 22469 -12062 22845 -12028
rect 23105 -12062 23481 -12028
rect 22469 -12330 22845 -12296
rect 23105 -12330 23481 -12296
rect 22376 -13088 22410 -12396
rect 22904 -13088 22938 -12396
rect 23012 -13088 23046 -12396
rect 23540 -13088 23574 -12396
rect 22469 -13188 22845 -13154
rect 23105 -13188 23481 -13154
rect 22413 -13322 23537 -13288
rect 24069 -11804 24445 -11770
rect 24705 -11804 25081 -11770
rect 23976 -11975 24010 -11857
rect 24504 -11975 24538 -11857
rect 24612 -11975 24646 -11857
rect 25140 -11975 25174 -11857
rect 24069 -12062 24445 -12028
rect 24705 -12062 25081 -12028
rect 24069 -12330 24445 -12296
rect 24705 -12330 25081 -12296
rect 23976 -13088 24010 -12396
rect 24504 -13088 24538 -12396
rect 24612 -13088 24646 -12396
rect 25140 -13088 25174 -12396
rect 24069 -13188 24445 -13154
rect 24705 -13188 25081 -13154
rect 24013 -13322 25137 -13288
rect 25669 -11804 26045 -11770
rect 26305 -11804 26681 -11770
rect 25576 -11975 25610 -11857
rect 26104 -11975 26138 -11857
rect 26212 -11975 26246 -11857
rect 26740 -11975 26774 -11857
rect 25669 -12062 26045 -12028
rect 26305 -12062 26681 -12028
rect 25669 -12330 26045 -12296
rect 26305 -12330 26681 -12296
rect 25576 -13088 25610 -12396
rect 26104 -13088 26138 -12396
rect 26212 -13088 26246 -12396
rect 26740 -13088 26774 -12396
rect 25669 -13188 26045 -13154
rect 26305 -13188 26681 -13154
rect 25613 -13322 26737 -13288
rect 27269 -11804 27645 -11770
rect 27905 -11804 28281 -11770
rect 27176 -11975 27210 -11857
rect 27704 -11975 27738 -11857
rect 27812 -11975 27846 -11857
rect 28340 -11975 28374 -11857
rect 27269 -12062 27645 -12028
rect 27905 -12062 28281 -12028
rect 27269 -12330 27645 -12296
rect 27905 -12330 28281 -12296
rect 27176 -13088 27210 -12396
rect 27704 -13088 27738 -12396
rect 27812 -13088 27846 -12396
rect 28340 -13088 28374 -12396
rect 27269 -13188 27645 -13154
rect 27905 -13188 28281 -13154
rect 27213 -13322 28337 -13288
rect 28869 -11804 29245 -11770
rect 29505 -11804 29881 -11770
rect 28776 -11975 28810 -11857
rect 29304 -11975 29338 -11857
rect 29412 -11975 29446 -11857
rect 29940 -11975 29974 -11857
rect 28869 -12062 29245 -12028
rect 29505 -12062 29881 -12028
rect 28869 -12330 29245 -12296
rect 29505 -12330 29881 -12296
rect 28776 -13088 28810 -12396
rect 29304 -13088 29338 -12396
rect 29412 -13088 29446 -12396
rect 29940 -13088 29974 -12396
rect 28869 -13188 29245 -13154
rect 29505 -13188 29881 -13154
rect 28813 -13322 29937 -13288
rect 30469 -11804 30845 -11770
rect 31105 -11804 31481 -11770
rect 30376 -11975 30410 -11857
rect 30904 -11975 30938 -11857
rect 31012 -11975 31046 -11857
rect 31540 -11975 31574 -11857
rect 30469 -12062 30845 -12028
rect 31105 -12062 31481 -12028
rect 30469 -12330 30845 -12296
rect 31105 -12330 31481 -12296
rect 30376 -13088 30410 -12396
rect 30904 -13088 30938 -12396
rect 31012 -13088 31046 -12396
rect 31540 -13088 31574 -12396
rect 30469 -13188 30845 -13154
rect 31105 -13188 31481 -13154
rect 30413 -13322 31537 -13288
rect 32069 -11804 32445 -11770
rect 32705 -11804 33081 -11770
rect 31976 -11975 32010 -11857
rect 32504 -11975 32538 -11857
rect 32612 -11975 32646 -11857
rect 33140 -11975 33174 -11857
rect 32069 -12062 32445 -12028
rect 32705 -12062 33081 -12028
rect 32069 -12330 32445 -12296
rect 32705 -12330 33081 -12296
rect 31976 -13088 32010 -12396
rect 32504 -13088 32538 -12396
rect 32612 -13088 32646 -12396
rect 33140 -13088 33174 -12396
rect 32069 -13188 32445 -13154
rect 32705 -13188 33081 -13154
rect 32013 -13322 33137 -13288
rect 33669 -11804 34045 -11770
rect 34305 -11804 34681 -11770
rect 33576 -11975 33610 -11857
rect 34104 -11975 34138 -11857
rect 34212 -11975 34246 -11857
rect 34740 -11975 34774 -11857
rect 33669 -12062 34045 -12028
rect 34305 -12062 34681 -12028
rect 33669 -12330 34045 -12296
rect 34305 -12330 34681 -12296
rect 33576 -13088 33610 -12396
rect 34104 -13088 34138 -12396
rect 34212 -13088 34246 -12396
rect 34740 -13088 34774 -12396
rect 33669 -13188 34045 -13154
rect 34305 -13188 34681 -13154
rect 33613 -13322 34737 -13288
rect 35269 -11804 35645 -11770
rect 35905 -11804 36281 -11770
rect 35176 -11975 35210 -11857
rect 35704 -11975 35738 -11857
rect 35812 -11975 35846 -11857
rect 36340 -11975 36374 -11857
rect 35269 -12062 35645 -12028
rect 35905 -12062 36281 -12028
rect 36869 -11804 37245 -11770
rect 37505 -11804 37881 -11770
rect 36776 -11975 36810 -11857
rect 37304 -11975 37338 -11857
rect 37412 -11975 37446 -11857
rect 37940 -11975 37974 -11857
rect 36869 -12062 37245 -12028
rect 37505 -12062 37881 -12028
rect 35269 -12330 35645 -12296
rect 35905 -12330 36281 -12296
rect 35176 -13088 35210 -12396
rect 35704 -13088 35738 -12396
rect 35812 -13088 35846 -12396
rect 36340 -13088 36374 -12396
rect 35269 -13188 35645 -13154
rect 35905 -13188 36281 -13154
rect 36869 -12330 37245 -12296
rect 37505 -12330 37881 -12296
rect 36776 -13088 36810 -12396
rect 37304 -13088 37338 -12396
rect 37412 -13088 37446 -12396
rect 37940 -13088 37974 -12396
rect 36869 -13188 37245 -13154
rect 37505 -13188 37881 -13154
rect 35213 -13322 36337 -13288
rect 36813 -13322 37937 -13288
rect 69 -13604 445 -13570
rect 705 -13604 1081 -13570
rect -24 -13775 10 -13657
rect 504 -13775 538 -13657
rect 612 -13775 646 -13657
rect 1140 -13775 1174 -13657
rect 69 -13862 445 -13828
rect 705 -13862 1081 -13828
rect 1669 -13604 2045 -13570
rect 2305 -13604 2681 -13570
rect 1576 -13775 1610 -13657
rect 2104 -13775 2138 -13657
rect 2212 -13775 2246 -13657
rect 2740 -13775 2774 -13657
rect 1669 -13862 2045 -13828
rect 2305 -13862 2681 -13828
rect 69 -14130 445 -14096
rect 705 -14130 1081 -14096
rect -24 -14888 10 -14196
rect 504 -14888 538 -14196
rect 612 -14888 646 -14196
rect 1140 -14888 1174 -14196
rect 69 -14988 445 -14954
rect 705 -14988 1081 -14954
rect 1669 -14130 2045 -14096
rect 2305 -14130 2681 -14096
rect 1576 -14888 1610 -14196
rect 2104 -14888 2138 -14196
rect 2212 -14888 2246 -14196
rect 2740 -14888 2774 -14196
rect 1669 -14988 2045 -14954
rect 2305 -14988 2681 -14954
rect 13 -15122 1137 -15088
rect 1613 -15122 2737 -15088
rect 3269 -13604 3645 -13570
rect 3905 -13604 4281 -13570
rect 3176 -13775 3210 -13657
rect 3704 -13775 3738 -13657
rect 3812 -13775 3846 -13657
rect 4340 -13775 4374 -13657
rect 3269 -13862 3645 -13828
rect 3905 -13862 4281 -13828
rect 3269 -14130 3645 -14096
rect 3905 -14130 4281 -14096
rect 3176 -14888 3210 -14196
rect 3704 -14888 3738 -14196
rect 3812 -14888 3846 -14196
rect 4340 -14888 4374 -14196
rect 3269 -14988 3645 -14954
rect 3905 -14988 4281 -14954
rect 3213 -15122 4337 -15088
rect 4869 -13604 5245 -13570
rect 5505 -13604 5881 -13570
rect 4776 -13775 4810 -13657
rect 5304 -13775 5338 -13657
rect 5412 -13775 5446 -13657
rect 5940 -13775 5974 -13657
rect 4869 -13862 5245 -13828
rect 5505 -13862 5881 -13828
rect 4869 -14130 5245 -14096
rect 5505 -14130 5881 -14096
rect 4776 -14888 4810 -14196
rect 5304 -14888 5338 -14196
rect 5412 -14888 5446 -14196
rect 5940 -14888 5974 -14196
rect 4869 -14988 5245 -14954
rect 5505 -14988 5881 -14954
rect 4813 -15122 5937 -15088
rect 6469 -13604 6845 -13570
rect 7105 -13604 7481 -13570
rect 6376 -13775 6410 -13657
rect 6904 -13775 6938 -13657
rect 7012 -13775 7046 -13657
rect 7540 -13775 7574 -13657
rect 6469 -13862 6845 -13828
rect 7105 -13862 7481 -13828
rect 6469 -14130 6845 -14096
rect 7105 -14130 7481 -14096
rect 6376 -14888 6410 -14196
rect 6904 -14888 6938 -14196
rect 7012 -14888 7046 -14196
rect 7540 -14888 7574 -14196
rect 6469 -14988 6845 -14954
rect 7105 -14988 7481 -14954
rect 6413 -15122 7537 -15088
rect 8069 -13604 8445 -13570
rect 8705 -13604 9081 -13570
rect 7976 -13775 8010 -13657
rect 8504 -13775 8538 -13657
rect 8612 -13775 8646 -13657
rect 9140 -13775 9174 -13657
rect 8069 -13862 8445 -13828
rect 8705 -13862 9081 -13828
rect 8069 -14130 8445 -14096
rect 8705 -14130 9081 -14096
rect 7976 -14888 8010 -14196
rect 8504 -14888 8538 -14196
rect 8612 -14888 8646 -14196
rect 9140 -14888 9174 -14196
rect 8069 -14988 8445 -14954
rect 8705 -14988 9081 -14954
rect 8013 -15122 9137 -15088
rect 9669 -13604 10045 -13570
rect 10305 -13604 10681 -13570
rect 9576 -13775 9610 -13657
rect 10104 -13775 10138 -13657
rect 10212 -13775 10246 -13657
rect 10740 -13775 10774 -13657
rect 9669 -13862 10045 -13828
rect 10305 -13862 10681 -13828
rect 9669 -14130 10045 -14096
rect 10305 -14130 10681 -14096
rect 9576 -14888 9610 -14196
rect 10104 -14888 10138 -14196
rect 10212 -14888 10246 -14196
rect 10740 -14888 10774 -14196
rect 9669 -14988 10045 -14954
rect 10305 -14988 10681 -14954
rect 9613 -15122 10737 -15088
rect 11269 -13604 11645 -13570
rect 11905 -13604 12281 -13570
rect 11176 -13775 11210 -13657
rect 11704 -13775 11738 -13657
rect 11812 -13775 11846 -13657
rect 12340 -13775 12374 -13657
rect 11269 -13862 11645 -13828
rect 11905 -13862 12281 -13828
rect 11269 -14130 11645 -14096
rect 11905 -14130 12281 -14096
rect 11176 -14888 11210 -14196
rect 11704 -14888 11738 -14196
rect 11812 -14888 11846 -14196
rect 12340 -14888 12374 -14196
rect 11269 -14988 11645 -14954
rect 11905 -14988 12281 -14954
rect 11213 -15122 12337 -15088
rect 12869 -13604 13245 -13570
rect 13505 -13604 13881 -13570
rect 12776 -13775 12810 -13657
rect 13304 -13775 13338 -13657
rect 13412 -13775 13446 -13657
rect 13940 -13775 13974 -13657
rect 12869 -13862 13245 -13828
rect 13505 -13862 13881 -13828
rect 12869 -14130 13245 -14096
rect 13505 -14130 13881 -14096
rect 12776 -14888 12810 -14196
rect 13304 -14888 13338 -14196
rect 13412 -14888 13446 -14196
rect 13940 -14888 13974 -14196
rect 12869 -14988 13245 -14954
rect 13505 -14988 13881 -14954
rect 12813 -15122 13937 -15088
rect 14469 -13604 14845 -13570
rect 15105 -13604 15481 -13570
rect 14376 -13775 14410 -13657
rect 14904 -13775 14938 -13657
rect 15012 -13775 15046 -13657
rect 15540 -13775 15574 -13657
rect 14469 -13862 14845 -13828
rect 15105 -13862 15481 -13828
rect 14469 -14130 14845 -14096
rect 15105 -14130 15481 -14096
rect 14376 -14888 14410 -14196
rect 14904 -14888 14938 -14196
rect 15012 -14888 15046 -14196
rect 15540 -14888 15574 -14196
rect 14469 -14988 14845 -14954
rect 15105 -14988 15481 -14954
rect 14413 -15122 15537 -15088
rect 16069 -13604 16445 -13570
rect 16705 -13604 17081 -13570
rect 15976 -13775 16010 -13657
rect 16504 -13775 16538 -13657
rect 16612 -13775 16646 -13657
rect 17140 -13775 17174 -13657
rect 16069 -13862 16445 -13828
rect 16705 -13862 17081 -13828
rect 16069 -14130 16445 -14096
rect 16705 -14130 17081 -14096
rect 15976 -14888 16010 -14196
rect 16504 -14888 16538 -14196
rect 16612 -14888 16646 -14196
rect 17140 -14888 17174 -14196
rect 16069 -14988 16445 -14954
rect 16705 -14988 17081 -14954
rect 16013 -15122 17137 -15088
rect 17669 -13604 18045 -13570
rect 18305 -13604 18681 -13570
rect 17576 -13775 17610 -13657
rect 18104 -13775 18138 -13657
rect 18212 -13775 18246 -13657
rect 18740 -13775 18774 -13657
rect 17669 -13862 18045 -13828
rect 18305 -13862 18681 -13828
rect 17669 -14130 18045 -14096
rect 18305 -14130 18681 -14096
rect 17576 -14888 17610 -14196
rect 18104 -14888 18138 -14196
rect 18212 -14888 18246 -14196
rect 18740 -14888 18774 -14196
rect 17669 -14988 18045 -14954
rect 18305 -14988 18681 -14954
rect 17613 -15122 18737 -15088
rect 19269 -13604 19645 -13570
rect 19905 -13604 20281 -13570
rect 19176 -13775 19210 -13657
rect 19704 -13775 19738 -13657
rect 19812 -13775 19846 -13657
rect 20340 -13775 20374 -13657
rect 19269 -13862 19645 -13828
rect 19905 -13862 20281 -13828
rect 19269 -14130 19645 -14096
rect 19905 -14130 20281 -14096
rect 19176 -14888 19210 -14196
rect 19704 -14888 19738 -14196
rect 19812 -14888 19846 -14196
rect 20340 -14888 20374 -14196
rect 19269 -14988 19645 -14954
rect 19905 -14988 20281 -14954
rect 19213 -15122 20337 -15088
rect 20869 -13604 21245 -13570
rect 21505 -13604 21881 -13570
rect 20776 -13775 20810 -13657
rect 21304 -13775 21338 -13657
rect 21412 -13775 21446 -13657
rect 21940 -13775 21974 -13657
rect 20869 -13862 21245 -13828
rect 21505 -13862 21881 -13828
rect 20869 -14130 21245 -14096
rect 21505 -14130 21881 -14096
rect 20776 -14888 20810 -14196
rect 21304 -14888 21338 -14196
rect 21412 -14888 21446 -14196
rect 21940 -14888 21974 -14196
rect 20869 -14988 21245 -14954
rect 21505 -14988 21881 -14954
rect 20813 -15122 21937 -15088
rect 22469 -13604 22845 -13570
rect 23105 -13604 23481 -13570
rect 22376 -13775 22410 -13657
rect 22904 -13775 22938 -13657
rect 23012 -13775 23046 -13657
rect 23540 -13775 23574 -13657
rect 22469 -13862 22845 -13828
rect 23105 -13862 23481 -13828
rect 22469 -14130 22845 -14096
rect 23105 -14130 23481 -14096
rect 22376 -14888 22410 -14196
rect 22904 -14888 22938 -14196
rect 23012 -14888 23046 -14196
rect 23540 -14888 23574 -14196
rect 22469 -14988 22845 -14954
rect 23105 -14988 23481 -14954
rect 22413 -15122 23537 -15088
rect 24069 -13604 24445 -13570
rect 24705 -13604 25081 -13570
rect 23976 -13775 24010 -13657
rect 24504 -13775 24538 -13657
rect 24612 -13775 24646 -13657
rect 25140 -13775 25174 -13657
rect 24069 -13862 24445 -13828
rect 24705 -13862 25081 -13828
rect 24069 -14130 24445 -14096
rect 24705 -14130 25081 -14096
rect 23976 -14888 24010 -14196
rect 24504 -14888 24538 -14196
rect 24612 -14888 24646 -14196
rect 25140 -14888 25174 -14196
rect 24069 -14988 24445 -14954
rect 24705 -14988 25081 -14954
rect 24013 -15122 25137 -15088
rect 25669 -13604 26045 -13570
rect 26305 -13604 26681 -13570
rect 25576 -13775 25610 -13657
rect 26104 -13775 26138 -13657
rect 26212 -13775 26246 -13657
rect 26740 -13775 26774 -13657
rect 25669 -13862 26045 -13828
rect 26305 -13862 26681 -13828
rect 25669 -14130 26045 -14096
rect 26305 -14130 26681 -14096
rect 25576 -14888 25610 -14196
rect 26104 -14888 26138 -14196
rect 26212 -14888 26246 -14196
rect 26740 -14888 26774 -14196
rect 25669 -14988 26045 -14954
rect 26305 -14988 26681 -14954
rect 25613 -15122 26737 -15088
rect 27269 -13604 27645 -13570
rect 27905 -13604 28281 -13570
rect 27176 -13775 27210 -13657
rect 27704 -13775 27738 -13657
rect 27812 -13775 27846 -13657
rect 28340 -13775 28374 -13657
rect 27269 -13862 27645 -13828
rect 27905 -13862 28281 -13828
rect 27269 -14130 27645 -14096
rect 27905 -14130 28281 -14096
rect 27176 -14888 27210 -14196
rect 27704 -14888 27738 -14196
rect 27812 -14888 27846 -14196
rect 28340 -14888 28374 -14196
rect 27269 -14988 27645 -14954
rect 27905 -14988 28281 -14954
rect 27213 -15122 28337 -15088
rect 28869 -13604 29245 -13570
rect 29505 -13604 29881 -13570
rect 28776 -13775 28810 -13657
rect 29304 -13775 29338 -13657
rect 29412 -13775 29446 -13657
rect 29940 -13775 29974 -13657
rect 28869 -13862 29245 -13828
rect 29505 -13862 29881 -13828
rect 28869 -14130 29245 -14096
rect 29505 -14130 29881 -14096
rect 28776 -14888 28810 -14196
rect 29304 -14888 29338 -14196
rect 29412 -14888 29446 -14196
rect 29940 -14888 29974 -14196
rect 28869 -14988 29245 -14954
rect 29505 -14988 29881 -14954
rect 28813 -15122 29937 -15088
rect 30469 -13604 30845 -13570
rect 31105 -13604 31481 -13570
rect 30376 -13775 30410 -13657
rect 30904 -13775 30938 -13657
rect 31012 -13775 31046 -13657
rect 31540 -13775 31574 -13657
rect 30469 -13862 30845 -13828
rect 31105 -13862 31481 -13828
rect 30469 -14130 30845 -14096
rect 31105 -14130 31481 -14096
rect 30376 -14888 30410 -14196
rect 30904 -14888 30938 -14196
rect 31012 -14888 31046 -14196
rect 31540 -14888 31574 -14196
rect 30469 -14988 30845 -14954
rect 31105 -14988 31481 -14954
rect 30413 -15122 31537 -15088
rect 32069 -13604 32445 -13570
rect 32705 -13604 33081 -13570
rect 31976 -13775 32010 -13657
rect 32504 -13775 32538 -13657
rect 32612 -13775 32646 -13657
rect 33140 -13775 33174 -13657
rect 32069 -13862 32445 -13828
rect 32705 -13862 33081 -13828
rect 32069 -14130 32445 -14096
rect 32705 -14130 33081 -14096
rect 31976 -14888 32010 -14196
rect 32504 -14888 32538 -14196
rect 32612 -14888 32646 -14196
rect 33140 -14888 33174 -14196
rect 32069 -14988 32445 -14954
rect 32705 -14988 33081 -14954
rect 32013 -15122 33137 -15088
rect 33669 -13604 34045 -13570
rect 34305 -13604 34681 -13570
rect 33576 -13775 33610 -13657
rect 34104 -13775 34138 -13657
rect 34212 -13775 34246 -13657
rect 34740 -13775 34774 -13657
rect 33669 -13862 34045 -13828
rect 34305 -13862 34681 -13828
rect 33669 -14130 34045 -14096
rect 34305 -14130 34681 -14096
rect 33576 -14888 33610 -14196
rect 34104 -14888 34138 -14196
rect 34212 -14888 34246 -14196
rect 34740 -14888 34774 -14196
rect 33669 -14988 34045 -14954
rect 34305 -14988 34681 -14954
rect 33613 -15122 34737 -15088
rect 35269 -13604 35645 -13570
rect 35905 -13604 36281 -13570
rect 35176 -13775 35210 -13657
rect 35704 -13775 35738 -13657
rect 35812 -13775 35846 -13657
rect 36340 -13775 36374 -13657
rect 35269 -13862 35645 -13828
rect 35905 -13862 36281 -13828
rect 36869 -13604 37245 -13570
rect 37505 -13604 37881 -13570
rect 36776 -13775 36810 -13657
rect 37304 -13775 37338 -13657
rect 37412 -13775 37446 -13657
rect 37940 -13775 37974 -13657
rect 36869 -13862 37245 -13828
rect 37505 -13862 37881 -13828
rect 35269 -14130 35645 -14096
rect 35905 -14130 36281 -14096
rect 35176 -14888 35210 -14196
rect 35704 -14888 35738 -14196
rect 35812 -14888 35846 -14196
rect 36340 -14888 36374 -14196
rect 35269 -14988 35645 -14954
rect 35905 -14988 36281 -14954
rect 36869 -14130 37245 -14096
rect 37505 -14130 37881 -14096
rect 36776 -14888 36810 -14196
rect 37304 -14888 37338 -14196
rect 37412 -14888 37446 -14196
rect 37940 -14888 37974 -14196
rect 36869 -14988 37245 -14954
rect 37505 -14988 37881 -14954
rect 35213 -15122 36337 -15088
rect 36813 -15122 37937 -15088
rect 69 -15404 445 -15370
rect 705 -15404 1081 -15370
rect -24 -15575 10 -15457
rect 504 -15575 538 -15457
rect 612 -15575 646 -15457
rect 1140 -15575 1174 -15457
rect 69 -15662 445 -15628
rect 705 -15662 1081 -15628
rect 1669 -15404 2045 -15370
rect 2305 -15404 2681 -15370
rect 1576 -15575 1610 -15457
rect 2104 -15575 2138 -15457
rect 2212 -15575 2246 -15457
rect 2740 -15575 2774 -15457
rect 1669 -15662 2045 -15628
rect 2305 -15662 2681 -15628
rect 69 -15930 445 -15896
rect 705 -15930 1081 -15896
rect -24 -16688 10 -15996
rect 504 -16688 538 -15996
rect 612 -16688 646 -15996
rect 1140 -16688 1174 -15996
rect 69 -16788 445 -16754
rect 705 -16788 1081 -16754
rect 1669 -15930 2045 -15896
rect 2305 -15930 2681 -15896
rect 1576 -16688 1610 -15996
rect 2104 -16688 2138 -15996
rect 2212 -16688 2246 -15996
rect 2740 -16688 2774 -15996
rect 1669 -16788 2045 -16754
rect 2305 -16788 2681 -16754
rect 13 -16922 1137 -16888
rect 1613 -16922 2737 -16888
rect 3269 -15404 3645 -15370
rect 3905 -15404 4281 -15370
rect 3176 -15575 3210 -15457
rect 3704 -15575 3738 -15457
rect 3812 -15575 3846 -15457
rect 4340 -15575 4374 -15457
rect 3269 -15662 3645 -15628
rect 3905 -15662 4281 -15628
rect 3269 -15930 3645 -15896
rect 3905 -15930 4281 -15896
rect 3176 -16688 3210 -15996
rect 3704 -16688 3738 -15996
rect 3812 -16688 3846 -15996
rect 4340 -16688 4374 -15996
rect 3269 -16788 3645 -16754
rect 3905 -16788 4281 -16754
rect 3213 -16922 4337 -16888
rect 4869 -15404 5245 -15370
rect 5505 -15404 5881 -15370
rect 4776 -15575 4810 -15457
rect 5304 -15575 5338 -15457
rect 5412 -15575 5446 -15457
rect 5940 -15575 5974 -15457
rect 4869 -15662 5245 -15628
rect 5505 -15662 5881 -15628
rect 4869 -15930 5245 -15896
rect 5505 -15930 5881 -15896
rect 4776 -16688 4810 -15996
rect 5304 -16688 5338 -15996
rect 5412 -16688 5446 -15996
rect 5940 -16688 5974 -15996
rect 4869 -16788 5245 -16754
rect 5505 -16788 5881 -16754
rect 4813 -16922 5937 -16888
rect 6469 -15404 6845 -15370
rect 7105 -15404 7481 -15370
rect 6376 -15575 6410 -15457
rect 6904 -15575 6938 -15457
rect 7012 -15575 7046 -15457
rect 7540 -15575 7574 -15457
rect 6469 -15662 6845 -15628
rect 7105 -15662 7481 -15628
rect 6469 -15930 6845 -15896
rect 7105 -15930 7481 -15896
rect 6376 -16688 6410 -15996
rect 6904 -16688 6938 -15996
rect 7012 -16688 7046 -15996
rect 7540 -16688 7574 -15996
rect 6469 -16788 6845 -16754
rect 7105 -16788 7481 -16754
rect 6413 -16922 7537 -16888
rect 8069 -15404 8445 -15370
rect 8705 -15404 9081 -15370
rect 7976 -15575 8010 -15457
rect 8504 -15575 8538 -15457
rect 8612 -15575 8646 -15457
rect 9140 -15575 9174 -15457
rect 8069 -15662 8445 -15628
rect 8705 -15662 9081 -15628
rect 8069 -15930 8445 -15896
rect 8705 -15930 9081 -15896
rect 7976 -16688 8010 -15996
rect 8504 -16688 8538 -15996
rect 8612 -16688 8646 -15996
rect 9140 -16688 9174 -15996
rect 8069 -16788 8445 -16754
rect 8705 -16788 9081 -16754
rect 8013 -16922 9137 -16888
rect 9669 -15404 10045 -15370
rect 10305 -15404 10681 -15370
rect 9576 -15575 9610 -15457
rect 10104 -15575 10138 -15457
rect 10212 -15575 10246 -15457
rect 10740 -15575 10774 -15457
rect 9669 -15662 10045 -15628
rect 10305 -15662 10681 -15628
rect 9669 -15930 10045 -15896
rect 10305 -15930 10681 -15896
rect 9576 -16688 9610 -15996
rect 10104 -16688 10138 -15996
rect 10212 -16688 10246 -15996
rect 10740 -16688 10774 -15996
rect 9669 -16788 10045 -16754
rect 10305 -16788 10681 -16754
rect 9613 -16922 10737 -16888
rect 11269 -15404 11645 -15370
rect 11905 -15404 12281 -15370
rect 11176 -15575 11210 -15457
rect 11704 -15575 11738 -15457
rect 11812 -15575 11846 -15457
rect 12340 -15575 12374 -15457
rect 11269 -15662 11645 -15628
rect 11905 -15662 12281 -15628
rect 11269 -15930 11645 -15896
rect 11905 -15930 12281 -15896
rect 11176 -16688 11210 -15996
rect 11704 -16688 11738 -15996
rect 11812 -16688 11846 -15996
rect 12340 -16688 12374 -15996
rect 11269 -16788 11645 -16754
rect 11905 -16788 12281 -16754
rect 11213 -16922 12337 -16888
rect 12869 -15404 13245 -15370
rect 13505 -15404 13881 -15370
rect 12776 -15575 12810 -15457
rect 13304 -15575 13338 -15457
rect 13412 -15575 13446 -15457
rect 13940 -15575 13974 -15457
rect 12869 -15662 13245 -15628
rect 13505 -15662 13881 -15628
rect 12869 -15930 13245 -15896
rect 13505 -15930 13881 -15896
rect 12776 -16688 12810 -15996
rect 13304 -16688 13338 -15996
rect 13412 -16688 13446 -15996
rect 13940 -16688 13974 -15996
rect 12869 -16788 13245 -16754
rect 13505 -16788 13881 -16754
rect 12813 -16922 13937 -16888
rect 14469 -15404 14845 -15370
rect 15105 -15404 15481 -15370
rect 14376 -15575 14410 -15457
rect 14904 -15575 14938 -15457
rect 15012 -15575 15046 -15457
rect 15540 -15575 15574 -15457
rect 14469 -15662 14845 -15628
rect 15105 -15662 15481 -15628
rect 14469 -15930 14845 -15896
rect 15105 -15930 15481 -15896
rect 14376 -16688 14410 -15996
rect 14904 -16688 14938 -15996
rect 15012 -16688 15046 -15996
rect 15540 -16688 15574 -15996
rect 14469 -16788 14845 -16754
rect 15105 -16788 15481 -16754
rect 14413 -16922 15537 -16888
rect 16069 -15404 16445 -15370
rect 16705 -15404 17081 -15370
rect 15976 -15575 16010 -15457
rect 16504 -15575 16538 -15457
rect 16612 -15575 16646 -15457
rect 17140 -15575 17174 -15457
rect 16069 -15662 16445 -15628
rect 16705 -15662 17081 -15628
rect 16069 -15930 16445 -15896
rect 16705 -15930 17081 -15896
rect 15976 -16688 16010 -15996
rect 16504 -16688 16538 -15996
rect 16612 -16688 16646 -15996
rect 17140 -16688 17174 -15996
rect 16069 -16788 16445 -16754
rect 16705 -16788 17081 -16754
rect 16013 -16922 17137 -16888
rect 17669 -15404 18045 -15370
rect 18305 -15404 18681 -15370
rect 17576 -15575 17610 -15457
rect 18104 -15575 18138 -15457
rect 18212 -15575 18246 -15457
rect 18740 -15575 18774 -15457
rect 17669 -15662 18045 -15628
rect 18305 -15662 18681 -15628
rect 17669 -15930 18045 -15896
rect 18305 -15930 18681 -15896
rect 17576 -16688 17610 -15996
rect 18104 -16688 18138 -15996
rect 18212 -16688 18246 -15996
rect 18740 -16688 18774 -15996
rect 17669 -16788 18045 -16754
rect 18305 -16788 18681 -16754
rect 17613 -16922 18737 -16888
rect 19269 -15404 19645 -15370
rect 19905 -15404 20281 -15370
rect 19176 -15575 19210 -15457
rect 19704 -15575 19738 -15457
rect 19812 -15575 19846 -15457
rect 20340 -15575 20374 -15457
rect 19269 -15662 19645 -15628
rect 19905 -15662 20281 -15628
rect 19269 -15930 19645 -15896
rect 19905 -15930 20281 -15896
rect 19176 -16688 19210 -15996
rect 19704 -16688 19738 -15996
rect 19812 -16688 19846 -15996
rect 20340 -16688 20374 -15996
rect 19269 -16788 19645 -16754
rect 19905 -16788 20281 -16754
rect 19213 -16922 20337 -16888
rect 20869 -15404 21245 -15370
rect 21505 -15404 21881 -15370
rect 20776 -15575 20810 -15457
rect 21304 -15575 21338 -15457
rect 21412 -15575 21446 -15457
rect 21940 -15575 21974 -15457
rect 20869 -15662 21245 -15628
rect 21505 -15662 21881 -15628
rect 20869 -15930 21245 -15896
rect 21505 -15930 21881 -15896
rect 20776 -16688 20810 -15996
rect 21304 -16688 21338 -15996
rect 21412 -16688 21446 -15996
rect 21940 -16688 21974 -15996
rect 20869 -16788 21245 -16754
rect 21505 -16788 21881 -16754
rect 20813 -16922 21937 -16888
rect 22469 -15404 22845 -15370
rect 23105 -15404 23481 -15370
rect 22376 -15575 22410 -15457
rect 22904 -15575 22938 -15457
rect 23012 -15575 23046 -15457
rect 23540 -15575 23574 -15457
rect 22469 -15662 22845 -15628
rect 23105 -15662 23481 -15628
rect 22469 -15930 22845 -15896
rect 23105 -15930 23481 -15896
rect 22376 -16688 22410 -15996
rect 22904 -16688 22938 -15996
rect 23012 -16688 23046 -15996
rect 23540 -16688 23574 -15996
rect 22469 -16788 22845 -16754
rect 23105 -16788 23481 -16754
rect 22413 -16922 23537 -16888
rect 24069 -15404 24445 -15370
rect 24705 -15404 25081 -15370
rect 23976 -15575 24010 -15457
rect 24504 -15575 24538 -15457
rect 24612 -15575 24646 -15457
rect 25140 -15575 25174 -15457
rect 24069 -15662 24445 -15628
rect 24705 -15662 25081 -15628
rect 24069 -15930 24445 -15896
rect 24705 -15930 25081 -15896
rect 23976 -16688 24010 -15996
rect 24504 -16688 24538 -15996
rect 24612 -16688 24646 -15996
rect 25140 -16688 25174 -15996
rect 24069 -16788 24445 -16754
rect 24705 -16788 25081 -16754
rect 24013 -16922 25137 -16888
rect 25669 -15404 26045 -15370
rect 26305 -15404 26681 -15370
rect 25576 -15575 25610 -15457
rect 26104 -15575 26138 -15457
rect 26212 -15575 26246 -15457
rect 26740 -15575 26774 -15457
rect 25669 -15662 26045 -15628
rect 26305 -15662 26681 -15628
rect 25669 -15930 26045 -15896
rect 26305 -15930 26681 -15896
rect 25576 -16688 25610 -15996
rect 26104 -16688 26138 -15996
rect 26212 -16688 26246 -15996
rect 26740 -16688 26774 -15996
rect 25669 -16788 26045 -16754
rect 26305 -16788 26681 -16754
rect 25613 -16922 26737 -16888
rect 27269 -15404 27645 -15370
rect 27905 -15404 28281 -15370
rect 27176 -15575 27210 -15457
rect 27704 -15575 27738 -15457
rect 27812 -15575 27846 -15457
rect 28340 -15575 28374 -15457
rect 27269 -15662 27645 -15628
rect 27905 -15662 28281 -15628
rect 27269 -15930 27645 -15896
rect 27905 -15930 28281 -15896
rect 27176 -16688 27210 -15996
rect 27704 -16688 27738 -15996
rect 27812 -16688 27846 -15996
rect 28340 -16688 28374 -15996
rect 27269 -16788 27645 -16754
rect 27905 -16788 28281 -16754
rect 27213 -16922 28337 -16888
rect 28869 -15404 29245 -15370
rect 29505 -15404 29881 -15370
rect 28776 -15575 28810 -15457
rect 29304 -15575 29338 -15457
rect 29412 -15575 29446 -15457
rect 29940 -15575 29974 -15457
rect 28869 -15662 29245 -15628
rect 29505 -15662 29881 -15628
rect 28869 -15930 29245 -15896
rect 29505 -15930 29881 -15896
rect 28776 -16688 28810 -15996
rect 29304 -16688 29338 -15996
rect 29412 -16688 29446 -15996
rect 29940 -16688 29974 -15996
rect 28869 -16788 29245 -16754
rect 29505 -16788 29881 -16754
rect 28813 -16922 29937 -16888
rect 30469 -15404 30845 -15370
rect 31105 -15404 31481 -15370
rect 30376 -15575 30410 -15457
rect 30904 -15575 30938 -15457
rect 31012 -15575 31046 -15457
rect 31540 -15575 31574 -15457
rect 30469 -15662 30845 -15628
rect 31105 -15662 31481 -15628
rect 30469 -15930 30845 -15896
rect 31105 -15930 31481 -15896
rect 30376 -16688 30410 -15996
rect 30904 -16688 30938 -15996
rect 31012 -16688 31046 -15996
rect 31540 -16688 31574 -15996
rect 30469 -16788 30845 -16754
rect 31105 -16788 31481 -16754
rect 30413 -16922 31537 -16888
rect 32069 -15404 32445 -15370
rect 32705 -15404 33081 -15370
rect 31976 -15575 32010 -15457
rect 32504 -15575 32538 -15457
rect 32612 -15575 32646 -15457
rect 33140 -15575 33174 -15457
rect 32069 -15662 32445 -15628
rect 32705 -15662 33081 -15628
rect 32069 -15930 32445 -15896
rect 32705 -15930 33081 -15896
rect 31976 -16688 32010 -15996
rect 32504 -16688 32538 -15996
rect 32612 -16688 32646 -15996
rect 33140 -16688 33174 -15996
rect 32069 -16788 32445 -16754
rect 32705 -16788 33081 -16754
rect 32013 -16922 33137 -16888
rect 33669 -15404 34045 -15370
rect 34305 -15404 34681 -15370
rect 33576 -15575 33610 -15457
rect 34104 -15575 34138 -15457
rect 34212 -15575 34246 -15457
rect 34740 -15575 34774 -15457
rect 33669 -15662 34045 -15628
rect 34305 -15662 34681 -15628
rect 33669 -15930 34045 -15896
rect 34305 -15930 34681 -15896
rect 33576 -16688 33610 -15996
rect 34104 -16688 34138 -15996
rect 34212 -16688 34246 -15996
rect 34740 -16688 34774 -15996
rect 33669 -16788 34045 -16754
rect 34305 -16788 34681 -16754
rect 33613 -16922 34737 -16888
rect 35269 -15404 35645 -15370
rect 35905 -15404 36281 -15370
rect 35176 -15575 35210 -15457
rect 35704 -15575 35738 -15457
rect 35812 -15575 35846 -15457
rect 36340 -15575 36374 -15457
rect 35269 -15662 35645 -15628
rect 35905 -15662 36281 -15628
rect 36869 -15404 37245 -15370
rect 37505 -15404 37881 -15370
rect 36776 -15575 36810 -15457
rect 37304 -15575 37338 -15457
rect 37412 -15575 37446 -15457
rect 37940 -15575 37974 -15457
rect 36869 -15662 37245 -15628
rect 37505 -15662 37881 -15628
rect 35269 -15930 35645 -15896
rect 35905 -15930 36281 -15896
rect 35176 -16688 35210 -15996
rect 35704 -16688 35738 -15996
rect 35812 -16688 35846 -15996
rect 36340 -16688 36374 -15996
rect 35269 -16788 35645 -16754
rect 35905 -16788 36281 -16754
rect 36869 -15930 37245 -15896
rect 37505 -15930 37881 -15896
rect 36776 -16688 36810 -15996
rect 37304 -16688 37338 -15996
rect 37412 -16688 37446 -15996
rect 37940 -16688 37974 -15996
rect 36869 -16788 37245 -16754
rect 37505 -16788 37881 -16754
rect 35213 -16922 36337 -16888
rect 36813 -16922 37937 -16888
rect 69 -17204 445 -17170
rect 705 -17204 1081 -17170
rect -24 -17375 10 -17257
rect 504 -17375 538 -17257
rect 612 -17375 646 -17257
rect 1140 -17375 1174 -17257
rect 69 -17462 445 -17428
rect 705 -17462 1081 -17428
rect 1669 -17204 2045 -17170
rect 2305 -17204 2681 -17170
rect 1576 -17375 1610 -17257
rect 2104 -17375 2138 -17257
rect 2212 -17375 2246 -17257
rect 2740 -17375 2774 -17257
rect 1669 -17462 2045 -17428
rect 2305 -17462 2681 -17428
rect 69 -17730 445 -17696
rect 705 -17730 1081 -17696
rect -24 -18488 10 -17796
rect 504 -18488 538 -17796
rect 612 -18488 646 -17796
rect 1140 -18488 1174 -17796
rect 69 -18588 445 -18554
rect 705 -18588 1081 -18554
rect 1669 -17730 2045 -17696
rect 2305 -17730 2681 -17696
rect 1576 -18488 1610 -17796
rect 2104 -18488 2138 -17796
rect 2212 -18488 2246 -17796
rect 2740 -18488 2774 -17796
rect 1669 -18588 2045 -18554
rect 2305 -18588 2681 -18554
rect 13 -18722 1137 -18688
rect 1613 -18722 2737 -18688
rect 3269 -17204 3645 -17170
rect 3905 -17204 4281 -17170
rect 3176 -17375 3210 -17257
rect 3704 -17375 3738 -17257
rect 3812 -17375 3846 -17257
rect 4340 -17375 4374 -17257
rect 3269 -17462 3645 -17428
rect 3905 -17462 4281 -17428
rect 3269 -17730 3645 -17696
rect 3905 -17730 4281 -17696
rect 3176 -18488 3210 -17796
rect 3704 -18488 3738 -17796
rect 3812 -18488 3846 -17796
rect 4340 -18488 4374 -17796
rect 3269 -18588 3645 -18554
rect 3905 -18588 4281 -18554
rect 3213 -18722 4337 -18688
rect 4869 -17204 5245 -17170
rect 5505 -17204 5881 -17170
rect 4776 -17375 4810 -17257
rect 5304 -17375 5338 -17257
rect 5412 -17375 5446 -17257
rect 5940 -17375 5974 -17257
rect 4869 -17462 5245 -17428
rect 5505 -17462 5881 -17428
rect 4869 -17730 5245 -17696
rect 5505 -17730 5881 -17696
rect 4776 -18488 4810 -17796
rect 5304 -18488 5338 -17796
rect 5412 -18488 5446 -17796
rect 5940 -18488 5974 -17796
rect 4869 -18588 5245 -18554
rect 5505 -18588 5881 -18554
rect 4813 -18722 5937 -18688
rect 6469 -17204 6845 -17170
rect 7105 -17204 7481 -17170
rect 6376 -17375 6410 -17257
rect 6904 -17375 6938 -17257
rect 7012 -17375 7046 -17257
rect 7540 -17375 7574 -17257
rect 6469 -17462 6845 -17428
rect 7105 -17462 7481 -17428
rect 6469 -17730 6845 -17696
rect 7105 -17730 7481 -17696
rect 6376 -18488 6410 -17796
rect 6904 -18488 6938 -17796
rect 7012 -18488 7046 -17796
rect 7540 -18488 7574 -17796
rect 6469 -18588 6845 -18554
rect 7105 -18588 7481 -18554
rect 6413 -18722 7537 -18688
rect 8069 -17204 8445 -17170
rect 8705 -17204 9081 -17170
rect 7976 -17375 8010 -17257
rect 8504 -17375 8538 -17257
rect 8612 -17375 8646 -17257
rect 9140 -17375 9174 -17257
rect 8069 -17462 8445 -17428
rect 8705 -17462 9081 -17428
rect 8069 -17730 8445 -17696
rect 8705 -17730 9081 -17696
rect 7976 -18488 8010 -17796
rect 8504 -18488 8538 -17796
rect 8612 -18488 8646 -17796
rect 9140 -18488 9174 -17796
rect 8069 -18588 8445 -18554
rect 8705 -18588 9081 -18554
rect 8013 -18722 9137 -18688
rect 9669 -17204 10045 -17170
rect 10305 -17204 10681 -17170
rect 9576 -17375 9610 -17257
rect 10104 -17375 10138 -17257
rect 10212 -17375 10246 -17257
rect 10740 -17375 10774 -17257
rect 9669 -17462 10045 -17428
rect 10305 -17462 10681 -17428
rect 9669 -17730 10045 -17696
rect 10305 -17730 10681 -17696
rect 9576 -18488 9610 -17796
rect 10104 -18488 10138 -17796
rect 10212 -18488 10246 -17796
rect 10740 -18488 10774 -17796
rect 9669 -18588 10045 -18554
rect 10305 -18588 10681 -18554
rect 9613 -18722 10737 -18688
rect 11269 -17204 11645 -17170
rect 11905 -17204 12281 -17170
rect 11176 -17375 11210 -17257
rect 11704 -17375 11738 -17257
rect 11812 -17375 11846 -17257
rect 12340 -17375 12374 -17257
rect 11269 -17462 11645 -17428
rect 11905 -17462 12281 -17428
rect 11269 -17730 11645 -17696
rect 11905 -17730 12281 -17696
rect 11176 -18488 11210 -17796
rect 11704 -18488 11738 -17796
rect 11812 -18488 11846 -17796
rect 12340 -18488 12374 -17796
rect 11269 -18588 11645 -18554
rect 11905 -18588 12281 -18554
rect 11213 -18722 12337 -18688
rect 12869 -17204 13245 -17170
rect 13505 -17204 13881 -17170
rect 12776 -17375 12810 -17257
rect 13304 -17375 13338 -17257
rect 13412 -17375 13446 -17257
rect 13940 -17375 13974 -17257
rect 12869 -17462 13245 -17428
rect 13505 -17462 13881 -17428
rect 12869 -17730 13245 -17696
rect 13505 -17730 13881 -17696
rect 12776 -18488 12810 -17796
rect 13304 -18488 13338 -17796
rect 13412 -18488 13446 -17796
rect 13940 -18488 13974 -17796
rect 12869 -18588 13245 -18554
rect 13505 -18588 13881 -18554
rect 12813 -18722 13937 -18688
rect 14469 -17204 14845 -17170
rect 15105 -17204 15481 -17170
rect 14376 -17375 14410 -17257
rect 14904 -17375 14938 -17257
rect 15012 -17375 15046 -17257
rect 15540 -17375 15574 -17257
rect 14469 -17462 14845 -17428
rect 15105 -17462 15481 -17428
rect 14469 -17730 14845 -17696
rect 15105 -17730 15481 -17696
rect 14376 -18488 14410 -17796
rect 14904 -18488 14938 -17796
rect 15012 -18488 15046 -17796
rect 15540 -18488 15574 -17796
rect 14469 -18588 14845 -18554
rect 15105 -18588 15481 -18554
rect 14413 -18722 15537 -18688
rect 16069 -17204 16445 -17170
rect 16705 -17204 17081 -17170
rect 15976 -17375 16010 -17257
rect 16504 -17375 16538 -17257
rect 16612 -17375 16646 -17257
rect 17140 -17375 17174 -17257
rect 16069 -17462 16445 -17428
rect 16705 -17462 17081 -17428
rect 16069 -17730 16445 -17696
rect 16705 -17730 17081 -17696
rect 15976 -18488 16010 -17796
rect 16504 -18488 16538 -17796
rect 16612 -18488 16646 -17796
rect 17140 -18488 17174 -17796
rect 16069 -18588 16445 -18554
rect 16705 -18588 17081 -18554
rect 16013 -18722 17137 -18688
rect 17669 -17204 18045 -17170
rect 18305 -17204 18681 -17170
rect 17576 -17375 17610 -17257
rect 18104 -17375 18138 -17257
rect 18212 -17375 18246 -17257
rect 18740 -17375 18774 -17257
rect 17669 -17462 18045 -17428
rect 18305 -17462 18681 -17428
rect 17669 -17730 18045 -17696
rect 18305 -17730 18681 -17696
rect 17576 -18488 17610 -17796
rect 18104 -18488 18138 -17796
rect 18212 -18488 18246 -17796
rect 18740 -18488 18774 -17796
rect 17669 -18588 18045 -18554
rect 18305 -18588 18681 -18554
rect 17613 -18722 18737 -18688
rect 19269 -17204 19645 -17170
rect 19905 -17204 20281 -17170
rect 19176 -17375 19210 -17257
rect 19704 -17375 19738 -17257
rect 19812 -17375 19846 -17257
rect 20340 -17375 20374 -17257
rect 19269 -17462 19645 -17428
rect 19905 -17462 20281 -17428
rect 19269 -17730 19645 -17696
rect 19905 -17730 20281 -17696
rect 19176 -18488 19210 -17796
rect 19704 -18488 19738 -17796
rect 19812 -18488 19846 -17796
rect 20340 -18488 20374 -17796
rect 19269 -18588 19645 -18554
rect 19905 -18588 20281 -18554
rect 19213 -18722 20337 -18688
rect 20869 -17204 21245 -17170
rect 21505 -17204 21881 -17170
rect 20776 -17375 20810 -17257
rect 21304 -17375 21338 -17257
rect 21412 -17375 21446 -17257
rect 21940 -17375 21974 -17257
rect 20869 -17462 21245 -17428
rect 21505 -17462 21881 -17428
rect 20869 -17730 21245 -17696
rect 21505 -17730 21881 -17696
rect 20776 -18488 20810 -17796
rect 21304 -18488 21338 -17796
rect 21412 -18488 21446 -17796
rect 21940 -18488 21974 -17796
rect 20869 -18588 21245 -18554
rect 21505 -18588 21881 -18554
rect 20813 -18722 21937 -18688
rect 22469 -17204 22845 -17170
rect 23105 -17204 23481 -17170
rect 22376 -17375 22410 -17257
rect 22904 -17375 22938 -17257
rect 23012 -17375 23046 -17257
rect 23540 -17375 23574 -17257
rect 22469 -17462 22845 -17428
rect 23105 -17462 23481 -17428
rect 22469 -17730 22845 -17696
rect 23105 -17730 23481 -17696
rect 22376 -18488 22410 -17796
rect 22904 -18488 22938 -17796
rect 23012 -18488 23046 -17796
rect 23540 -18488 23574 -17796
rect 22469 -18588 22845 -18554
rect 23105 -18588 23481 -18554
rect 22413 -18722 23537 -18688
rect 24069 -17204 24445 -17170
rect 24705 -17204 25081 -17170
rect 23976 -17375 24010 -17257
rect 24504 -17375 24538 -17257
rect 24612 -17375 24646 -17257
rect 25140 -17375 25174 -17257
rect 24069 -17462 24445 -17428
rect 24705 -17462 25081 -17428
rect 24069 -17730 24445 -17696
rect 24705 -17730 25081 -17696
rect 23976 -18488 24010 -17796
rect 24504 -18488 24538 -17796
rect 24612 -18488 24646 -17796
rect 25140 -18488 25174 -17796
rect 24069 -18588 24445 -18554
rect 24705 -18588 25081 -18554
rect 24013 -18722 25137 -18688
rect 25669 -17204 26045 -17170
rect 26305 -17204 26681 -17170
rect 25576 -17375 25610 -17257
rect 26104 -17375 26138 -17257
rect 26212 -17375 26246 -17257
rect 26740 -17375 26774 -17257
rect 25669 -17462 26045 -17428
rect 26305 -17462 26681 -17428
rect 25669 -17730 26045 -17696
rect 26305 -17730 26681 -17696
rect 25576 -18488 25610 -17796
rect 26104 -18488 26138 -17796
rect 26212 -18488 26246 -17796
rect 26740 -18488 26774 -17796
rect 25669 -18588 26045 -18554
rect 26305 -18588 26681 -18554
rect 25613 -18722 26737 -18688
rect 27269 -17204 27645 -17170
rect 27905 -17204 28281 -17170
rect 27176 -17375 27210 -17257
rect 27704 -17375 27738 -17257
rect 27812 -17375 27846 -17257
rect 28340 -17375 28374 -17257
rect 27269 -17462 27645 -17428
rect 27905 -17462 28281 -17428
rect 27269 -17730 27645 -17696
rect 27905 -17730 28281 -17696
rect 27176 -18488 27210 -17796
rect 27704 -18488 27738 -17796
rect 27812 -18488 27846 -17796
rect 28340 -18488 28374 -17796
rect 27269 -18588 27645 -18554
rect 27905 -18588 28281 -18554
rect 27213 -18722 28337 -18688
rect 28869 -17204 29245 -17170
rect 29505 -17204 29881 -17170
rect 28776 -17375 28810 -17257
rect 29304 -17375 29338 -17257
rect 29412 -17375 29446 -17257
rect 29940 -17375 29974 -17257
rect 28869 -17462 29245 -17428
rect 29505 -17462 29881 -17428
rect 28869 -17730 29245 -17696
rect 29505 -17730 29881 -17696
rect 28776 -18488 28810 -17796
rect 29304 -18488 29338 -17796
rect 29412 -18488 29446 -17796
rect 29940 -18488 29974 -17796
rect 28869 -18588 29245 -18554
rect 29505 -18588 29881 -18554
rect 28813 -18722 29937 -18688
rect 30469 -17204 30845 -17170
rect 31105 -17204 31481 -17170
rect 30376 -17375 30410 -17257
rect 30904 -17375 30938 -17257
rect 31012 -17375 31046 -17257
rect 31540 -17375 31574 -17257
rect 30469 -17462 30845 -17428
rect 31105 -17462 31481 -17428
rect 30469 -17730 30845 -17696
rect 31105 -17730 31481 -17696
rect 30376 -18488 30410 -17796
rect 30904 -18488 30938 -17796
rect 31012 -18488 31046 -17796
rect 31540 -18488 31574 -17796
rect 30469 -18588 30845 -18554
rect 31105 -18588 31481 -18554
rect 30413 -18722 31537 -18688
rect 32069 -17204 32445 -17170
rect 32705 -17204 33081 -17170
rect 31976 -17375 32010 -17257
rect 32504 -17375 32538 -17257
rect 32612 -17375 32646 -17257
rect 33140 -17375 33174 -17257
rect 32069 -17462 32445 -17428
rect 32705 -17462 33081 -17428
rect 32069 -17730 32445 -17696
rect 32705 -17730 33081 -17696
rect 31976 -18488 32010 -17796
rect 32504 -18488 32538 -17796
rect 32612 -18488 32646 -17796
rect 33140 -18488 33174 -17796
rect 32069 -18588 32445 -18554
rect 32705 -18588 33081 -18554
rect 32013 -18722 33137 -18688
rect 33669 -17204 34045 -17170
rect 34305 -17204 34681 -17170
rect 33576 -17375 33610 -17257
rect 34104 -17375 34138 -17257
rect 34212 -17375 34246 -17257
rect 34740 -17375 34774 -17257
rect 33669 -17462 34045 -17428
rect 34305 -17462 34681 -17428
rect 33669 -17730 34045 -17696
rect 34305 -17730 34681 -17696
rect 33576 -18488 33610 -17796
rect 34104 -18488 34138 -17796
rect 34212 -18488 34246 -17796
rect 34740 -18488 34774 -17796
rect 33669 -18588 34045 -18554
rect 34305 -18588 34681 -18554
rect 33613 -18722 34737 -18688
rect 35269 -17204 35645 -17170
rect 35905 -17204 36281 -17170
rect 35176 -17375 35210 -17257
rect 35704 -17375 35738 -17257
rect 35812 -17375 35846 -17257
rect 36340 -17375 36374 -17257
rect 35269 -17462 35645 -17428
rect 35905 -17462 36281 -17428
rect 36869 -17204 37245 -17170
rect 37505 -17204 37881 -17170
rect 36776 -17375 36810 -17257
rect 37304 -17375 37338 -17257
rect 37412 -17375 37446 -17257
rect 37940 -17375 37974 -17257
rect 36869 -17462 37245 -17428
rect 37505 -17462 37881 -17428
rect 35269 -17730 35645 -17696
rect 35905 -17730 36281 -17696
rect 35176 -18488 35210 -17796
rect 35704 -18488 35738 -17796
rect 35812 -18488 35846 -17796
rect 36340 -18488 36374 -17796
rect 35269 -18588 35645 -18554
rect 35905 -18588 36281 -18554
rect 36869 -17730 37245 -17696
rect 37505 -17730 37881 -17696
rect 36776 -18488 36810 -17796
rect 37304 -18488 37338 -17796
rect 37412 -18488 37446 -17796
rect 37940 -18488 37974 -17796
rect 36869 -18588 37245 -18554
rect 37505 -18588 37881 -18554
rect 35213 -18722 36337 -18688
rect 36813 -18722 37937 -18688
rect 69 -19004 445 -18970
rect 705 -19004 1081 -18970
rect -24 -19175 10 -19057
rect 504 -19175 538 -19057
rect 612 -19175 646 -19057
rect 1140 -19175 1174 -19057
rect 69 -19262 445 -19228
rect 705 -19262 1081 -19228
rect 1669 -19004 2045 -18970
rect 2305 -19004 2681 -18970
rect 1576 -19175 1610 -19057
rect 2104 -19175 2138 -19057
rect 2212 -19175 2246 -19057
rect 2740 -19175 2774 -19057
rect 1669 -19262 2045 -19228
rect 2305 -19262 2681 -19228
rect 69 -19530 445 -19496
rect 705 -19530 1081 -19496
rect -24 -20288 10 -19596
rect 504 -20288 538 -19596
rect 612 -20288 646 -19596
rect 1140 -20288 1174 -19596
rect 69 -20388 445 -20354
rect 705 -20388 1081 -20354
rect 1669 -19530 2045 -19496
rect 2305 -19530 2681 -19496
rect 1576 -20288 1610 -19596
rect 2104 -20288 2138 -19596
rect 2212 -20288 2246 -19596
rect 2740 -20288 2774 -19596
rect 1669 -20388 2045 -20354
rect 2305 -20388 2681 -20354
rect 13 -20522 1137 -20488
rect 1613 -20522 2737 -20488
rect 3269 -19004 3645 -18970
rect 3905 -19004 4281 -18970
rect 3176 -19175 3210 -19057
rect 3704 -19175 3738 -19057
rect 3812 -19175 3846 -19057
rect 4340 -19175 4374 -19057
rect 3269 -19262 3645 -19228
rect 3905 -19262 4281 -19228
rect 3269 -19530 3645 -19496
rect 3905 -19530 4281 -19496
rect 3176 -20288 3210 -19596
rect 3704 -20288 3738 -19596
rect 3812 -20288 3846 -19596
rect 4340 -20288 4374 -19596
rect 3269 -20388 3645 -20354
rect 3905 -20388 4281 -20354
rect 3213 -20522 4337 -20488
rect 4869 -19004 5245 -18970
rect 5505 -19004 5881 -18970
rect 4776 -19175 4810 -19057
rect 5304 -19175 5338 -19057
rect 5412 -19175 5446 -19057
rect 5940 -19175 5974 -19057
rect 4869 -19262 5245 -19228
rect 5505 -19262 5881 -19228
rect 4869 -19530 5245 -19496
rect 5505 -19530 5881 -19496
rect 4776 -20288 4810 -19596
rect 5304 -20288 5338 -19596
rect 5412 -20288 5446 -19596
rect 5940 -20288 5974 -19596
rect 4869 -20388 5245 -20354
rect 5505 -20388 5881 -20354
rect 4813 -20522 5937 -20488
rect 6469 -19004 6845 -18970
rect 7105 -19004 7481 -18970
rect 6376 -19175 6410 -19057
rect 6904 -19175 6938 -19057
rect 7012 -19175 7046 -19057
rect 7540 -19175 7574 -19057
rect 6469 -19262 6845 -19228
rect 7105 -19262 7481 -19228
rect 6469 -19530 6845 -19496
rect 7105 -19530 7481 -19496
rect 6376 -20288 6410 -19596
rect 6904 -20288 6938 -19596
rect 7012 -20288 7046 -19596
rect 7540 -20288 7574 -19596
rect 6469 -20388 6845 -20354
rect 7105 -20388 7481 -20354
rect 6413 -20522 7537 -20488
rect 8069 -19004 8445 -18970
rect 8705 -19004 9081 -18970
rect 7976 -19175 8010 -19057
rect 8504 -19175 8538 -19057
rect 8612 -19175 8646 -19057
rect 9140 -19175 9174 -19057
rect 8069 -19262 8445 -19228
rect 8705 -19262 9081 -19228
rect 8069 -19530 8445 -19496
rect 8705 -19530 9081 -19496
rect 7976 -20288 8010 -19596
rect 8504 -20288 8538 -19596
rect 8612 -20288 8646 -19596
rect 9140 -20288 9174 -19596
rect 8069 -20388 8445 -20354
rect 8705 -20388 9081 -20354
rect 8013 -20522 9137 -20488
rect 9669 -19004 10045 -18970
rect 10305 -19004 10681 -18970
rect 9576 -19175 9610 -19057
rect 10104 -19175 10138 -19057
rect 10212 -19175 10246 -19057
rect 10740 -19175 10774 -19057
rect 9669 -19262 10045 -19228
rect 10305 -19262 10681 -19228
rect 9669 -19530 10045 -19496
rect 10305 -19530 10681 -19496
rect 9576 -20288 9610 -19596
rect 10104 -20288 10138 -19596
rect 10212 -20288 10246 -19596
rect 10740 -20288 10774 -19596
rect 9669 -20388 10045 -20354
rect 10305 -20388 10681 -20354
rect 9613 -20522 10737 -20488
rect 11269 -19004 11645 -18970
rect 11905 -19004 12281 -18970
rect 11176 -19175 11210 -19057
rect 11704 -19175 11738 -19057
rect 11812 -19175 11846 -19057
rect 12340 -19175 12374 -19057
rect 11269 -19262 11645 -19228
rect 11905 -19262 12281 -19228
rect 11269 -19530 11645 -19496
rect 11905 -19530 12281 -19496
rect 11176 -20288 11210 -19596
rect 11704 -20288 11738 -19596
rect 11812 -20288 11846 -19596
rect 12340 -20288 12374 -19596
rect 11269 -20388 11645 -20354
rect 11905 -20388 12281 -20354
rect 11213 -20522 12337 -20488
rect 12869 -19004 13245 -18970
rect 13505 -19004 13881 -18970
rect 12776 -19175 12810 -19057
rect 13304 -19175 13338 -19057
rect 13412 -19175 13446 -19057
rect 13940 -19175 13974 -19057
rect 12869 -19262 13245 -19228
rect 13505 -19262 13881 -19228
rect 12869 -19530 13245 -19496
rect 13505 -19530 13881 -19496
rect 12776 -20288 12810 -19596
rect 13304 -20288 13338 -19596
rect 13412 -20288 13446 -19596
rect 13940 -20288 13974 -19596
rect 12869 -20388 13245 -20354
rect 13505 -20388 13881 -20354
rect 12813 -20522 13937 -20488
rect 14469 -19004 14845 -18970
rect 15105 -19004 15481 -18970
rect 14376 -19175 14410 -19057
rect 14904 -19175 14938 -19057
rect 15012 -19175 15046 -19057
rect 15540 -19175 15574 -19057
rect 14469 -19262 14845 -19228
rect 15105 -19262 15481 -19228
rect 14469 -19530 14845 -19496
rect 15105 -19530 15481 -19496
rect 14376 -20288 14410 -19596
rect 14904 -20288 14938 -19596
rect 15012 -20288 15046 -19596
rect 15540 -20288 15574 -19596
rect 14469 -20388 14845 -20354
rect 15105 -20388 15481 -20354
rect 14413 -20522 15537 -20488
rect 16069 -19004 16445 -18970
rect 16705 -19004 17081 -18970
rect 15976 -19175 16010 -19057
rect 16504 -19175 16538 -19057
rect 16612 -19175 16646 -19057
rect 17140 -19175 17174 -19057
rect 16069 -19262 16445 -19228
rect 16705 -19262 17081 -19228
rect 16069 -19530 16445 -19496
rect 16705 -19530 17081 -19496
rect 15976 -20288 16010 -19596
rect 16504 -20288 16538 -19596
rect 16612 -20288 16646 -19596
rect 17140 -20288 17174 -19596
rect 16069 -20388 16445 -20354
rect 16705 -20388 17081 -20354
rect 16013 -20522 17137 -20488
rect 17669 -19004 18045 -18970
rect 18305 -19004 18681 -18970
rect 17576 -19175 17610 -19057
rect 18104 -19175 18138 -19057
rect 18212 -19175 18246 -19057
rect 18740 -19175 18774 -19057
rect 17669 -19262 18045 -19228
rect 18305 -19262 18681 -19228
rect 17669 -19530 18045 -19496
rect 18305 -19530 18681 -19496
rect 17576 -20288 17610 -19596
rect 18104 -20288 18138 -19596
rect 18212 -20288 18246 -19596
rect 18740 -20288 18774 -19596
rect 17669 -20388 18045 -20354
rect 18305 -20388 18681 -20354
rect 17613 -20522 18737 -20488
rect 19269 -19004 19645 -18970
rect 19905 -19004 20281 -18970
rect 19176 -19175 19210 -19057
rect 19704 -19175 19738 -19057
rect 19812 -19175 19846 -19057
rect 20340 -19175 20374 -19057
rect 19269 -19262 19645 -19228
rect 19905 -19262 20281 -19228
rect 19269 -19530 19645 -19496
rect 19905 -19530 20281 -19496
rect 19176 -20288 19210 -19596
rect 19704 -20288 19738 -19596
rect 19812 -20288 19846 -19596
rect 20340 -20288 20374 -19596
rect 19269 -20388 19645 -20354
rect 19905 -20388 20281 -20354
rect 19213 -20522 20337 -20488
rect 20869 -19004 21245 -18970
rect 21505 -19004 21881 -18970
rect 20776 -19175 20810 -19057
rect 21304 -19175 21338 -19057
rect 21412 -19175 21446 -19057
rect 21940 -19175 21974 -19057
rect 20869 -19262 21245 -19228
rect 21505 -19262 21881 -19228
rect 20869 -19530 21245 -19496
rect 21505 -19530 21881 -19496
rect 20776 -20288 20810 -19596
rect 21304 -20288 21338 -19596
rect 21412 -20288 21446 -19596
rect 21940 -20288 21974 -19596
rect 20869 -20388 21245 -20354
rect 21505 -20388 21881 -20354
rect 20813 -20522 21937 -20488
rect 22469 -19004 22845 -18970
rect 23105 -19004 23481 -18970
rect 22376 -19175 22410 -19057
rect 22904 -19175 22938 -19057
rect 23012 -19175 23046 -19057
rect 23540 -19175 23574 -19057
rect 22469 -19262 22845 -19228
rect 23105 -19262 23481 -19228
rect 22469 -19530 22845 -19496
rect 23105 -19530 23481 -19496
rect 22376 -20288 22410 -19596
rect 22904 -20288 22938 -19596
rect 23012 -20288 23046 -19596
rect 23540 -20288 23574 -19596
rect 22469 -20388 22845 -20354
rect 23105 -20388 23481 -20354
rect 22413 -20522 23537 -20488
rect 24069 -19004 24445 -18970
rect 24705 -19004 25081 -18970
rect 23976 -19175 24010 -19057
rect 24504 -19175 24538 -19057
rect 24612 -19175 24646 -19057
rect 25140 -19175 25174 -19057
rect 24069 -19262 24445 -19228
rect 24705 -19262 25081 -19228
rect 24069 -19530 24445 -19496
rect 24705 -19530 25081 -19496
rect 23976 -20288 24010 -19596
rect 24504 -20288 24538 -19596
rect 24612 -20288 24646 -19596
rect 25140 -20288 25174 -19596
rect 24069 -20388 24445 -20354
rect 24705 -20388 25081 -20354
rect 24013 -20522 25137 -20488
rect 25669 -19004 26045 -18970
rect 26305 -19004 26681 -18970
rect 25576 -19175 25610 -19057
rect 26104 -19175 26138 -19057
rect 26212 -19175 26246 -19057
rect 26740 -19175 26774 -19057
rect 25669 -19262 26045 -19228
rect 26305 -19262 26681 -19228
rect 25669 -19530 26045 -19496
rect 26305 -19530 26681 -19496
rect 25576 -20288 25610 -19596
rect 26104 -20288 26138 -19596
rect 26212 -20288 26246 -19596
rect 26740 -20288 26774 -19596
rect 25669 -20388 26045 -20354
rect 26305 -20388 26681 -20354
rect 25613 -20522 26737 -20488
rect 27269 -19004 27645 -18970
rect 27905 -19004 28281 -18970
rect 27176 -19175 27210 -19057
rect 27704 -19175 27738 -19057
rect 27812 -19175 27846 -19057
rect 28340 -19175 28374 -19057
rect 27269 -19262 27645 -19228
rect 27905 -19262 28281 -19228
rect 27269 -19530 27645 -19496
rect 27905 -19530 28281 -19496
rect 27176 -20288 27210 -19596
rect 27704 -20288 27738 -19596
rect 27812 -20288 27846 -19596
rect 28340 -20288 28374 -19596
rect 27269 -20388 27645 -20354
rect 27905 -20388 28281 -20354
rect 27213 -20522 28337 -20488
rect 28869 -19004 29245 -18970
rect 29505 -19004 29881 -18970
rect 28776 -19175 28810 -19057
rect 29304 -19175 29338 -19057
rect 29412 -19175 29446 -19057
rect 29940 -19175 29974 -19057
rect 28869 -19262 29245 -19228
rect 29505 -19262 29881 -19228
rect 28869 -19530 29245 -19496
rect 29505 -19530 29881 -19496
rect 28776 -20288 28810 -19596
rect 29304 -20288 29338 -19596
rect 29412 -20288 29446 -19596
rect 29940 -20288 29974 -19596
rect 28869 -20388 29245 -20354
rect 29505 -20388 29881 -20354
rect 28813 -20522 29937 -20488
rect 30469 -19004 30845 -18970
rect 31105 -19004 31481 -18970
rect 30376 -19175 30410 -19057
rect 30904 -19175 30938 -19057
rect 31012 -19175 31046 -19057
rect 31540 -19175 31574 -19057
rect 30469 -19262 30845 -19228
rect 31105 -19262 31481 -19228
rect 30469 -19530 30845 -19496
rect 31105 -19530 31481 -19496
rect 30376 -20288 30410 -19596
rect 30904 -20288 30938 -19596
rect 31012 -20288 31046 -19596
rect 31540 -20288 31574 -19596
rect 30469 -20388 30845 -20354
rect 31105 -20388 31481 -20354
rect 30413 -20522 31537 -20488
rect 32069 -19004 32445 -18970
rect 32705 -19004 33081 -18970
rect 31976 -19175 32010 -19057
rect 32504 -19175 32538 -19057
rect 32612 -19175 32646 -19057
rect 33140 -19175 33174 -19057
rect 32069 -19262 32445 -19228
rect 32705 -19262 33081 -19228
rect 32069 -19530 32445 -19496
rect 32705 -19530 33081 -19496
rect 31976 -20288 32010 -19596
rect 32504 -20288 32538 -19596
rect 32612 -20288 32646 -19596
rect 33140 -20288 33174 -19596
rect 32069 -20388 32445 -20354
rect 32705 -20388 33081 -20354
rect 32013 -20522 33137 -20488
rect 33669 -19004 34045 -18970
rect 34305 -19004 34681 -18970
rect 33576 -19175 33610 -19057
rect 34104 -19175 34138 -19057
rect 34212 -19175 34246 -19057
rect 34740 -19175 34774 -19057
rect 33669 -19262 34045 -19228
rect 34305 -19262 34681 -19228
rect 33669 -19530 34045 -19496
rect 34305 -19530 34681 -19496
rect 33576 -20288 33610 -19596
rect 34104 -20288 34138 -19596
rect 34212 -20288 34246 -19596
rect 34740 -20288 34774 -19596
rect 33669 -20388 34045 -20354
rect 34305 -20388 34681 -20354
rect 33613 -20522 34737 -20488
rect 35269 -19004 35645 -18970
rect 35905 -19004 36281 -18970
rect 35176 -19175 35210 -19057
rect 35704 -19175 35738 -19057
rect 35812 -19175 35846 -19057
rect 36340 -19175 36374 -19057
rect 35269 -19262 35645 -19228
rect 35905 -19262 36281 -19228
rect 36869 -19004 37245 -18970
rect 37505 -19004 37881 -18970
rect 36776 -19175 36810 -19057
rect 37304 -19175 37338 -19057
rect 37412 -19175 37446 -19057
rect 37940 -19175 37974 -19057
rect 36869 -19262 37245 -19228
rect 37505 -19262 37881 -19228
rect 35269 -19530 35645 -19496
rect 35905 -19530 36281 -19496
rect 35176 -20288 35210 -19596
rect 35704 -20288 35738 -19596
rect 35812 -20288 35846 -19596
rect 36340 -20288 36374 -19596
rect 35269 -20388 35645 -20354
rect 35905 -20388 36281 -20354
rect 36869 -19530 37245 -19496
rect 37505 -19530 37881 -19496
rect 36776 -20288 36810 -19596
rect 37304 -20288 37338 -19596
rect 37412 -20288 37446 -19596
rect 37940 -20288 37974 -19596
rect 36869 -20388 37245 -20354
rect 37505 -20388 37881 -20354
rect 35213 -20522 36337 -20488
rect 36813 -20522 37937 -20488
rect 69 -20804 445 -20770
rect 705 -20804 1081 -20770
rect -24 -20975 10 -20857
rect 504 -20975 538 -20857
rect 612 -20975 646 -20857
rect 1140 -20975 1174 -20857
rect 69 -21062 445 -21028
rect 705 -21062 1081 -21028
rect 1669 -20804 2045 -20770
rect 2305 -20804 2681 -20770
rect 1576 -20975 1610 -20857
rect 2104 -20975 2138 -20857
rect 2212 -20975 2246 -20857
rect 2740 -20975 2774 -20857
rect 1669 -21062 2045 -21028
rect 2305 -21062 2681 -21028
rect 69 -21330 445 -21296
rect 705 -21330 1081 -21296
rect -24 -22088 10 -21396
rect 504 -22088 538 -21396
rect 612 -22088 646 -21396
rect 1140 -22088 1174 -21396
rect 69 -22188 445 -22154
rect 705 -22188 1081 -22154
rect 1669 -21330 2045 -21296
rect 2305 -21330 2681 -21296
rect 1576 -22088 1610 -21396
rect 2104 -22088 2138 -21396
rect 2212 -22088 2246 -21396
rect 2740 -22088 2774 -21396
rect 1669 -22188 2045 -22154
rect 2305 -22188 2681 -22154
rect 13 -22322 1137 -22288
rect 1613 -22322 2737 -22288
rect 3269 -20804 3645 -20770
rect 3905 -20804 4281 -20770
rect 3176 -20975 3210 -20857
rect 3704 -20975 3738 -20857
rect 3812 -20975 3846 -20857
rect 4340 -20975 4374 -20857
rect 3269 -21062 3645 -21028
rect 3905 -21062 4281 -21028
rect 3269 -21330 3645 -21296
rect 3905 -21330 4281 -21296
rect 3176 -22088 3210 -21396
rect 3704 -22088 3738 -21396
rect 3812 -22088 3846 -21396
rect 4340 -22088 4374 -21396
rect 3269 -22188 3645 -22154
rect 3905 -22188 4281 -22154
rect 4869 -20804 5245 -20770
rect 5505 -20804 5881 -20770
rect 4776 -20975 4810 -20857
rect 5304 -20975 5338 -20857
rect 5412 -20975 5446 -20857
rect 5940 -20975 5974 -20857
rect 4869 -21062 5245 -21028
rect 5505 -21062 5881 -21028
rect 4869 -21330 5245 -21296
rect 5505 -21330 5881 -21296
rect 4776 -22088 4810 -21396
rect 5304 -22088 5338 -21396
rect 5412 -22088 5446 -21396
rect 5940 -22088 5974 -21396
rect 4869 -22188 5245 -22154
rect 5505 -22188 5881 -22154
rect 6469 -20804 6845 -20770
rect 7105 -20804 7481 -20770
rect 6376 -20975 6410 -20857
rect 6904 -20975 6938 -20857
rect 7012 -20975 7046 -20857
rect 7540 -20975 7574 -20857
rect 6469 -21062 6845 -21028
rect 7105 -21062 7481 -21028
rect 6469 -21330 6845 -21296
rect 7105 -21330 7481 -21296
rect 6376 -22088 6410 -21396
rect 6904 -22088 6938 -21396
rect 7012 -22088 7046 -21396
rect 7540 -22088 7574 -21396
rect 6469 -22188 6845 -22154
rect 7105 -22188 7481 -22154
rect 8069 -20804 8445 -20770
rect 8705 -20804 9081 -20770
rect 7976 -20975 8010 -20857
rect 8504 -20975 8538 -20857
rect 8612 -20975 8646 -20857
rect 9140 -20975 9174 -20857
rect 8069 -21062 8445 -21028
rect 8705 -21062 9081 -21028
rect 8069 -21330 8445 -21296
rect 8705 -21330 9081 -21296
rect 7976 -22088 8010 -21396
rect 8504 -22088 8538 -21396
rect 8612 -22088 8646 -21396
rect 9140 -22088 9174 -21396
rect 8069 -22188 8445 -22154
rect 8705 -22188 9081 -22154
rect 9669 -20804 10045 -20770
rect 10305 -20804 10681 -20770
rect 9576 -20975 9610 -20857
rect 10104 -20975 10138 -20857
rect 10212 -20975 10246 -20857
rect 10740 -20975 10774 -20857
rect 9669 -21062 10045 -21028
rect 10305 -21062 10681 -21028
rect 9669 -21330 10045 -21296
rect 10305 -21330 10681 -21296
rect 9576 -22088 9610 -21396
rect 10104 -22088 10138 -21396
rect 10212 -22088 10246 -21396
rect 10740 -22088 10774 -21396
rect 9669 -22188 10045 -22154
rect 10305 -22188 10681 -22154
rect 11269 -20804 11645 -20770
rect 11905 -20804 12281 -20770
rect 11176 -20975 11210 -20857
rect 11704 -20975 11738 -20857
rect 11812 -20975 11846 -20857
rect 12340 -20975 12374 -20857
rect 11269 -21062 11645 -21028
rect 11905 -21062 12281 -21028
rect 11269 -21330 11645 -21296
rect 11905 -21330 12281 -21296
rect 11176 -22088 11210 -21396
rect 11704 -22088 11738 -21396
rect 11812 -22088 11846 -21396
rect 12340 -22088 12374 -21396
rect 11269 -22188 11645 -22154
rect 11905 -22188 12281 -22154
rect 12869 -20804 13245 -20770
rect 13505 -20804 13881 -20770
rect 12776 -20975 12810 -20857
rect 13304 -20975 13338 -20857
rect 13412 -20975 13446 -20857
rect 13940 -20975 13974 -20857
rect 12869 -21062 13245 -21028
rect 13505 -21062 13881 -21028
rect 12869 -21330 13245 -21296
rect 13505 -21330 13881 -21296
rect 12776 -22088 12810 -21396
rect 13304 -22088 13338 -21396
rect 13412 -22088 13446 -21396
rect 13940 -22088 13974 -21396
rect 12869 -22188 13245 -22154
rect 13505 -22188 13881 -22154
rect 14469 -20804 14845 -20770
rect 15105 -20804 15481 -20770
rect 14376 -20975 14410 -20857
rect 14904 -20975 14938 -20857
rect 15012 -20975 15046 -20857
rect 15540 -20975 15574 -20857
rect 14469 -21062 14845 -21028
rect 15105 -21062 15481 -21028
rect 14469 -21330 14845 -21296
rect 15105 -21330 15481 -21296
rect 14376 -22088 14410 -21396
rect 14904 -22088 14938 -21396
rect 15012 -22088 15046 -21396
rect 15540 -22088 15574 -21396
rect 14469 -22188 14845 -22154
rect 15105 -22188 15481 -22154
rect 16069 -20804 16445 -20770
rect 16705 -20804 17081 -20770
rect 15976 -20975 16010 -20857
rect 16504 -20975 16538 -20857
rect 16612 -20975 16646 -20857
rect 17140 -20975 17174 -20857
rect 16069 -21062 16445 -21028
rect 16705 -21062 17081 -21028
rect 16069 -21330 16445 -21296
rect 16705 -21330 17081 -21296
rect 15976 -22088 16010 -21396
rect 16504 -22088 16538 -21396
rect 16612 -22088 16646 -21396
rect 17140 -22088 17174 -21396
rect 16069 -22188 16445 -22154
rect 16705 -22188 17081 -22154
rect 17669 -20804 18045 -20770
rect 18305 -20804 18681 -20770
rect 17576 -20975 17610 -20857
rect 18104 -20975 18138 -20857
rect 18212 -20975 18246 -20857
rect 18740 -20975 18774 -20857
rect 17669 -21062 18045 -21028
rect 18305 -21062 18681 -21028
rect 17669 -21330 18045 -21296
rect 18305 -21330 18681 -21296
rect 17576 -22088 17610 -21396
rect 18104 -22088 18138 -21396
rect 18212 -22088 18246 -21396
rect 18740 -22088 18774 -21396
rect 17669 -22188 18045 -22154
rect 18305 -22188 18681 -22154
rect 19269 -20804 19645 -20770
rect 19905 -20804 20281 -20770
rect 19176 -20975 19210 -20857
rect 19704 -20975 19738 -20857
rect 19812 -20975 19846 -20857
rect 20340 -20975 20374 -20857
rect 19269 -21062 19645 -21028
rect 19905 -21062 20281 -21028
rect 19269 -21330 19645 -21296
rect 19905 -21330 20281 -21296
rect 19176 -22088 19210 -21396
rect 19704 -22088 19738 -21396
rect 19812 -22088 19846 -21396
rect 20340 -22088 20374 -21396
rect 19269 -22188 19645 -22154
rect 19905 -22188 20281 -22154
rect 20869 -20804 21245 -20770
rect 21505 -20804 21881 -20770
rect 20776 -20975 20810 -20857
rect 21304 -20975 21338 -20857
rect 21412 -20975 21446 -20857
rect 21940 -20975 21974 -20857
rect 20869 -21062 21245 -21028
rect 21505 -21062 21881 -21028
rect 20869 -21330 21245 -21296
rect 21505 -21330 21881 -21296
rect 20776 -22088 20810 -21396
rect 21304 -22088 21338 -21396
rect 21412 -22088 21446 -21396
rect 21940 -22088 21974 -21396
rect 20869 -22188 21245 -22154
rect 21505 -22188 21881 -22154
rect 3213 -22322 4337 -22288
rect 4813 -22322 5937 -22288
rect 6413 -22322 7537 -22288
rect 8013 -22322 9137 -22288
rect 9613 -22322 10737 -22288
rect 11213 -22322 12337 -22288
rect 12813 -22322 13937 -22288
rect 14413 -22322 15537 -22288
rect 16013 -22322 17137 -22288
rect 17613 -22322 18737 -22288
rect 19213 -22322 20337 -22288
rect 20813 -22322 21937 -22288
rect 22469 -20804 22845 -20770
rect 23105 -20804 23481 -20770
rect 22376 -20975 22410 -20857
rect 22904 -20975 22938 -20857
rect 23012 -20975 23046 -20857
rect 23540 -20975 23574 -20857
rect 22469 -21062 22845 -21028
rect 23105 -21062 23481 -21028
rect 22469 -21330 22845 -21296
rect 23105 -21330 23481 -21296
rect 22376 -22088 22410 -21396
rect 22904 -22088 22938 -21396
rect 23012 -22088 23046 -21396
rect 23540 -22088 23574 -21396
rect 22469 -22188 22845 -22154
rect 23105 -22188 23481 -22154
rect 22413 -22322 23537 -22288
rect 24069 -20804 24445 -20770
rect 24705 -20804 25081 -20770
rect 23976 -20975 24010 -20857
rect 24504 -20975 24538 -20857
rect 24612 -20975 24646 -20857
rect 25140 -20975 25174 -20857
rect 24069 -21062 24445 -21028
rect 24705 -21062 25081 -21028
rect 24069 -21330 24445 -21296
rect 24705 -21330 25081 -21296
rect 23976 -22088 24010 -21396
rect 24504 -22088 24538 -21396
rect 24612 -22088 24646 -21396
rect 25140 -22088 25174 -21396
rect 24069 -22188 24445 -22154
rect 24705 -22188 25081 -22154
rect 24013 -22322 25137 -22288
rect 25669 -20804 26045 -20770
rect 26305 -20804 26681 -20770
rect 25576 -20975 25610 -20857
rect 26104 -20975 26138 -20857
rect 26212 -20975 26246 -20857
rect 26740 -20975 26774 -20857
rect 25669 -21062 26045 -21028
rect 26305 -21062 26681 -21028
rect 25669 -21330 26045 -21296
rect 26305 -21330 26681 -21296
rect 25576 -22088 25610 -21396
rect 26104 -22088 26138 -21396
rect 26212 -22088 26246 -21396
rect 26740 -22088 26774 -21396
rect 25669 -22188 26045 -22154
rect 26305 -22188 26681 -22154
rect 25613 -22322 26737 -22288
rect 27269 -20804 27645 -20770
rect 27905 -20804 28281 -20770
rect 27176 -20975 27210 -20857
rect 27704 -20975 27738 -20857
rect 27812 -20975 27846 -20857
rect 28340 -20975 28374 -20857
rect 27269 -21062 27645 -21028
rect 27905 -21062 28281 -21028
rect 27269 -21330 27645 -21296
rect 27905 -21330 28281 -21296
rect 27176 -22088 27210 -21396
rect 27704 -22088 27738 -21396
rect 27812 -22088 27846 -21396
rect 28340 -22088 28374 -21396
rect 27269 -22188 27645 -22154
rect 27905 -22188 28281 -22154
rect 27213 -22322 28337 -22288
rect 28869 -20804 29245 -20770
rect 29505 -20804 29881 -20770
rect 28776 -20975 28810 -20857
rect 29304 -20975 29338 -20857
rect 29412 -20975 29446 -20857
rect 29940 -20975 29974 -20857
rect 28869 -21062 29245 -21028
rect 29505 -21062 29881 -21028
rect 28869 -21330 29245 -21296
rect 29505 -21330 29881 -21296
rect 28776 -22088 28810 -21396
rect 29304 -22088 29338 -21396
rect 29412 -22088 29446 -21396
rect 29940 -22088 29974 -21396
rect 28869 -22188 29245 -22154
rect 29505 -22188 29881 -22154
rect 28813 -22322 29937 -22288
rect 30469 -20804 30845 -20770
rect 31105 -20804 31481 -20770
rect 30376 -20975 30410 -20857
rect 30904 -20975 30938 -20857
rect 31012 -20975 31046 -20857
rect 31540 -20975 31574 -20857
rect 30469 -21062 30845 -21028
rect 31105 -21062 31481 -21028
rect 30469 -21330 30845 -21296
rect 31105 -21330 31481 -21296
rect 30376 -22088 30410 -21396
rect 30904 -22088 30938 -21396
rect 31012 -22088 31046 -21396
rect 31540 -22088 31574 -21396
rect 30469 -22188 30845 -22154
rect 31105 -22188 31481 -22154
rect 30413 -22322 31537 -22288
rect 32069 -20804 32445 -20770
rect 32705 -20804 33081 -20770
rect 31976 -20975 32010 -20857
rect 32504 -20975 32538 -20857
rect 32612 -20975 32646 -20857
rect 33140 -20975 33174 -20857
rect 32069 -21062 32445 -21028
rect 32705 -21062 33081 -21028
rect 32069 -21330 32445 -21296
rect 32705 -21330 33081 -21296
rect 31976 -22088 32010 -21396
rect 32504 -22088 32538 -21396
rect 32612 -22088 32646 -21396
rect 33140 -22088 33174 -21396
rect 32069 -22188 32445 -22154
rect 32705 -22188 33081 -22154
rect 32013 -22322 33137 -22288
rect 33669 -20804 34045 -20770
rect 34305 -20804 34681 -20770
rect 33576 -20975 33610 -20857
rect 34104 -20975 34138 -20857
rect 34212 -20975 34246 -20857
rect 34740 -20975 34774 -20857
rect 33669 -21062 34045 -21028
rect 34305 -21062 34681 -21028
rect 33669 -21330 34045 -21296
rect 34305 -21330 34681 -21296
rect 33576 -22088 33610 -21396
rect 34104 -22088 34138 -21396
rect 34212 -22088 34246 -21396
rect 34740 -22088 34774 -21396
rect 33669 -22188 34045 -22154
rect 34305 -22188 34681 -22154
rect 33613 -22322 34737 -22288
rect 35269 -20804 35645 -20770
rect 35905 -20804 36281 -20770
rect 35176 -20975 35210 -20857
rect 35704 -20975 35738 -20857
rect 35812 -20975 35846 -20857
rect 36340 -20975 36374 -20857
rect 35269 -21062 35645 -21028
rect 35905 -21062 36281 -21028
rect 36869 -20804 37245 -20770
rect 37505 -20804 37881 -20770
rect 36776 -20975 36810 -20857
rect 37304 -20975 37338 -20857
rect 37412 -20975 37446 -20857
rect 37940 -20975 37974 -20857
rect 36869 -21062 37245 -21028
rect 37505 -21062 37881 -21028
rect 35269 -21330 35645 -21296
rect 35905 -21330 36281 -21296
rect 35176 -22088 35210 -21396
rect 35704 -22088 35738 -21396
rect 35812 -22088 35846 -21396
rect 36340 -22088 36374 -21396
rect 35269 -22188 35645 -22154
rect 35905 -22188 36281 -22154
rect 36869 -21330 37245 -21296
rect 37505 -21330 37881 -21296
rect 36776 -22088 36810 -21396
rect 37304 -22088 37338 -21396
rect 37412 -22088 37446 -21396
rect 37940 -22088 37974 -21396
rect 36869 -22188 37245 -22154
rect 37505 -22188 37881 -22154
rect 35213 -22322 36337 -22288
rect 36813 -22322 37937 -22288
rect 28352 -23460 28386 -22684
rect 28510 -23460 28544 -22684
rect 28668 -23460 28702 -22684
rect 28826 -23460 28860 -22684
rect 28984 -23460 29018 -22684
rect 28414 -23553 28482 -23519
rect 28572 -23553 28640 -23519
rect 28730 -23553 28798 -23519
rect 28888 -23553 28956 -23519
rect 32498 -23131 32532 -22515
rect 32711 -22576 32745 -22542
rect 32869 -22576 32903 -22542
rect 33027 -22576 33061 -22542
rect 33185 -22576 33219 -22542
rect 32632 -23011 32666 -22635
rect 32790 -23011 32824 -22635
rect 32948 -23011 32982 -22635
rect 33106 -23011 33140 -22635
rect 33264 -23011 33298 -22635
rect 32711 -23104 32745 -23070
rect 32869 -23104 32903 -23070
rect 33027 -23104 33061 -23070
rect 33185 -23104 33219 -23070
rect 33398 -23131 33432 -22515
rect 33868 -23151 33902 -22535
rect 34081 -22596 34115 -22562
rect 34239 -22596 34273 -22562
rect 34002 -23031 34036 -22655
rect 34160 -23031 34194 -22655
rect 34318 -23031 34352 -22655
rect 34081 -23124 34115 -23090
rect 34239 -23124 34273 -23090
rect 32619 -23242 33311 -23208
rect 34452 -23151 34486 -22535
rect 33957 -23262 33964 -23228
rect 33964 -23262 34390 -23228
rect 34390 -23262 34397 -23228
rect 33036 -24273 33070 -23657
rect 33249 -23718 33283 -23684
rect 33407 -23718 33441 -23684
rect 33565 -23718 33599 -23684
rect 33723 -23718 33757 -23684
rect 33881 -23718 33915 -23684
rect 34039 -23718 34073 -23684
rect 33170 -24153 33204 -23777
rect 33328 -24153 33362 -23777
rect 33486 -24153 33520 -23777
rect 33644 -24153 33678 -23777
rect 33802 -24153 33836 -23777
rect 33960 -24153 33994 -23777
rect 34118 -24153 34152 -23777
rect 33249 -24246 33283 -24212
rect 33407 -24246 33441 -24212
rect 33565 -24246 33599 -24212
rect 33723 -24246 33757 -24212
rect 33881 -24246 33915 -24212
rect 34039 -24246 34073 -24212
rect 22470 -24548 26790 -24514
rect 2479 -25140 4055 -25106
rect 2386 -25436 2420 -25168
rect 4114 -25436 4148 -25168
rect 2479 -25498 4055 -25464
rect 4679 -25140 6255 -25106
rect 4586 -25436 4620 -25168
rect 6314 -25436 6348 -25168
rect 4679 -25498 6255 -25464
rect 6879 -25140 8455 -25106
rect 6786 -25436 6820 -25168
rect 8514 -25436 8548 -25168
rect 6879 -25498 8455 -25464
rect 9079 -25140 10655 -25106
rect 8986 -25436 9020 -25168
rect 10714 -25436 10748 -25168
rect 9079 -25498 10655 -25464
rect 11279 -25140 12855 -25106
rect 11186 -25436 11220 -25168
rect 12914 -25436 12948 -25168
rect 11279 -25498 12855 -25464
rect 13479 -25140 15055 -25106
rect 13386 -25436 13420 -25168
rect 15114 -25436 15148 -25168
rect 13479 -25498 15055 -25464
rect 15679 -25140 17255 -25106
rect 15586 -25436 15620 -25168
rect 17314 -25436 17348 -25168
rect 15679 -25498 17255 -25464
rect 17879 -25140 19455 -25106
rect 17786 -25436 17820 -25168
rect 19514 -25436 19548 -25168
rect 17879 -25498 19455 -25464
rect 2479 -25940 4055 -25906
rect 2386 -26236 2420 -25968
rect 4114 -26236 4148 -25968
rect 2479 -26298 4055 -26264
rect 4679 -25940 6255 -25906
rect 4586 -26236 4620 -25968
rect 6314 -26236 6348 -25968
rect 4679 -26298 6255 -26264
rect 6879 -25940 8455 -25906
rect 6786 -26236 6820 -25968
rect 8514 -26236 8548 -25968
rect 6879 -26298 8455 -26264
rect 9079 -25940 10655 -25906
rect 8986 -26236 9020 -25968
rect 10714 -26236 10748 -25968
rect 9079 -26298 10655 -26264
rect 11279 -25940 12855 -25906
rect 11186 -26236 11220 -25968
rect 12914 -26236 12948 -25968
rect 11279 -26298 12855 -26264
rect 13479 -25940 15055 -25906
rect 13386 -26236 13420 -25968
rect 15114 -26236 15148 -25968
rect 13479 -26298 15055 -26264
rect 15679 -25940 17255 -25906
rect 15586 -26236 15620 -25968
rect 17314 -26236 17348 -25968
rect 15679 -26298 17255 -26264
rect 17879 -25940 19455 -25906
rect 17786 -26236 17820 -25968
rect 19514 -26236 19548 -25968
rect 17879 -26298 19455 -26264
rect 2479 -26740 4055 -26706
rect 2386 -27036 2420 -26768
rect 4114 -27036 4148 -26768
rect 2479 -27098 4055 -27064
rect 4679 -26740 6255 -26706
rect 4586 -27036 4620 -26768
rect 6314 -27036 6348 -26768
rect 4679 -27098 6255 -27064
rect 6879 -26740 8455 -26706
rect 6786 -27036 6820 -26768
rect 8514 -27036 8548 -26768
rect 6879 -27098 8455 -27064
rect 9079 -26740 10655 -26706
rect 8986 -27036 9020 -26768
rect 10714 -27036 10748 -26768
rect 9079 -27098 10655 -27064
rect 11279 -26740 12855 -26706
rect 11186 -27036 11220 -26768
rect 12914 -27036 12948 -26768
rect 11279 -27098 12855 -27064
rect 13479 -26740 15055 -26706
rect 13386 -27036 13420 -26768
rect 15114 -27036 15148 -26768
rect 13479 -27098 15055 -27064
rect 15679 -26740 17255 -26706
rect 15586 -27036 15620 -26768
rect 17314 -27036 17348 -26768
rect 15679 -27098 17255 -27064
rect 17879 -26740 19455 -26706
rect 17786 -27036 17820 -26768
rect 19514 -27036 19548 -26768
rect 17879 -27098 19455 -27064
rect 2479 -27540 4055 -27506
rect 2386 -27836 2420 -27568
rect 4114 -27836 4148 -27568
rect 2479 -27898 4055 -27864
rect 4679 -27540 6255 -27506
rect 4586 -27836 4620 -27568
rect 6314 -27836 6348 -27568
rect 4679 -27898 6255 -27864
rect 6879 -27540 8455 -27506
rect 6786 -27836 6820 -27568
rect 8514 -27836 8548 -27568
rect 6879 -27898 8455 -27864
rect 9079 -27540 10655 -27506
rect 8986 -27836 9020 -27568
rect 10714 -27836 10748 -27568
rect 9079 -27898 10655 -27864
rect 11279 -27540 12855 -27506
rect 11186 -27836 11220 -27568
rect 12914 -27836 12948 -27568
rect 11279 -27898 12855 -27864
rect 13479 -27540 15055 -27506
rect 13386 -27836 13420 -27568
rect 15114 -27836 15148 -27568
rect 13479 -27898 15055 -27864
rect 15679 -27540 17255 -27506
rect 15586 -27836 15620 -27568
rect 17314 -27836 17348 -27568
rect 15679 -27898 17255 -27864
rect 17879 -27540 19455 -27506
rect 17786 -27836 17820 -27568
rect 19514 -27836 19548 -27568
rect 17879 -27898 19455 -27864
rect 2479 -28340 4055 -28306
rect 2386 -28636 2420 -28368
rect 4114 -28636 4148 -28368
rect 2479 -28698 4055 -28664
rect 4679 -28340 6255 -28306
rect 4586 -28636 4620 -28368
rect 6314 -28636 6348 -28368
rect 4679 -28698 6255 -28664
rect 6879 -28340 8455 -28306
rect 6786 -28636 6820 -28368
rect 8514 -28636 8548 -28368
rect 6879 -28698 8455 -28664
rect 9079 -28340 10655 -28306
rect 8986 -28636 9020 -28368
rect 10714 -28636 10748 -28368
rect 9079 -28698 10655 -28664
rect 11279 -28340 12855 -28306
rect 11186 -28636 11220 -28368
rect 12914 -28636 12948 -28368
rect 11279 -28698 12855 -28664
rect 13479 -28340 15055 -28306
rect 13386 -28636 13420 -28368
rect 15114 -28636 15148 -28368
rect 13479 -28698 15055 -28664
rect 15679 -28340 17255 -28306
rect 15586 -28636 15620 -28368
rect 17314 -28636 17348 -28368
rect 15679 -28698 17255 -28664
rect 17879 -28340 19455 -28306
rect 17786 -28636 17820 -28368
rect 19514 -28636 19548 -28368
rect 17879 -28698 19455 -28664
rect 2479 -29140 4055 -29106
rect 2386 -29436 2420 -29168
rect 4114 -29436 4148 -29168
rect 2479 -29498 4055 -29464
rect 4679 -29140 6255 -29106
rect 4586 -29436 4620 -29168
rect 6314 -29436 6348 -29168
rect 4679 -29498 6255 -29464
rect 6879 -29140 8455 -29106
rect 6786 -29436 6820 -29168
rect 8514 -29436 8548 -29168
rect 6879 -29498 8455 -29464
rect 9079 -29140 10655 -29106
rect 8986 -29436 9020 -29168
rect 10714 -29436 10748 -29168
rect 9079 -29498 10655 -29464
rect 11279 -29140 12855 -29106
rect 11186 -29436 11220 -29168
rect 12914 -29436 12948 -29168
rect 11279 -29498 12855 -29464
rect 13479 -29140 15055 -29106
rect 13386 -29436 13420 -29168
rect 15114 -29436 15148 -29168
rect 13479 -29498 15055 -29464
rect 15679 -29140 17255 -29106
rect 15586 -29436 15620 -29168
rect 17314 -29436 17348 -29168
rect 15679 -29498 17255 -29464
rect 17879 -29140 19455 -29106
rect 17786 -29436 17820 -29168
rect 19514 -29436 19548 -29168
rect 17879 -29498 19455 -29464
rect 2479 -29940 4055 -29906
rect 2386 -30236 2420 -29968
rect 4114 -30236 4148 -29968
rect 2479 -30298 4055 -30264
rect 4679 -29940 6255 -29906
rect 4586 -30236 4620 -29968
rect 6314 -30236 6348 -29968
rect 4679 -30298 6255 -30264
rect 6879 -29940 8455 -29906
rect 6786 -30236 6820 -29968
rect 8514 -30236 8548 -29968
rect 6879 -30298 8455 -30264
rect 9079 -29940 10655 -29906
rect 8986 -30236 9020 -29968
rect 10714 -30236 10748 -29968
rect 9079 -30298 10655 -30264
rect 11279 -29940 12855 -29906
rect 11186 -30236 11220 -29968
rect 12914 -30236 12948 -29968
rect 11279 -30298 12855 -30264
rect 13479 -29940 15055 -29906
rect 13386 -30236 13420 -29968
rect 15114 -30236 15148 -29968
rect 13479 -30298 15055 -30264
rect 15679 -29940 17255 -29906
rect 15586 -30236 15620 -29968
rect 17314 -30236 17348 -29968
rect 15679 -30298 17255 -30264
rect 17879 -29940 19455 -29906
rect 17786 -30236 17820 -29968
rect 19514 -30236 19548 -29968
rect 17879 -30298 19455 -30264
rect 2479 -30740 4055 -30706
rect 2386 -31036 2420 -30768
rect 4114 -31036 4148 -30768
rect 2479 -31098 4055 -31064
rect 4679 -30740 6255 -30706
rect 4586 -31036 4620 -30768
rect 6314 -31036 6348 -30768
rect 4679 -31098 6255 -31064
rect 6879 -30740 8455 -30706
rect 6786 -31036 6820 -30768
rect 8514 -31036 8548 -30768
rect 6879 -31098 8455 -31064
rect 9079 -30740 10655 -30706
rect 8986 -31036 9020 -30768
rect 10714 -31036 10748 -30768
rect 9079 -31098 10655 -31064
rect 11279 -30740 12855 -30706
rect 11186 -31036 11220 -30768
rect 12914 -31036 12948 -30768
rect 11279 -31098 12855 -31064
rect 13479 -30740 15055 -30706
rect 13386 -31036 13420 -30768
rect 15114 -31036 15148 -30768
rect 13479 -31098 15055 -31064
rect 15679 -30740 17255 -30706
rect 15586 -31036 15620 -30768
rect 17314 -31036 17348 -30768
rect 15679 -31098 17255 -31064
rect 17879 -30740 19455 -30706
rect 17786 -31036 17820 -30768
rect 19514 -31036 19548 -30768
rect 17879 -31098 19455 -31064
rect 22196 -31656 22230 -24922
rect 22363 -25080 22901 -24683
rect 23029 -25080 23567 -24683
rect 23695 -25080 24233 -24683
rect 24361 -25080 24899 -24683
rect 25027 -25080 25565 -24683
rect 25693 -25080 26231 -24683
rect 26359 -25080 26897 -24683
rect 22363 -31895 22901 -31498
rect 23029 -31895 23567 -31498
rect 23695 -31895 24233 -31498
rect 24361 -31895 24899 -31498
rect 25027 -31895 25565 -31498
rect 25693 -31895 26231 -31498
rect 26359 -31895 26897 -31498
rect 27030 -31656 27064 -24922
rect 22470 -32064 26790 -32030
rect 34252 -24273 34286 -23657
rect 33188 -24384 34134 -24350
rect 34408 -24271 34442 -23655
rect 34621 -23716 34655 -23682
rect 34779 -23716 34813 -23682
rect 34937 -23716 34971 -23682
rect 35095 -23716 35129 -23682
rect 35253 -23716 35287 -23682
rect 35411 -23716 35445 -23682
rect 35569 -23716 35603 -23682
rect 35727 -23716 35761 -23682
rect 35885 -23716 35919 -23682
rect 36043 -23716 36077 -23682
rect 36201 -23716 36235 -23682
rect 36359 -23716 36393 -23682
rect 36517 -23716 36551 -23682
rect 36675 -23716 36709 -23682
rect 36833 -23716 36867 -23682
rect 36991 -23716 37025 -23682
rect 34542 -24151 34576 -23775
rect 34700 -24151 34734 -23775
rect 34858 -24151 34892 -23775
rect 35016 -24151 35050 -23775
rect 35174 -24151 35208 -23775
rect 35332 -24151 35366 -23775
rect 35490 -24151 35524 -23775
rect 35648 -24151 35682 -23775
rect 35806 -24151 35840 -23775
rect 35964 -24151 35998 -23775
rect 36122 -24151 36156 -23775
rect 36280 -24151 36314 -23775
rect 36438 -24151 36472 -23775
rect 36596 -24151 36630 -23775
rect 36754 -24151 36788 -23775
rect 36912 -24151 36946 -23775
rect 37070 -24151 37104 -23775
rect 34621 -24244 34655 -24210
rect 34779 -24244 34813 -24210
rect 34937 -24244 34971 -24210
rect 35095 -24244 35129 -24210
rect 35253 -24244 35287 -24210
rect 35411 -24244 35445 -24210
rect 35569 -24244 35603 -24210
rect 35727 -24244 35761 -24210
rect 35885 -24244 35919 -24210
rect 36043 -24244 36077 -24210
rect 36201 -24244 36235 -24210
rect 36359 -24244 36393 -24210
rect 36517 -24244 36551 -24210
rect 36675 -24244 36709 -24210
rect 36833 -24244 36867 -24210
rect 36991 -24244 37025 -24210
rect 37204 -24271 37238 -23655
rect 34718 -24382 36928 -24348
rect 27931 -24536 28805 -24502
rect 27984 -24674 28752 -24640
rect 27922 -25100 27956 -24724
rect 28780 -25100 28814 -24724
rect 27984 -25184 28752 -25150
rect 28914 -25213 28948 -24611
rect 27931 -25322 28805 -25288
rect 27931 -25442 28803 -25408
rect 27948 -25576 28724 -25542
rect 28774 -25665 28808 -25611
rect 27948 -25734 28724 -25700
rect 28774 -25823 28808 -25769
rect 27948 -25892 28724 -25858
rect 28774 -25981 28808 -25927
rect 27948 -26050 28724 -26016
rect 28774 -26139 28808 -26085
rect 27948 -26208 28724 -26174
rect 27931 -26342 28803 -26308
rect 27931 -26482 28803 -26448
rect 27948 -26616 28724 -26582
rect 28774 -26705 28808 -26651
rect 27948 -26774 28724 -26740
rect 28774 -26863 28808 -26809
rect 27948 -26932 28724 -26898
rect 28774 -27021 28808 -26967
rect 27948 -27090 28724 -27056
rect 28774 -27179 28808 -27125
rect 27948 -27248 28724 -27214
rect 34989 -24864 35765 -24830
rect 34896 -25043 34930 -24909
rect 35824 -25043 35858 -24909
rect 34989 -25122 35765 -25088
rect 34896 -25301 34930 -25167
rect 35824 -25301 35858 -25167
rect 34989 -25380 35765 -25346
rect 34896 -25559 34930 -25425
rect 35824 -25559 35858 -25425
rect 34989 -25638 35765 -25604
rect 34896 -25817 34930 -25683
rect 35824 -25817 35858 -25683
rect 34989 -25896 35765 -25862
rect 34896 -26075 34930 -25941
rect 35824 -26075 35858 -25941
rect 34989 -26154 35765 -26120
rect 34896 -26333 34930 -26199
rect 35824 -26333 35858 -26199
rect 34989 -26412 35765 -26378
rect 34896 -26591 34930 -26457
rect 35824 -26591 35858 -26457
rect 34989 -26670 35765 -26636
rect 34896 -26849 34930 -26715
rect 35824 -26849 35858 -26715
rect 34989 -26928 35765 -26894
rect 36329 -24864 37105 -24830
rect 36236 -25043 36270 -24909
rect 37164 -25043 37198 -24909
rect 36329 -25122 37105 -25088
rect 36236 -25301 36270 -25167
rect 37164 -25301 37198 -25167
rect 36329 -25380 37105 -25346
rect 36236 -25559 36270 -25425
rect 37164 -25559 37198 -25425
rect 36329 -25638 37105 -25604
rect 36236 -25817 36270 -25683
rect 37164 -25817 37198 -25683
rect 36329 -25896 37105 -25862
rect 36236 -26075 36270 -25941
rect 37164 -26075 37198 -25941
rect 36329 -26154 37105 -26120
rect 36236 -26333 36270 -26199
rect 37164 -26333 37198 -26199
rect 36329 -26412 37105 -26378
rect 36236 -26591 36270 -26457
rect 37164 -26591 37198 -26457
rect 36329 -26670 37105 -26636
rect 36236 -26849 36270 -26715
rect 37164 -26849 37198 -26715
rect 36329 -26928 37105 -26894
rect 27931 -27382 28803 -27348
rect 27931 -27522 28803 -27488
rect 27948 -27656 28724 -27622
rect 28774 -27745 28808 -27691
rect 27948 -27814 28724 -27780
rect 28774 -27903 28808 -27849
rect 27948 -27972 28724 -27938
rect 28774 -28061 28808 -28007
rect 27948 -28130 28724 -28096
rect 28774 -28219 28808 -28165
rect 27948 -28288 28724 -28254
rect 27931 -28422 28803 -28388
rect 27931 -28562 28803 -28528
rect 27948 -28696 28724 -28662
rect 28774 -28785 28808 -28731
rect 27948 -28854 28724 -28820
rect 28774 -28943 28808 -28889
rect 27948 -29012 28724 -28978
rect 28774 -29101 28808 -29047
rect 27948 -29170 28724 -29136
rect 28774 -29259 28808 -29205
rect 27948 -29328 28724 -29294
rect 31712 -28336 31774 -28302
rect 31774 -28336 32042 -28302
rect 32042 -28336 32104 -28302
rect 32152 -28336 32214 -28302
rect 32214 -28336 32482 -28302
rect 32482 -28336 32544 -28302
rect 31888 -28474 31928 -28440
rect 31812 -28909 31846 -28533
rect 31970 -28909 32004 -28533
rect 31888 -29002 31928 -28968
rect 32328 -28474 32368 -28440
rect 32252 -28909 32286 -28533
rect 32410 -28909 32444 -28533
rect 32328 -29002 32368 -28968
rect 32592 -28336 32654 -28302
rect 32654 -28336 32922 -28302
rect 32922 -28336 32984 -28302
rect 32768 -28474 32808 -28440
rect 32692 -28909 32726 -28533
rect 32850 -28909 32884 -28533
rect 33912 -28336 33974 -28302
rect 33974 -28336 34242 -28302
rect 34242 -28336 34304 -28302
rect 33075 -28636 33629 -28602
rect 32972 -28698 33006 -28683
rect 32768 -29002 32808 -28968
rect 32972 -29044 33006 -28698
rect 32972 -29059 33006 -29044
rect 33242 -28774 33462 -28740
rect 33106 -28909 33140 -28833
rect 33564 -28909 33598 -28833
rect 33242 -29002 33462 -28968
rect 34352 -28336 34414 -28302
rect 34414 -28336 34682 -28302
rect 34682 -28336 34744 -28302
rect 34088 -28474 34128 -28440
rect 34012 -28909 34046 -28533
rect 34170 -28909 34204 -28533
rect 34088 -29002 34128 -28968
rect 34528 -28474 34568 -28440
rect 34452 -28909 34486 -28533
rect 34610 -28909 34644 -28533
rect 34528 -29002 34568 -28968
rect 34792 -28336 34854 -28302
rect 34854 -28336 35122 -28302
rect 35122 -28336 35184 -28302
rect 34968 -28474 35008 -28440
rect 34892 -28909 34926 -28533
rect 35050 -28909 35084 -28533
rect 36112 -28336 36174 -28302
rect 36174 -28336 36442 -28302
rect 36442 -28336 36504 -28302
rect 35275 -28636 35829 -28602
rect 35172 -28698 35206 -28683
rect 34968 -29002 35008 -28968
rect 35172 -29044 35206 -28698
rect 35172 -29059 35206 -29044
rect 35442 -28774 35662 -28740
rect 35306 -28909 35340 -28833
rect 35764 -28909 35798 -28833
rect 35442 -29002 35662 -28968
rect 36552 -28336 36614 -28302
rect 36614 -28336 36882 -28302
rect 36882 -28336 36944 -28302
rect 36288 -28474 36328 -28440
rect 36212 -28909 36246 -28533
rect 36370 -28909 36404 -28533
rect 36288 -29002 36328 -28968
rect 36728 -28474 36768 -28440
rect 36652 -28909 36686 -28533
rect 36810 -28909 36844 -28533
rect 36728 -29002 36768 -28968
rect 36992 -28336 37054 -28302
rect 37054 -28336 37322 -28302
rect 37322 -28336 37384 -28302
rect 37168 -28474 37208 -28440
rect 37092 -28909 37126 -28533
rect 37250 -28909 37284 -28533
rect 37475 -28636 38029 -28602
rect 37372 -28698 37406 -28683
rect 37168 -29002 37208 -28968
rect 37372 -29044 37406 -28698
rect 37372 -29059 37406 -29044
rect 37642 -28774 37862 -28740
rect 37506 -28909 37540 -28833
rect 37964 -28909 37998 -28833
rect 37642 -29002 37862 -28968
rect 27931 -29462 28803 -29428
rect 27931 -29602 28803 -29568
rect 27948 -29736 28724 -29702
rect 28774 -29825 28808 -29771
rect 27948 -29894 28724 -29860
rect 28774 -29983 28808 -29929
rect 27948 -30052 28724 -30018
rect 28774 -30141 28808 -30087
rect 27948 -30210 28724 -30176
rect 28774 -30299 28808 -30245
rect 27948 -30368 28724 -30334
rect 27931 -30502 28803 -30468
rect 27931 -30642 28803 -30608
rect 27948 -30776 28724 -30742
rect 28774 -30865 28808 -30811
rect 27948 -30934 28724 -30900
rect 28774 -31023 28808 -30969
rect 27948 -31092 28724 -31058
rect 28774 -31181 28808 -31127
rect 27948 -31250 28724 -31216
rect 28774 -31339 28808 -31285
rect 27948 -31408 28724 -31374
rect 32119 -29427 32153 -29420
rect 31875 -29503 31943 -29469
rect 31813 -29729 31847 -29553
rect 31971 -29729 32005 -29553
rect 31875 -29813 31943 -29779
rect 32119 -29855 32139 -29427
rect 32139 -29855 32153 -29427
rect 32315 -29503 32383 -29469
rect 32253 -29729 32287 -29553
rect 32411 -29729 32445 -29553
rect 32315 -29813 32383 -29779
rect 32119 -29862 32153 -29855
rect 32769 -29503 32809 -29469
rect 32693 -29729 32727 -29553
rect 32851 -29729 32885 -29553
rect 32769 -29813 32809 -29779
rect 32998 -29427 33032 -29420
rect 32998 -29855 33032 -29427
rect 33208 -29503 33248 -29469
rect 33366 -29503 33406 -29469
rect 33524 -29503 33564 -29469
rect 33132 -29729 33166 -29553
rect 33290 -29729 33324 -29553
rect 33448 -29729 33482 -29553
rect 33606 -29729 33640 -29553
rect 33208 -29813 33248 -29779
rect 33366 -29813 33406 -29779
rect 33524 -29813 33564 -29779
rect 32998 -29862 33032 -29855
rect 34319 -29427 34353 -29420
rect 34075 -29503 34143 -29469
rect 34013 -29729 34047 -29553
rect 34171 -29729 34205 -29553
rect 34075 -29813 34143 -29779
rect 34319 -29855 34339 -29427
rect 34339 -29855 34353 -29427
rect 34515 -29503 34583 -29469
rect 34453 -29729 34487 -29553
rect 34611 -29729 34645 -29553
rect 34515 -29813 34583 -29779
rect 34319 -29862 34353 -29855
rect 34969 -29503 35009 -29469
rect 34893 -29729 34927 -29553
rect 35051 -29729 35085 -29553
rect 34969 -29813 35009 -29779
rect 35198 -29427 35232 -29420
rect 35198 -29855 35232 -29427
rect 35408 -29503 35448 -29469
rect 35566 -29503 35606 -29469
rect 35724 -29503 35764 -29469
rect 35332 -29729 35366 -29553
rect 35490 -29729 35524 -29553
rect 35648 -29729 35682 -29553
rect 35806 -29729 35840 -29553
rect 35408 -29813 35448 -29779
rect 35566 -29813 35606 -29779
rect 35724 -29813 35764 -29779
rect 35198 -29862 35232 -29855
rect 36519 -29427 36553 -29420
rect 36275 -29503 36343 -29469
rect 36213 -29729 36247 -29553
rect 36371 -29729 36405 -29553
rect 36275 -29813 36343 -29779
rect 36519 -29855 36539 -29427
rect 36539 -29855 36553 -29427
rect 36715 -29503 36783 -29469
rect 36653 -29729 36687 -29553
rect 36811 -29729 36845 -29553
rect 36715 -29813 36783 -29779
rect 36519 -29862 36553 -29855
rect 37169 -29503 37209 -29469
rect 37093 -29729 37127 -29553
rect 37251 -29729 37285 -29553
rect 37169 -29813 37209 -29779
rect 37398 -29427 37432 -29420
rect 37398 -29855 37432 -29427
rect 37608 -29503 37648 -29469
rect 37766 -29503 37806 -29469
rect 37924 -29503 37964 -29469
rect 37532 -29729 37566 -29553
rect 37690 -29729 37724 -29553
rect 37848 -29729 37882 -29553
rect 38006 -29729 38040 -29553
rect 37608 -29813 37648 -29779
rect 37766 -29813 37806 -29779
rect 37924 -29813 37964 -29779
rect 37398 -29862 37432 -29855
rect 31713 -29951 31775 -29917
rect 31775 -29951 32043 -29917
rect 32043 -29951 32105 -29917
rect 32192 -29951 32215 -29917
rect 32215 -29951 32483 -29917
rect 32483 -29951 32506 -29917
rect 32593 -29951 32655 -29917
rect 32655 -29951 32923 -29917
rect 32923 -29951 32985 -29917
rect 33103 -29951 33669 -29917
rect 33913 -29951 33975 -29917
rect 33975 -29951 34243 -29917
rect 34243 -29951 34305 -29917
rect 34392 -29951 34415 -29917
rect 34415 -29951 34683 -29917
rect 34683 -29951 34706 -29917
rect 34793 -29951 34855 -29917
rect 34855 -29951 35123 -29917
rect 35123 -29951 35185 -29917
rect 35303 -29951 35869 -29917
rect 36113 -29951 36175 -29917
rect 36175 -29951 36443 -29917
rect 36443 -29951 36505 -29917
rect 36592 -29951 36615 -29917
rect 36615 -29951 36883 -29917
rect 36883 -29951 36906 -29917
rect 36993 -29951 37055 -29917
rect 37055 -29951 37323 -29917
rect 37323 -29951 37385 -29917
rect 37503 -29951 38069 -29917
rect 31753 -30107 32319 -30073
rect 32437 -30107 32499 -30073
rect 32499 -30107 32767 -30073
rect 32767 -30107 32829 -30073
rect 32916 -30107 32939 -30073
rect 32939 -30107 33207 -30073
rect 33207 -30107 33230 -30073
rect 33317 -30107 33379 -30073
rect 33379 -30107 33647 -30073
rect 33647 -30107 33709 -30073
rect 33953 -30107 34519 -30073
rect 34637 -30107 34699 -30073
rect 34699 -30107 34967 -30073
rect 34967 -30107 35029 -30073
rect 35116 -30107 35139 -30073
rect 35139 -30107 35407 -30073
rect 35407 -30107 35430 -30073
rect 35517 -30107 35579 -30073
rect 35579 -30107 35847 -30073
rect 35847 -30107 35909 -30073
rect 36153 -30107 36719 -30073
rect 36837 -30107 36899 -30073
rect 36899 -30107 37167 -30073
rect 37167 -30107 37229 -30073
rect 37316 -30107 37339 -30073
rect 37339 -30107 37607 -30073
rect 37607 -30107 37630 -30073
rect 37717 -30107 37779 -30073
rect 37779 -30107 38047 -30073
rect 38047 -30107 38109 -30073
rect 32390 -30169 32424 -30162
rect 31858 -30245 31898 -30211
rect 32016 -30245 32056 -30211
rect 32174 -30245 32214 -30211
rect 31782 -30471 31816 -30295
rect 31940 -30471 31974 -30295
rect 32098 -30471 32132 -30295
rect 32256 -30471 32290 -30295
rect 31858 -30555 31898 -30521
rect 32016 -30555 32056 -30521
rect 32174 -30555 32214 -30521
rect 32390 -30597 32424 -30169
rect 32390 -30604 32424 -30597
rect 32613 -30245 32653 -30211
rect 32537 -30471 32571 -30295
rect 32695 -30471 32729 -30295
rect 32613 -30555 32653 -30521
rect 33269 -30169 33303 -30162
rect 33039 -30245 33107 -30211
rect 32977 -30471 33011 -30295
rect 33135 -30471 33169 -30295
rect 33039 -30555 33107 -30521
rect 33269 -30597 33283 -30169
rect 33283 -30597 33303 -30169
rect 33479 -30245 33547 -30211
rect 33417 -30471 33451 -30295
rect 33575 -30471 33609 -30295
rect 33479 -30555 33547 -30521
rect 33269 -30604 33303 -30597
rect 34590 -30169 34624 -30162
rect 34058 -30245 34098 -30211
rect 34216 -30245 34256 -30211
rect 34374 -30245 34414 -30211
rect 33982 -30471 34016 -30295
rect 34140 -30471 34174 -30295
rect 34298 -30471 34332 -30295
rect 34456 -30471 34490 -30295
rect 34058 -30555 34098 -30521
rect 34216 -30555 34256 -30521
rect 34374 -30555 34414 -30521
rect 34590 -30597 34624 -30169
rect 34590 -30604 34624 -30597
rect 34813 -30245 34853 -30211
rect 34737 -30471 34771 -30295
rect 34895 -30471 34929 -30295
rect 34813 -30555 34853 -30521
rect 35469 -30169 35503 -30162
rect 35239 -30245 35307 -30211
rect 35177 -30471 35211 -30295
rect 35335 -30471 35369 -30295
rect 35239 -30555 35307 -30521
rect 35469 -30597 35483 -30169
rect 35483 -30597 35503 -30169
rect 35679 -30245 35747 -30211
rect 35617 -30471 35651 -30295
rect 35775 -30471 35809 -30295
rect 35679 -30555 35747 -30521
rect 35469 -30604 35503 -30597
rect 36790 -30169 36824 -30162
rect 36258 -30245 36298 -30211
rect 36416 -30245 36456 -30211
rect 36574 -30245 36614 -30211
rect 36182 -30471 36216 -30295
rect 36340 -30471 36374 -30295
rect 36498 -30471 36532 -30295
rect 36656 -30471 36690 -30295
rect 36258 -30555 36298 -30521
rect 36416 -30555 36456 -30521
rect 36574 -30555 36614 -30521
rect 36790 -30597 36824 -30169
rect 36790 -30604 36824 -30597
rect 37013 -30245 37053 -30211
rect 36937 -30471 36971 -30295
rect 37095 -30471 37129 -30295
rect 37013 -30555 37053 -30521
rect 37669 -30169 37703 -30162
rect 37439 -30245 37507 -30211
rect 37377 -30471 37411 -30295
rect 37535 -30471 37569 -30295
rect 37439 -30555 37507 -30521
rect 37669 -30597 37683 -30169
rect 37683 -30597 37703 -30169
rect 37879 -30245 37947 -30211
rect 37817 -30471 37851 -30295
rect 37975 -30471 38009 -30295
rect 37879 -30555 37947 -30521
rect 37669 -30604 37703 -30597
rect 31960 -31056 32180 -31022
rect 31824 -31191 31858 -31115
rect 32282 -31191 32316 -31115
rect 31960 -31284 32180 -31250
rect 32416 -30980 32450 -30965
rect 32416 -31326 32450 -30980
rect 32614 -31056 32654 -31022
rect 32416 -31341 32450 -31326
rect 31793 -31422 32347 -31388
rect 27931 -31542 28803 -31508
rect 32538 -31491 32572 -31115
rect 32696 -31491 32730 -31115
rect 32614 -31584 32654 -31550
rect 32438 -31722 32500 -31688
rect 32500 -31722 32768 -31688
rect 32768 -31722 32830 -31688
rect 33054 -31056 33094 -31022
rect 32978 -31491 33012 -31115
rect 33136 -31491 33170 -31115
rect 33054 -31584 33094 -31550
rect 33494 -31056 33534 -31022
rect 33418 -31491 33452 -31115
rect 33576 -31491 33610 -31115
rect 33494 -31584 33534 -31550
rect 32878 -31722 32940 -31688
rect 32940 -31722 33208 -31688
rect 33208 -31722 33270 -31688
rect 34160 -31056 34380 -31022
rect 34024 -31191 34058 -31115
rect 34482 -31191 34516 -31115
rect 34160 -31284 34380 -31250
rect 34616 -30980 34650 -30965
rect 34616 -31326 34650 -30980
rect 34814 -31056 34854 -31022
rect 34616 -31341 34650 -31326
rect 33993 -31422 34547 -31388
rect 33318 -31722 33380 -31688
rect 33380 -31722 33648 -31688
rect 33648 -31722 33710 -31688
rect 34738 -31491 34772 -31115
rect 34896 -31491 34930 -31115
rect 34814 -31584 34854 -31550
rect 34638 -31722 34700 -31688
rect 34700 -31722 34968 -31688
rect 34968 -31722 35030 -31688
rect 35254 -31056 35294 -31022
rect 35178 -31491 35212 -31115
rect 35336 -31491 35370 -31115
rect 35254 -31584 35294 -31550
rect 35694 -31056 35734 -31022
rect 35618 -31491 35652 -31115
rect 35776 -31491 35810 -31115
rect 35694 -31584 35734 -31550
rect 35078 -31722 35140 -31688
rect 35140 -31722 35408 -31688
rect 35408 -31722 35470 -31688
rect 36360 -31056 36580 -31022
rect 36224 -31191 36258 -31115
rect 36682 -31191 36716 -31115
rect 36360 -31284 36580 -31250
rect 36816 -30980 36850 -30965
rect 36816 -31326 36850 -30980
rect 37014 -31056 37054 -31022
rect 36816 -31341 36850 -31326
rect 36193 -31422 36747 -31388
rect 35518 -31722 35580 -31688
rect 35580 -31722 35848 -31688
rect 35848 -31722 35910 -31688
rect 36938 -31491 36972 -31115
rect 37096 -31491 37130 -31115
rect 37014 -31584 37054 -31550
rect 36838 -31722 36900 -31688
rect 36900 -31722 37168 -31688
rect 37168 -31722 37230 -31688
rect 37454 -31056 37494 -31022
rect 37378 -31491 37412 -31115
rect 37536 -31491 37570 -31115
rect 37454 -31584 37494 -31550
rect 37894 -31056 37934 -31022
rect 37818 -31491 37852 -31115
rect 37976 -31491 38010 -31115
rect 37894 -31584 37934 -31550
rect 37278 -31722 37340 -31688
rect 37340 -31722 37608 -31688
rect 37608 -31722 37670 -31688
rect 37718 -31722 37780 -31688
rect 37780 -31722 38048 -31688
rect 38048 -31722 38110 -31688
<< metal1 >>
rect 29990 11986 36820 11990
rect 29986 11980 36820 11986
rect 22496 11944 26802 11950
rect 22496 11910 22508 11944
rect 26790 11910 26802 11944
rect 22496 11904 26802 11910
rect 29986 11937 36480 11980
rect 29986 11903 30073 11937
rect 30639 11903 30757 11937
rect 31149 11903 31236 11937
rect 31550 11903 31637 11937
rect 32029 11903 32273 11937
rect 32839 11903 32957 11937
rect 33349 11903 33436 11937
rect 33750 11903 33837 11937
rect 34229 11903 34473 11937
rect 35039 11903 35157 11937
rect 35549 11903 35636 11937
rect 35950 11903 36037 11937
rect 36429 11903 36480 11937
rect 29986 11890 36480 11903
rect 29986 11886 32112 11890
rect 32186 11886 34312 11890
rect 34386 11886 36480 11890
rect 22370 11796 22932 11802
rect 22230 11538 22276 11550
rect 2500 11180 2510 11240
rect 2690 11180 2700 11240
rect 2500 10980 2700 11180
rect 3160 11180 3170 11240
rect 3350 11180 3360 11240
rect 3160 10980 3360 11180
rect 3820 11180 3830 11240
rect 4010 11180 4020 11240
rect 3820 10980 4020 11180
rect 4700 11180 4710 11240
rect 4890 11180 4900 11240
rect 4700 10980 4900 11180
rect 5360 11180 5370 11240
rect 5550 11180 5560 11240
rect 5360 10980 5560 11180
rect 6020 11180 6030 11240
rect 6210 11180 6220 11240
rect 6020 10980 6220 11180
rect 6900 11100 7100 11240
rect 6900 11040 6910 11100
rect 7090 11040 7100 11100
rect 6900 10980 7100 11040
rect 7560 11100 7760 11240
rect 7560 11040 7570 11100
rect 7750 11040 7760 11100
rect 7560 10980 7760 11040
rect 8220 11100 8420 11240
rect 8220 11040 8230 11100
rect 8410 11040 8420 11100
rect 8220 10980 8420 11040
rect 9100 11100 9300 11240
rect 9100 11040 9110 11100
rect 9290 11040 9300 11100
rect 9100 10980 9300 11040
rect 9760 11100 9960 11240
rect 9760 11040 9770 11100
rect 9950 11040 9960 11100
rect 9760 10980 9960 11040
rect 10420 11100 10620 11240
rect 10420 11040 10430 11100
rect 10610 11040 10620 11100
rect 10420 10980 10620 11040
rect 11300 11100 11500 11240
rect 11300 11040 11310 11100
rect 11490 11040 11500 11100
rect 11300 10980 11500 11040
rect 11960 11100 12160 11240
rect 11960 11040 11970 11100
rect 12150 11040 12160 11100
rect 11960 10980 12160 11040
rect 12620 11100 12820 11240
rect 12620 11040 12630 11100
rect 12810 11040 12820 11100
rect 12620 10980 12820 11040
rect 13500 11100 13700 11240
rect 13500 11040 13510 11100
rect 13690 11040 13700 11100
rect 13500 10980 13700 11040
rect 14160 11100 14360 11240
rect 14160 11040 14170 11100
rect 14350 11040 14360 11100
rect 14160 10980 14360 11040
rect 14820 11100 15020 11240
rect 14820 11040 14830 11100
rect 15010 11040 15020 11100
rect 14820 10980 15020 11040
rect 15700 11180 15710 11240
rect 15890 11180 15900 11240
rect 15700 10980 15900 11180
rect 16360 11180 16370 11240
rect 16550 11180 16560 11240
rect 16360 10980 16560 11180
rect 17020 11180 17030 11240
rect 17210 11180 17220 11240
rect 17020 10980 17220 11180
rect 17900 11180 17910 11240
rect 18090 11180 18100 11240
rect 17900 10980 18100 11180
rect 18560 11180 18570 11240
rect 18750 11180 18760 11240
rect 18560 10980 18760 11180
rect 19220 11180 19230 11240
rect 19410 11180 19420 11240
rect 19220 10980 19420 11180
rect 2458 10974 4058 10980
rect 2458 10940 2470 10974
rect 4046 10940 4058 10974
rect 4658 10974 6258 10980
rect 4658 10940 4670 10974
rect 6246 10940 6258 10974
rect 6858 10974 8458 10980
rect 6858 10940 6870 10974
rect 8446 10940 8458 10974
rect 9058 10974 10658 10980
rect 9058 10940 9070 10974
rect 10646 10940 10658 10974
rect 11258 10974 12858 10980
rect 11258 10940 11270 10974
rect 12846 10940 12858 10974
rect 13458 10974 15058 10980
rect 13458 10940 13470 10974
rect 15046 10940 15058 10974
rect 15658 10974 17258 10980
rect 15658 10940 15670 10974
rect 17246 10940 17258 10974
rect 17858 10974 19458 10980
rect 17858 10940 17870 10974
rect 19446 10940 19458 10974
rect -90 10930 10 10940
rect -90 10870 -70 10930
rect -10 10870 10 10930
rect -90 10860 10 10870
rect 2110 10930 2210 10940
rect 2458 10934 4058 10940
rect 2110 10870 2130 10930
rect 2190 10870 2210 10930
rect 4310 10930 4410 10940
rect 4658 10934 6258 10940
rect 2110 10860 2210 10870
rect 2380 10912 2426 10924
rect 2380 10710 2386 10912
rect 2010 10650 2020 10710
rect 2080 10650 2386 10710
rect 2380 10644 2386 10650
rect 2420 10644 2426 10912
rect 2380 10632 2426 10644
rect 4090 10912 4136 10924
rect 4090 10644 4096 10912
rect 4130 10820 4136 10912
rect 4310 10870 4330 10930
rect 4390 10870 4410 10930
rect 6510 10930 6610 10940
rect 6858 10934 8458 10940
rect 4310 10860 4410 10870
rect 4580 10912 4626 10924
rect 4130 10760 4220 10820
rect 4280 10760 4510 10820
rect 4130 10644 4136 10760
rect 4580 10710 4586 10912
rect 4210 10650 4220 10710
rect 4280 10650 4586 10710
rect 4090 10632 4136 10644
rect 4580 10644 4586 10650
rect 4620 10644 4626 10912
rect 4580 10632 4626 10644
rect 6290 10912 6336 10924
rect 6290 10644 6296 10912
rect 6330 10820 6336 10912
rect 6510 10870 6530 10930
rect 6590 10870 6610 10930
rect 8710 10930 8810 10940
rect 9058 10934 10658 10940
rect 6510 10860 6610 10870
rect 6780 10912 6826 10924
rect 6330 10760 6420 10820
rect 6480 10760 6710 10820
rect 6330 10644 6336 10760
rect 6780 10710 6786 10912
rect 6410 10650 6640 10710
rect 6700 10650 6786 10710
rect 6290 10632 6336 10644
rect 6780 10644 6786 10650
rect 6820 10644 6826 10912
rect 6780 10632 6826 10644
rect 8490 10912 8536 10924
rect 8490 10644 8496 10912
rect 8530 10820 8536 10912
rect 8710 10870 8730 10930
rect 8790 10870 8810 10930
rect 10910 10930 11010 10940
rect 11258 10934 12858 10940
rect 8710 10860 8810 10870
rect 8980 10912 9026 10924
rect 8530 10760 8840 10820
rect 8900 10760 8910 10820
rect 8530 10644 8536 10760
rect 8980 10710 8986 10912
rect 8610 10650 8840 10710
rect 8900 10650 8986 10710
rect 8490 10632 8536 10644
rect 8980 10644 8986 10650
rect 9020 10644 9026 10912
rect 8980 10632 9026 10644
rect 10690 10912 10736 10924
rect 10690 10644 10696 10912
rect 10730 10820 10736 10912
rect 10910 10870 10930 10930
rect 10990 10870 11010 10930
rect 13110 10930 13210 10940
rect 13458 10934 15058 10940
rect 10910 10860 11010 10870
rect 11180 10912 11226 10924
rect 10730 10760 11040 10820
rect 11100 10760 11110 10820
rect 10730 10644 10736 10760
rect 11180 10710 11186 10912
rect 10810 10650 11040 10710
rect 11100 10650 11186 10710
rect 10690 10632 10736 10644
rect 11180 10644 11186 10650
rect 11220 10644 11226 10912
rect 11180 10632 11226 10644
rect 12890 10912 12936 10924
rect 12890 10644 12896 10912
rect 12930 10820 12936 10912
rect 13110 10870 13130 10930
rect 13190 10870 13210 10930
rect 15310 10930 15410 10940
rect 15658 10934 17258 10940
rect 13110 10860 13210 10870
rect 13380 10912 13426 10924
rect 12930 10760 13240 10820
rect 13300 10760 13310 10820
rect 12930 10644 12936 10760
rect 13380 10710 13386 10912
rect 13010 10650 13240 10710
rect 13300 10650 13386 10710
rect 12890 10632 12936 10644
rect 13380 10644 13386 10650
rect 13420 10644 13426 10912
rect 13380 10632 13426 10644
rect 15090 10912 15136 10924
rect 15090 10644 15096 10912
rect 15130 10820 15136 10912
rect 15310 10870 15330 10930
rect 15390 10870 15410 10930
rect 17510 10930 17610 10940
rect 17858 10934 19458 10940
rect 15310 10860 15410 10870
rect 15580 10912 15626 10924
rect 15130 10760 15440 10820
rect 15500 10760 15510 10820
rect 15130 10644 15136 10760
rect 15580 10710 15586 10912
rect 15210 10650 15220 10710
rect 15280 10650 15586 10710
rect 15090 10632 15136 10644
rect 15580 10644 15586 10650
rect 15620 10644 15626 10912
rect 15580 10632 15626 10644
rect 17290 10912 17336 10924
rect 17290 10644 17296 10912
rect 17330 10820 17336 10912
rect 17510 10870 17530 10930
rect 17590 10870 17610 10930
rect 19710 10930 19810 10940
rect 17510 10860 17610 10870
rect 17780 10912 17826 10924
rect 17330 10760 17420 10820
rect 17480 10760 17710 10820
rect 17330 10644 17336 10760
rect 17780 10710 17786 10912
rect 17410 10650 17420 10710
rect 17480 10650 17786 10710
rect 17290 10632 17336 10644
rect 17780 10644 17786 10650
rect 17820 10644 17826 10912
rect 17780 10632 17826 10644
rect 19490 10912 19536 10924
rect 19490 10644 19496 10912
rect 19530 10800 19536 10912
rect 19710 10870 19730 10930
rect 19790 10870 19810 10930
rect 19710 10860 19810 10870
rect 21910 10930 22010 10940
rect 21910 10870 21930 10930
rect 21990 10870 22010 10930
rect 21910 10860 22010 10870
rect 19530 10740 19620 10800
rect 19680 10740 19910 10800
rect 19530 10644 19536 10740
rect 19490 10632 19536 10644
rect 2458 10616 4058 10622
rect 2458 10582 2470 10616
rect 4046 10582 4058 10616
rect 2458 10576 2510 10582
rect 2500 10550 2510 10576
rect 4010 10576 4058 10582
rect 4658 10616 6258 10622
rect 4658 10582 4670 10616
rect 6246 10582 6258 10616
rect 4658 10576 4710 10582
rect 4010 10550 4020 10576
rect 2500 10540 4020 10550
rect 4700 10550 4710 10576
rect 6210 10576 6258 10582
rect 6858 10616 8458 10622
rect 6858 10582 6870 10616
rect 8446 10582 8458 10616
rect 6858 10576 6910 10582
rect 6210 10550 6220 10576
rect 4700 10540 6220 10550
rect 6900 10550 6910 10576
rect 8410 10576 8458 10582
rect 9058 10616 10658 10622
rect 9058 10582 9070 10616
rect 10646 10582 10658 10616
rect 9058 10576 9110 10582
rect 8410 10550 8420 10576
rect 6900 10540 8420 10550
rect 9100 10550 9110 10576
rect 10610 10576 10658 10582
rect 11258 10616 12858 10622
rect 11258 10582 11270 10616
rect 12846 10582 12858 10616
rect 11258 10576 11310 10582
rect 10610 10550 10620 10576
rect 9100 10540 10620 10550
rect 11300 10550 11310 10576
rect 12810 10576 12858 10582
rect 13458 10616 15058 10622
rect 13458 10582 13470 10616
rect 15046 10582 15058 10616
rect 13458 10576 13510 10582
rect 12810 10550 12820 10576
rect 11300 10540 12820 10550
rect 13500 10550 13510 10576
rect 15010 10576 15058 10582
rect 15658 10616 17258 10622
rect 15658 10582 15670 10616
rect 17246 10582 17258 10616
rect 15658 10576 15710 10582
rect 15010 10550 15020 10576
rect 13500 10540 15020 10550
rect 15700 10550 15710 10576
rect 17210 10576 17258 10582
rect 17858 10616 19458 10622
rect 17858 10582 17870 10616
rect 19446 10582 19458 10616
rect 17858 10576 17910 10582
rect 17210 10550 17220 10576
rect 15700 10540 17220 10550
rect 17900 10550 17910 10576
rect 19410 10576 19458 10582
rect 19410 10550 19420 10576
rect 17900 10540 19420 10550
rect 2500 10300 2700 10440
rect 2500 10240 2510 10300
rect 2690 10240 2700 10300
rect 2500 10180 2700 10240
rect 3160 10300 3360 10440
rect 3160 10240 3170 10300
rect 3350 10240 3360 10300
rect 3160 10180 3360 10240
rect 3820 10300 4020 10440
rect 3820 10240 3830 10300
rect 4010 10240 4020 10300
rect 3820 10180 4020 10240
rect 4700 10300 4900 10440
rect 4700 10240 4710 10300
rect 4890 10240 4900 10300
rect 4700 10180 4900 10240
rect 5360 10300 5560 10440
rect 5360 10240 5370 10300
rect 5550 10240 5560 10300
rect 5360 10180 5560 10240
rect 6020 10300 6220 10440
rect 6020 10240 6030 10300
rect 6210 10240 6220 10300
rect 6020 10180 6220 10240
rect 6900 10380 6910 10440
rect 7090 10380 7100 10440
rect 6900 10180 7100 10380
rect 7560 10380 7570 10440
rect 7750 10380 7760 10440
rect 7560 10180 7760 10380
rect 8220 10380 8230 10440
rect 8410 10380 8420 10440
rect 8220 10180 8420 10380
rect 9100 10380 9110 10440
rect 9290 10380 9300 10440
rect 9100 10180 9300 10380
rect 9760 10380 9770 10440
rect 9950 10380 9960 10440
rect 9760 10180 9960 10380
rect 10420 10380 10430 10440
rect 10610 10380 10620 10440
rect 10420 10180 10620 10380
rect 11300 10380 11310 10440
rect 11490 10380 11500 10440
rect 11300 10180 11500 10380
rect 11960 10380 11970 10440
rect 12150 10380 12160 10440
rect 11960 10180 12160 10380
rect 12620 10380 12630 10440
rect 12810 10380 12820 10440
rect 12620 10180 12820 10380
rect 13500 10380 13510 10440
rect 13690 10380 13700 10440
rect 13500 10180 13700 10380
rect 14160 10380 14170 10440
rect 14350 10380 14360 10440
rect 14160 10180 14360 10380
rect 14820 10380 14830 10440
rect 15010 10380 15020 10440
rect 14820 10180 15020 10380
rect 15700 10300 15900 10440
rect 15700 10240 15710 10300
rect 15890 10240 15900 10300
rect 15700 10180 15900 10240
rect 16360 10300 16560 10440
rect 16360 10240 16370 10300
rect 16550 10240 16560 10300
rect 16360 10180 16560 10240
rect 17020 10300 17220 10440
rect 17020 10240 17030 10300
rect 17210 10240 17220 10300
rect 17020 10180 17220 10240
rect 17900 10300 18100 10440
rect 17900 10240 17910 10300
rect 18090 10240 18100 10300
rect 17900 10180 18100 10240
rect 18560 10300 18760 10440
rect 18560 10240 18570 10300
rect 18750 10240 18760 10300
rect 18560 10180 18760 10240
rect 19220 10300 19420 10440
rect 19220 10240 19230 10300
rect 19410 10240 19420 10300
rect 19220 10180 19420 10240
rect 2458 10174 4058 10180
rect 2458 10140 2470 10174
rect 4046 10140 4058 10174
rect 4658 10174 6258 10180
rect 4658 10140 4670 10174
rect 6246 10140 6258 10174
rect 6858 10174 8458 10180
rect 6858 10140 6870 10174
rect 8446 10140 8458 10174
rect 9058 10174 10658 10180
rect 9058 10140 9070 10174
rect 10646 10140 10658 10174
rect 11258 10174 12858 10180
rect 11258 10140 11270 10174
rect 12846 10140 12858 10174
rect 13458 10174 15058 10180
rect 13458 10140 13470 10174
rect 15046 10140 15058 10174
rect 15658 10174 17258 10180
rect 15658 10140 15670 10174
rect 17246 10140 17258 10174
rect 17858 10174 19458 10180
rect 17858 10140 17870 10174
rect 19446 10140 19458 10174
rect -90 10130 10 10140
rect -90 10070 -70 10130
rect -10 10070 10 10130
rect -90 10060 10 10070
rect 2110 10130 2210 10140
rect 2458 10134 4058 10140
rect 2110 10070 2130 10130
rect 2190 10070 2210 10130
rect 4310 10130 4410 10140
rect 4658 10134 6258 10140
rect 2110 10060 2210 10070
rect 2380 10112 2426 10124
rect 2380 9910 2386 10112
rect 2010 9850 2240 9910
rect 2300 9850 2386 9910
rect 2380 9844 2386 9850
rect 2420 9844 2426 10112
rect 2380 9832 2426 9844
rect 4090 10112 4136 10124
rect 4090 9844 4096 10112
rect 4130 10020 4136 10112
rect 4310 10070 4330 10130
rect 4390 10070 4410 10130
rect 6510 10130 6610 10140
rect 6858 10134 8458 10140
rect 4310 10060 4410 10070
rect 4580 10112 4626 10124
rect 4130 9960 4440 10020
rect 4500 9960 4510 10020
rect 4130 9844 4136 9960
rect 4580 9910 4586 10112
rect 4210 9850 4440 9910
rect 4500 9850 4586 9910
rect 4090 9832 4136 9844
rect 4580 9844 4586 9850
rect 4620 9844 4626 10112
rect 4580 9832 4626 9844
rect 6290 10112 6336 10124
rect 6290 9844 6296 10112
rect 6330 10020 6336 10112
rect 6510 10070 6530 10130
rect 6590 10070 6610 10130
rect 8710 10130 8810 10140
rect 9058 10134 10658 10140
rect 6510 10060 6610 10070
rect 6780 10112 6826 10124
rect 6330 9960 6640 10020
rect 6700 9960 6710 10020
rect 6330 9844 6336 9960
rect 6780 9910 6786 10112
rect 6410 9850 6420 9910
rect 6480 9850 6786 9910
rect 6290 9832 6336 9844
rect 6780 9844 6786 9850
rect 6820 9844 6826 10112
rect 6780 9832 6826 9844
rect 8490 10112 8536 10124
rect 8490 9844 8496 10112
rect 8530 10020 8536 10112
rect 8710 10070 8730 10130
rect 8790 10070 8810 10130
rect 10910 10130 11010 10140
rect 11258 10134 12858 10140
rect 8710 10060 8810 10070
rect 8980 10112 9026 10124
rect 8530 9960 8620 10020
rect 8680 9960 8910 10020
rect 8530 9844 8536 9960
rect 8980 9910 8986 10112
rect 8610 9850 8620 9910
rect 8680 9850 8986 9910
rect 8490 9832 8536 9844
rect 8980 9844 8986 9850
rect 9020 9844 9026 10112
rect 8980 9832 9026 9844
rect 10690 10112 10736 10124
rect 10690 9844 10696 10112
rect 10730 10020 10736 10112
rect 10910 10070 10930 10130
rect 10990 10070 11010 10130
rect 13110 10130 13210 10140
rect 13458 10134 15058 10140
rect 10910 10060 11010 10070
rect 11180 10112 11226 10124
rect 10730 9960 10820 10020
rect 10880 9960 11110 10020
rect 10730 9844 10736 9960
rect 11180 9910 11186 10112
rect 10810 9850 10820 9910
rect 10880 9850 11186 9910
rect 10690 9832 10736 9844
rect 11180 9844 11186 9850
rect 11220 9844 11226 10112
rect 11180 9832 11226 9844
rect 12890 10112 12936 10124
rect 12890 9844 12896 10112
rect 12930 10020 12936 10112
rect 13110 10070 13130 10130
rect 13190 10070 13210 10130
rect 15310 10130 15410 10140
rect 15658 10134 17258 10140
rect 13110 10060 13210 10070
rect 13380 10112 13426 10124
rect 12930 9960 13020 10020
rect 13080 9960 13310 10020
rect 12930 9844 12936 9960
rect 13380 9910 13386 10112
rect 13010 9850 13020 9910
rect 13080 9850 13386 9910
rect 12890 9832 12936 9844
rect 13380 9844 13386 9850
rect 13420 9844 13426 10112
rect 13380 9832 13426 9844
rect 15090 10112 15136 10124
rect 15090 9844 15096 10112
rect 15130 10020 15136 10112
rect 15310 10070 15330 10130
rect 15390 10070 15410 10130
rect 17510 10130 17610 10140
rect 17858 10134 19458 10140
rect 15310 10060 15410 10070
rect 15580 10112 15626 10124
rect 15130 9960 15220 10020
rect 15280 9960 15510 10020
rect 15130 9844 15136 9960
rect 15580 9910 15586 10112
rect 15210 9850 15440 9910
rect 15500 9850 15586 9910
rect 15090 9832 15136 9844
rect 15580 9844 15586 9850
rect 15620 9844 15626 10112
rect 15580 9832 15626 9844
rect 17290 10112 17336 10124
rect 17290 9844 17296 10112
rect 17330 10020 17336 10112
rect 17510 10070 17530 10130
rect 17590 10070 17610 10130
rect 19710 10130 19810 10140
rect 17510 10060 17610 10070
rect 17780 10112 17826 10124
rect 17330 9960 17640 10020
rect 17700 9960 17710 10020
rect 17330 9844 17336 9960
rect 17780 9910 17786 10112
rect 17410 9850 17640 9910
rect 17700 9850 17786 9910
rect 17290 9832 17336 9844
rect 17780 9844 17786 9850
rect 17820 9844 17826 10112
rect 17780 9832 17826 9844
rect 19490 10112 19536 10124
rect 19490 9844 19496 10112
rect 19530 10000 19536 10112
rect 19710 10070 19730 10130
rect 19790 10070 19810 10130
rect 19710 10060 19810 10070
rect 21910 10130 22010 10140
rect 21910 10070 21930 10130
rect 21990 10070 22010 10130
rect 21910 10060 22010 10070
rect 19530 9940 19840 10000
rect 19900 9940 19910 10000
rect 19530 9844 19536 9940
rect 19490 9832 19536 9844
rect 2458 9816 4058 9822
rect 2458 9782 2470 9816
rect 4046 9782 4058 9816
rect 2458 9776 2510 9782
rect 2500 9750 2510 9776
rect 4010 9776 4058 9782
rect 4658 9816 6258 9822
rect 4658 9782 4670 9816
rect 6246 9782 6258 9816
rect 4658 9776 4710 9782
rect 4010 9750 4020 9776
rect 2500 9740 4020 9750
rect 4700 9750 4710 9776
rect 6210 9776 6258 9782
rect 6858 9816 8458 9822
rect 6858 9782 6870 9816
rect 8446 9782 8458 9816
rect 6858 9776 6910 9782
rect 6210 9750 6220 9776
rect 4700 9740 6220 9750
rect 6900 9750 6910 9776
rect 8410 9776 8458 9782
rect 9058 9816 10658 9822
rect 9058 9782 9070 9816
rect 10646 9782 10658 9816
rect 9058 9776 9110 9782
rect 8410 9750 8420 9776
rect 6900 9740 8420 9750
rect 9100 9750 9110 9776
rect 10610 9776 10658 9782
rect 11258 9816 12858 9822
rect 11258 9782 11270 9816
rect 12846 9782 12858 9816
rect 11258 9776 11310 9782
rect 10610 9750 10620 9776
rect 9100 9740 10620 9750
rect 11300 9750 11310 9776
rect 12810 9776 12858 9782
rect 13458 9816 15058 9822
rect 13458 9782 13470 9816
rect 15046 9782 15058 9816
rect 13458 9776 13510 9782
rect 12810 9750 12820 9776
rect 11300 9740 12820 9750
rect 13500 9750 13510 9776
rect 15010 9776 15058 9782
rect 15658 9816 17258 9822
rect 15658 9782 15670 9816
rect 17246 9782 17258 9816
rect 15658 9776 15710 9782
rect 15010 9750 15020 9776
rect 13500 9740 15020 9750
rect 15700 9750 15710 9776
rect 17210 9776 17258 9782
rect 17858 9816 19458 9822
rect 17858 9782 17870 9816
rect 19446 9782 19458 9816
rect 17858 9776 17910 9782
rect 17210 9750 17220 9776
rect 15700 9740 17220 9750
rect 17900 9750 17910 9776
rect 19410 9776 19458 9782
rect 19410 9750 19420 9776
rect 17900 9740 19420 9750
rect 2500 9580 2510 9640
rect 2690 9580 2700 9640
rect 2500 9380 2700 9580
rect 3160 9580 3170 9640
rect 3350 9580 3360 9640
rect 3160 9380 3360 9580
rect 3820 9580 3830 9640
rect 4010 9580 4020 9640
rect 3820 9380 4020 9580
rect 4700 9580 4710 9640
rect 4890 9580 4900 9640
rect 4700 9380 4900 9580
rect 5360 9580 5370 9640
rect 5550 9580 5560 9640
rect 5360 9380 5560 9580
rect 6020 9580 6030 9640
rect 6210 9580 6220 9640
rect 6020 9380 6220 9580
rect 6900 9500 7100 9640
rect 6900 9440 6910 9500
rect 7090 9440 7100 9500
rect 6900 9380 7100 9440
rect 7560 9500 7760 9640
rect 7560 9440 7570 9500
rect 7750 9440 7760 9500
rect 7560 9380 7760 9440
rect 8220 9500 8420 9640
rect 8220 9440 8230 9500
rect 8410 9440 8420 9500
rect 8220 9380 8420 9440
rect 9100 9500 9300 9640
rect 9100 9440 9110 9500
rect 9290 9440 9300 9500
rect 9100 9380 9300 9440
rect 9760 9500 9960 9640
rect 9760 9440 9770 9500
rect 9950 9440 9960 9500
rect 9760 9380 9960 9440
rect 10420 9500 10620 9640
rect 10420 9440 10430 9500
rect 10610 9440 10620 9500
rect 10420 9380 10620 9440
rect 11300 9500 11500 9640
rect 11300 9440 11310 9500
rect 11490 9440 11500 9500
rect 11300 9380 11500 9440
rect 11960 9500 12160 9640
rect 11960 9440 11970 9500
rect 12150 9440 12160 9500
rect 11960 9380 12160 9440
rect 12620 9500 12820 9640
rect 12620 9440 12630 9500
rect 12810 9440 12820 9500
rect 12620 9380 12820 9440
rect 13500 9500 13700 9640
rect 13500 9440 13510 9500
rect 13690 9440 13700 9500
rect 13500 9380 13700 9440
rect 14160 9500 14360 9640
rect 14160 9440 14170 9500
rect 14350 9440 14360 9500
rect 14160 9380 14360 9440
rect 14820 9500 15020 9640
rect 14820 9440 14830 9500
rect 15010 9440 15020 9500
rect 14820 9380 15020 9440
rect 15700 9580 15710 9640
rect 15890 9580 15900 9640
rect 15700 9380 15900 9580
rect 16360 9580 16370 9640
rect 16550 9580 16560 9640
rect 16360 9380 16560 9580
rect 17020 9580 17030 9640
rect 17210 9580 17220 9640
rect 17020 9380 17220 9580
rect 17900 9580 17910 9640
rect 18090 9580 18100 9640
rect 17900 9380 18100 9580
rect 18560 9580 18570 9640
rect 18750 9580 18760 9640
rect 18560 9380 18760 9580
rect 19220 9580 19230 9640
rect 19410 9580 19420 9640
rect 19220 9380 19420 9580
rect 2458 9374 4058 9380
rect 2458 9340 2470 9374
rect 4046 9340 4058 9374
rect 4658 9374 6258 9380
rect 4658 9340 4670 9374
rect 6246 9340 6258 9374
rect 6858 9374 8458 9380
rect 6858 9340 6870 9374
rect 8446 9340 8458 9374
rect 9058 9374 10658 9380
rect 9058 9340 9070 9374
rect 10646 9340 10658 9374
rect 11258 9374 12858 9380
rect 11258 9340 11270 9374
rect 12846 9340 12858 9374
rect 13458 9374 15058 9380
rect 13458 9340 13470 9374
rect 15046 9340 15058 9374
rect 15658 9374 17258 9380
rect 15658 9340 15670 9374
rect 17246 9340 17258 9374
rect 17858 9374 19458 9380
rect 17858 9340 17870 9374
rect 19446 9340 19458 9374
rect -90 9330 10 9340
rect -90 9270 -70 9330
rect -10 9270 10 9330
rect -90 9260 10 9270
rect 2110 9330 2210 9340
rect 2458 9334 4058 9340
rect 2110 9270 2130 9330
rect 2190 9270 2210 9330
rect 4310 9330 4410 9340
rect 4658 9334 6258 9340
rect 2110 9260 2210 9270
rect 2380 9312 2426 9324
rect 1410 9210 1490 9220
rect 1410 9060 1420 9210
rect 1480 9110 1490 9210
rect 2380 9110 2386 9312
rect 1480 9060 2386 9110
rect 1410 9050 2386 9060
rect 2380 9044 2386 9050
rect 2420 9044 2426 9312
rect 2380 9032 2426 9044
rect 4090 9312 4136 9324
rect 4090 9044 4096 9312
rect 4130 9220 4136 9312
rect 4310 9270 4330 9330
rect 4390 9270 4410 9330
rect 6510 9330 6610 9340
rect 6858 9334 8458 9340
rect 4310 9260 4410 9270
rect 4580 9312 4626 9324
rect 4130 9160 4510 9220
rect 4130 9044 4136 9160
rect 4580 9110 4586 9312
rect 4210 9050 4220 9110
rect 4280 9050 4586 9110
rect 4090 9032 4136 9044
rect 4580 9044 4586 9050
rect 4620 9044 4626 9312
rect 4580 9032 4626 9044
rect 6290 9312 6336 9324
rect 6290 9044 6296 9312
rect 6330 9220 6336 9312
rect 6510 9270 6530 9330
rect 6590 9270 6610 9330
rect 8710 9330 8810 9340
rect 9058 9334 10658 9340
rect 6510 9260 6610 9270
rect 6780 9312 6826 9324
rect 6330 9160 6420 9220
rect 6480 9160 6710 9220
rect 6330 9044 6336 9160
rect 6780 9110 6786 9312
rect 6410 9050 6640 9110
rect 6700 9050 6786 9110
rect 6290 9032 6336 9044
rect 6780 9044 6786 9050
rect 6820 9044 6826 9312
rect 6780 9032 6826 9044
rect 8490 9312 8536 9324
rect 8490 9044 8496 9312
rect 8530 9220 8536 9312
rect 8710 9270 8730 9330
rect 8790 9270 8810 9330
rect 10910 9330 11010 9340
rect 11258 9334 12858 9340
rect 8710 9260 8810 9270
rect 8980 9312 9026 9324
rect 8530 9160 8840 9220
rect 8900 9160 8910 9220
rect 8530 9044 8536 9160
rect 8980 9110 8986 9312
rect 8610 9050 8840 9110
rect 8900 9050 8986 9110
rect 8490 9032 8536 9044
rect 8980 9044 8986 9050
rect 9020 9044 9026 9312
rect 8980 9032 9026 9044
rect 10690 9312 10736 9324
rect 10690 9044 10696 9312
rect 10730 9220 10736 9312
rect 10910 9270 10930 9330
rect 10990 9270 11010 9330
rect 13110 9330 13210 9340
rect 13458 9334 15058 9340
rect 10910 9260 11010 9270
rect 11180 9312 11226 9324
rect 10730 9160 11040 9220
rect 11100 9160 11110 9220
rect 10730 9044 10736 9160
rect 11180 9110 11186 9312
rect 10810 9050 11040 9110
rect 11100 9050 11186 9110
rect 10690 9032 10736 9044
rect 11180 9044 11186 9050
rect 11220 9044 11226 9312
rect 11180 9032 11226 9044
rect 12890 9312 12936 9324
rect 12890 9044 12896 9312
rect 12930 9220 12936 9312
rect 13110 9270 13130 9330
rect 13190 9270 13210 9330
rect 15310 9330 15410 9340
rect 15658 9334 17258 9340
rect 13110 9260 13210 9270
rect 13380 9312 13426 9324
rect 12930 9160 13240 9220
rect 13300 9160 13310 9220
rect 12930 9044 12936 9160
rect 13380 9110 13386 9312
rect 13010 9050 13240 9110
rect 13300 9050 13386 9110
rect 12890 9032 12936 9044
rect 13380 9044 13386 9050
rect 13420 9044 13426 9312
rect 13380 9032 13426 9044
rect 15090 9312 15136 9324
rect 15090 9044 15096 9312
rect 15130 9220 15136 9312
rect 15310 9270 15330 9330
rect 15390 9270 15410 9330
rect 17510 9330 17610 9340
rect 17858 9334 19458 9340
rect 15310 9260 15410 9270
rect 15580 9312 15626 9324
rect 15130 9160 15440 9220
rect 15500 9160 15510 9220
rect 15130 9044 15136 9160
rect 15580 9110 15586 9312
rect 15210 9050 15220 9110
rect 15280 9050 15586 9110
rect 15090 9032 15136 9044
rect 15580 9044 15586 9050
rect 15620 9044 15626 9312
rect 15580 9032 15626 9044
rect 17290 9312 17336 9324
rect 17290 9044 17296 9312
rect 17330 9220 17336 9312
rect 17510 9270 17530 9330
rect 17590 9270 17610 9330
rect 19710 9330 19810 9340
rect 17510 9260 17610 9270
rect 17780 9312 17826 9324
rect 17330 9160 17420 9220
rect 17480 9160 17710 9220
rect 17330 9044 17336 9160
rect 17780 9110 17786 9312
rect 17410 9050 17786 9110
rect 17290 9032 17336 9044
rect 17780 9044 17786 9050
rect 17820 9044 17826 9312
rect 17780 9032 17826 9044
rect 19490 9312 19536 9324
rect 19490 9044 19496 9312
rect 19530 9200 19536 9312
rect 19710 9270 19730 9330
rect 19790 9270 19810 9330
rect 21910 9330 22010 9340
rect 19710 9260 19810 9270
rect 20230 9300 20310 9310
rect 20230 9200 20240 9300
rect 19530 9150 20240 9200
rect 20300 9150 20310 9300
rect 21910 9270 21930 9330
rect 21990 9270 22010 9330
rect 21910 9260 22010 9270
rect 19530 9140 20310 9150
rect 19530 9044 19536 9140
rect 19490 9032 19536 9044
rect 2458 9016 4058 9022
rect 420 8990 620 9000
rect 420 8910 430 8990
rect 610 8980 620 8990
rect 2458 8982 2470 9016
rect 4046 8982 4058 9016
rect 2458 8980 4058 8982
rect 610 8976 4058 8980
rect 4658 9016 6258 9022
rect 4658 8982 4670 9016
rect 6246 8982 6258 9016
rect 4658 8976 4710 8982
rect 610 8920 4040 8976
rect 4700 8950 4710 8976
rect 6210 8976 6258 8982
rect 6858 9016 8458 9022
rect 6858 8982 6870 9016
rect 8446 8982 8458 9016
rect 6858 8976 6910 8982
rect 6210 8950 6220 8976
rect 4700 8940 6220 8950
rect 6900 8950 6910 8976
rect 8410 8976 8458 8982
rect 9058 9016 10658 9022
rect 9058 8982 9070 9016
rect 10646 8982 10658 9016
rect 9058 8976 9110 8982
rect 8410 8950 8420 8976
rect 6900 8940 8420 8950
rect 9100 8950 9110 8976
rect 10610 8976 10658 8982
rect 11258 9016 12858 9022
rect 11258 8982 11270 9016
rect 12846 8982 12858 9016
rect 11258 8976 11310 8982
rect 10610 8950 10620 8976
rect 9100 8940 10620 8950
rect 11300 8950 11310 8976
rect 12810 8976 12858 8982
rect 13458 9016 15058 9022
rect 13458 8982 13470 9016
rect 15046 8982 15058 9016
rect 13458 8976 13510 8982
rect 12810 8950 12820 8976
rect 11300 8940 12820 8950
rect 13500 8950 13510 8976
rect 15010 8976 15058 8982
rect 15658 9016 17258 9022
rect 15658 8982 15670 9016
rect 17246 8982 17258 9016
rect 15658 8976 15710 8982
rect 15010 8950 15020 8976
rect 13500 8940 15020 8950
rect 15700 8950 15710 8976
rect 17210 8976 17258 8982
rect 17858 9016 19458 9022
rect 17858 8982 17870 9016
rect 19446 8982 19458 9016
rect 17858 8980 19458 8982
rect 21300 8990 21500 9000
rect 21300 8980 21310 8990
rect 17858 8976 21310 8980
rect 17210 8950 17220 8976
rect 15700 8940 17220 8950
rect 17880 8920 21310 8976
rect 610 8910 620 8920
rect 420 8900 620 8910
rect 21300 8910 21310 8920
rect 21490 8910 21500 8990
rect 21300 8900 21500 8910
rect 2500 8700 2700 8840
rect 2500 8640 2510 8700
rect 2690 8640 2700 8700
rect 2500 8580 2700 8640
rect 3160 8700 3360 8840
rect 3160 8640 3170 8700
rect 3350 8640 3360 8700
rect 3160 8580 3360 8640
rect 3820 8700 4020 8840
rect 3820 8640 3830 8700
rect 4010 8640 4020 8700
rect 3820 8580 4020 8640
rect 4700 8700 4900 8840
rect 4700 8640 4710 8700
rect 4890 8640 4900 8700
rect 4700 8580 4900 8640
rect 5360 8700 5560 8840
rect 5360 8640 5370 8700
rect 5550 8640 5560 8700
rect 5360 8580 5560 8640
rect 6020 8700 6220 8840
rect 6020 8640 6030 8700
rect 6210 8640 6220 8700
rect 6020 8580 6220 8640
rect 6900 8780 6910 8840
rect 7090 8780 7100 8840
rect 6900 8580 7100 8780
rect 7560 8780 7570 8840
rect 7750 8780 7760 8840
rect 7560 8580 7760 8780
rect 8220 8780 8230 8840
rect 8410 8780 8420 8840
rect 8220 8580 8420 8780
rect 9100 8780 9110 8840
rect 9290 8780 9300 8840
rect 9100 8580 9300 8780
rect 9760 8780 9770 8840
rect 9950 8780 9960 8840
rect 9760 8580 9960 8780
rect 10420 8780 10430 8840
rect 10610 8780 10620 8840
rect 10420 8580 10620 8780
rect 11300 8780 11310 8840
rect 11490 8780 11500 8840
rect 11300 8580 11500 8780
rect 11960 8780 11970 8840
rect 12150 8780 12160 8840
rect 11960 8580 12160 8780
rect 12620 8780 12630 8840
rect 12810 8780 12820 8840
rect 12620 8580 12820 8780
rect 13500 8780 13510 8840
rect 13690 8780 13700 8840
rect 13500 8580 13700 8780
rect 14160 8780 14170 8840
rect 14350 8780 14360 8840
rect 14160 8580 14360 8780
rect 14820 8780 14830 8840
rect 15010 8780 15020 8840
rect 14820 8580 15020 8780
rect 15700 8700 15900 8840
rect 15700 8640 15710 8700
rect 15890 8640 15900 8700
rect 15700 8580 15900 8640
rect 16360 8700 16560 8840
rect 16360 8640 16370 8700
rect 16550 8640 16560 8700
rect 16360 8580 16560 8640
rect 17020 8700 17220 8840
rect 17020 8640 17030 8700
rect 17210 8640 17220 8700
rect 17020 8580 17220 8640
rect 17900 8700 18100 8840
rect 17900 8640 17910 8700
rect 18090 8640 18100 8700
rect 17900 8580 18100 8640
rect 18560 8700 18760 8840
rect 18560 8640 18570 8700
rect 18750 8640 18760 8700
rect 18560 8580 18760 8640
rect 19220 8700 19420 8840
rect 19220 8640 19230 8700
rect 19410 8640 19420 8700
rect 19220 8580 19420 8640
rect 2458 8574 4058 8580
rect 2458 8540 2470 8574
rect 4046 8540 4058 8574
rect 4658 8574 6258 8580
rect 4658 8540 4670 8574
rect 6246 8540 6258 8574
rect 6858 8574 8458 8580
rect 6858 8540 6870 8574
rect 8446 8540 8458 8574
rect 9058 8574 10658 8580
rect 9058 8540 9070 8574
rect 10646 8540 10658 8574
rect 11258 8574 12858 8580
rect 11258 8540 11270 8574
rect 12846 8540 12858 8574
rect 13458 8574 15058 8580
rect 13458 8540 13470 8574
rect 15046 8540 15058 8574
rect 15658 8574 17258 8580
rect 15658 8540 15670 8574
rect 17246 8540 17258 8574
rect 17858 8574 19458 8580
rect 17858 8540 17870 8574
rect 19446 8540 19458 8574
rect -90 8530 10 8540
rect -90 8470 -70 8530
rect -10 8470 10 8530
rect -90 8460 10 8470
rect 2110 8530 2210 8540
rect 2458 8534 4058 8540
rect 2110 8470 2130 8530
rect 2190 8470 2210 8530
rect 4310 8530 4410 8540
rect 4658 8534 6258 8540
rect 2110 8460 2210 8470
rect 2380 8512 2426 8524
rect 1610 8410 1690 8420
rect 1610 8260 1620 8410
rect 1680 8310 1690 8410
rect 2380 8310 2386 8512
rect 1680 8260 2386 8310
rect 1610 8250 2386 8260
rect 2380 8244 2386 8250
rect 2420 8244 2426 8512
rect 2380 8232 2426 8244
rect 4090 8512 4136 8524
rect 4090 8244 4096 8512
rect 4130 8420 4136 8512
rect 4310 8470 4330 8530
rect 4390 8470 4410 8530
rect 6510 8530 6610 8540
rect 6858 8534 8458 8540
rect 4310 8460 4410 8470
rect 4580 8512 4626 8524
rect 4130 8360 4510 8420
rect 4130 8244 4136 8360
rect 4580 8310 4586 8512
rect 4210 8250 4440 8310
rect 4500 8250 4586 8310
rect 4090 8232 4136 8244
rect 4580 8244 4586 8250
rect 4620 8244 4626 8512
rect 4580 8232 4626 8244
rect 6290 8512 6336 8524
rect 6290 8244 6296 8512
rect 6330 8420 6336 8512
rect 6510 8470 6530 8530
rect 6590 8470 6610 8530
rect 8710 8530 8810 8540
rect 9058 8534 10658 8540
rect 6510 8460 6610 8470
rect 6780 8512 6826 8524
rect 6330 8360 6640 8420
rect 6700 8360 6710 8420
rect 6330 8244 6336 8360
rect 6780 8310 6786 8512
rect 6410 8250 6420 8310
rect 6480 8250 6786 8310
rect 6290 8232 6336 8244
rect 6780 8244 6786 8250
rect 6820 8244 6826 8512
rect 6780 8232 6826 8244
rect 8490 8512 8536 8524
rect 8490 8244 8496 8512
rect 8530 8420 8536 8512
rect 8710 8470 8730 8530
rect 8790 8470 8810 8530
rect 10910 8530 11010 8540
rect 11258 8534 12858 8540
rect 8710 8460 8810 8470
rect 8980 8512 9026 8524
rect 8530 8360 8620 8420
rect 8680 8360 8910 8420
rect 8530 8244 8536 8360
rect 8980 8310 8986 8512
rect 8610 8250 8620 8310
rect 8680 8250 8986 8310
rect 8490 8232 8536 8244
rect 8980 8244 8986 8250
rect 9020 8244 9026 8512
rect 8980 8232 9026 8244
rect 10690 8512 10736 8524
rect 10690 8244 10696 8512
rect 10730 8420 10736 8512
rect 10910 8470 10930 8530
rect 10990 8470 11010 8530
rect 13110 8530 13210 8540
rect 13458 8534 15058 8540
rect 10910 8460 11010 8470
rect 11180 8512 11226 8524
rect 10730 8360 10820 8420
rect 10880 8360 11110 8420
rect 10730 8244 10736 8360
rect 11180 8310 11186 8512
rect 10810 8250 10820 8310
rect 10880 8250 11186 8310
rect 10690 8232 10736 8244
rect 11180 8244 11186 8250
rect 11220 8244 11226 8512
rect 11180 8232 11226 8244
rect 12890 8512 12936 8524
rect 12890 8244 12896 8512
rect 12930 8420 12936 8512
rect 13110 8470 13130 8530
rect 13190 8470 13210 8530
rect 15310 8530 15410 8540
rect 15658 8534 17258 8540
rect 13110 8460 13210 8470
rect 13380 8512 13426 8524
rect 12930 8360 13020 8420
rect 13080 8360 13310 8420
rect 12930 8244 12936 8360
rect 13380 8310 13386 8512
rect 13010 8250 13020 8310
rect 13080 8250 13386 8310
rect 12890 8232 12936 8244
rect 13380 8244 13386 8250
rect 13420 8244 13426 8512
rect 13380 8232 13426 8244
rect 15090 8512 15136 8524
rect 15090 8244 15096 8512
rect 15130 8420 15136 8512
rect 15310 8470 15330 8530
rect 15390 8470 15410 8530
rect 17510 8530 17610 8540
rect 17858 8534 19458 8540
rect 15310 8460 15410 8470
rect 15580 8512 15626 8524
rect 15130 8360 15220 8420
rect 15280 8360 15510 8420
rect 15130 8244 15136 8360
rect 15580 8310 15586 8512
rect 15210 8250 15440 8310
rect 15500 8250 15586 8310
rect 15090 8232 15136 8244
rect 15580 8244 15586 8250
rect 15620 8244 15626 8512
rect 15580 8232 15626 8244
rect 17290 8512 17336 8524
rect 17290 8244 17296 8512
rect 17330 8420 17336 8512
rect 17510 8470 17530 8530
rect 17590 8470 17610 8530
rect 19710 8530 19810 8540
rect 17510 8460 17610 8470
rect 17780 8512 17826 8524
rect 17330 8360 17640 8420
rect 17700 8360 17710 8420
rect 17330 8244 17336 8360
rect 17780 8310 17786 8512
rect 17410 8250 17786 8310
rect 17290 8232 17336 8244
rect 17780 8244 17786 8250
rect 17820 8244 17826 8512
rect 17780 8232 17826 8244
rect 19490 8512 19536 8524
rect 19490 8244 19496 8512
rect 19530 8400 19536 8512
rect 19710 8470 19730 8530
rect 19790 8470 19810 8530
rect 21910 8530 22010 8540
rect 19710 8460 19810 8470
rect 20430 8500 20510 8510
rect 20430 8400 20440 8500
rect 19530 8350 20440 8400
rect 20500 8350 20510 8500
rect 21910 8470 21930 8530
rect 21990 8470 22010 8530
rect 21910 8460 22010 8470
rect 19530 8340 20510 8350
rect 19530 8244 19536 8340
rect 19490 8232 19536 8244
rect 2458 8216 4058 8222
rect 420 8190 620 8200
rect 420 8110 430 8190
rect 610 8180 620 8190
rect 2458 8182 2470 8216
rect 4046 8182 4058 8216
rect 2458 8180 4058 8182
rect 610 8176 4058 8180
rect 4658 8216 6258 8222
rect 4658 8182 4670 8216
rect 6246 8182 6258 8216
rect 4658 8176 4710 8182
rect 610 8120 4040 8176
rect 4700 8150 4710 8176
rect 6210 8176 6258 8182
rect 6858 8216 8458 8222
rect 6858 8182 6870 8216
rect 8446 8182 8458 8216
rect 6858 8176 6910 8182
rect 6210 8150 6220 8176
rect 4700 8140 6220 8150
rect 6900 8150 6910 8176
rect 8410 8176 8458 8182
rect 9058 8216 10658 8222
rect 9058 8182 9070 8216
rect 10646 8182 10658 8216
rect 9058 8176 9110 8182
rect 8410 8150 8420 8176
rect 6900 8140 8420 8150
rect 9100 8150 9110 8176
rect 10610 8176 10658 8182
rect 11258 8216 12858 8222
rect 11258 8182 11270 8216
rect 12846 8182 12858 8216
rect 11258 8176 11310 8182
rect 10610 8150 10620 8176
rect 9100 8140 10620 8150
rect 11300 8150 11310 8176
rect 12810 8176 12858 8182
rect 13458 8216 15058 8222
rect 13458 8182 13470 8216
rect 15046 8182 15058 8216
rect 13458 8176 13510 8182
rect 12810 8150 12820 8176
rect 11300 8140 12820 8150
rect 13500 8150 13510 8176
rect 15010 8176 15058 8182
rect 15658 8216 17258 8222
rect 15658 8182 15670 8216
rect 17246 8182 17258 8216
rect 15658 8176 15710 8182
rect 15010 8150 15020 8176
rect 13500 8140 15020 8150
rect 15700 8150 15710 8176
rect 17210 8176 17258 8182
rect 17858 8216 19458 8222
rect 17858 8182 17870 8216
rect 19446 8182 19458 8216
rect 17858 8180 19458 8182
rect 21300 8190 21500 8200
rect 21300 8180 21310 8190
rect 17858 8176 21310 8180
rect 17210 8150 17220 8176
rect 15700 8140 17220 8150
rect 17880 8120 21310 8176
rect 610 8110 620 8120
rect 420 8100 620 8110
rect 21300 8110 21310 8120
rect 21490 8110 21500 8190
rect 21300 8100 21500 8110
rect 2500 7900 2700 8040
rect 2500 7840 2510 7900
rect 2690 7840 2700 7900
rect 2500 7780 2700 7840
rect 3160 7900 3360 8040
rect 3160 7840 3170 7900
rect 3350 7840 3360 7900
rect 3160 7780 3360 7840
rect 3820 7900 4020 8040
rect 3820 7840 3830 7900
rect 4010 7840 4020 7900
rect 3820 7780 4020 7840
rect 4700 7900 4900 8040
rect 4700 7840 4710 7900
rect 4890 7840 4900 7900
rect 4700 7780 4900 7840
rect 5360 7900 5560 8040
rect 5360 7840 5370 7900
rect 5550 7840 5560 7900
rect 5360 7780 5560 7840
rect 6020 7900 6220 8040
rect 6020 7840 6030 7900
rect 6210 7840 6220 7900
rect 6020 7780 6220 7840
rect 6900 7980 6910 8040
rect 7090 7980 7100 8040
rect 6900 7780 7100 7980
rect 7560 7980 7570 8040
rect 7750 7980 7760 8040
rect 7560 7780 7760 7980
rect 8220 7980 8230 8040
rect 8410 7980 8420 8040
rect 8220 7780 8420 7980
rect 9100 7980 9110 8040
rect 9290 7980 9300 8040
rect 9100 7780 9300 7980
rect 9760 7980 9770 8040
rect 9950 7980 9960 8040
rect 9760 7780 9960 7980
rect 10420 7980 10430 8040
rect 10610 7980 10620 8040
rect 10420 7780 10620 7980
rect 11300 7980 11310 8040
rect 11490 7980 11500 8040
rect 11300 7780 11500 7980
rect 11960 7980 11970 8040
rect 12150 7980 12160 8040
rect 11960 7780 12160 7980
rect 12620 7980 12630 8040
rect 12810 7980 12820 8040
rect 12620 7780 12820 7980
rect 13500 7980 13510 8040
rect 13690 7980 13700 8040
rect 13500 7780 13700 7980
rect 14160 7980 14170 8040
rect 14350 7980 14360 8040
rect 14160 7780 14360 7980
rect 14820 7980 14830 8040
rect 15010 7980 15020 8040
rect 14820 7780 15020 7980
rect 15700 7900 15900 8040
rect 15700 7840 15710 7900
rect 15890 7840 15900 7900
rect 15700 7780 15900 7840
rect 16360 7900 16560 8040
rect 16360 7840 16370 7900
rect 16550 7840 16560 7900
rect 16360 7780 16560 7840
rect 17020 7900 17220 8040
rect 17020 7840 17030 7900
rect 17210 7840 17220 7900
rect 17020 7780 17220 7840
rect 17900 7900 18100 8040
rect 17900 7840 17910 7900
rect 18090 7840 18100 7900
rect 17900 7780 18100 7840
rect 18560 7900 18760 8040
rect 18560 7840 18570 7900
rect 18750 7840 18760 7900
rect 18560 7780 18760 7840
rect 19220 7900 19420 8040
rect 19220 7840 19230 7900
rect 19410 7840 19420 7900
rect 19220 7780 19420 7840
rect 2458 7774 4058 7780
rect 2458 7740 2470 7774
rect 4046 7740 4058 7774
rect 4658 7774 6258 7780
rect 4658 7740 4670 7774
rect 6246 7740 6258 7774
rect 6858 7774 8458 7780
rect 6858 7740 6870 7774
rect 8446 7740 8458 7774
rect 9058 7774 10658 7780
rect 9058 7740 9070 7774
rect 10646 7740 10658 7774
rect 11258 7774 12858 7780
rect 11258 7740 11270 7774
rect 12846 7740 12858 7774
rect 13458 7774 15058 7780
rect 13458 7740 13470 7774
rect 15046 7740 15058 7774
rect 15658 7774 17258 7780
rect 15658 7740 15670 7774
rect 17246 7740 17258 7774
rect 17858 7774 19458 7780
rect 17858 7740 17870 7774
rect 19446 7740 19458 7774
rect -90 7730 10 7740
rect -90 7670 -70 7730
rect -10 7670 10 7730
rect -90 7660 10 7670
rect 2110 7730 2210 7740
rect 2458 7734 4058 7740
rect 2110 7670 2130 7730
rect 2190 7670 2210 7730
rect 4310 7730 4410 7740
rect 4658 7734 6258 7740
rect 2110 7660 2210 7670
rect 2380 7712 2426 7724
rect 1610 7610 1690 7620
rect 1610 7460 1620 7610
rect 1680 7510 1690 7610
rect 2380 7510 2386 7712
rect 1680 7460 2386 7510
rect 1610 7450 2386 7460
rect 2380 7444 2386 7450
rect 2420 7444 2426 7712
rect 2380 7432 2426 7444
rect 4090 7712 4136 7724
rect 4090 7444 4096 7712
rect 4130 7620 4136 7712
rect 4310 7670 4330 7730
rect 4390 7670 4410 7730
rect 6510 7730 6610 7740
rect 6858 7734 8458 7740
rect 4310 7660 4410 7670
rect 4580 7712 4626 7724
rect 4130 7560 4510 7620
rect 4130 7444 4136 7560
rect 4580 7510 4586 7712
rect 4210 7450 4440 7510
rect 4500 7450 4586 7510
rect 4090 7432 4136 7444
rect 4580 7444 4586 7450
rect 4620 7444 4626 7712
rect 4580 7432 4626 7444
rect 6290 7712 6336 7724
rect 6290 7444 6296 7712
rect 6330 7620 6336 7712
rect 6510 7670 6530 7730
rect 6590 7670 6610 7730
rect 8710 7730 8810 7740
rect 9058 7734 10658 7740
rect 6510 7660 6610 7670
rect 6780 7712 6826 7724
rect 6330 7560 6640 7620
rect 6700 7560 6710 7620
rect 6330 7444 6336 7560
rect 6780 7510 6786 7712
rect 6410 7450 6420 7510
rect 6480 7450 6786 7510
rect 6290 7432 6336 7444
rect 6780 7444 6786 7450
rect 6820 7444 6826 7712
rect 6780 7432 6826 7444
rect 8490 7712 8536 7724
rect 8490 7444 8496 7712
rect 8530 7620 8536 7712
rect 8710 7670 8730 7730
rect 8790 7670 8810 7730
rect 10910 7730 11010 7740
rect 11258 7734 12858 7740
rect 8710 7660 8810 7670
rect 8980 7712 9026 7724
rect 8530 7560 8620 7620
rect 8680 7560 8910 7620
rect 8530 7444 8536 7560
rect 8980 7510 8986 7712
rect 8610 7450 8620 7510
rect 8680 7450 8986 7510
rect 8490 7432 8536 7444
rect 8980 7444 8986 7450
rect 9020 7444 9026 7712
rect 8980 7432 9026 7444
rect 10690 7712 10736 7724
rect 10690 7444 10696 7712
rect 10730 7620 10736 7712
rect 10910 7670 10930 7730
rect 10990 7670 11010 7730
rect 13110 7730 13210 7740
rect 13458 7734 15058 7740
rect 10910 7660 11010 7670
rect 11180 7712 11226 7724
rect 10730 7560 10820 7620
rect 10880 7560 11110 7620
rect 10730 7444 10736 7560
rect 11180 7510 11186 7712
rect 10810 7450 10820 7510
rect 10880 7450 11186 7510
rect 10690 7432 10736 7444
rect 11180 7444 11186 7450
rect 11220 7444 11226 7712
rect 11180 7432 11226 7444
rect 12890 7712 12936 7724
rect 12890 7444 12896 7712
rect 12930 7620 12936 7712
rect 13110 7670 13130 7730
rect 13190 7670 13210 7730
rect 15310 7730 15410 7740
rect 15658 7734 17258 7740
rect 13110 7660 13210 7670
rect 13380 7712 13426 7724
rect 12930 7560 13020 7620
rect 13080 7560 13310 7620
rect 12930 7444 12936 7560
rect 13380 7510 13386 7712
rect 13010 7450 13020 7510
rect 13080 7450 13386 7510
rect 12890 7432 12936 7444
rect 13380 7444 13386 7450
rect 13420 7444 13426 7712
rect 13380 7432 13426 7444
rect 15090 7712 15136 7724
rect 15090 7444 15096 7712
rect 15130 7620 15136 7712
rect 15310 7670 15330 7730
rect 15390 7670 15410 7730
rect 17510 7730 17610 7740
rect 17858 7734 19458 7740
rect 15310 7660 15410 7670
rect 15580 7712 15626 7724
rect 15130 7560 15220 7620
rect 15280 7560 15510 7620
rect 15130 7444 15136 7560
rect 15580 7510 15586 7712
rect 15210 7450 15440 7510
rect 15500 7450 15586 7510
rect 15090 7432 15136 7444
rect 15580 7444 15586 7450
rect 15620 7444 15626 7712
rect 15580 7432 15626 7444
rect 17290 7712 17336 7724
rect 17290 7444 17296 7712
rect 17330 7620 17336 7712
rect 17510 7670 17530 7730
rect 17590 7670 17610 7730
rect 19710 7730 19810 7740
rect 17510 7660 17610 7670
rect 17780 7712 17826 7724
rect 17330 7560 17640 7620
rect 17700 7560 17710 7620
rect 17330 7444 17336 7560
rect 17780 7510 17786 7712
rect 17410 7450 17786 7510
rect 17290 7432 17336 7444
rect 17780 7444 17786 7450
rect 17820 7444 17826 7712
rect 17780 7432 17826 7444
rect 19490 7712 19536 7724
rect 19490 7444 19496 7712
rect 19530 7600 19536 7712
rect 19710 7670 19730 7730
rect 19790 7670 19810 7730
rect 21910 7730 22010 7740
rect 19710 7660 19810 7670
rect 20430 7700 20510 7710
rect 20430 7600 20440 7700
rect 19530 7550 20440 7600
rect 20500 7550 20510 7700
rect 21910 7670 21930 7730
rect 21990 7670 22010 7730
rect 21910 7660 22010 7670
rect 19530 7540 20510 7550
rect 19530 7444 19536 7540
rect 19490 7432 19536 7444
rect 2458 7416 4058 7422
rect 420 7390 620 7400
rect 420 7310 430 7390
rect 610 7380 620 7390
rect 2458 7382 2470 7416
rect 4046 7382 4058 7416
rect 2458 7380 4058 7382
rect 610 7376 4058 7380
rect 4658 7416 6258 7422
rect 4658 7382 4670 7416
rect 6246 7382 6258 7416
rect 4658 7376 4710 7382
rect 610 7320 4040 7376
rect 4700 7350 4710 7376
rect 6210 7376 6258 7382
rect 6858 7416 8458 7422
rect 6858 7382 6870 7416
rect 8446 7382 8458 7416
rect 6858 7376 6910 7382
rect 6210 7350 6220 7376
rect 4700 7340 6220 7350
rect 6900 7350 6910 7376
rect 8410 7376 8458 7382
rect 9058 7416 10658 7422
rect 9058 7382 9070 7416
rect 10646 7382 10658 7416
rect 9058 7376 9110 7382
rect 8410 7350 8420 7376
rect 6900 7340 8420 7350
rect 9100 7350 9110 7376
rect 10610 7376 10658 7382
rect 11258 7416 12858 7422
rect 11258 7382 11270 7416
rect 12846 7382 12858 7416
rect 11258 7376 11310 7382
rect 10610 7350 10620 7376
rect 9100 7340 10620 7350
rect 11300 7350 11310 7376
rect 12810 7376 12858 7382
rect 13458 7416 15058 7422
rect 13458 7382 13470 7416
rect 15046 7382 15058 7416
rect 13458 7376 13510 7382
rect 12810 7350 12820 7376
rect 11300 7340 12820 7350
rect 13500 7350 13510 7376
rect 15010 7376 15058 7382
rect 15658 7416 17258 7422
rect 15658 7382 15670 7416
rect 17246 7382 17258 7416
rect 15658 7376 15710 7382
rect 15010 7350 15020 7376
rect 13500 7340 15020 7350
rect 15700 7350 15710 7376
rect 17210 7376 17258 7382
rect 17858 7416 19458 7422
rect 17858 7382 17870 7416
rect 19446 7382 19458 7416
rect 17858 7380 19458 7382
rect 21300 7390 21500 7400
rect 21300 7380 21310 7390
rect 17858 7376 21310 7380
rect 17210 7350 17220 7376
rect 15700 7340 17220 7350
rect 17880 7320 21310 7376
rect 610 7310 620 7320
rect 420 7300 620 7310
rect 21300 7310 21310 7320
rect 21490 7310 21500 7390
rect 21300 7300 21500 7310
rect 2500 7180 2510 7240
rect 2690 7180 2700 7240
rect 2500 6980 2700 7180
rect 3160 7180 3170 7240
rect 3350 7180 3360 7240
rect 3160 6980 3360 7180
rect 3820 7180 3830 7240
rect 4010 7180 4020 7240
rect 3820 6980 4020 7180
rect 4700 7180 4710 7240
rect 4890 7180 4900 7240
rect 4700 6980 4900 7180
rect 5360 7180 5370 7240
rect 5550 7180 5560 7240
rect 5360 6980 5560 7180
rect 6020 7180 6030 7240
rect 6210 7180 6220 7240
rect 6020 6980 6220 7180
rect 6900 7100 7100 7240
rect 6900 7040 6910 7100
rect 7090 7040 7100 7100
rect 6900 6980 7100 7040
rect 7560 7100 7760 7240
rect 7560 7040 7570 7100
rect 7750 7040 7760 7100
rect 7560 6980 7760 7040
rect 8220 7100 8420 7240
rect 8220 7040 8230 7100
rect 8410 7040 8420 7100
rect 8220 6980 8420 7040
rect 9100 7100 9300 7240
rect 9100 7040 9110 7100
rect 9290 7040 9300 7100
rect 9100 6980 9300 7040
rect 9760 7100 9960 7240
rect 9760 7040 9770 7100
rect 9950 7040 9960 7100
rect 9760 6980 9960 7040
rect 10420 7100 10620 7240
rect 10420 7040 10430 7100
rect 10610 7040 10620 7100
rect 10420 6980 10620 7040
rect 11300 7100 11500 7240
rect 11300 7040 11310 7100
rect 11490 7040 11500 7100
rect 11300 6980 11500 7040
rect 11960 7100 12160 7240
rect 11960 7040 11970 7100
rect 12150 7040 12160 7100
rect 11960 6980 12160 7040
rect 12620 7100 12820 7240
rect 12620 7040 12630 7100
rect 12810 7040 12820 7100
rect 12620 6980 12820 7040
rect 13500 7100 13700 7240
rect 13500 7040 13510 7100
rect 13690 7040 13700 7100
rect 13500 6980 13700 7040
rect 14160 7100 14360 7240
rect 14160 7040 14170 7100
rect 14350 7040 14360 7100
rect 14160 6980 14360 7040
rect 14820 7100 15020 7240
rect 14820 7040 14830 7100
rect 15010 7040 15020 7100
rect 14820 6980 15020 7040
rect 15700 7180 15710 7240
rect 15890 7180 15900 7240
rect 15700 6980 15900 7180
rect 16360 7180 16370 7240
rect 16550 7180 16560 7240
rect 16360 6980 16560 7180
rect 17020 7180 17030 7240
rect 17210 7180 17220 7240
rect 17020 6980 17220 7180
rect 17900 7180 17910 7240
rect 18090 7180 18100 7240
rect 17900 6980 18100 7180
rect 18560 7180 18570 7240
rect 18750 7180 18760 7240
rect 18560 6980 18760 7180
rect 19220 7180 19230 7240
rect 19410 7180 19420 7240
rect 19220 6980 19420 7180
rect 2458 6974 4058 6980
rect 2458 6940 2470 6974
rect 4046 6940 4058 6974
rect 4658 6974 6258 6980
rect 4658 6940 4670 6974
rect 6246 6940 6258 6974
rect 6858 6974 8458 6980
rect 6858 6940 6870 6974
rect 8446 6940 8458 6974
rect 9058 6974 10658 6980
rect 9058 6940 9070 6974
rect 10646 6940 10658 6974
rect 11258 6974 12858 6980
rect 11258 6940 11270 6974
rect 12846 6940 12858 6974
rect 13458 6974 15058 6980
rect 13458 6940 13470 6974
rect 15046 6940 15058 6974
rect 15658 6974 17258 6980
rect 15658 6940 15670 6974
rect 17246 6940 17258 6974
rect 17858 6974 19458 6980
rect 17858 6940 17870 6974
rect 19446 6940 19458 6974
rect -90 6930 10 6940
rect -90 6870 -70 6930
rect -10 6870 10 6930
rect -90 6860 10 6870
rect 2110 6930 2210 6940
rect 2458 6934 4058 6940
rect 2110 6870 2130 6930
rect 2190 6870 2210 6930
rect 4310 6930 4410 6940
rect 4658 6934 6258 6940
rect 2110 6860 2210 6870
rect 2380 6912 2426 6924
rect 1410 6810 1490 6820
rect 1410 6660 1420 6810
rect 1480 6710 1490 6810
rect 2380 6710 2386 6912
rect 1480 6660 2386 6710
rect 1410 6650 2386 6660
rect 2380 6644 2386 6650
rect 2420 6644 2426 6912
rect 2380 6632 2426 6644
rect 4090 6912 4136 6924
rect 4090 6644 4096 6912
rect 4130 6820 4136 6912
rect 4310 6870 4330 6930
rect 4390 6870 4410 6930
rect 6510 6930 6610 6940
rect 6858 6934 8458 6940
rect 4310 6860 4410 6870
rect 4580 6912 4626 6924
rect 4130 6760 4510 6820
rect 4130 6644 4136 6760
rect 4580 6710 4586 6912
rect 4210 6650 4220 6710
rect 4280 6650 4586 6710
rect 4090 6632 4136 6644
rect 4580 6644 4586 6650
rect 4620 6644 4626 6912
rect 4580 6632 4626 6644
rect 6290 6912 6336 6924
rect 6290 6644 6296 6912
rect 6330 6820 6336 6912
rect 6510 6870 6530 6930
rect 6590 6870 6610 6930
rect 8710 6930 8810 6940
rect 9058 6934 10658 6940
rect 6510 6860 6610 6870
rect 6780 6912 6826 6924
rect 6330 6760 6420 6820
rect 6480 6760 6710 6820
rect 6330 6644 6336 6760
rect 6780 6710 6786 6912
rect 6410 6650 6640 6710
rect 6700 6650 6786 6710
rect 6290 6632 6336 6644
rect 6780 6644 6786 6650
rect 6820 6644 6826 6912
rect 6780 6632 6826 6644
rect 8490 6912 8536 6924
rect 8490 6644 8496 6912
rect 8530 6820 8536 6912
rect 8710 6870 8730 6930
rect 8790 6870 8810 6930
rect 10910 6930 11010 6940
rect 11258 6934 12858 6940
rect 8710 6860 8810 6870
rect 8980 6912 9026 6924
rect 8530 6760 8840 6820
rect 8900 6760 8910 6820
rect 8530 6644 8536 6760
rect 8980 6710 8986 6912
rect 8610 6650 8840 6710
rect 8900 6650 8986 6710
rect 8490 6632 8536 6644
rect 8980 6644 8986 6650
rect 9020 6644 9026 6912
rect 8980 6632 9026 6644
rect 10690 6912 10736 6924
rect 10690 6644 10696 6912
rect 10730 6820 10736 6912
rect 10910 6870 10930 6930
rect 10990 6870 11010 6930
rect 13110 6930 13210 6940
rect 13458 6934 15058 6940
rect 10910 6860 11010 6870
rect 11180 6912 11226 6924
rect 10730 6760 11040 6820
rect 11100 6760 11110 6820
rect 10730 6644 10736 6760
rect 11180 6710 11186 6912
rect 10810 6650 11040 6710
rect 11100 6650 11186 6710
rect 10690 6632 10736 6644
rect 11180 6644 11186 6650
rect 11220 6644 11226 6912
rect 11180 6632 11226 6644
rect 12890 6912 12936 6924
rect 12890 6644 12896 6912
rect 12930 6820 12936 6912
rect 13110 6870 13130 6930
rect 13190 6870 13210 6930
rect 15310 6930 15410 6940
rect 15658 6934 17258 6940
rect 13110 6860 13210 6870
rect 13380 6912 13426 6924
rect 12930 6760 13240 6820
rect 13300 6760 13310 6820
rect 12930 6644 12936 6760
rect 13380 6710 13386 6912
rect 13010 6650 13240 6710
rect 13300 6650 13386 6710
rect 12890 6632 12936 6644
rect 13380 6644 13386 6650
rect 13420 6644 13426 6912
rect 13380 6632 13426 6644
rect 15090 6912 15136 6924
rect 15090 6644 15096 6912
rect 15130 6820 15136 6912
rect 15310 6870 15330 6930
rect 15390 6870 15410 6930
rect 17510 6930 17610 6940
rect 17858 6934 19458 6940
rect 15310 6860 15410 6870
rect 15580 6912 15626 6924
rect 15130 6760 15440 6820
rect 15500 6760 15510 6820
rect 15130 6644 15136 6760
rect 15580 6710 15586 6912
rect 15210 6650 15220 6710
rect 15280 6650 15586 6710
rect 15090 6632 15136 6644
rect 15580 6644 15586 6650
rect 15620 6644 15626 6912
rect 15580 6632 15626 6644
rect 17290 6912 17336 6924
rect 17290 6644 17296 6912
rect 17330 6820 17336 6912
rect 17510 6870 17530 6930
rect 17590 6870 17610 6930
rect 19710 6930 19810 6940
rect 17510 6860 17610 6870
rect 17780 6912 17826 6924
rect 17330 6760 17420 6820
rect 17480 6760 17710 6820
rect 17330 6644 17336 6760
rect 17780 6710 17786 6912
rect 17410 6650 17786 6710
rect 17290 6632 17336 6644
rect 17780 6644 17786 6650
rect 17820 6644 17826 6912
rect 17780 6632 17826 6644
rect 19490 6912 19536 6924
rect 19490 6644 19496 6912
rect 19530 6800 19536 6912
rect 19710 6870 19730 6930
rect 19790 6870 19810 6930
rect 21910 6930 22010 6940
rect 19710 6860 19810 6870
rect 20230 6900 20310 6910
rect 20230 6800 20240 6900
rect 19530 6750 20240 6800
rect 20300 6750 20310 6900
rect 21910 6870 21930 6930
rect 21990 6870 22010 6930
rect 21910 6860 22010 6870
rect 19530 6740 20310 6750
rect 19530 6644 19536 6740
rect 19490 6632 19536 6644
rect 2458 6616 4058 6622
rect 420 6590 620 6600
rect 420 6510 430 6590
rect 610 6580 620 6590
rect 2458 6582 2470 6616
rect 4046 6582 4058 6616
rect 2458 6580 4058 6582
rect 610 6576 4058 6580
rect 4658 6616 6258 6622
rect 4658 6582 4670 6616
rect 6246 6582 6258 6616
rect 4658 6576 4710 6582
rect 610 6520 4040 6576
rect 4700 6550 4710 6576
rect 6210 6576 6258 6582
rect 6858 6616 8458 6622
rect 6858 6582 6870 6616
rect 8446 6582 8458 6616
rect 6858 6576 6910 6582
rect 6210 6550 6220 6576
rect 4700 6540 6220 6550
rect 6900 6550 6910 6576
rect 8410 6576 8458 6582
rect 9058 6616 10658 6622
rect 9058 6582 9070 6616
rect 10646 6582 10658 6616
rect 9058 6576 9110 6582
rect 8410 6550 8420 6576
rect 6900 6540 8420 6550
rect 9100 6550 9110 6576
rect 10610 6576 10658 6582
rect 11258 6616 12858 6622
rect 11258 6582 11270 6616
rect 12846 6582 12858 6616
rect 11258 6576 11310 6582
rect 10610 6550 10620 6576
rect 9100 6540 10620 6550
rect 11300 6550 11310 6576
rect 12810 6576 12858 6582
rect 13458 6616 15058 6622
rect 13458 6582 13470 6616
rect 15046 6582 15058 6616
rect 13458 6576 13510 6582
rect 12810 6550 12820 6576
rect 11300 6540 12820 6550
rect 13500 6550 13510 6576
rect 15010 6576 15058 6582
rect 15658 6616 17258 6622
rect 15658 6582 15670 6616
rect 17246 6582 17258 6616
rect 15658 6576 15710 6582
rect 15010 6550 15020 6576
rect 13500 6540 15020 6550
rect 15700 6550 15710 6576
rect 17210 6576 17258 6582
rect 17858 6616 19458 6622
rect 17858 6582 17870 6616
rect 19446 6582 19458 6616
rect 17858 6580 19458 6582
rect 21300 6590 21500 6600
rect 21300 6580 21310 6590
rect 17858 6576 21310 6580
rect 17210 6550 17220 6576
rect 15700 6540 17220 6550
rect 17880 6520 21310 6576
rect 610 6510 620 6520
rect 420 6500 620 6510
rect 21300 6510 21310 6520
rect 21490 6510 21500 6590
rect 21300 6500 21500 6510
rect 2500 6300 2700 6440
rect 2500 6240 2510 6300
rect 2690 6240 2700 6300
rect 2500 6180 2700 6240
rect 3160 6300 3360 6440
rect 3160 6240 3170 6300
rect 3350 6240 3360 6300
rect 3160 6180 3360 6240
rect 3820 6300 4020 6440
rect 3820 6240 3830 6300
rect 4010 6240 4020 6300
rect 3820 6180 4020 6240
rect 4700 6300 4900 6440
rect 4700 6240 4710 6300
rect 4890 6240 4900 6300
rect 4700 6180 4900 6240
rect 5360 6300 5560 6440
rect 5360 6240 5370 6300
rect 5550 6240 5560 6300
rect 5360 6180 5560 6240
rect 6020 6300 6220 6440
rect 6020 6240 6030 6300
rect 6210 6240 6220 6300
rect 6020 6180 6220 6240
rect 6900 6380 6910 6440
rect 7090 6380 7100 6440
rect 6900 6180 7100 6380
rect 7560 6380 7570 6440
rect 7750 6380 7760 6440
rect 7560 6180 7760 6380
rect 8220 6380 8230 6440
rect 8410 6380 8420 6440
rect 8220 6180 8420 6380
rect 9100 6380 9110 6440
rect 9290 6380 9300 6440
rect 9100 6180 9300 6380
rect 9760 6380 9770 6440
rect 9950 6380 9960 6440
rect 9760 6180 9960 6380
rect 10420 6380 10430 6440
rect 10610 6380 10620 6440
rect 10420 6180 10620 6380
rect 11300 6380 11310 6440
rect 11490 6380 11500 6440
rect 11300 6180 11500 6380
rect 11960 6380 11970 6440
rect 12150 6380 12160 6440
rect 11960 6180 12160 6380
rect 12620 6380 12630 6440
rect 12810 6380 12820 6440
rect 12620 6180 12820 6380
rect 13500 6380 13510 6440
rect 13690 6380 13700 6440
rect 13500 6180 13700 6380
rect 14160 6380 14170 6440
rect 14350 6380 14360 6440
rect 14160 6180 14360 6380
rect 14820 6380 14830 6440
rect 15010 6380 15020 6440
rect 14820 6180 15020 6380
rect 15700 6300 15900 6440
rect 15700 6240 15710 6300
rect 15890 6240 15900 6300
rect 15700 6180 15900 6240
rect 16360 6300 16560 6440
rect 16360 6240 16370 6300
rect 16550 6240 16560 6300
rect 16360 6180 16560 6240
rect 17020 6300 17220 6440
rect 17020 6240 17030 6300
rect 17210 6240 17220 6300
rect 17020 6180 17220 6240
rect 17900 6300 18100 6440
rect 17900 6240 17910 6300
rect 18090 6240 18100 6300
rect 17900 6180 18100 6240
rect 18560 6300 18760 6440
rect 18560 6240 18570 6300
rect 18750 6240 18760 6300
rect 18560 6180 18760 6240
rect 19220 6300 19420 6440
rect 19220 6240 19230 6300
rect 19410 6240 19420 6300
rect 19220 6180 19420 6240
rect 2458 6174 4058 6180
rect 2458 6140 2470 6174
rect 4046 6140 4058 6174
rect 4658 6174 6258 6180
rect 4658 6140 4670 6174
rect 6246 6140 6258 6174
rect 6858 6174 8458 6180
rect 6858 6140 6870 6174
rect 8446 6140 8458 6174
rect 9058 6174 10658 6180
rect 9058 6140 9070 6174
rect 10646 6140 10658 6174
rect 11258 6174 12858 6180
rect 11258 6140 11270 6174
rect 12846 6140 12858 6174
rect 13458 6174 15058 6180
rect 13458 6140 13470 6174
rect 15046 6140 15058 6174
rect 15658 6174 17258 6180
rect 15658 6140 15670 6174
rect 17246 6140 17258 6174
rect 17858 6174 19458 6180
rect 17858 6140 17870 6174
rect 19446 6140 19458 6174
rect -90 6130 10 6140
rect -90 6070 -70 6130
rect -10 6070 10 6130
rect -90 6060 10 6070
rect 2110 6130 2210 6140
rect 2458 6134 4058 6140
rect 2110 6070 2130 6130
rect 2190 6070 2210 6130
rect 4310 6130 4410 6140
rect 4658 6134 6258 6140
rect 2110 6060 2210 6070
rect 2380 6112 2426 6124
rect 2380 5910 2386 6112
rect 2010 5850 2240 5910
rect 2300 5850 2386 5910
rect 2380 5844 2386 5850
rect 2420 5844 2426 6112
rect 2380 5832 2426 5844
rect 4090 6112 4136 6124
rect 4090 5844 4096 6112
rect 4130 6020 4136 6112
rect 4310 6070 4330 6130
rect 4390 6070 4410 6130
rect 6510 6130 6610 6140
rect 6858 6134 8458 6140
rect 4310 6060 4410 6070
rect 4580 6112 4626 6124
rect 4130 5960 4440 6020
rect 4500 5960 4510 6020
rect 4130 5844 4136 5960
rect 4580 5910 4586 6112
rect 4210 5850 4440 5910
rect 4500 5850 4586 5910
rect 4090 5832 4136 5844
rect 4580 5844 4586 5850
rect 4620 5844 4626 6112
rect 4580 5832 4626 5844
rect 6290 6112 6336 6124
rect 6290 5844 6296 6112
rect 6330 6020 6336 6112
rect 6510 6070 6530 6130
rect 6590 6070 6610 6130
rect 8710 6130 8810 6140
rect 9058 6134 10658 6140
rect 6510 6060 6610 6070
rect 6780 6112 6826 6124
rect 6330 5960 6640 6020
rect 6700 5960 6710 6020
rect 6330 5844 6336 5960
rect 6780 5910 6786 6112
rect 6410 5850 6420 5910
rect 6480 5850 6786 5910
rect 6290 5832 6336 5844
rect 6780 5844 6786 5850
rect 6820 5844 6826 6112
rect 6780 5832 6826 5844
rect 8490 6112 8536 6124
rect 8490 5844 8496 6112
rect 8530 6020 8536 6112
rect 8710 6070 8730 6130
rect 8790 6070 8810 6130
rect 10910 6130 11010 6140
rect 11258 6134 12858 6140
rect 8710 6060 8810 6070
rect 8980 6112 9026 6124
rect 8530 5960 8620 6020
rect 8680 5960 8910 6020
rect 8530 5844 8536 5960
rect 8980 5910 8986 6112
rect 8610 5850 8620 5910
rect 8680 5850 8986 5910
rect 8490 5832 8536 5844
rect 8980 5844 8986 5850
rect 9020 5844 9026 6112
rect 8980 5832 9026 5844
rect 10690 6112 10736 6124
rect 10690 5844 10696 6112
rect 10730 6020 10736 6112
rect 10910 6070 10930 6130
rect 10990 6070 11010 6130
rect 13110 6130 13210 6140
rect 13458 6134 15058 6140
rect 10910 6060 11010 6070
rect 11180 6112 11226 6124
rect 10730 5960 10820 6020
rect 10880 5960 11110 6020
rect 10730 5844 10736 5960
rect 11180 5910 11186 6112
rect 10810 5850 10820 5910
rect 10880 5850 11186 5910
rect 10690 5832 10736 5844
rect 11180 5844 11186 5850
rect 11220 5844 11226 6112
rect 11180 5832 11226 5844
rect 12890 6112 12936 6124
rect 12890 5844 12896 6112
rect 12930 6020 12936 6112
rect 13110 6070 13130 6130
rect 13190 6070 13210 6130
rect 15310 6130 15410 6140
rect 15658 6134 17258 6140
rect 13110 6060 13210 6070
rect 13380 6112 13426 6124
rect 12930 5960 13020 6020
rect 13080 5960 13310 6020
rect 12930 5844 12936 5960
rect 13380 5910 13386 6112
rect 13010 5850 13020 5910
rect 13080 5850 13386 5910
rect 12890 5832 12936 5844
rect 13380 5844 13386 5850
rect 13420 5844 13426 6112
rect 13380 5832 13426 5844
rect 15090 6112 15136 6124
rect 15090 5844 15096 6112
rect 15130 6020 15136 6112
rect 15310 6070 15330 6130
rect 15390 6070 15410 6130
rect 17510 6130 17610 6140
rect 17858 6134 19458 6140
rect 15310 6060 15410 6070
rect 15580 6112 15626 6124
rect 15130 5960 15220 6020
rect 15280 5960 15510 6020
rect 15130 5844 15136 5960
rect 15580 5910 15586 6112
rect 15210 5850 15440 5910
rect 15500 5850 15586 5910
rect 15090 5832 15136 5844
rect 15580 5844 15586 5850
rect 15620 5844 15626 6112
rect 15580 5832 15626 5844
rect 17290 6112 17336 6124
rect 17290 5844 17296 6112
rect 17330 6020 17336 6112
rect 17510 6070 17530 6130
rect 17590 6070 17610 6130
rect 19710 6130 19810 6140
rect 17510 6060 17610 6070
rect 17780 6112 17826 6124
rect 17330 5960 17640 6020
rect 17700 5960 17710 6020
rect 17330 5844 17336 5960
rect 17780 5910 17786 6112
rect 17410 5850 17640 5910
rect 17700 5850 17786 5910
rect 17290 5832 17336 5844
rect 17780 5844 17786 5850
rect 17820 5844 17826 6112
rect 17780 5832 17826 5844
rect 19490 6112 19536 6124
rect 19490 5844 19496 6112
rect 19530 6000 19536 6112
rect 19710 6070 19730 6130
rect 19790 6070 19810 6130
rect 19710 6060 19810 6070
rect 21910 6130 22010 6140
rect 21910 6070 21930 6130
rect 21990 6070 22010 6130
rect 21910 6060 22010 6070
rect 19530 5940 19840 6000
rect 19900 5940 19910 6000
rect 19530 5844 19536 5940
rect 19490 5832 19536 5844
rect 2458 5816 4058 5822
rect 2458 5782 2470 5816
rect 4046 5782 4058 5816
rect 2458 5776 2510 5782
rect 2500 5750 2510 5776
rect 4010 5776 4058 5782
rect 4658 5816 6258 5822
rect 4658 5782 4670 5816
rect 6246 5782 6258 5816
rect 4658 5776 4710 5782
rect 4010 5750 4020 5776
rect 2500 5740 4020 5750
rect 4700 5750 4710 5776
rect 6210 5776 6258 5782
rect 6858 5816 8458 5822
rect 6858 5782 6870 5816
rect 8446 5782 8458 5816
rect 6858 5776 6910 5782
rect 6210 5750 6220 5776
rect 4700 5740 6220 5750
rect 6900 5750 6910 5776
rect 8410 5776 8458 5782
rect 9058 5816 10658 5822
rect 9058 5782 9070 5816
rect 10646 5782 10658 5816
rect 9058 5776 9110 5782
rect 8410 5750 8420 5776
rect 6900 5740 8420 5750
rect 9100 5750 9110 5776
rect 10610 5776 10658 5782
rect 11258 5816 12858 5822
rect 11258 5782 11270 5816
rect 12846 5782 12858 5816
rect 11258 5776 11310 5782
rect 10610 5750 10620 5776
rect 9100 5740 10620 5750
rect 11300 5750 11310 5776
rect 12810 5776 12858 5782
rect 13458 5816 15058 5822
rect 13458 5782 13470 5816
rect 15046 5782 15058 5816
rect 13458 5776 13510 5782
rect 12810 5750 12820 5776
rect 11300 5740 12820 5750
rect 13500 5750 13510 5776
rect 15010 5776 15058 5782
rect 15658 5816 17258 5822
rect 15658 5782 15670 5816
rect 17246 5782 17258 5816
rect 15658 5776 15710 5782
rect 15010 5750 15020 5776
rect 13500 5740 15020 5750
rect 15700 5750 15710 5776
rect 17210 5776 17258 5782
rect 17858 5816 19458 5822
rect 17858 5782 17870 5816
rect 19446 5782 19458 5816
rect 17858 5776 17910 5782
rect 17210 5750 17220 5776
rect 15700 5740 17220 5750
rect 17900 5750 17910 5776
rect 19410 5776 19458 5782
rect 19410 5750 19420 5776
rect 17900 5740 19420 5750
rect 2500 5580 2510 5640
rect 2690 5580 2700 5640
rect 2500 5380 2700 5580
rect 3160 5580 3170 5640
rect 3350 5580 3360 5640
rect 3160 5380 3360 5580
rect 3820 5580 3830 5640
rect 4010 5580 4020 5640
rect 3820 5380 4020 5580
rect 4700 5580 4710 5640
rect 4890 5580 4900 5640
rect 4700 5380 4900 5580
rect 5360 5580 5370 5640
rect 5550 5580 5560 5640
rect 5360 5380 5560 5580
rect 6020 5580 6030 5640
rect 6210 5580 6220 5640
rect 6020 5380 6220 5580
rect 6900 5500 7100 5640
rect 6900 5440 6910 5500
rect 7090 5440 7100 5500
rect 6900 5380 7100 5440
rect 7560 5500 7760 5640
rect 7560 5440 7570 5500
rect 7750 5440 7760 5500
rect 7560 5380 7760 5440
rect 8220 5500 8420 5640
rect 8220 5440 8230 5500
rect 8410 5440 8420 5500
rect 8220 5380 8420 5440
rect 9100 5500 9300 5640
rect 9100 5440 9110 5500
rect 9290 5440 9300 5500
rect 9100 5380 9300 5440
rect 9760 5500 9960 5640
rect 9760 5440 9770 5500
rect 9950 5440 9960 5500
rect 9760 5380 9960 5440
rect 10420 5500 10620 5640
rect 10420 5440 10430 5500
rect 10610 5440 10620 5500
rect 10420 5380 10620 5440
rect 11300 5500 11500 5640
rect 11300 5440 11310 5500
rect 11490 5440 11500 5500
rect 11300 5380 11500 5440
rect 11960 5500 12160 5640
rect 11960 5440 11970 5500
rect 12150 5440 12160 5500
rect 11960 5380 12160 5440
rect 12620 5500 12820 5640
rect 12620 5440 12630 5500
rect 12810 5440 12820 5500
rect 12620 5380 12820 5440
rect 13500 5500 13700 5640
rect 13500 5440 13510 5500
rect 13690 5440 13700 5500
rect 13500 5380 13700 5440
rect 14160 5500 14360 5640
rect 14160 5440 14170 5500
rect 14350 5440 14360 5500
rect 14160 5380 14360 5440
rect 14820 5500 15020 5640
rect 14820 5440 14830 5500
rect 15010 5440 15020 5500
rect 14820 5380 15020 5440
rect 15700 5580 15710 5640
rect 15890 5580 15900 5640
rect 15700 5380 15900 5580
rect 16360 5580 16370 5640
rect 16550 5580 16560 5640
rect 16360 5380 16560 5580
rect 17020 5580 17030 5640
rect 17210 5580 17220 5640
rect 17020 5380 17220 5580
rect 17900 5580 17910 5640
rect 18090 5580 18100 5640
rect 17900 5380 18100 5580
rect 18560 5580 18570 5640
rect 18750 5580 18760 5640
rect 18560 5380 18760 5580
rect 19220 5580 19230 5640
rect 19410 5580 19420 5640
rect 19220 5380 19420 5580
rect 2458 5374 4058 5380
rect 2458 5340 2470 5374
rect 4046 5340 4058 5374
rect 4658 5374 6258 5380
rect 4658 5340 4670 5374
rect 6246 5340 6258 5374
rect 6858 5374 8458 5380
rect 6858 5340 6870 5374
rect 8446 5340 8458 5374
rect 9058 5374 10658 5380
rect 9058 5340 9070 5374
rect 10646 5340 10658 5374
rect 11258 5374 12858 5380
rect 11258 5340 11270 5374
rect 12846 5340 12858 5374
rect 13458 5374 15058 5380
rect 13458 5340 13470 5374
rect 15046 5340 15058 5374
rect 15658 5374 17258 5380
rect 15658 5340 15670 5374
rect 17246 5340 17258 5374
rect 17858 5374 19458 5380
rect 17858 5340 17870 5374
rect 19446 5340 19458 5374
rect -90 5330 10 5340
rect -90 5270 -70 5330
rect -10 5270 10 5330
rect -90 5260 10 5270
rect 2110 5330 2210 5340
rect 2458 5334 4058 5340
rect 2110 5270 2130 5330
rect 2190 5270 2210 5330
rect 4310 5330 4410 5340
rect 4658 5334 6258 5340
rect 2110 5260 2210 5270
rect 2380 5312 2426 5324
rect 2380 5110 2386 5312
rect 2010 5050 2020 5110
rect 2080 5050 2386 5110
rect 2380 5044 2386 5050
rect 2420 5044 2426 5312
rect 2380 5032 2426 5044
rect 4090 5312 4136 5324
rect 4090 5044 4096 5312
rect 4130 5220 4136 5312
rect 4310 5270 4330 5330
rect 4390 5270 4410 5330
rect 6510 5330 6610 5340
rect 6858 5334 8458 5340
rect 4310 5260 4410 5270
rect 4580 5312 4626 5324
rect 4130 5160 4220 5220
rect 4280 5160 4510 5220
rect 4130 5044 4136 5160
rect 4580 5110 4586 5312
rect 4210 5050 4220 5110
rect 4280 5050 4586 5110
rect 4090 5032 4136 5044
rect 4580 5044 4586 5050
rect 4620 5044 4626 5312
rect 4580 5032 4626 5044
rect 6290 5312 6336 5324
rect 6290 5044 6296 5312
rect 6330 5220 6336 5312
rect 6510 5270 6530 5330
rect 6590 5270 6610 5330
rect 8710 5330 8810 5340
rect 9058 5334 10658 5340
rect 6510 5260 6610 5270
rect 6780 5312 6826 5324
rect 6330 5160 6420 5220
rect 6480 5160 6710 5220
rect 6330 5044 6336 5160
rect 6780 5110 6786 5312
rect 6410 5050 6640 5110
rect 6700 5050 6786 5110
rect 6290 5032 6336 5044
rect 6780 5044 6786 5050
rect 6820 5044 6826 5312
rect 6780 5032 6826 5044
rect 8490 5312 8536 5324
rect 8490 5044 8496 5312
rect 8530 5220 8536 5312
rect 8710 5270 8730 5330
rect 8790 5270 8810 5330
rect 10910 5330 11010 5340
rect 11258 5334 12858 5340
rect 8710 5260 8810 5270
rect 8980 5312 9026 5324
rect 8530 5160 8840 5220
rect 8900 5160 8910 5220
rect 8530 5044 8536 5160
rect 8980 5110 8986 5312
rect 8610 5050 8840 5110
rect 8900 5050 8986 5110
rect 8490 5032 8536 5044
rect 8980 5044 8986 5050
rect 9020 5044 9026 5312
rect 8980 5032 9026 5044
rect 10690 5312 10736 5324
rect 10690 5044 10696 5312
rect 10730 5220 10736 5312
rect 10910 5270 10930 5330
rect 10990 5270 11010 5330
rect 13110 5330 13210 5340
rect 13458 5334 15058 5340
rect 10910 5260 11010 5270
rect 11180 5312 11226 5324
rect 10730 5160 11040 5220
rect 11100 5160 11110 5220
rect 10730 5044 10736 5160
rect 11180 5110 11186 5312
rect 10810 5050 11040 5110
rect 11100 5050 11186 5110
rect 10690 5032 10736 5044
rect 11180 5044 11186 5050
rect 11220 5044 11226 5312
rect 11180 5032 11226 5044
rect 12890 5312 12936 5324
rect 12890 5044 12896 5312
rect 12930 5220 12936 5312
rect 13110 5270 13130 5330
rect 13190 5270 13210 5330
rect 15310 5330 15410 5340
rect 15658 5334 17258 5340
rect 13110 5260 13210 5270
rect 13380 5312 13426 5324
rect 12930 5160 13240 5220
rect 13300 5160 13310 5220
rect 12930 5044 12936 5160
rect 13380 5110 13386 5312
rect 13010 5050 13240 5110
rect 13300 5050 13386 5110
rect 12890 5032 12936 5044
rect 13380 5044 13386 5050
rect 13420 5044 13426 5312
rect 13380 5032 13426 5044
rect 15090 5312 15136 5324
rect 15090 5044 15096 5312
rect 15130 5220 15136 5312
rect 15310 5270 15330 5330
rect 15390 5270 15410 5330
rect 17510 5330 17610 5340
rect 17858 5334 19458 5340
rect 15310 5260 15410 5270
rect 15580 5312 15626 5324
rect 15130 5160 15440 5220
rect 15500 5160 15510 5220
rect 15130 5044 15136 5160
rect 15580 5110 15586 5312
rect 15210 5050 15220 5110
rect 15280 5050 15586 5110
rect 15090 5032 15136 5044
rect 15580 5044 15586 5050
rect 15620 5044 15626 5312
rect 15580 5032 15626 5044
rect 17290 5312 17336 5324
rect 17290 5044 17296 5312
rect 17330 5220 17336 5312
rect 17510 5270 17530 5330
rect 17590 5270 17610 5330
rect 19710 5330 19810 5340
rect 17510 5260 17610 5270
rect 17780 5312 17826 5324
rect 17330 5160 17420 5220
rect 17480 5160 17710 5220
rect 17330 5044 17336 5160
rect 17780 5110 17786 5312
rect 17410 5050 17420 5110
rect 17480 5050 17786 5110
rect 17290 5032 17336 5044
rect 17780 5044 17786 5050
rect 17820 5044 17826 5312
rect 17780 5032 17826 5044
rect 19490 5312 19536 5324
rect 19490 5044 19496 5312
rect 19530 5200 19536 5312
rect 19710 5270 19730 5330
rect 19790 5270 19810 5330
rect 19710 5260 19810 5270
rect 21910 5330 22010 5340
rect 21910 5270 21930 5330
rect 21990 5270 22010 5330
rect 21910 5260 22010 5270
rect 19530 5140 19620 5200
rect 19680 5140 19910 5200
rect 19530 5044 19536 5140
rect 19490 5032 19536 5044
rect 2458 5016 4058 5022
rect 2458 4982 2470 5016
rect 4046 4982 4058 5016
rect 2458 4976 2510 4982
rect 2500 4950 2510 4976
rect 4010 4976 4058 4982
rect 4658 5016 6258 5022
rect 4658 4982 4670 5016
rect 6246 4982 6258 5016
rect 4658 4976 4710 4982
rect 4010 4950 4020 4976
rect 2500 4940 4020 4950
rect 4700 4950 4710 4976
rect 6210 4976 6258 4982
rect 6858 5016 8458 5022
rect 6858 4982 6870 5016
rect 8446 4982 8458 5016
rect 6858 4976 6910 4982
rect 6210 4950 6220 4976
rect 4700 4940 6220 4950
rect 6900 4950 6910 4976
rect 8410 4976 8458 4982
rect 9058 5016 10658 5022
rect 9058 4982 9070 5016
rect 10646 4982 10658 5016
rect 9058 4976 9110 4982
rect 8410 4950 8420 4976
rect 6900 4940 8420 4950
rect 9100 4950 9110 4976
rect 10610 4976 10658 4982
rect 11258 5016 12858 5022
rect 11258 4982 11270 5016
rect 12846 4982 12858 5016
rect 11258 4976 11310 4982
rect 10610 4950 10620 4976
rect 9100 4940 10620 4950
rect 11300 4950 11310 4976
rect 12810 4976 12858 4982
rect 13458 5016 15058 5022
rect 13458 4982 13470 5016
rect 15046 4982 15058 5016
rect 13458 4976 13510 4982
rect 12810 4950 12820 4976
rect 11300 4940 12820 4950
rect 13500 4950 13510 4976
rect 15010 4976 15058 4982
rect 15658 5016 17258 5022
rect 15658 4982 15670 5016
rect 17246 4982 17258 5016
rect 15658 4976 15710 4982
rect 15010 4950 15020 4976
rect 13500 4940 15020 4950
rect 15700 4950 15710 4976
rect 17210 4976 17258 4982
rect 17858 5016 19458 5022
rect 17858 4982 17870 5016
rect 19446 4982 19458 5016
rect 17858 4976 17910 4982
rect 17210 4950 17220 4976
rect 15700 4940 17220 4950
rect 17900 4950 17910 4976
rect 19410 4976 19458 4982
rect 19410 4950 19420 4976
rect 17900 4940 19420 4950
rect 22230 4842 22236 11538
rect 22270 4842 22276 11538
rect 22370 11399 22382 11796
rect 22920 11399 22932 11796
rect 22370 11393 22932 11399
rect 23036 11796 23598 11802
rect 23036 11399 23048 11796
rect 23586 11790 23598 11796
rect 23702 11796 24264 11802
rect 23702 11790 23714 11796
rect 23586 11400 23714 11790
rect 23586 11399 23598 11400
rect 23036 11393 23598 11399
rect 23702 11399 23714 11400
rect 24252 11399 24264 11796
rect 23702 11393 24264 11399
rect 24368 11796 24930 11802
rect 24368 11399 24380 11796
rect 24918 11790 24930 11796
rect 25034 11796 25596 11802
rect 25034 11790 25046 11796
rect 24918 11400 25046 11790
rect 24918 11399 24930 11400
rect 24368 11393 24930 11399
rect 25034 11399 25046 11400
rect 25584 11399 25596 11796
rect 25034 11393 25596 11399
rect 25700 11796 26262 11802
rect 25700 11399 25712 11796
rect 26250 11399 26262 11796
rect 25700 11393 26262 11399
rect 26366 11796 26928 11802
rect 26366 11399 26378 11796
rect 26916 11399 26928 11796
rect 30084 11727 30130 11886
rect 30166 11800 30230 11805
rect 30324 11800 30388 11805
rect 30166 11799 30388 11800
rect 30166 11765 30178 11799
rect 30218 11765 30336 11799
rect 30376 11765 30388 11799
rect 30166 11760 30388 11765
rect 30166 11759 30230 11760
rect 30324 11759 30388 11760
rect 30084 11715 30142 11727
rect 27910 11592 28814 11598
rect 27910 11558 27922 11592
rect 28802 11558 28814 11592
rect 27910 11552 28814 11558
rect 26366 11393 26928 11399
rect 27022 11538 27068 11550
rect 22230 4830 22276 4842
rect 22370 4981 22932 4987
rect 7790 4680 7950 4690
rect 7790 4540 7800 4680
rect 7940 4660 7950 4680
rect 7940 4582 12840 4660
rect 22370 4584 22382 4981
rect 22920 4584 22932 4981
rect 7940 4576 12860 4582
rect 22370 4578 22932 4584
rect 23036 4981 23598 4987
rect 23036 4584 23048 4981
rect 23586 4584 23598 4981
rect 23036 4578 23598 4584
rect 23702 4981 24264 4987
rect 23702 4584 23714 4981
rect 24252 4980 24264 4981
rect 24368 4981 24930 4987
rect 24368 4980 24380 4981
rect 24252 4590 24380 4980
rect 24252 4584 24264 4590
rect 23702 4578 24264 4584
rect 24368 4584 24380 4590
rect 24918 4584 24930 4981
rect 24368 4578 24930 4584
rect 25034 4981 25596 4987
rect 25034 4584 25046 4981
rect 25584 4980 25596 4981
rect 25700 4981 26262 4987
rect 25700 4980 25712 4981
rect 25584 4590 25712 4980
rect 25584 4584 25596 4590
rect 25034 4578 25596 4584
rect 25700 4584 25712 4590
rect 26250 4584 26262 4981
rect 25700 4578 26262 4584
rect 26366 4981 26928 4987
rect 26366 4584 26378 4981
rect 26916 4584 26928 4981
rect 27022 4842 27028 11538
rect 27062 4842 27068 11538
rect 30084 11539 30102 11715
rect 30136 11539 30142 11715
rect 30084 11528 30142 11539
rect 30096 11527 30142 11528
rect 27250 11490 27330 11500
rect 30178 11495 30218 11759
rect 30254 11715 30300 11727
rect 30254 11539 30260 11715
rect 30294 11539 30300 11715
rect 30254 11527 30300 11539
rect 27250 11400 27260 11490
rect 27320 11464 27330 11490
rect 30166 11489 30230 11495
rect 27320 11458 28726 11464
rect 27320 11424 27938 11458
rect 28714 11424 28726 11458
rect 30166 11455 30178 11489
rect 30218 11455 30230 11489
rect 30166 11449 30230 11455
rect 30178 11448 30218 11449
rect 27320 11418 28726 11424
rect 30260 11418 30294 11527
rect 30336 11495 30376 11759
rect 30416 11727 30454 11886
rect 30704 11848 30756 11886
rect 30482 11799 30546 11805
rect 30482 11765 30494 11799
rect 30534 11765 30546 11799
rect 30482 11759 30546 11765
rect 30412 11715 30458 11727
rect 30412 11539 30418 11715
rect 30452 11539 30458 11715
rect 30412 11527 30458 11539
rect 30494 11495 30534 11759
rect 30570 11722 30670 11728
rect 30570 11532 30576 11722
rect 30664 11532 30670 11722
rect 30570 11526 30670 11532
rect 30324 11494 30388 11495
rect 30482 11494 30546 11495
rect 30324 11489 30546 11494
rect 30324 11455 30336 11489
rect 30376 11455 30494 11489
rect 30534 11455 30546 11489
rect 30324 11450 30546 11455
rect 30324 11449 30388 11450
rect 30482 11449 30546 11450
rect 27320 11400 27330 11418
rect 30148 11416 30294 11418
rect 27250 11390 27330 11400
rect 28767 11389 28813 11401
rect 27730 11330 27810 11340
rect 27730 11306 27740 11330
rect 27260 11260 27740 11306
rect 27730 11240 27740 11260
rect 27800 11306 27810 11330
rect 28767 11335 28773 11389
rect 28807 11335 28813 11389
rect 30148 11364 30154 11416
rect 30288 11364 30294 11416
rect 30148 11362 30294 11364
rect 28767 11323 28813 11335
rect 27800 11300 28726 11306
rect 27800 11266 27938 11300
rect 28714 11266 28726 11300
rect 27800 11260 28726 11266
rect 28770 11270 28810 11323
rect 30336 11280 30376 11449
rect 30494 11432 30534 11449
rect 30594 11326 30638 11526
rect 30704 11406 30710 11848
rect 30744 11406 30756 11848
rect 30830 11727 30874 11886
rect 30934 11805 30974 11806
rect 30921 11799 30985 11805
rect 30921 11765 30933 11799
rect 30973 11765 30985 11799
rect 30921 11759 30985 11765
rect 30830 11715 30897 11727
rect 30830 11539 30857 11715
rect 30891 11539 30897 11715
rect 30830 11527 30897 11539
rect 30830 11524 30874 11527
rect 30934 11495 30974 11759
rect 31034 11727 31078 11728
rect 31009 11715 31078 11727
rect 31009 11539 31015 11715
rect 31049 11539 31078 11715
rect 31009 11527 31078 11539
rect 30921 11489 30985 11495
rect 30921 11455 30933 11489
rect 30973 11455 30985 11489
rect 30921 11449 30985 11455
rect 30704 11394 30756 11406
rect 30594 11320 30744 11326
rect 30180 11270 30400 11280
rect 28770 11260 28850 11270
rect 27800 11240 27810 11260
rect 28770 11243 28780 11260
rect 27730 11230 27810 11240
rect 28767 11231 28780 11243
rect 27250 11170 27330 11180
rect 27250 11080 27260 11170
rect 27320 11148 27330 11170
rect 28767 11177 28773 11231
rect 28767 11165 28780 11177
rect 27320 11142 28726 11148
rect 27320 11108 27938 11142
rect 28714 11108 28726 11142
rect 27320 11102 28726 11108
rect 27320 11080 27330 11102
rect 28770 11085 28780 11165
rect 27250 11070 27330 11080
rect 28767 11073 28780 11085
rect 27730 11015 27810 11025
rect 27730 10990 27740 11015
rect 27260 10944 27740 10990
rect 27730 10925 27740 10944
rect 27800 10990 27810 11015
rect 28767 11019 28773 11073
rect 28840 11040 28850 11260
rect 30180 11190 30190 11270
rect 30390 11190 30400 11270
rect 30180 11180 30400 11190
rect 30594 11262 30600 11320
rect 30738 11262 30744 11320
rect 30594 11256 30744 11262
rect 30594 11198 30638 11256
rect 30934 11198 30974 11449
rect 28807 11030 28850 11040
rect 28807 11019 28813 11030
rect 28767 11007 28813 11019
rect 27800 10984 28726 10990
rect 27800 10950 27938 10984
rect 28714 10950 28726 10984
rect 27800 10944 28726 10950
rect 27800 10925 27810 10944
rect 28770 10927 28810 11007
rect 30336 10994 30376 11180
rect 30594 11138 30974 11198
rect 30268 10988 30512 10994
rect 30268 10954 30280 10988
rect 30500 10954 30512 10988
rect 27730 10915 27810 10925
rect 28767 10915 28813 10927
rect 27250 10855 27330 10865
rect 27250 10765 27260 10855
rect 27320 10832 27330 10855
rect 28767 10861 28773 10915
rect 28807 10861 28813 10915
rect 28767 10849 28813 10861
rect 30138 10895 30184 10907
rect 27320 10826 28726 10832
rect 27320 10792 27938 10826
rect 28714 10792 28726 10826
rect 27320 10786 28726 10792
rect 30138 10819 30144 10895
rect 30178 10819 30184 10895
rect 27320 10765 27330 10786
rect 27250 10755 27330 10765
rect 27910 10692 28814 10698
rect 27910 10658 27922 10692
rect 28802 10658 28814 10692
rect 27910 10652 28814 10658
rect 30138 10628 30184 10819
rect 30268 10760 30512 10954
rect 30620 10907 30664 11138
rect 30596 10895 30664 10907
rect 30596 10819 30602 10895
rect 30636 10819 30664 10895
rect 30596 10808 30664 10819
rect 30730 11045 30776 11104
rect 30596 10807 30642 10808
rect 30268 10726 30280 10760
rect 30500 10726 30512 10760
rect 30268 10720 30512 10726
rect 30730 10669 30736 11045
rect 30770 10669 30776 11045
rect 30934 10994 30974 11138
rect 31034 11198 31078 11527
rect 31270 11727 31314 11886
rect 31582 11848 31640 11886
rect 31374 11805 31414 11806
rect 31347 11799 31439 11805
rect 31347 11765 31359 11799
rect 31427 11765 31439 11799
rect 31347 11759 31439 11765
rect 31270 11715 31337 11727
rect 31270 11539 31297 11715
rect 31331 11539 31337 11715
rect 31270 11527 31337 11539
rect 31270 11524 31314 11527
rect 31374 11495 31414 11759
rect 31472 11727 31542 11728
rect 31449 11722 31542 11727
rect 31449 11715 31478 11722
rect 31449 11539 31455 11715
rect 31449 11536 31478 11539
rect 31536 11536 31542 11722
rect 31449 11530 31542 11536
rect 31449 11528 31516 11530
rect 31449 11527 31495 11528
rect 31347 11489 31439 11495
rect 31347 11455 31359 11489
rect 31427 11455 31439 11489
rect 31347 11449 31439 11455
rect 31374 11326 31414 11449
rect 31582 11406 31589 11848
rect 31623 11406 31640 11848
rect 31814 11805 31854 11806
rect 31787 11799 31879 11805
rect 31787 11765 31799 11799
rect 31867 11765 31879 11799
rect 31787 11759 31879 11765
rect 31731 11726 31777 11727
rect 31684 11720 31777 11726
rect 31684 11534 31690 11720
rect 31748 11715 31777 11720
rect 31771 11539 31777 11715
rect 31748 11534 31777 11539
rect 31684 11528 31777 11534
rect 31731 11527 31777 11528
rect 31814 11495 31854 11759
rect 31912 11727 31956 11886
rect 31889 11715 31956 11727
rect 31889 11539 31895 11715
rect 31929 11539 31956 11715
rect 31889 11527 31956 11539
rect 32284 11727 32330 11886
rect 32366 11800 32430 11805
rect 32524 11800 32588 11805
rect 32366 11799 32588 11800
rect 32366 11765 32378 11799
rect 32418 11765 32536 11799
rect 32576 11765 32588 11799
rect 32366 11760 32588 11765
rect 32366 11759 32430 11760
rect 32524 11759 32588 11760
rect 32284 11715 32342 11727
rect 32284 11539 32302 11715
rect 32336 11539 32342 11715
rect 32284 11528 32342 11539
rect 32296 11527 32342 11528
rect 31912 11524 31956 11527
rect 32378 11495 32418 11759
rect 32454 11715 32500 11727
rect 32454 11539 32460 11715
rect 32494 11539 32500 11715
rect 32454 11527 32500 11539
rect 31787 11489 31879 11495
rect 31787 11455 31799 11489
rect 31867 11455 31879 11489
rect 31787 11449 31879 11455
rect 32366 11489 32430 11495
rect 32366 11455 32378 11489
rect 32418 11455 32430 11489
rect 32366 11449 32430 11455
rect 31582 11394 31640 11406
rect 31264 11320 31414 11326
rect 31264 11262 31270 11320
rect 31408 11262 31414 11320
rect 31264 11256 31414 11262
rect 31814 11198 31854 11449
rect 32378 11448 32418 11449
rect 32460 11418 32494 11527
rect 32536 11495 32576 11759
rect 32616 11727 32654 11886
rect 32904 11848 32956 11886
rect 32682 11799 32746 11805
rect 32682 11765 32694 11799
rect 32734 11765 32746 11799
rect 32682 11759 32746 11765
rect 32612 11715 32658 11727
rect 32612 11539 32618 11715
rect 32652 11539 32658 11715
rect 32612 11527 32658 11539
rect 32694 11495 32734 11759
rect 32770 11722 32870 11728
rect 32770 11532 32776 11722
rect 32864 11532 32870 11722
rect 32770 11526 32870 11532
rect 32524 11494 32588 11495
rect 32682 11494 32746 11495
rect 32524 11489 32746 11494
rect 32524 11455 32536 11489
rect 32576 11455 32694 11489
rect 32734 11455 32746 11489
rect 32524 11450 32746 11455
rect 32524 11449 32588 11450
rect 32682 11449 32746 11450
rect 32348 11416 32494 11418
rect 32348 11364 32354 11416
rect 32488 11364 32494 11416
rect 32348 11362 32494 11364
rect 32536 11280 32576 11449
rect 32694 11432 32734 11449
rect 32794 11326 32838 11526
rect 32904 11406 32910 11848
rect 32944 11406 32956 11848
rect 33030 11727 33074 11886
rect 33134 11805 33174 11806
rect 33121 11799 33185 11805
rect 33121 11765 33133 11799
rect 33173 11765 33185 11799
rect 33121 11759 33185 11765
rect 33030 11715 33097 11727
rect 33030 11539 33057 11715
rect 33091 11539 33097 11715
rect 33030 11527 33097 11539
rect 33030 11524 33074 11527
rect 33134 11495 33174 11759
rect 33234 11727 33278 11728
rect 33209 11715 33278 11727
rect 33209 11539 33215 11715
rect 33249 11539 33278 11715
rect 33209 11527 33278 11539
rect 33121 11489 33185 11495
rect 33121 11455 33133 11489
rect 33173 11455 33185 11489
rect 33121 11449 33185 11455
rect 32904 11394 32956 11406
rect 32794 11320 32944 11326
rect 31034 11138 31854 11198
rect 32380 11270 32600 11280
rect 32380 11190 32390 11270
rect 32590 11190 32600 11270
rect 32380 11180 32600 11190
rect 32794 11262 32800 11320
rect 32938 11262 32944 11320
rect 32794 11256 32944 11262
rect 32794 11198 32838 11256
rect 33134 11198 33174 11449
rect 30922 10988 30986 10994
rect 30922 10954 30934 10988
rect 30974 10954 30986 10988
rect 30922 10948 30986 10954
rect 30852 10906 30898 10907
rect 30730 10628 30776 10669
rect 30032 10622 30776 10628
rect 30032 10588 30113 10622
rect 30667 10594 30776 10622
rect 30832 10895 30898 10906
rect 30667 10588 30748 10594
rect 27910 10552 28814 10558
rect 27910 10518 27922 10552
rect 28802 10518 28814 10552
rect 27910 10512 28814 10518
rect 27730 10450 27810 10460
rect 27730 10424 27740 10450
rect 27260 10378 27740 10424
rect 27730 10360 27740 10378
rect 27800 10424 27810 10450
rect 27800 10418 28726 10424
rect 27800 10384 27938 10418
rect 28714 10384 28726 10418
rect 27800 10378 28726 10384
rect 27800 10360 27810 10378
rect 27730 10350 27810 10360
rect 28767 10360 28813 10361
rect 28767 10349 28820 10360
rect 27370 10290 27450 10300
rect 27370 10266 27380 10290
rect 27260 10220 27380 10266
rect 27370 10200 27380 10220
rect 27440 10266 27450 10290
rect 28767 10295 28773 10349
rect 28807 10295 28820 10349
rect 30032 10346 30748 10588
rect 30832 10519 30858 10895
rect 30892 10519 30898 10895
rect 30832 10507 30898 10519
rect 30832 10346 30876 10507
rect 30934 10466 30974 10948
rect 31034 10907 31078 11138
rect 31374 10994 31414 11006
rect 31814 10994 31854 11006
rect 32536 10994 32576 11180
rect 32794 11138 33174 11198
rect 31362 10988 31638 10994
rect 31362 10954 31374 10988
rect 31414 10954 31638 10988
rect 31362 10948 31638 10954
rect 31802 10988 31866 10994
rect 31802 10954 31814 10988
rect 31854 10954 31866 10988
rect 31802 10948 31866 10954
rect 32468 10988 32712 10994
rect 32468 10954 32480 10988
rect 32700 10954 32712 10988
rect 31010 10895 31078 10907
rect 31292 10906 31338 10907
rect 31010 10519 31016 10895
rect 31050 10519 31078 10895
rect 31010 10508 31078 10519
rect 31270 10895 31338 10906
rect 31270 10519 31298 10895
rect 31332 10519 31338 10895
rect 31010 10507 31056 10508
rect 31270 10507 31338 10519
rect 30922 10460 30986 10466
rect 30922 10426 30934 10460
rect 30974 10426 30986 10460
rect 30922 10420 30986 10426
rect 31270 10346 31314 10507
rect 31374 10466 31414 10948
rect 31450 10906 31496 10907
rect 31590 10906 31638 10948
rect 31732 10906 31778 10907
rect 31450 10900 31542 10906
rect 31450 10895 31478 10900
rect 31450 10519 31456 10895
rect 31536 10556 31542 10900
rect 31590 10900 31778 10906
rect 31590 10860 31690 10900
rect 31748 10895 31778 10900
rect 31450 10514 31478 10519
rect 31536 10514 31638 10556
rect 31450 10510 31638 10514
rect 31450 10508 31542 10510
rect 31450 10507 31496 10508
rect 31590 10466 31638 10510
rect 31684 10514 31690 10860
rect 31772 10519 31778 10895
rect 31748 10514 31778 10519
rect 31684 10508 31778 10514
rect 31732 10507 31778 10508
rect 31814 10466 31854 10948
rect 31890 10906 31936 10907
rect 31890 10895 31958 10906
rect 31890 10519 31896 10895
rect 31930 10519 31958 10895
rect 32338 10895 32384 10907
rect 32338 10819 32344 10895
rect 32378 10819 32384 10895
rect 32338 10628 32384 10819
rect 32468 10760 32712 10954
rect 32820 10907 32864 11138
rect 32796 10895 32864 10907
rect 32796 10819 32802 10895
rect 32836 10819 32864 10895
rect 32796 10808 32864 10819
rect 32930 11045 32976 11104
rect 32796 10807 32842 10808
rect 32468 10726 32480 10760
rect 32700 10726 32712 10760
rect 32468 10720 32712 10726
rect 32930 10669 32936 11045
rect 32970 10669 32976 11045
rect 33134 10994 33174 11138
rect 33234 11198 33278 11527
rect 33470 11727 33514 11886
rect 33782 11848 33840 11886
rect 33574 11805 33614 11806
rect 33547 11799 33639 11805
rect 33547 11765 33559 11799
rect 33627 11765 33639 11799
rect 33547 11759 33639 11765
rect 33470 11715 33537 11727
rect 33470 11539 33497 11715
rect 33531 11539 33537 11715
rect 33470 11527 33537 11539
rect 33470 11524 33514 11527
rect 33574 11495 33614 11759
rect 33672 11727 33742 11728
rect 33649 11722 33742 11727
rect 33649 11715 33678 11722
rect 33649 11539 33655 11715
rect 33649 11536 33678 11539
rect 33736 11536 33742 11722
rect 33649 11530 33742 11536
rect 33649 11528 33716 11530
rect 33649 11527 33695 11528
rect 33547 11489 33639 11495
rect 33547 11455 33559 11489
rect 33627 11455 33639 11489
rect 33547 11449 33639 11455
rect 33574 11326 33614 11449
rect 33782 11406 33789 11848
rect 33823 11406 33840 11848
rect 34014 11805 34054 11806
rect 33987 11799 34079 11805
rect 33987 11765 33999 11799
rect 34067 11765 34079 11799
rect 33987 11759 34079 11765
rect 33931 11726 33977 11727
rect 33884 11720 33977 11726
rect 33884 11534 33890 11720
rect 33948 11715 33977 11720
rect 33971 11539 33977 11715
rect 33948 11534 33977 11539
rect 33884 11528 33977 11534
rect 33931 11527 33977 11528
rect 34014 11495 34054 11759
rect 34112 11727 34156 11886
rect 34089 11715 34156 11727
rect 34089 11539 34095 11715
rect 34129 11539 34156 11715
rect 34089 11527 34156 11539
rect 34484 11727 34530 11886
rect 34566 11800 34630 11805
rect 34724 11800 34788 11805
rect 34566 11799 34788 11800
rect 34566 11765 34578 11799
rect 34618 11765 34736 11799
rect 34776 11765 34788 11799
rect 34566 11760 34788 11765
rect 34566 11759 34630 11760
rect 34724 11759 34788 11760
rect 34484 11715 34542 11727
rect 34484 11539 34502 11715
rect 34536 11539 34542 11715
rect 34484 11528 34542 11539
rect 34496 11527 34542 11528
rect 34112 11524 34156 11527
rect 34578 11495 34618 11759
rect 34654 11715 34700 11727
rect 34654 11539 34660 11715
rect 34694 11539 34700 11715
rect 34654 11527 34700 11539
rect 33987 11489 34079 11495
rect 33987 11455 33999 11489
rect 34067 11455 34079 11489
rect 33987 11449 34079 11455
rect 34566 11489 34630 11495
rect 34566 11455 34578 11489
rect 34618 11455 34630 11489
rect 34566 11449 34630 11455
rect 33782 11394 33840 11406
rect 33464 11320 33614 11326
rect 33464 11262 33470 11320
rect 33608 11262 33614 11320
rect 33464 11256 33614 11262
rect 34014 11198 34054 11449
rect 34578 11448 34618 11449
rect 34660 11418 34694 11527
rect 34736 11495 34776 11759
rect 34816 11727 34854 11886
rect 35104 11848 35156 11886
rect 34882 11799 34946 11805
rect 34882 11765 34894 11799
rect 34934 11765 34946 11799
rect 34882 11759 34946 11765
rect 34812 11715 34858 11727
rect 34812 11539 34818 11715
rect 34852 11539 34858 11715
rect 34812 11527 34858 11539
rect 34894 11495 34934 11759
rect 34970 11722 35070 11728
rect 34970 11532 34976 11722
rect 35064 11532 35070 11722
rect 34970 11526 35070 11532
rect 34724 11494 34788 11495
rect 34882 11494 34946 11495
rect 34724 11489 34946 11494
rect 34724 11455 34736 11489
rect 34776 11455 34894 11489
rect 34934 11455 34946 11489
rect 34724 11450 34946 11455
rect 34724 11449 34788 11450
rect 34882 11449 34946 11450
rect 34548 11416 34694 11418
rect 34548 11364 34554 11416
rect 34688 11364 34694 11416
rect 34548 11362 34694 11364
rect 34736 11280 34776 11449
rect 34894 11432 34934 11449
rect 34994 11326 35038 11526
rect 35104 11406 35110 11848
rect 35144 11406 35156 11848
rect 35230 11727 35274 11886
rect 35334 11805 35374 11806
rect 35321 11799 35385 11805
rect 35321 11765 35333 11799
rect 35373 11765 35385 11799
rect 35321 11759 35385 11765
rect 35230 11715 35297 11727
rect 35230 11539 35257 11715
rect 35291 11539 35297 11715
rect 35230 11527 35297 11539
rect 35230 11524 35274 11527
rect 35334 11495 35374 11759
rect 35434 11727 35478 11728
rect 35409 11715 35478 11727
rect 35409 11539 35415 11715
rect 35449 11539 35478 11715
rect 35409 11527 35478 11539
rect 35321 11489 35385 11495
rect 35321 11455 35333 11489
rect 35373 11455 35385 11489
rect 35321 11449 35385 11455
rect 35104 11394 35156 11406
rect 34994 11320 35144 11326
rect 33234 11138 34054 11198
rect 34560 11270 34780 11280
rect 34560 11190 34570 11270
rect 34770 11190 34780 11270
rect 34560 11180 34780 11190
rect 34994 11262 35000 11320
rect 35138 11262 35144 11320
rect 34994 11256 35144 11262
rect 34994 11198 35038 11256
rect 35334 11198 35374 11449
rect 33122 10988 33186 10994
rect 33122 10954 33134 10988
rect 33174 10954 33186 10988
rect 33122 10948 33186 10954
rect 33052 10906 33098 10907
rect 32930 10628 32976 10669
rect 31890 10507 31958 10519
rect 31362 10460 31426 10466
rect 31362 10426 31374 10460
rect 31414 10426 31426 10460
rect 31362 10420 31426 10426
rect 31590 10460 31866 10466
rect 31590 10426 31814 10460
rect 31854 10426 31866 10460
rect 31590 10420 31866 10426
rect 31914 10346 31958 10507
rect 32232 10622 32976 10628
rect 32232 10588 32313 10622
rect 32867 10594 32976 10622
rect 33032 10895 33098 10906
rect 32867 10588 32948 10594
rect 32232 10346 32948 10588
rect 33032 10519 33058 10895
rect 33092 10519 33098 10895
rect 33032 10507 33098 10519
rect 33032 10346 33076 10507
rect 33134 10466 33174 10948
rect 33234 10907 33278 11138
rect 33574 10994 33614 11006
rect 34014 10994 34054 11006
rect 34736 10994 34776 11180
rect 34994 11138 35374 11198
rect 33562 10988 33838 10994
rect 33562 10954 33574 10988
rect 33614 10954 33838 10988
rect 33562 10948 33838 10954
rect 34002 10988 34066 10994
rect 34002 10954 34014 10988
rect 34054 10954 34066 10988
rect 34002 10948 34066 10954
rect 34668 10988 34912 10994
rect 34668 10954 34680 10988
rect 34900 10954 34912 10988
rect 33210 10895 33278 10907
rect 33492 10906 33538 10907
rect 33210 10519 33216 10895
rect 33250 10519 33278 10895
rect 33210 10508 33278 10519
rect 33470 10895 33538 10906
rect 33470 10519 33498 10895
rect 33532 10519 33538 10895
rect 33210 10507 33256 10508
rect 33470 10507 33538 10519
rect 33122 10460 33186 10466
rect 33122 10426 33134 10460
rect 33174 10426 33186 10460
rect 33122 10420 33186 10426
rect 33470 10346 33514 10507
rect 33574 10466 33614 10948
rect 33650 10906 33696 10907
rect 33790 10906 33838 10948
rect 33932 10906 33978 10907
rect 33650 10900 33742 10906
rect 33650 10895 33678 10900
rect 33650 10519 33656 10895
rect 33736 10556 33742 10900
rect 33790 10900 33978 10906
rect 33790 10860 33890 10900
rect 33948 10895 33978 10900
rect 33650 10514 33678 10519
rect 33736 10514 33838 10556
rect 33650 10510 33838 10514
rect 33650 10508 33742 10510
rect 33650 10507 33696 10508
rect 33790 10466 33838 10510
rect 33884 10514 33890 10860
rect 33972 10519 33978 10895
rect 33948 10514 33978 10519
rect 33884 10508 33978 10514
rect 33932 10507 33978 10508
rect 34014 10466 34054 10948
rect 34090 10906 34136 10907
rect 34090 10895 34158 10906
rect 34090 10519 34096 10895
rect 34130 10519 34158 10895
rect 34538 10895 34584 10907
rect 34538 10819 34544 10895
rect 34578 10819 34584 10895
rect 34538 10628 34584 10819
rect 34668 10760 34912 10954
rect 35020 10907 35064 11138
rect 34996 10895 35064 10907
rect 34996 10819 35002 10895
rect 35036 10819 35064 10895
rect 34996 10808 35064 10819
rect 35130 11045 35176 11104
rect 34996 10807 35042 10808
rect 34668 10726 34680 10760
rect 34900 10726 34912 10760
rect 34668 10720 34912 10726
rect 35130 10669 35136 11045
rect 35170 10669 35176 11045
rect 35334 10994 35374 11138
rect 35434 11198 35478 11527
rect 35670 11727 35714 11886
rect 35982 11848 36040 11886
rect 35774 11805 35814 11806
rect 35747 11799 35839 11805
rect 35747 11765 35759 11799
rect 35827 11765 35839 11799
rect 35747 11759 35839 11765
rect 35670 11715 35737 11727
rect 35670 11539 35697 11715
rect 35731 11539 35737 11715
rect 35670 11527 35737 11539
rect 35670 11524 35714 11527
rect 35774 11495 35814 11759
rect 35872 11727 35942 11728
rect 35849 11722 35942 11727
rect 35849 11715 35878 11722
rect 35849 11539 35855 11715
rect 35849 11536 35878 11539
rect 35936 11536 35942 11722
rect 35849 11530 35942 11536
rect 35849 11528 35916 11530
rect 35849 11527 35895 11528
rect 35747 11489 35839 11495
rect 35747 11455 35759 11489
rect 35827 11455 35839 11489
rect 35747 11449 35839 11455
rect 35774 11326 35814 11449
rect 35982 11406 35989 11848
rect 36023 11406 36040 11848
rect 36214 11805 36254 11806
rect 36187 11799 36279 11805
rect 36187 11765 36199 11799
rect 36267 11765 36279 11799
rect 36187 11759 36279 11765
rect 36131 11726 36177 11727
rect 36084 11720 36177 11726
rect 36084 11534 36090 11720
rect 36148 11715 36177 11720
rect 36171 11539 36177 11715
rect 36148 11534 36177 11539
rect 36084 11528 36177 11534
rect 36131 11527 36177 11528
rect 36214 11495 36254 11759
rect 36312 11727 36356 11886
rect 36289 11715 36356 11727
rect 36289 11539 36295 11715
rect 36329 11539 36356 11715
rect 36289 11527 36356 11539
rect 36312 11524 36356 11527
rect 36470 11510 36480 11886
rect 36810 11510 36820 11980
rect 36470 11500 36820 11510
rect 36187 11489 36279 11495
rect 36187 11455 36199 11489
rect 36267 11455 36279 11489
rect 36187 11449 36279 11455
rect 35982 11394 36040 11406
rect 35664 11320 35814 11326
rect 35664 11262 35670 11320
rect 35808 11262 35814 11320
rect 35664 11256 35814 11262
rect 36214 11198 36254 11449
rect 35434 11138 36254 11198
rect 35322 10988 35386 10994
rect 35322 10954 35334 10988
rect 35374 10954 35386 10988
rect 35322 10948 35386 10954
rect 35252 10906 35298 10907
rect 35130 10628 35176 10669
rect 34090 10507 34158 10519
rect 33562 10460 33626 10466
rect 33562 10426 33574 10460
rect 33614 10426 33626 10460
rect 33562 10420 33626 10426
rect 33790 10460 34066 10466
rect 33790 10426 34014 10460
rect 34054 10426 34066 10460
rect 33790 10420 34066 10426
rect 34114 10346 34158 10507
rect 34432 10622 35176 10628
rect 34432 10588 34513 10622
rect 35067 10594 35176 10622
rect 35232 10895 35298 10906
rect 35067 10588 35148 10594
rect 34432 10346 35148 10588
rect 35232 10519 35258 10895
rect 35292 10519 35298 10895
rect 35232 10507 35298 10519
rect 35232 10346 35276 10507
rect 35334 10466 35374 10948
rect 35434 10907 35478 11138
rect 35774 10994 35814 11006
rect 36214 10994 36254 11006
rect 35762 10988 36038 10994
rect 35762 10954 35774 10988
rect 35814 10954 36038 10988
rect 35762 10948 36038 10954
rect 36202 10988 36266 10994
rect 36202 10954 36214 10988
rect 36254 10954 36266 10988
rect 36202 10948 36266 10954
rect 35410 10895 35478 10907
rect 35692 10906 35738 10907
rect 35410 10519 35416 10895
rect 35450 10519 35478 10895
rect 35410 10508 35478 10519
rect 35670 10895 35738 10906
rect 35670 10519 35698 10895
rect 35732 10519 35738 10895
rect 35410 10507 35456 10508
rect 35670 10507 35738 10519
rect 35322 10460 35386 10466
rect 35322 10426 35334 10460
rect 35374 10426 35386 10460
rect 35322 10420 35386 10426
rect 35670 10346 35714 10507
rect 35774 10466 35814 10948
rect 35850 10906 35896 10907
rect 35990 10906 36038 10948
rect 36132 10906 36178 10907
rect 35850 10900 35942 10906
rect 35850 10895 35878 10900
rect 35850 10519 35856 10895
rect 35936 10556 35942 10900
rect 35990 10900 36178 10906
rect 35990 10860 36090 10900
rect 36148 10895 36178 10900
rect 35850 10514 35878 10519
rect 35936 10514 36038 10556
rect 35850 10510 36038 10514
rect 35850 10508 35942 10510
rect 35850 10507 35896 10508
rect 35990 10466 36038 10510
rect 36084 10514 36090 10860
rect 36172 10519 36178 10895
rect 36148 10514 36178 10519
rect 36084 10508 36178 10514
rect 36132 10507 36178 10508
rect 36214 10466 36254 10948
rect 36290 10906 36336 10907
rect 36290 10895 36358 10906
rect 36290 10519 36296 10895
rect 36330 10519 36358 10895
rect 36290 10507 36358 10519
rect 35762 10460 35826 10466
rect 35762 10426 35774 10460
rect 35814 10426 35826 10460
rect 35762 10420 35826 10426
rect 35990 10460 36266 10466
rect 35990 10426 36214 10460
rect 36254 10426 36266 10460
rect 35990 10420 36266 10426
rect 36314 10346 36358 10507
rect 30032 10330 32112 10346
rect 32232 10330 34312 10346
rect 34432 10330 36512 10346
rect 28767 10283 28820 10295
rect 27440 10260 28726 10266
rect 27440 10226 27938 10260
rect 28714 10226 28726 10260
rect 27440 10220 28726 10226
rect 27440 10200 27450 10220
rect 28770 10203 28820 10283
rect 27370 10190 27450 10200
rect 28767 10191 28820 10203
rect 29930 10322 36512 10330
rect 29930 10288 30758 10322
rect 31150 10288 31198 10322
rect 31590 10288 31638 10322
rect 32030 10288 32958 10322
rect 33350 10288 33398 10322
rect 33790 10288 33838 10322
rect 34230 10288 35158 10322
rect 35550 10288 35598 10322
rect 35990 10288 36038 10322
rect 36430 10288 36512 10322
rect 29930 10246 36512 10288
rect 27730 10130 27810 10140
rect 27730 10108 27740 10130
rect 27260 10062 27740 10108
rect 27730 10040 27740 10062
rect 27800 10108 27810 10130
rect 28767 10137 28773 10191
rect 28807 10137 28820 10191
rect 28767 10125 28820 10137
rect 28770 10120 28820 10125
rect 29130 10190 29210 10200
rect 29930 10190 36510 10246
rect 29130 10120 29140 10190
rect 27800 10102 28726 10108
rect 27800 10068 27938 10102
rect 28714 10068 28726 10102
rect 27800 10062 28726 10068
rect 27800 10040 27810 10062
rect 28770 10045 29140 10120
rect 27730 10030 27810 10040
rect 28767 10040 29140 10045
rect 28767 10033 28820 10040
rect 27370 9975 27450 9985
rect 27370 9950 27380 9975
rect 27260 9904 27380 9950
rect 27370 9885 27380 9904
rect 27440 9950 27450 9975
rect 28767 9979 28773 10033
rect 28807 9979 28820 10033
rect 28767 9967 28820 9979
rect 27440 9944 28726 9950
rect 27440 9910 27938 9944
rect 28714 9910 28726 9944
rect 27440 9904 28726 9910
rect 27440 9885 27450 9904
rect 28770 9887 28820 9967
rect 29130 9970 29140 10040
rect 29200 9970 29210 10190
rect 29130 9960 29210 9970
rect 29560 10020 36510 10190
rect 27370 9875 27450 9885
rect 28767 9875 28820 9887
rect 27730 9815 27810 9825
rect 27730 9792 27740 9815
rect 27260 9746 27740 9792
rect 27730 9725 27740 9746
rect 27800 9792 27810 9815
rect 28767 9821 28773 9875
rect 28807 9821 28820 9875
rect 28767 9810 28820 9821
rect 29560 9816 31680 10020
rect 28767 9809 28813 9810
rect 29560 9800 29827 9816
rect 27800 9786 28726 9792
rect 27800 9752 27938 9786
rect 28714 9752 28726 9786
rect 27800 9746 28726 9752
rect 27800 9725 27810 9746
rect 27730 9715 27810 9725
rect 27910 9652 28814 9658
rect 27910 9618 27922 9652
rect 28802 9618 28814 9652
rect 27910 9612 28814 9618
rect 29560 9597 29750 9800
rect 29815 9782 29827 9800
rect 31387 9800 31680 9816
rect 31387 9782 31399 9800
rect 29815 9776 31399 9782
rect 29782 9678 30574 9684
rect 29782 9644 29794 9678
rect 30562 9644 30574 9678
rect 29782 9638 30574 9644
rect 30640 9678 31432 9684
rect 30640 9644 30652 9678
rect 31420 9644 31432 9678
rect 30640 9638 31432 9644
rect 29560 9585 29772 9597
rect 29560 9551 29732 9585
rect 27910 9512 28814 9518
rect 27910 9478 27922 9512
rect 28802 9478 28814 9512
rect 27910 9472 28814 9478
rect 27250 9405 27330 9415
rect 27250 9315 27260 9405
rect 27320 9384 27330 9405
rect 27320 9378 28726 9384
rect 27320 9344 27938 9378
rect 28714 9344 28726 9378
rect 27320 9338 28726 9344
rect 27320 9315 27330 9338
rect 27250 9305 27330 9315
rect 28767 9309 28813 9321
rect 27490 9250 27570 9260
rect 27490 9226 27500 9250
rect 27260 9180 27500 9226
rect 27490 9160 27500 9180
rect 27560 9226 27570 9250
rect 28767 9255 28773 9309
rect 28807 9255 28813 9309
rect 28767 9243 28813 9255
rect 29560 9243 29598 9551
rect 29632 9243 29732 9551
rect 27560 9220 28726 9226
rect 27560 9186 27938 9220
rect 28714 9186 28726 9220
rect 27560 9180 28726 9186
rect 27560 9160 27570 9180
rect 28770 9163 28810 9243
rect 29560 9220 29732 9243
rect 29726 9209 29732 9220
rect 29766 9209 29772 9585
rect 29726 9197 29772 9209
rect 27490 9150 27570 9160
rect 28767 9151 28813 9163
rect 27250 9090 27330 9100
rect 27250 9000 27260 9090
rect 27320 9068 27330 9090
rect 28767 9097 28773 9151
rect 28807 9100 28813 9151
rect 28870 9160 28950 9170
rect 28870 9100 28880 9160
rect 28807 9097 28880 9100
rect 28767 9085 28880 9097
rect 27320 9062 28726 9068
rect 27320 9028 27938 9062
rect 28714 9028 28726 9062
rect 27320 9022 28726 9028
rect 27320 9000 27330 9022
rect 28770 9005 28880 9085
rect 27250 8990 27330 9000
rect 28767 9000 28880 9005
rect 28767 8993 28813 9000
rect 27490 8935 27570 8945
rect 27490 8910 27500 8935
rect 27260 8864 27500 8910
rect 27490 8845 27500 8864
rect 27560 8910 27570 8935
rect 28767 8939 28773 8993
rect 28807 8939 28813 8993
rect 28767 8927 28813 8939
rect 28870 8940 28880 9000
rect 28940 8940 28950 9160
rect 30120 9156 30230 9638
rect 30560 9585 30650 9600
rect 30560 9209 30590 9585
rect 30624 9209 30650 9585
rect 30560 9156 30650 9209
rect 30970 9156 31080 9638
rect 31460 9597 31680 9800
rect 31442 9585 31680 9597
rect 31442 9209 31448 9585
rect 31482 9551 31680 9585
rect 31482 9410 31582 9551
rect 31616 9410 31680 9551
rect 31670 9220 31680 9410
rect 31482 9210 31680 9220
rect 31482 9209 31488 9210
rect 31442 9197 31488 9209
rect 29782 9150 31432 9156
rect 29520 9116 29794 9150
rect 30562 9116 30652 9150
rect 31420 9120 32210 9150
rect 31420 9116 32070 9120
rect 29520 9070 32070 9116
rect 29815 9012 31399 9018
rect 29815 9010 29827 9012
rect 28870 8930 28950 8940
rect 29590 8978 29827 9010
rect 31387 9010 31399 9012
rect 31387 8990 31750 9010
rect 31387 8978 31450 8990
rect 27560 8904 28726 8910
rect 27560 8870 27938 8904
rect 28714 8870 28726 8904
rect 27560 8864 28726 8870
rect 27560 8845 27570 8864
rect 28770 8847 28810 8927
rect 27490 8835 27570 8845
rect 28767 8835 28813 8847
rect 27250 8775 27330 8785
rect 27250 8685 27260 8775
rect 27320 8752 27330 8775
rect 28767 8781 28773 8835
rect 28807 8781 28813 8835
rect 28767 8769 28813 8781
rect 29590 8812 31450 8978
rect 29590 8790 29827 8812
rect 27320 8746 28726 8752
rect 27320 8712 27938 8746
rect 28714 8712 28726 8746
rect 27320 8706 28726 8712
rect 27320 8685 27330 8706
rect 27250 8675 27330 8685
rect 29590 8637 29740 8790
rect 29815 8778 29827 8790
rect 31387 8780 31450 8812
rect 31680 8780 31750 8990
rect 32060 8990 32070 9070
rect 32200 8990 32210 9120
rect 32810 9042 35710 9300
rect 32810 9020 32830 9042
rect 32818 9008 32830 9020
rect 33540 9020 33670 9042
rect 33540 9008 33552 9020
rect 32818 9002 33552 9008
rect 33658 9008 33670 9020
rect 34380 9030 35710 9042
rect 34380 9020 37110 9030
rect 34380 9008 34392 9020
rect 33658 9002 34392 9008
rect 32060 8980 32210 8990
rect 31387 8778 31750 8780
rect 29815 8772 31750 8778
rect 31380 8770 31750 8772
rect 32904 8940 33118 8946
rect 32904 8906 33006 8940
rect 33106 8906 33120 8940
rect 32904 8900 33120 8906
rect 32904 8847 32950 8900
rect 27910 8612 28814 8618
rect 27910 8578 27922 8612
rect 28802 8578 28814 8612
rect 27910 8572 28814 8578
rect 27910 8472 28814 8478
rect 27910 8438 27922 8472
rect 28802 8438 28814 8472
rect 27910 8432 28814 8438
rect 27250 8370 27330 8380
rect 27250 8280 27260 8370
rect 27320 8344 27330 8370
rect 27320 8338 28726 8344
rect 27320 8304 27938 8338
rect 28714 8304 28726 8338
rect 27320 8298 28726 8304
rect 27320 8280 27330 8298
rect 27250 8270 27330 8280
rect 28767 8269 28813 8281
rect 27610 8210 27690 8220
rect 27610 8186 27620 8210
rect 27260 8140 27620 8186
rect 27610 8120 27620 8140
rect 27680 8186 27690 8210
rect 28767 8215 28773 8269
rect 28807 8215 28813 8269
rect 28767 8203 28813 8215
rect 27680 8180 28726 8186
rect 27680 8146 27938 8180
rect 28714 8146 28726 8180
rect 27680 8140 28726 8146
rect 27680 8120 27690 8140
rect 28770 8123 28810 8203
rect 27610 8110 27690 8120
rect 28767 8111 28813 8123
rect 27250 8050 27330 8060
rect 27250 7960 27260 8050
rect 27320 8028 27330 8050
rect 28767 8057 28773 8111
rect 28807 8057 28813 8111
rect 28767 8050 28813 8057
rect 29000 8110 29080 8120
rect 29000 8050 29010 8110
rect 28767 8045 29010 8050
rect 27320 8022 28726 8028
rect 27320 7988 27938 8022
rect 28714 7988 28726 8022
rect 27320 7982 28726 7988
rect 27320 7960 27330 7982
rect 28770 7965 29010 8045
rect 27250 7950 27330 7960
rect 28767 7960 29010 7965
rect 28767 7953 28813 7960
rect 27610 7890 27690 7900
rect 27610 7870 27620 7890
rect 27260 7824 27620 7870
rect 27610 7800 27620 7824
rect 27680 7870 27690 7890
rect 28767 7899 28773 7953
rect 28807 7899 28813 7953
rect 28767 7887 28813 7899
rect 29000 7890 29010 7960
rect 29070 7890 29080 8110
rect 27680 7864 28726 7870
rect 27680 7830 27938 7864
rect 28714 7830 28726 7864
rect 27680 7824 28726 7830
rect 27680 7800 27690 7824
rect 28770 7807 28810 7887
rect 29000 7880 29080 7890
rect 27610 7790 27690 7800
rect 28767 7795 28813 7807
rect 27250 7740 27330 7750
rect 27250 7650 27260 7740
rect 27320 7712 27330 7740
rect 28767 7741 28773 7795
rect 28807 7741 28813 7795
rect 28767 7729 28813 7741
rect 27320 7706 28726 7712
rect 27320 7672 27938 7706
rect 28714 7672 28726 7706
rect 27320 7666 28726 7672
rect 27320 7650 27330 7666
rect 27250 7640 27330 7650
rect 27910 7572 28814 7578
rect 27910 7538 27922 7572
rect 28802 7538 28814 7572
rect 27910 7532 28814 7538
rect 29590 7513 29598 8637
rect 29632 8593 29740 8637
rect 29782 8674 30574 8680
rect 29782 8640 29794 8674
rect 30562 8640 30574 8674
rect 29782 8634 30574 8640
rect 30640 8674 31432 8680
rect 30640 8640 30652 8674
rect 31420 8640 31432 8674
rect 30640 8634 31432 8640
rect 31480 8637 31630 8770
rect 29632 8581 29772 8593
rect 29632 8205 29732 8581
rect 29766 8205 29772 8581
rect 29632 8193 29772 8205
rect 29632 7957 29740 8193
rect 30080 8152 30280 8634
rect 30584 8590 30630 8593
rect 30560 8581 30650 8590
rect 30560 8580 30590 8581
rect 30624 8580 30650 8581
rect 30560 8210 30570 8580
rect 30640 8210 30650 8580
rect 30560 8205 30590 8210
rect 30624 8205 30650 8210
rect 30560 8200 30650 8205
rect 30584 8193 30630 8200
rect 30900 8152 31100 8634
rect 31480 8593 31582 8637
rect 31442 8581 31582 8593
rect 31442 8205 31448 8581
rect 31482 8205 31582 8581
rect 31442 8193 31582 8205
rect 29782 8146 30574 8152
rect 29782 8112 29794 8146
rect 30562 8130 30574 8146
rect 30640 8146 31432 8152
rect 30640 8130 30652 8146
rect 30562 8112 30652 8130
rect 31420 8112 31432 8146
rect 29782 8106 30890 8112
rect 29800 8044 30890 8106
rect 29782 8038 30890 8044
rect 31280 8106 31432 8112
rect 31280 8044 31420 8106
rect 31280 8038 31432 8044
rect 29782 8004 29794 8038
rect 30562 8020 30652 8038
rect 30562 8004 30574 8020
rect 29782 7998 30574 8004
rect 30640 8004 30652 8020
rect 31420 8004 31432 8038
rect 30640 7998 31432 8004
rect 29632 7945 29772 7957
rect 29632 7569 29732 7945
rect 29766 7569 29772 7945
rect 29632 7557 29772 7569
rect 29632 7513 29740 7557
rect 30080 7516 30280 7998
rect 30584 7950 30630 7957
rect 30560 7945 30650 7950
rect 30560 7940 30590 7945
rect 30624 7940 30650 7945
rect 30560 7570 30570 7940
rect 30640 7570 30650 7940
rect 30560 7569 30590 7570
rect 30624 7569 30650 7570
rect 30560 7560 30650 7569
rect 30584 7557 30630 7560
rect 30900 7516 31100 7998
rect 31480 7957 31582 8193
rect 31442 7945 31582 7957
rect 31442 7569 31448 7945
rect 31482 7569 31582 7945
rect 31442 7557 31582 7569
rect 29590 7510 29740 7513
rect 29782 7510 30574 7516
rect 29592 7501 29638 7510
rect 29782 7476 29794 7510
rect 30562 7476 30574 7510
rect 29782 7470 30574 7476
rect 30640 7510 31432 7516
rect 30640 7476 30652 7510
rect 31420 7476 31432 7510
rect 30640 7470 31432 7476
rect 31480 7513 31582 7557
rect 31616 7513 31630 8637
rect 32904 8071 32910 8847
rect 32944 8071 32950 8847
rect 32904 8018 32950 8071
rect 33000 8018 33120 8900
rect 33170 8859 33200 9002
rect 33252 8940 33466 8946
rect 33252 8906 33264 8940
rect 33364 8906 33466 8940
rect 33252 8900 33466 8906
rect 33834 8940 33958 8946
rect 33834 8906 33846 8940
rect 33946 8906 33958 8940
rect 33834 8900 33958 8906
rect 33162 8847 33208 8859
rect 33162 8071 33168 8847
rect 33202 8071 33208 8847
rect 33162 8059 33208 8071
rect 33260 8018 33380 8900
rect 33420 8847 33466 8900
rect 33420 8071 33426 8847
rect 33460 8071 33466 8847
rect 33744 8847 33790 8859
rect 33744 8840 33750 8847
rect 33420 8018 33466 8071
rect 33660 8830 33750 8840
rect 33660 8030 33670 8830
rect 33784 8071 33790 8847
rect 33770 8059 33790 8071
rect 33770 8030 33780 8059
rect 33660 8020 33780 8030
rect 33860 8018 33920 8900
rect 34010 8859 34040 9002
rect 34092 8940 34216 8946
rect 34092 8906 34104 8940
rect 34204 8906 34216 8940
rect 34092 8900 34216 8906
rect 34450 8940 37110 9020
rect 34002 8847 34048 8859
rect 34002 8071 34008 8847
rect 34042 8071 34048 8847
rect 34002 8059 34048 8071
rect 34120 8018 34180 8900
rect 34450 8880 34500 8940
rect 35520 8880 37110 8940
rect 34260 8847 34306 8859
rect 34260 8071 34266 8847
rect 34300 8840 34306 8847
rect 34300 8730 34340 8840
rect 34450 8822 37110 8880
rect 34450 8800 34510 8822
rect 34498 8788 34510 8800
rect 34792 8800 34930 8822
rect 34792 8788 34804 8800
rect 34498 8782 34804 8788
rect 34918 8788 34930 8800
rect 35212 8800 35350 8822
rect 35212 8788 35224 8800
rect 34918 8782 35224 8788
rect 35338 8788 35350 8800
rect 35632 8800 37110 8822
rect 35632 8788 35644 8800
rect 35338 8782 35644 8788
rect 34300 8726 34670 8730
rect 34300 8720 34680 8726
rect 34300 8686 34634 8720
rect 34668 8686 34680 8720
rect 34300 8680 34680 8686
rect 34710 8720 35100 8730
rect 34710 8686 35054 8720
rect 35088 8686 35100 8720
rect 34710 8680 35100 8686
rect 35130 8720 35520 8730
rect 35130 8686 35474 8720
rect 35508 8686 35520 8720
rect 35130 8680 35520 8686
rect 34300 8071 34340 8680
rect 34710 8639 34790 8680
rect 35130 8639 35210 8680
rect 34584 8627 34630 8639
rect 34584 8610 34590 8627
rect 34500 8600 34590 8610
rect 34500 8440 34510 8600
rect 34500 8430 34590 8440
rect 34584 8251 34590 8430
rect 34624 8251 34630 8627
rect 34584 8239 34630 8251
rect 34672 8627 34790 8639
rect 34672 8251 34678 8627
rect 34712 8620 34790 8627
rect 35004 8627 35050 8639
rect 34712 8251 34800 8620
rect 35004 8610 35010 8627
rect 34920 8600 35010 8610
rect 34920 8440 34930 8600
rect 34920 8430 35010 8440
rect 34672 8239 34800 8251
rect 35004 8251 35010 8430
rect 35044 8251 35050 8627
rect 35004 8239 35050 8251
rect 35092 8627 35210 8639
rect 35092 8251 35098 8627
rect 35132 8620 35210 8627
rect 35424 8627 35470 8639
rect 35424 8620 35430 8627
rect 35132 8251 35220 8620
rect 35340 8610 35430 8620
rect 35340 8450 35350 8610
rect 35340 8440 35430 8450
rect 35092 8239 35220 8251
rect 35424 8251 35430 8440
rect 35464 8251 35470 8627
rect 35424 8239 35470 8251
rect 35512 8627 35558 8639
rect 35512 8251 35518 8627
rect 35552 8620 35558 8627
rect 35552 8251 35640 8620
rect 35512 8239 35640 8251
rect 34680 8238 34800 8239
rect 35100 8238 35220 8239
rect 35520 8238 35640 8239
rect 34260 8059 34340 8071
rect 32904 8012 33120 8018
rect 32904 8000 33006 8012
rect 32900 7980 33006 8000
rect 32290 7978 33006 7980
rect 33106 8000 33120 8012
rect 33252 8012 33466 8018
rect 33252 8000 33264 8012
rect 33106 7978 33264 8000
rect 33364 7990 33466 8012
rect 33834 8012 33958 8018
rect 33834 7990 33846 8012
rect 33364 7978 33846 7990
rect 33946 7990 33958 8012
rect 34092 8012 34216 8018
rect 34092 7990 34104 8012
rect 33946 7978 34104 7990
rect 34204 7978 34216 8012
rect 32290 7972 34216 7978
rect 34280 8000 34340 8059
rect 34620 8192 34680 8200
rect 34620 8158 34634 8192
rect 34668 8158 34680 8192
rect 34280 7990 34370 8000
rect 32290 7970 34210 7972
rect 32290 7890 32300 7970
rect 32460 7890 34210 7970
rect 32290 7880 34210 7890
rect 34280 7790 34290 7990
rect 34360 7940 34370 7990
rect 34620 7940 34680 8158
rect 34360 7930 34680 7940
rect 34610 7850 34680 7930
rect 34360 7840 34680 7850
rect 34360 7790 34370 7840
rect 34280 7780 34370 7790
rect 32250 7770 32320 7780
rect 32250 7570 32260 7770
rect 32320 7660 32330 7680
rect 34280 7660 34340 7780
rect 32320 7570 34340 7660
rect 32250 7560 34340 7570
rect 31480 7460 31630 7513
rect 33470 7550 34340 7560
rect 33470 7438 33500 7550
rect 33536 7510 33600 7516
rect 33536 7476 33548 7510
rect 33588 7476 33600 7510
rect 33536 7470 33600 7476
rect 33694 7510 33758 7516
rect 33694 7476 33706 7510
rect 33746 7476 33758 7510
rect 33694 7470 33758 7476
rect 27910 7432 28814 7438
rect 27910 7398 27922 7432
rect 28802 7398 28814 7432
rect 27910 7392 28814 7398
rect 33466 7426 33512 7438
rect 27370 7330 27450 7340
rect 27370 7304 27380 7330
rect 27260 7258 27380 7304
rect 27370 7240 27380 7258
rect 27440 7304 27450 7330
rect 27440 7298 28726 7304
rect 27440 7264 27938 7298
rect 28714 7264 28726 7298
rect 27440 7258 28726 7264
rect 27440 7240 27450 7258
rect 27370 7230 27450 7240
rect 28767 7229 28813 7241
rect 27610 7170 27690 7180
rect 27610 7146 27620 7170
rect 27260 7100 27620 7146
rect 27610 7080 27620 7100
rect 27680 7146 27690 7170
rect 28767 7175 28773 7229
rect 28807 7175 28813 7229
rect 28767 7163 28813 7175
rect 27680 7140 28726 7146
rect 27680 7106 27938 7140
rect 28714 7106 28726 7140
rect 27680 7100 28726 7106
rect 27680 7080 27690 7100
rect 28770 7083 28810 7163
rect 29770 7150 31890 7160
rect 29532 7115 29578 7127
rect 27610 7070 27690 7080
rect 28767 7071 28813 7083
rect 27370 7015 27450 7025
rect 27370 6988 27380 7015
rect 27260 6942 27380 6988
rect 27370 6925 27380 6942
rect 27440 6988 27450 7015
rect 28767 7017 28773 7071
rect 28807 7020 28813 7071
rect 28870 7080 28950 7090
rect 28870 7020 28880 7080
rect 28807 7017 28880 7020
rect 28767 7005 28880 7017
rect 27440 6982 28726 6988
rect 27440 6948 27938 6982
rect 28714 6948 28726 6982
rect 27440 6942 28726 6948
rect 27440 6925 27450 6942
rect 28770 6925 28880 7005
rect 27370 6915 27450 6925
rect 28767 6913 28880 6925
rect 27610 6855 27690 6865
rect 27610 6830 27620 6855
rect 27260 6784 27620 6830
rect 27610 6765 27620 6784
rect 27680 6830 27690 6855
rect 28767 6859 28773 6913
rect 28807 6910 28880 6913
rect 28807 6859 28813 6910
rect 28767 6847 28813 6859
rect 28870 6860 28880 6910
rect 28940 6860 28950 7080
rect 28870 6850 28950 6860
rect 27680 6824 28726 6830
rect 27680 6790 27938 6824
rect 28714 6790 28726 6824
rect 27680 6784 28726 6790
rect 27680 6765 27690 6784
rect 28770 6767 28810 6847
rect 27610 6755 27690 6765
rect 28767 6755 28813 6767
rect 27370 6700 27450 6710
rect 27370 6672 27380 6700
rect 27260 6626 27380 6672
rect 27370 6610 27380 6626
rect 27440 6672 27450 6700
rect 28767 6701 28773 6755
rect 28807 6701 28813 6755
rect 29532 6721 29538 7115
rect 29572 6721 29578 7115
rect 29770 7070 30470 7150
rect 29757 7064 30470 7070
rect 30850 7070 31890 7150
rect 30850 7064 31897 7070
rect 29757 7030 29769 7064
rect 30850 7050 31109 7064
rect 30545 7040 31109 7050
rect 30545 7030 30557 7040
rect 29757 7024 30557 7030
rect 31097 7030 31109 7040
rect 31885 7030 31897 7064
rect 33466 7050 33472 7426
rect 33506 7050 33512 7426
rect 33466 7038 33512 7050
rect 31097 7024 31897 7030
rect 33550 7006 33590 7470
rect 33624 7426 33670 7438
rect 33624 7050 33630 7426
rect 33664 7050 33670 7426
rect 33624 7038 33670 7050
rect 33536 7000 33600 7006
rect 33450 6990 33548 7000
rect 33588 6990 33600 7000
rect 29670 6970 29716 6980
rect 30598 6970 30644 6980
rect 31010 6970 31056 6980
rect 31938 6970 31984 6980
rect 29670 6968 30790 6970
rect 29670 6868 29676 6968
rect 29710 6870 30604 6968
rect 29710 6868 29716 6870
rect 29670 6856 29716 6868
rect 30598 6868 30604 6870
rect 30638 6870 30790 6968
rect 30638 6868 30644 6870
rect 30598 6856 30644 6868
rect 29757 6806 30557 6812
rect 29757 6772 29769 6806
rect 30545 6772 30557 6806
rect 29757 6766 30557 6772
rect 29532 6709 29578 6721
rect 28767 6689 28813 6701
rect 29780 6680 30550 6766
rect 27440 6666 28726 6672
rect 27440 6632 27938 6666
rect 28714 6632 28726 6666
rect 27440 6626 28726 6632
rect 27440 6610 27450 6626
rect 27370 6600 27450 6610
rect 27910 6532 28814 6538
rect 27910 6498 27922 6532
rect 28802 6498 28814 6532
rect 27910 6492 28814 6498
rect 30090 6480 30210 6680
rect 30090 6470 30430 6480
rect 30090 6410 30120 6470
rect 30420 6410 30430 6470
rect 30090 6400 30430 6410
rect 27910 6392 28814 6398
rect 27910 6358 27922 6392
rect 28802 6358 28814 6392
rect 27910 6352 28814 6358
rect 30090 6330 30210 6400
rect 27370 6290 27450 6300
rect 27370 6264 27380 6290
rect 27260 6218 27380 6264
rect 27370 6200 27380 6218
rect 27440 6264 27450 6290
rect 27440 6258 28726 6264
rect 27440 6224 27938 6258
rect 28714 6224 28726 6258
rect 29770 6240 30680 6330
rect 27440 6218 28726 6224
rect 29758 6234 30680 6240
rect 27440 6200 27450 6218
rect 27370 6190 27450 6200
rect 28767 6189 28813 6201
rect 29758 6200 29770 6234
rect 30546 6200 30680 6234
rect 29758 6194 30680 6200
rect 27490 6130 27570 6140
rect 27490 6106 27500 6130
rect 27260 6060 27500 6106
rect 27490 6040 27500 6060
rect 27560 6106 27570 6130
rect 28767 6135 28773 6189
rect 28807 6135 28813 6189
rect 28767 6123 28813 6135
rect 29680 6155 29726 6167
rect 27560 6100 28726 6106
rect 27560 6066 27938 6100
rect 28714 6066 28726 6100
rect 27560 6060 28726 6066
rect 27560 6040 27570 6060
rect 28770 6043 28810 6123
rect 27490 6030 27570 6040
rect 28767 6031 28813 6043
rect 27370 5975 27450 5985
rect 27370 5948 27380 5975
rect 27260 5902 27380 5948
rect 27370 5885 27380 5902
rect 27440 5948 27450 5975
rect 28767 5977 28773 6031
rect 28807 5977 28813 6031
rect 28767 5970 28813 5977
rect 29000 6040 29080 6050
rect 29000 5970 29010 6040
rect 27440 5942 28726 5948
rect 27440 5908 27938 5942
rect 28714 5908 28726 5942
rect 27440 5902 28726 5908
rect 27440 5885 27450 5902
rect 27370 5875 27450 5885
rect 28760 5873 29010 5970
rect 28760 5860 28773 5873
rect 27490 5815 27570 5825
rect 27490 5790 27500 5815
rect 27260 5744 27500 5790
rect 27490 5725 27500 5744
rect 27560 5790 27570 5815
rect 28767 5819 28773 5860
rect 28807 5860 29010 5873
rect 28807 5819 28813 5860
rect 28767 5807 28813 5819
rect 29000 5820 29010 5860
rect 29070 5820 29080 6040
rect 29680 6021 29686 6155
rect 29720 6150 29726 6155
rect 30550 6155 30680 6194
rect 30550 6150 30596 6155
rect 29720 6030 30596 6150
rect 29720 6021 29726 6030
rect 29680 6009 29726 6021
rect 30590 6021 30596 6030
rect 30630 6021 30680 6155
rect 30590 6009 30680 6021
rect 29758 5976 30558 5982
rect 29758 5970 29770 5976
rect 29000 5810 29080 5820
rect 29630 5942 29770 5970
rect 30546 5942 30558 5976
rect 29630 5936 30558 5942
rect 29630 5820 30550 5936
rect 27560 5784 28726 5790
rect 27560 5750 27938 5784
rect 28714 5750 28726 5784
rect 27560 5744 28726 5750
rect 27560 5725 27570 5744
rect 28770 5727 28810 5807
rect 27490 5715 27570 5725
rect 28767 5715 28813 5727
rect 27370 5660 27450 5670
rect 27370 5632 27380 5660
rect 27260 5586 27380 5632
rect 27370 5570 27380 5586
rect 27440 5632 27450 5660
rect 28767 5661 28773 5715
rect 28807 5661 28813 5715
rect 28767 5649 28813 5661
rect 27440 5626 28726 5632
rect 27440 5592 27938 5626
rect 28714 5592 28726 5626
rect 27440 5586 28726 5592
rect 27440 5570 27450 5586
rect 27370 5560 27450 5570
rect 27910 5492 28814 5498
rect 27910 5458 27922 5492
rect 28802 5458 28814 5492
rect 27910 5452 28814 5458
rect 27909 5376 28807 5382
rect 27909 5342 27921 5376
rect 28795 5342 28807 5376
rect 27909 5336 28807 5342
rect 27170 5244 28750 5250
rect 27170 5240 28754 5244
rect 27170 5110 27180 5240
rect 27310 5238 28754 5240
rect 27310 5204 27974 5238
rect 28742 5204 28754 5238
rect 29630 5240 29800 5820
rect 30050 5730 30250 5740
rect 29880 5670 30060 5730
rect 30240 5670 30250 5730
rect 29880 5508 29940 5670
rect 30050 5660 30250 5670
rect 30600 5620 30680 6009
rect 29980 5586 30680 5620
rect 29972 5580 30680 5586
rect 29972 5546 29984 5580
rect 30352 5550 30680 5580
rect 30352 5546 30364 5550
rect 29972 5540 30364 5546
rect 29880 5496 29962 5508
rect 29880 5420 29922 5496
rect 29956 5420 29962 5496
rect 29916 5408 29962 5420
rect 30110 5376 30190 5540
rect 30400 5508 30460 5510
rect 30374 5496 30460 5508
rect 30374 5420 30380 5496
rect 30414 5420 30460 5496
rect 30374 5408 30460 5420
rect 29972 5370 30364 5376
rect 29972 5336 29984 5370
rect 30352 5336 30364 5370
rect 29972 5330 30364 5336
rect 30400 5240 30460 5408
rect 27310 5198 28754 5204
rect 28898 5225 28944 5237
rect 27310 5190 28750 5198
rect 27310 5157 27950 5190
rect 27310 5145 27952 5157
rect 27310 5110 27912 5145
rect 27170 5100 27912 5110
rect 27022 4830 27068 4842
rect 26366 4578 26928 4584
rect 7940 4560 9072 4576
rect 7940 4540 7950 4560
rect 7790 4530 7950 4540
rect 9060 4542 9072 4560
rect 10648 4560 11272 4576
rect 10648 4542 10660 4560
rect 9060 4536 10660 4542
rect 11260 4542 11272 4560
rect 12848 4542 12860 4576
rect 11260 4536 12860 4542
rect 8982 4487 9028 4499
rect 8982 4310 8988 4487
rect 8610 4250 8620 4310
rect 8680 4273 8988 4310
rect 9022 4273 9028 4487
rect 8680 4261 9028 4273
rect 10692 4487 10738 4499
rect 10692 4273 10698 4487
rect 10732 4420 10738 4487
rect 11182 4487 11228 4499
rect 10732 4360 10820 4420
rect 10880 4360 11110 4420
rect 10732 4273 10738 4360
rect 11182 4310 11188 4487
rect 10692 4261 10738 4273
rect 8680 4250 9026 4261
rect 10810 4250 11040 4310
rect 11100 4273 11188 4310
rect 11222 4273 11228 4487
rect 11100 4261 11228 4273
rect 12892 4487 12938 4499
rect 12892 4273 12898 4487
rect 12932 4420 12938 4487
rect 22496 4470 26802 4476
rect 22496 4436 22508 4470
rect 26790 4436 26802 4470
rect 22496 4430 26802 4436
rect 12932 4360 13240 4420
rect 13300 4360 13310 4420
rect 27880 4369 27912 5100
rect 27946 4369 27952 5145
rect 12932 4273 12938 4360
rect 12892 4261 12938 4273
rect 27880 4357 27952 4369
rect 28764 5150 28810 5157
rect 28898 5150 28904 5225
rect 28764 5145 28904 5150
rect 28764 4369 28770 5145
rect 28804 4369 28904 5145
rect 28764 4360 28904 4369
rect 28764 4357 28810 4360
rect 27880 4320 27950 4357
rect 27880 4316 28750 4320
rect 27880 4310 28754 4316
rect 27880 4276 27974 4310
rect 28742 4276 28754 4310
rect 28898 4289 28904 4360
rect 28938 4289 28944 5225
rect 29630 5170 30460 5240
rect 29630 5070 30040 5170
rect 30320 5070 30460 5170
rect 29980 4980 30460 5070
rect 29758 4974 30558 4980
rect 29758 4940 29770 4974
rect 30546 4940 30558 4974
rect 29758 4934 30558 4940
rect 30600 4907 30680 5550
rect 29680 4895 29726 4907
rect 29680 4761 29686 4895
rect 29720 4890 29726 4895
rect 30590 4895 30680 4907
rect 30590 4890 30596 4895
rect 29720 4770 30596 4890
rect 29720 4761 29726 4770
rect 29680 4749 29726 4761
rect 30590 4761 30596 4770
rect 30630 4770 30680 4895
rect 30630 4761 30636 4770
rect 30590 4749 30636 4761
rect 29758 4720 30558 4722
rect 29758 4716 30560 4720
rect 29758 4676 29770 4716
rect 30546 4710 30560 4716
rect 29760 4640 29770 4676
rect 30550 4640 30560 4710
rect 29760 4630 30560 4640
rect 30730 4610 30790 6870
rect 28898 4277 28944 4289
rect 30650 4530 30790 4610
rect 30860 6968 31984 6970
rect 30860 6870 31016 6968
rect 30860 4610 30920 6870
rect 31010 6868 31016 6870
rect 31050 6870 31944 6968
rect 31050 6868 31056 6870
rect 31010 6856 31056 6868
rect 31938 6868 31944 6870
rect 31978 6868 31984 6968
rect 33450 6930 33460 6990
rect 33590 6930 33600 6990
rect 33450 6920 33600 6930
rect 33630 6868 33660 7038
rect 33710 7006 33750 7470
rect 33790 7438 33820 7550
rect 33852 7510 33916 7516
rect 33852 7476 33864 7510
rect 33904 7476 33916 7510
rect 33852 7470 33916 7476
rect 34010 7510 34074 7516
rect 34010 7476 34022 7510
rect 34062 7476 34074 7510
rect 34010 7470 34074 7476
rect 33782 7426 33828 7438
rect 33782 7050 33788 7426
rect 33822 7050 33828 7426
rect 33782 7038 33828 7050
rect 33860 7006 33900 7470
rect 33940 7426 33986 7438
rect 33940 7050 33946 7426
rect 33980 7050 33986 7426
rect 33940 7038 33986 7050
rect 33694 7000 33758 7006
rect 33852 7000 33916 7006
rect 33690 6990 33706 7000
rect 33746 6990 33864 7000
rect 33904 6990 33920 7000
rect 33690 6930 33700 6990
rect 33910 6930 33920 6990
rect 33690 6920 33920 6930
rect 33950 6868 33980 7038
rect 34020 7006 34060 7470
rect 34110 7438 34140 7550
rect 34098 7426 34144 7438
rect 34098 7050 34104 7426
rect 34138 7050 34144 7426
rect 34280 7100 34340 7550
rect 34620 7402 34680 7840
rect 34620 7368 34634 7402
rect 34668 7368 34680 7402
rect 34620 7360 34680 7368
rect 34740 8190 34800 8238
rect 35040 8192 35100 8200
rect 34740 8180 34900 8190
rect 34740 7960 34750 8180
rect 34890 7960 34900 8180
rect 34740 7950 34900 7960
rect 35040 8158 35054 8192
rect 35088 8158 35100 8192
rect 34740 7620 34800 7950
rect 35040 7620 35100 8158
rect 34740 7560 35100 7620
rect 34740 7330 34800 7560
rect 35040 7402 35100 7560
rect 35040 7368 35054 7402
rect 35088 7368 35100 7402
rect 35040 7360 35100 7368
rect 35160 7990 35220 8238
rect 35460 8192 35520 8200
rect 35460 8158 35474 8192
rect 35508 8158 35520 8192
rect 35160 7980 35320 7990
rect 35160 7760 35170 7980
rect 35310 7760 35320 7980
rect 35160 7750 35320 7760
rect 35160 7620 35220 7750
rect 35460 7620 35520 8158
rect 35160 7560 35520 7620
rect 35160 7330 35220 7560
rect 35460 7402 35520 7560
rect 35460 7368 35474 7402
rect 35508 7368 35520 7402
rect 35460 7360 35520 7368
rect 35580 7680 35640 8238
rect 35580 7560 36610 7680
rect 35580 7330 35640 7560
rect 34584 7320 34630 7330
rect 34490 7318 34630 7320
rect 34490 7310 34590 7318
rect 34490 7150 34500 7310
rect 34490 7142 34590 7150
rect 34624 7142 34630 7318
rect 34490 7140 34630 7142
rect 34580 7130 34630 7140
rect 34672 7318 34800 7330
rect 35004 7320 35050 7330
rect 34672 7142 34678 7318
rect 34712 7142 34800 7318
rect 34672 7130 34800 7142
rect 34910 7318 35050 7320
rect 34910 7310 35010 7318
rect 34910 7150 34920 7310
rect 34910 7142 35010 7150
rect 35044 7142 35050 7318
rect 34910 7140 35050 7142
rect 35000 7130 35050 7140
rect 35092 7318 35220 7330
rect 35424 7320 35470 7330
rect 35092 7142 35098 7318
rect 35132 7142 35220 7318
rect 35092 7130 35220 7142
rect 35330 7318 35470 7320
rect 35330 7310 35430 7318
rect 35330 7150 35340 7310
rect 35330 7142 35430 7150
rect 35464 7142 35470 7318
rect 35330 7140 35470 7142
rect 35420 7130 35470 7140
rect 35512 7318 35640 7330
rect 35512 7142 35518 7318
rect 35552 7142 35640 7318
rect 35512 7140 35640 7142
rect 35512 7130 35558 7140
rect 34710 7100 34800 7130
rect 35130 7100 35220 7130
rect 34280 7092 34680 7100
rect 34280 7058 34634 7092
rect 34668 7058 34680 7092
rect 34280 7050 34680 7058
rect 34710 7092 35100 7100
rect 34710 7058 35054 7092
rect 35088 7058 35100 7092
rect 34710 7050 35100 7058
rect 35130 7092 35520 7100
rect 35130 7058 35474 7092
rect 35508 7058 35520 7092
rect 35130 7050 35520 7058
rect 34098 7038 34144 7050
rect 34010 7000 34074 7006
rect 34010 6990 34022 7000
rect 34062 6990 34200 7000
rect 34010 6930 34020 6990
rect 34190 6930 34200 6990
rect 34498 6990 34804 6996
rect 34498 6980 34510 6990
rect 34010 6920 34200 6930
rect 34480 6956 34510 6980
rect 34792 6980 34804 6990
rect 34918 6990 35224 6996
rect 34918 6980 34930 6990
rect 34792 6956 34930 6980
rect 35212 6980 35224 6990
rect 35338 6990 35644 6996
rect 35338 6980 35350 6990
rect 35212 6956 35350 6980
rect 35632 6980 35644 6990
rect 35632 6956 36700 6980
rect 34480 6920 36700 6956
rect 31938 6856 31984 6868
rect 33360 6862 34250 6868
rect 33360 6850 33372 6862
rect 33330 6828 33372 6850
rect 34238 6850 34250 6862
rect 34238 6846 34410 6850
rect 34480 6846 34500 6920
rect 34238 6830 34500 6846
rect 35540 6830 36700 6920
rect 34238 6828 36700 6830
rect 31097 6806 31897 6812
rect 31097 6772 31109 6806
rect 31885 6772 31897 6806
rect 31097 6766 31897 6772
rect 31110 6680 31870 6766
rect 33330 6748 36700 6828
rect 33330 6700 35660 6748
rect 31410 6330 31530 6680
rect 33334 6630 35660 6700
rect 33330 6614 35554 6630
rect 30970 6310 31880 6330
rect 30970 6250 31080 6310
rect 31380 6250 31880 6310
rect 30970 6240 31880 6250
rect 30970 6234 31898 6240
rect 30970 6200 31110 6234
rect 31886 6200 31898 6234
rect 30970 6194 31898 6200
rect 30970 6155 31110 6194
rect 30970 6021 31026 6155
rect 31060 6150 31110 6155
rect 31930 6155 31976 6167
rect 31930 6150 31936 6155
rect 31060 6030 31936 6150
rect 31060 6021 31066 6030
rect 30970 6009 31066 6021
rect 31930 6021 31936 6030
rect 31970 6021 31976 6155
rect 31930 6009 31976 6021
rect 30970 5620 31050 6009
rect 31098 5976 31898 5982
rect 31098 5942 31110 5976
rect 31886 5970 31898 5976
rect 33330 5970 33560 6614
rect 36220 6260 36420 6270
rect 36220 6200 36230 6260
rect 36060 6080 36230 6200
rect 36410 6080 36420 6260
rect 36060 6000 36420 6080
rect 36520 6260 36720 6270
rect 36520 6080 36530 6260
rect 36710 6220 36720 6260
rect 36710 6110 38010 6220
rect 36710 6080 36720 6110
rect 36520 6070 36720 6080
rect 37420 6006 38010 6110
rect 36448 6000 36848 6006
rect 36060 5970 36460 6000
rect 31886 5942 33650 5970
rect 31098 5936 33650 5942
rect 31110 5820 33650 5936
rect 31370 5740 31570 5750
rect 31370 5680 31380 5740
rect 31560 5680 31770 5740
rect 31370 5670 31570 5680
rect 30970 5586 31650 5620
rect 30970 5580 31674 5586
rect 30970 5550 31294 5580
rect 30970 4907 31050 5550
rect 31282 5546 31294 5550
rect 31662 5546 31674 5580
rect 31282 5540 31674 5546
rect 31140 5508 31250 5510
rect 31140 5496 31272 5508
rect 31140 5420 31232 5496
rect 31266 5420 31272 5496
rect 31140 5408 31272 5420
rect 31140 5220 31250 5408
rect 31440 5376 31520 5540
rect 31710 5508 31770 5680
rect 31684 5496 31770 5508
rect 31684 5420 31690 5496
rect 31724 5420 31770 5496
rect 31684 5408 31730 5420
rect 31282 5370 31674 5376
rect 31282 5336 31294 5370
rect 31662 5336 31674 5370
rect 31282 5330 31674 5336
rect 33350 5300 33560 5820
rect 36060 5480 36140 5970
rect 36448 5966 36460 5970
rect 36836 5966 36848 6000
rect 36448 5960 36848 5966
rect 37234 6000 38010 6006
rect 37234 5966 37246 6000
rect 37622 5970 38010 6000
rect 37622 5966 37634 5970
rect 37234 5960 37634 5966
rect 36370 5921 36416 5933
rect 36370 5900 36376 5921
rect 36290 5890 36376 5900
rect 36410 5920 36416 5921
rect 36880 5921 36926 5933
rect 36880 5920 36886 5921
rect 36290 5820 36300 5890
rect 36290 5810 36376 5820
rect 36370 5787 36376 5810
rect 36410 5790 36886 5920
rect 36410 5787 36416 5790
rect 36370 5775 36416 5787
rect 36880 5787 36886 5790
rect 36920 5787 36926 5921
rect 36880 5775 36926 5787
rect 36448 5742 36848 5748
rect 36448 5708 36460 5742
rect 36836 5740 36848 5742
rect 37000 5740 37080 5960
rect 37156 5921 37202 5933
rect 37156 5787 37162 5921
rect 37196 5920 37202 5921
rect 37666 5921 37712 5933
rect 37666 5920 37672 5921
rect 37196 5790 37672 5920
rect 37706 5900 37712 5921
rect 37706 5890 37780 5900
rect 37770 5820 37780 5890
rect 37196 5787 37202 5790
rect 37156 5775 37202 5787
rect 37666 5787 37672 5790
rect 37706 5810 37780 5820
rect 37706 5787 37712 5810
rect 37666 5775 37712 5787
rect 37234 5742 37634 5748
rect 37234 5740 37246 5742
rect 36836 5710 37246 5740
rect 36836 5708 36848 5710
rect 36448 5702 36848 5708
rect 36370 5663 36416 5675
rect 36370 5640 36376 5663
rect 36290 5630 36376 5640
rect 36410 5660 36416 5663
rect 36880 5663 36926 5675
rect 36880 5660 36886 5663
rect 36290 5560 36300 5630
rect 36290 5550 36376 5560
rect 36370 5529 36376 5550
rect 36410 5530 36886 5660
rect 36410 5529 36416 5530
rect 36370 5517 36416 5529
rect 36880 5529 36886 5530
rect 36920 5529 36926 5663
rect 36880 5517 36926 5529
rect 36448 5484 36848 5490
rect 36448 5480 36460 5484
rect 36060 5450 36460 5480
rect 36836 5450 36848 5484
rect 33320 5290 33640 5300
rect 33320 5220 33330 5290
rect 31140 5100 33330 5220
rect 31140 4980 31670 5100
rect 33320 5020 33330 5100
rect 33630 5020 33640 5290
rect 33320 5010 33640 5020
rect 31098 4974 31898 4980
rect 31098 4940 31110 4974
rect 31886 4940 31898 4974
rect 31098 4934 31898 4940
rect 36060 4970 36140 5450
rect 36448 5444 36848 5450
rect 36370 5405 36416 5417
rect 36370 5380 36376 5405
rect 36290 5370 36376 5380
rect 36410 5400 36416 5405
rect 36880 5405 36926 5417
rect 36880 5400 36886 5405
rect 36290 5300 36300 5370
rect 36290 5290 36376 5300
rect 36370 5271 36376 5290
rect 36410 5271 36886 5400
rect 36920 5271 36926 5405
rect 36370 5270 36926 5271
rect 36370 5259 36416 5270
rect 36880 5259 36926 5270
rect 36448 5226 36848 5232
rect 36448 5192 36460 5226
rect 36836 5220 36848 5226
rect 37000 5220 37080 5710
rect 37234 5708 37246 5710
rect 37622 5708 37634 5742
rect 37234 5702 37634 5708
rect 37156 5663 37202 5675
rect 37156 5529 37162 5663
rect 37196 5660 37202 5663
rect 37666 5663 37712 5675
rect 37666 5660 37672 5663
rect 37196 5530 37672 5660
rect 37706 5640 37712 5663
rect 37706 5630 37780 5640
rect 37770 5560 37780 5630
rect 37196 5529 37202 5530
rect 37156 5517 37202 5529
rect 37666 5529 37672 5530
rect 37706 5550 37780 5560
rect 37706 5529 37712 5550
rect 37666 5517 37712 5529
rect 37234 5484 37634 5490
rect 37234 5450 37246 5484
rect 37622 5480 37634 5484
rect 37930 5480 38010 5970
rect 37622 5450 38010 5480
rect 37234 5444 37634 5450
rect 37156 5405 37202 5417
rect 37156 5271 37162 5405
rect 37196 5400 37202 5405
rect 37666 5405 37712 5417
rect 37666 5400 37672 5405
rect 37196 5271 37672 5400
rect 37706 5380 37712 5405
rect 37706 5370 37780 5380
rect 37770 5300 37780 5370
rect 37706 5290 37780 5300
rect 37706 5271 37712 5290
rect 37156 5270 37712 5271
rect 37156 5259 37202 5270
rect 37666 5259 37712 5270
rect 37234 5226 37634 5232
rect 37234 5220 37246 5226
rect 36836 5192 37246 5220
rect 37622 5192 37634 5226
rect 36448 5190 37634 5192
rect 36448 5186 36848 5190
rect 36370 5147 36416 5159
rect 36370 5120 36376 5147
rect 36290 5110 36376 5120
rect 36410 5140 36416 5147
rect 36880 5147 36926 5159
rect 36880 5140 36886 5147
rect 36290 5040 36300 5110
rect 36290 5030 36376 5040
rect 36370 5013 36376 5030
rect 36410 5013 36886 5140
rect 36920 5013 36926 5147
rect 36370 5010 36926 5013
rect 36370 5001 36416 5010
rect 36880 5001 36926 5010
rect 36448 4970 36848 4974
rect 36060 4968 36850 4970
rect 36060 4940 36460 4968
rect 30970 4895 31066 4907
rect 30970 4770 31026 4895
rect 31020 4761 31026 4770
rect 31060 4890 31066 4895
rect 31930 4895 31976 4907
rect 31930 4890 31936 4895
rect 31060 4770 31936 4890
rect 31060 4761 31066 4770
rect 31020 4749 31066 4761
rect 31930 4761 31936 4770
rect 31970 4761 31976 4895
rect 31930 4749 31976 4761
rect 32250 4880 32330 4890
rect 31098 4716 31898 4722
rect 31098 4682 31110 4716
rect 31886 4700 31898 4716
rect 32250 4700 32260 4880
rect 31886 4682 32260 4700
rect 31098 4676 32260 4682
rect 31110 4650 32260 4676
rect 32320 4650 32330 4880
rect 31110 4640 32330 4650
rect 30860 4530 31000 4610
rect 27880 4270 28754 4276
rect 11100 4250 11226 4261
rect 27880 4260 28750 4270
rect 9060 4218 10660 4224
rect 9060 4184 9072 4218
rect 10648 4200 10660 4218
rect 11260 4218 12860 4224
rect 11260 4200 11272 4218
rect 10648 4184 11272 4200
rect 12848 4184 12860 4218
rect 9060 4178 12860 4184
rect 9080 4100 12840 4178
rect 27909 4172 28807 4178
rect 27909 4138 27921 4172
rect 28795 4138 28807 4172
rect 27909 4132 28807 4138
rect 10880 3960 10890 4100
rect 11030 3960 11040 4100
rect 10880 3950 11040 3960
rect 30070 4040 30270 4050
rect 30070 3860 30080 4040
rect 30260 4000 30270 4040
rect 30650 4000 30750 4530
rect 30260 3890 30750 4000
rect 30900 4000 31000 4530
rect 36060 4450 36140 4940
rect 36448 4934 36460 4940
rect 36836 4940 36850 4968
rect 36836 4934 36848 4940
rect 36448 4928 36848 4934
rect 36370 4890 36416 4901
rect 36880 4890 36926 4901
rect 36370 4889 36926 4890
rect 36370 4860 36376 4889
rect 36290 4850 36376 4860
rect 36290 4780 36300 4850
rect 36290 4770 36376 4780
rect 36370 4755 36376 4770
rect 36410 4760 36886 4889
rect 36410 4755 36416 4760
rect 36370 4743 36416 4755
rect 36880 4755 36886 4760
rect 36920 4755 36926 4889
rect 36880 4743 36926 4755
rect 36448 4710 36848 4716
rect 37000 4710 37080 5190
rect 37234 5186 37634 5190
rect 37156 5147 37202 5159
rect 37156 5013 37162 5147
rect 37196 5140 37202 5147
rect 37666 5147 37712 5159
rect 37666 5140 37672 5147
rect 37196 5013 37672 5140
rect 37706 5120 37712 5147
rect 37706 5110 37780 5120
rect 37770 5040 37780 5110
rect 37706 5030 37780 5040
rect 37706 5013 37712 5030
rect 37156 5010 37712 5013
rect 37156 5001 37202 5010
rect 37666 5001 37712 5010
rect 37234 4970 37634 4974
rect 37930 4970 38010 5450
rect 37234 4968 38010 4970
rect 37234 4934 37246 4968
rect 37622 4940 38010 4968
rect 37622 4934 37634 4940
rect 37234 4928 37634 4934
rect 37156 4890 37202 4901
rect 37666 4890 37712 4901
rect 37156 4889 37712 4890
rect 37156 4755 37162 4889
rect 37196 4760 37672 4889
rect 37706 4860 37712 4889
rect 37706 4850 37780 4860
rect 37770 4780 37780 4850
rect 37196 4755 37202 4760
rect 37156 4743 37202 4755
rect 37666 4755 37672 4760
rect 37706 4770 37780 4780
rect 37706 4755 37712 4770
rect 37666 4743 37712 4755
rect 37234 4710 37634 4716
rect 36448 4676 36460 4710
rect 36836 4680 37246 4710
rect 36836 4676 36848 4680
rect 36448 4670 36848 4676
rect 36370 4631 36416 4643
rect 36370 4600 36376 4631
rect 36290 4590 36376 4600
rect 36410 4630 36416 4631
rect 36880 4631 36926 4643
rect 36880 4630 36886 4631
rect 36290 4520 36300 4590
rect 36290 4510 36376 4520
rect 36370 4497 36376 4510
rect 36410 4500 36886 4630
rect 36410 4497 36416 4500
rect 36370 4485 36416 4497
rect 36880 4497 36886 4500
rect 36920 4497 36926 4631
rect 36880 4485 36926 4497
rect 36448 4452 36848 4458
rect 36448 4450 36460 4452
rect 36060 4420 36460 4450
rect 32240 4168 34160 4240
rect 32240 4134 32772 4168
rect 33970 4134 34160 4168
rect 32240 4128 34160 4134
rect 32240 4059 32760 4128
rect 31670 4040 31870 4050
rect 31670 4000 31680 4040
rect 30900 3890 31680 4000
rect 30260 3860 30270 3890
rect 30070 3850 30270 3860
rect 31670 3860 31680 3890
rect 31860 3860 31870 4040
rect 31670 3850 31870 3860
rect 32240 3457 32588 4059
rect 32622 3958 32760 4059
rect 32800 4070 32990 4080
rect 32800 4036 32810 4070
rect 32789 4030 32810 4036
rect 32980 4036 32990 4070
rect 32980 4030 33005 4036
rect 32789 3996 32801 4030
rect 32835 3996 32959 4010
rect 32993 3996 33005 4030
rect 32789 3990 33005 3996
rect 32622 3946 32762 3958
rect 32622 3570 32722 3946
rect 32756 3570 32762 3946
rect 32622 3558 32762 3570
rect 32622 3457 32760 3558
rect 32790 3526 32846 3990
rect 32874 3946 32920 3958
rect 32874 3570 32880 3946
rect 32914 3570 32920 3946
rect 32874 3558 32920 3570
rect 32789 3520 32847 3526
rect 32789 3486 32801 3520
rect 32835 3486 32847 3520
rect 32789 3480 32847 3486
rect 17150 3388 18160 3410
rect 17150 3360 17164 3388
rect 17152 3354 17164 3360
rect 17232 3360 17322 3388
rect 17232 3354 17244 3360
rect 17152 3348 17244 3354
rect 17310 3354 17322 3360
rect 17390 3360 17480 3388
rect 17390 3354 17402 3360
rect 17310 3348 17402 3354
rect 17468 3354 17480 3360
rect 17548 3360 17638 3388
rect 17548 3354 17560 3360
rect 17468 3348 17560 3354
rect 17626 3354 17638 3360
rect 17706 3360 18160 3388
rect 17706 3354 17718 3360
rect 17626 3348 17718 3354
rect 17096 3304 17142 3316
rect 7800 2500 7940 2900
rect 17096 2790 17102 3304
rect 16900 2780 17102 2790
rect 16900 2640 16910 2780
rect 16900 2630 17102 2640
rect 17096 2528 17102 2630
rect 17136 2528 17142 3304
rect 17096 2516 17142 2528
rect 17254 3304 17300 3316
rect 17254 2528 17260 3304
rect 17294 2528 17300 3304
rect 17412 3304 17458 3316
rect 17412 2790 17418 3304
rect 17370 2780 17418 2790
rect 17452 2790 17458 3304
rect 17570 3304 17616 3316
rect 17452 2780 17500 2790
rect 17370 2640 17380 2780
rect 17490 2640 17500 2780
rect 17370 2630 17418 2640
rect 17254 2516 17300 2528
rect 17412 2528 17418 2630
rect 17452 2630 17500 2640
rect 17452 2528 17458 2630
rect 17412 2516 17458 2528
rect 17570 2528 17576 3304
rect 17610 2528 17616 3304
rect 17570 2516 17616 2528
rect 17728 3304 17774 3316
rect 17728 2528 17734 3304
rect 17768 2790 17774 3304
rect 18110 3020 18160 3360
rect 32240 3280 32760 3457
rect 32880 3440 32914 3558
rect 32948 3526 33004 3990
rect 33038 3958 33072 4128
rect 33120 4070 33310 4080
rect 33120 4036 33130 4070
rect 33105 4030 33130 4036
rect 33300 4036 33310 4070
rect 33300 4030 33321 4036
rect 33105 3996 33117 4030
rect 33151 3996 33275 4010
rect 33309 3996 33321 4030
rect 33105 3990 33321 3996
rect 33032 3946 33078 3958
rect 33032 3570 33038 3946
rect 33072 3570 33078 3946
rect 33032 3558 33078 3570
rect 33106 3526 33162 3990
rect 33190 3946 33236 3958
rect 33190 3570 33196 3946
rect 33230 3570 33236 3946
rect 33190 3558 33236 3570
rect 32947 3520 33005 3526
rect 32947 3486 32959 3520
rect 32993 3486 33005 3520
rect 32947 3480 33005 3486
rect 33105 3520 33163 3526
rect 33105 3486 33117 3520
rect 33151 3486 33163 3520
rect 33105 3480 33163 3486
rect 33196 3440 33230 3558
rect 33264 3526 33320 3990
rect 33354 3958 33388 4128
rect 33430 4070 33620 4080
rect 33430 4036 33440 4070
rect 33421 4030 33440 4036
rect 33610 4036 33620 4070
rect 33610 4030 33637 4036
rect 33421 3996 33433 4030
rect 33467 3996 33591 4010
rect 33625 3996 33637 4030
rect 33421 3990 33637 3996
rect 33348 3946 33394 3958
rect 33348 3570 33354 3946
rect 33388 3570 33394 3946
rect 33348 3558 33394 3570
rect 33422 3526 33478 3990
rect 33506 3946 33552 3958
rect 33506 3570 33512 3946
rect 33546 3570 33552 3946
rect 33506 3558 33552 3570
rect 33263 3520 33321 3526
rect 33263 3486 33275 3520
rect 33309 3486 33321 3520
rect 33263 3480 33321 3486
rect 33421 3520 33479 3526
rect 33421 3486 33433 3520
rect 33467 3486 33479 3520
rect 33421 3480 33479 3486
rect 33512 3440 33546 3558
rect 33580 3526 33636 3990
rect 33670 3958 33704 4128
rect 33960 4120 34160 4128
rect 33750 4070 33940 4080
rect 33750 4036 33760 4070
rect 33737 4030 33760 4036
rect 33930 4036 33940 4070
rect 33990 4059 34160 4120
rect 33930 4030 33953 4036
rect 33737 3996 33749 4030
rect 33783 3996 33907 4010
rect 33941 3996 33953 4030
rect 33737 3990 33953 3996
rect 33664 3946 33710 3958
rect 33664 3570 33670 3946
rect 33704 3570 33710 3946
rect 33664 3558 33710 3570
rect 33738 3526 33794 3990
rect 33822 3946 33868 3958
rect 33822 3570 33828 3946
rect 33862 3570 33868 3946
rect 33822 3558 33868 3570
rect 33579 3520 33637 3526
rect 33579 3486 33591 3520
rect 33625 3486 33637 3520
rect 33579 3480 33637 3486
rect 33737 3520 33795 3526
rect 33737 3486 33749 3520
rect 33783 3486 33795 3520
rect 33737 3480 33795 3486
rect 33828 3440 33862 3558
rect 33896 3526 33952 3990
rect 33990 3958 34120 4059
rect 33980 3946 34120 3958
rect 33980 3570 33986 3946
rect 34020 3570 34120 3946
rect 33980 3558 34120 3570
rect 33895 3520 33953 3526
rect 33895 3486 33907 3520
rect 33941 3486 33953 3520
rect 33895 3480 33953 3486
rect 33990 3457 34120 3558
rect 34154 3560 34160 4059
rect 34740 4168 35740 4240
rect 34740 4140 34883 4168
rect 34740 4071 34800 4140
rect 34871 4134 34883 4140
rect 35449 4140 35740 4168
rect 35449 4134 35461 4140
rect 34871 4128 35461 4134
rect 34860 4090 35200 4100
rect 34740 4059 34818 4071
rect 34740 3560 34778 4059
rect 34154 3457 34778 3560
rect 34812 3958 34818 4059
rect 34860 4010 34870 4090
rect 35190 4010 35200 4090
rect 34860 4000 34991 4010
rect 34979 3996 34991 4000
rect 35025 3996 35149 4010
rect 35183 4000 35200 4010
rect 35183 3996 35195 4000
rect 34979 3992 35195 3996
rect 34979 3990 35037 3992
rect 35137 3990 35195 3992
rect 34812 3946 34952 3958
rect 34812 3570 34912 3946
rect 34946 3570 34952 3946
rect 34812 3558 34952 3570
rect 34812 3457 34818 3558
rect 34980 3526 35036 3990
rect 35064 3946 35110 3958
rect 35064 3570 35070 3946
rect 35104 3570 35110 3946
rect 35064 3558 35110 3570
rect 34979 3520 35037 3526
rect 34979 3486 34991 3520
rect 35025 3486 35037 3520
rect 34979 3480 35037 3486
rect 33990 3445 34818 3457
rect 32840 3430 33880 3440
rect 32840 3350 32850 3430
rect 33870 3350 33880 3430
rect 32840 3340 33880 3350
rect 32240 3244 32880 3280
rect 33990 3250 34800 3445
rect 35070 3440 35104 3558
rect 35138 3526 35194 3990
rect 35228 3958 35262 4128
rect 35540 4071 35740 4140
rect 35514 4059 35740 4071
rect 35295 4030 35353 4036
rect 35295 3996 35307 4030
rect 35341 3996 35353 4030
rect 35295 3990 35353 3996
rect 35222 3946 35268 3958
rect 35222 3570 35228 3946
rect 35262 3570 35268 3946
rect 35222 3558 35268 3570
rect 35296 3526 35352 3990
rect 35380 3946 35426 3958
rect 35380 3570 35386 3946
rect 35420 3570 35426 3946
rect 35380 3558 35426 3570
rect 35137 3520 35353 3526
rect 35137 3486 35149 3520
rect 35183 3486 35307 3520
rect 35341 3486 35353 3520
rect 35137 3480 35353 3486
rect 35386 3440 35420 3558
rect 35514 3457 35520 4059
rect 35554 3457 35740 4059
rect 36060 3930 36140 4420
rect 36448 4418 36460 4420
rect 36836 4450 36848 4452
rect 36836 4420 36850 4450
rect 36836 4418 36848 4420
rect 36448 4412 36848 4418
rect 36370 4373 36416 4385
rect 36370 4340 36376 4373
rect 36290 4330 36376 4340
rect 36410 4370 36416 4373
rect 36880 4373 36926 4385
rect 36880 4370 36886 4373
rect 36290 4260 36300 4330
rect 36290 4250 36376 4260
rect 36370 4239 36376 4250
rect 36410 4240 36886 4370
rect 36410 4239 36416 4240
rect 36370 4227 36416 4239
rect 36880 4239 36886 4240
rect 36920 4239 36926 4373
rect 36880 4227 36926 4239
rect 36448 4194 36848 4200
rect 36448 4160 36460 4194
rect 36836 4190 36848 4194
rect 37000 4190 37080 4680
rect 37234 4676 37246 4680
rect 37622 4676 37634 4710
rect 37234 4670 37634 4676
rect 37156 4631 37202 4643
rect 37156 4497 37162 4631
rect 37196 4630 37202 4631
rect 37666 4631 37712 4643
rect 37666 4630 37672 4631
rect 37196 4500 37672 4630
rect 37706 4600 37712 4631
rect 37706 4590 37780 4600
rect 37770 4520 37780 4590
rect 37196 4497 37202 4500
rect 37156 4485 37202 4497
rect 37666 4497 37672 4500
rect 37706 4510 37780 4520
rect 37706 4497 37712 4510
rect 37666 4485 37712 4497
rect 37234 4452 37634 4458
rect 37234 4418 37246 4452
rect 37622 4450 37634 4452
rect 37930 4450 38010 4940
rect 37622 4420 38010 4450
rect 37622 4418 37634 4420
rect 37234 4412 37634 4418
rect 37156 4373 37202 4385
rect 37156 4239 37162 4373
rect 37196 4370 37202 4373
rect 37666 4373 37712 4385
rect 37666 4370 37672 4373
rect 37196 4240 37672 4370
rect 37706 4340 37712 4373
rect 37706 4330 37780 4340
rect 37770 4260 37780 4330
rect 37196 4239 37202 4240
rect 37156 4227 37202 4239
rect 37666 4239 37672 4240
rect 37706 4250 37780 4260
rect 37706 4239 37712 4250
rect 37666 4227 37712 4239
rect 37234 4194 37634 4200
rect 37234 4190 37246 4194
rect 36836 4160 37246 4190
rect 37622 4160 37634 4194
rect 36448 4154 36848 4160
rect 36370 4115 36416 4127
rect 36370 4080 36376 4115
rect 36290 4070 36376 4080
rect 36410 4110 36416 4115
rect 36880 4115 36926 4127
rect 36880 4110 36886 4115
rect 36290 4000 36300 4070
rect 36290 3990 36376 4000
rect 36370 3981 36376 3990
rect 36410 3981 36886 4110
rect 36920 3981 36926 4115
rect 36370 3980 36926 3981
rect 36370 3969 36416 3980
rect 36880 3969 36926 3980
rect 36448 3936 36848 3942
rect 36448 3930 36460 3936
rect 36060 3902 36460 3930
rect 36836 3902 36848 3936
rect 36060 3900 36848 3902
rect 36060 3860 36140 3900
rect 36448 3896 36848 3900
rect 35514 3445 35740 3457
rect 35060 3430 35420 3440
rect 35060 3350 35070 3430
rect 35410 3350 35420 3430
rect 35060 3340 35420 3350
rect 35540 3340 35740 3445
rect 36370 3580 36530 3590
rect 36370 3440 36380 3580
rect 36520 3560 36530 3580
rect 37000 3560 37080 4160
rect 37234 4154 37634 4160
rect 37156 4115 37202 4127
rect 37156 3981 37162 4115
rect 37196 4110 37202 4115
rect 37666 4115 37712 4127
rect 37666 4110 37672 4115
rect 37196 3981 37672 4110
rect 37706 4080 37712 4115
rect 37706 4070 37780 4080
rect 37770 4000 37780 4070
rect 37706 3990 37780 4000
rect 37706 3981 37712 3990
rect 37156 3980 37712 3981
rect 37156 3969 37202 3980
rect 37666 3969 37712 3980
rect 37234 3936 37634 3942
rect 37234 3902 37246 3936
rect 37622 3930 37634 3936
rect 37930 3930 38010 4420
rect 37622 3902 38010 3930
rect 37234 3900 38010 3902
rect 37234 3896 37634 3900
rect 37930 3860 38010 3900
rect 36520 3460 37080 3560
rect 36520 3440 36530 3460
rect 36370 3430 36530 3440
rect 35540 3260 36200 3340
rect 33980 3244 34800 3250
rect 32240 3238 32882 3244
rect 32240 3204 32347 3238
rect 32787 3204 32882 3238
rect 32240 3198 32882 3204
rect 32240 3129 32348 3198
rect 18050 3010 18210 3020
rect 18050 2870 18060 3010
rect 18200 2870 18210 3010
rect 18050 2860 18210 2870
rect 17768 2780 17970 2790
rect 17960 2640 17970 2780
rect 17768 2630 17970 2640
rect 17768 2528 17774 2630
rect 17728 2516 17774 2528
rect 32240 2527 32258 3129
rect 32292 3028 32348 3129
rect 32460 3156 32674 3162
rect 32460 3106 32466 3156
rect 32459 3068 32466 3106
rect 32668 3106 32674 3156
rect 32786 3129 32882 3198
rect 32668 3068 32675 3106
rect 32459 3066 32471 3068
rect 32505 3066 32629 3068
rect 32663 3066 32675 3068
rect 32459 3062 32675 3066
rect 32459 3060 32517 3062
rect 32617 3060 32675 3062
rect 32292 3016 32432 3028
rect 32292 2640 32392 3016
rect 32426 2640 32432 3016
rect 32292 2628 32432 2640
rect 32292 2527 32392 2628
rect 32460 2596 32516 3060
rect 32544 3016 32590 3028
rect 32544 2640 32550 3016
rect 32584 2640 32590 3016
rect 32544 2628 32590 2640
rect 32459 2590 32517 2596
rect 32459 2556 32471 2590
rect 32505 2556 32517 2590
rect 32459 2550 32517 2556
rect -140 2480 14240 2500
rect 17260 2480 17300 2516
rect 17570 2480 17610 2516
rect 32240 2480 32392 2527
rect 32548 2520 32586 2628
rect 32618 2596 32674 3060
rect 32786 3028 32842 3129
rect 32702 3016 32842 3028
rect 32702 2640 32708 3016
rect 32742 2640 32842 3016
rect 32702 2628 32842 2640
rect 32617 2590 32675 2596
rect 32617 2556 32629 2590
rect 32663 2556 32675 2590
rect 32617 2550 32675 2556
rect 32742 2527 32842 2628
rect 32876 2760 32882 3129
rect 33852 3238 34800 3244
rect 33852 3204 33947 3238
rect 34387 3220 34800 3238
rect 35360 3238 36200 3260
rect 34387 3204 34680 3220
rect 33852 3198 34680 3204
rect 33852 3129 33948 3198
rect 33852 2760 33858 3129
rect 32876 2527 33858 2760
rect 33892 3028 33948 3129
rect 34060 3156 34274 3162
rect 34060 3106 34066 3156
rect 34059 3068 34066 3106
rect 34268 3106 34274 3156
rect 34386 3129 34680 3198
rect 34268 3068 34275 3106
rect 34059 3066 34071 3068
rect 34105 3066 34229 3068
rect 34263 3066 34275 3068
rect 34059 3062 34275 3066
rect 34059 3060 34117 3062
rect 34217 3060 34275 3062
rect 33892 3016 34032 3028
rect 33892 2640 33992 3016
rect 34026 2640 34032 3016
rect 33892 2628 34032 2640
rect 33892 2527 33992 2628
rect 34060 2596 34116 3060
rect 34144 3016 34190 3028
rect 34144 2640 34150 3016
rect 34184 2640 34190 3016
rect 34144 2628 34190 2640
rect 34059 2590 34117 2596
rect 34059 2556 34071 2590
rect 34105 2556 34117 2590
rect 34059 2550 34117 2556
rect -140 2380 32392 2480
rect 32440 2510 32700 2520
rect 32440 2430 32450 2510
rect 32690 2430 32700 2510
rect 32440 2420 32700 2430
rect 32742 2380 33992 2527
rect 34148 2520 34186 2628
rect 34218 2596 34274 3060
rect 34386 3028 34442 3129
rect 34302 3016 34442 3028
rect 34302 2640 34308 3016
rect 34342 2640 34442 3016
rect 34302 2628 34442 2640
rect 34217 2590 34275 2596
rect 34217 2556 34229 2590
rect 34263 2556 34275 2590
rect 34217 2550 34275 2556
rect 34342 2527 34442 2628
rect 34476 2527 34680 3129
rect 34040 2510 34300 2520
rect 34040 2430 34050 2510
rect 34290 2430 34300 2510
rect 34040 2420 34300 2430
rect 34342 2380 34680 2527
rect 35360 3204 35547 3238
rect 35987 3204 36200 3238
rect 35360 3198 36200 3204
rect 35360 3129 35548 3198
rect 35360 2527 35458 3129
rect 35492 3028 35548 3129
rect 35660 3156 35874 3162
rect 35660 3106 35666 3156
rect 35659 3068 35666 3106
rect 35868 3106 35874 3156
rect 35986 3129 36200 3198
rect 35868 3068 35875 3106
rect 35659 3066 35671 3068
rect 35705 3066 35829 3068
rect 35863 3066 35875 3068
rect 35659 3062 35875 3066
rect 35659 3060 35717 3062
rect 35817 3060 35875 3062
rect 35492 3016 35632 3028
rect 35492 2640 35592 3016
rect 35626 2640 35632 3016
rect 35492 2628 35632 2640
rect 35492 2527 35592 2628
rect 35660 2596 35716 3060
rect 35744 3016 35790 3028
rect 35744 2640 35750 3016
rect 35784 2640 35790 3016
rect 35744 2628 35790 2640
rect 35659 2590 35717 2596
rect 35659 2556 35671 2590
rect 35705 2556 35717 2590
rect 35659 2550 35717 2556
rect 35360 2380 35592 2527
rect 35748 2520 35786 2628
rect 35818 2596 35874 3060
rect 35986 3028 36042 3129
rect 35902 3016 36042 3028
rect 35902 2640 35908 3016
rect 35942 2640 36042 3016
rect 35902 2628 36042 2640
rect 35817 2590 35875 2596
rect 35817 2556 35829 2590
rect 35863 2556 35875 2590
rect 35817 2550 35875 2556
rect 35942 2527 36042 2628
rect 36076 2527 36200 3129
rect 35640 2510 35900 2520
rect 35640 2430 35650 2510
rect 35890 2430 35900 2510
rect 35640 2420 35900 2430
rect 35942 2380 36200 2527
rect -140 2235 37880 2380
rect -140 2229 38065 2235
rect -140 2195 -117 2229
rect 1253 2195 1483 2229
rect 2853 2195 3083 2229
rect 4453 2195 4683 2229
rect 6053 2195 6283 2229
rect 7653 2195 7883 2229
rect 9253 2195 9483 2229
rect 10853 2195 11083 2229
rect 12453 2195 12683 2229
rect 14053 2195 14283 2229
rect 15653 2195 15883 2229
rect 17253 2195 17483 2229
rect 18853 2195 19083 2229
rect 20453 2195 20683 2229
rect 22053 2195 22283 2229
rect 23653 2195 23883 2229
rect 25253 2195 25483 2229
rect 26853 2195 27083 2229
rect 28453 2195 28683 2229
rect 30053 2195 30283 2229
rect 31653 2195 31883 2229
rect 33253 2195 33483 2229
rect 34853 2195 35083 2229
rect 36453 2195 36683 2229
rect 38053 2195 38065 2229
rect -140 2095 480 2195
rect -140 2061 71 2095
rect 447 2061 480 2095
rect -140 2060 480 2061
rect -140 2007 0 2060
rect 59 2055 480 2060
rect -140 1995 27 2007
rect -140 1303 -13 1995
rect 21 1303 27 1995
rect -140 1291 27 1303
rect -140 882 0 1291
rect 440 1243 480 2055
rect 660 2189 38065 2195
rect 660 2180 37880 2189
rect 660 2095 11160 2180
rect 660 2061 689 2095
rect 1065 2061 1671 2095
rect 2047 2061 2289 2095
rect 2665 2061 3271 2095
rect 3647 2061 3889 2095
rect 4265 2061 4871 2095
rect 5247 2061 5489 2095
rect 5865 2061 6471 2095
rect 6847 2061 7089 2095
rect 7465 2061 8071 2095
rect 8447 2061 8689 2095
rect 9065 2061 9671 2095
rect 10047 2061 10289 2095
rect 10665 2061 11160 2095
rect 660 2060 11160 2061
rect 11240 2095 12300 2140
rect 11240 2061 11271 2095
rect 11647 2061 11889 2095
rect 12265 2061 12300 2095
rect 11240 2060 12300 2061
rect 12380 2060 12760 2180
rect 12840 2095 13900 2140
rect 12840 2061 12871 2095
rect 13247 2061 13489 2095
rect 13865 2061 13900 2095
rect 12840 2060 13900 2061
rect 13980 2100 31780 2180
rect 32060 2130 34680 2140
rect 32060 2101 32450 2130
rect 13980 2095 14870 2100
rect 13980 2061 14471 2095
rect 14847 2061 14870 2095
rect 13980 2060 14870 2061
rect 15070 2095 31780 2100
rect 15070 2061 15089 2095
rect 15465 2061 16071 2095
rect 16447 2061 16689 2095
rect 17065 2061 17671 2095
rect 18047 2061 18289 2095
rect 18665 2061 19271 2095
rect 19647 2061 19889 2095
rect 20265 2061 20871 2095
rect 21247 2061 21489 2095
rect 21865 2061 22471 2095
rect 22847 2061 23089 2095
rect 23465 2061 24071 2095
rect 24447 2061 24689 2095
rect 25065 2061 25671 2095
rect 26047 2061 26289 2095
rect 26665 2061 27271 2095
rect 27647 2061 27889 2095
rect 28265 2061 28871 2095
rect 29247 2061 29489 2095
rect 29865 2061 30471 2095
rect 30847 2061 31089 2095
rect 31465 2061 31780 2095
rect 15070 2060 31780 2061
rect 32059 2095 32450 2101
rect 32690 2095 34050 2130
rect 34290 2095 34680 2130
rect 35270 2130 36270 2140
rect 35270 2101 35650 2130
rect 32059 2061 32071 2095
rect 32447 2070 32450 2095
rect 32447 2061 32689 2070
rect 33065 2061 33671 2095
rect 34047 2070 34050 2095
rect 34047 2061 34289 2070
rect 34665 2061 34680 2095
rect 32059 2060 34680 2061
rect 35259 2095 35650 2101
rect 35890 2101 36270 2130
rect 35890 2095 36277 2101
rect 35259 2061 35271 2095
rect 35647 2070 35650 2095
rect 35647 2061 35889 2070
rect 36265 2061 36277 2095
rect 35259 2060 36277 2061
rect 36760 2095 37880 2180
rect 36760 2061 36871 2095
rect 37247 2061 37489 2095
rect 37865 2061 37880 2095
rect 36760 2060 37880 2061
rect 660 2055 1077 2060
rect 1659 2055 2059 2060
rect 2277 2055 2677 2060
rect 3259 2055 3659 2060
rect 3877 2055 4277 2060
rect 4859 2055 5259 2060
rect 5477 2055 5877 2060
rect 6459 2055 6859 2060
rect 7077 2055 7477 2060
rect 8059 2055 8459 2060
rect 8677 2055 9077 2060
rect 9659 2055 10059 2060
rect 10277 2055 10677 2060
rect 11259 2055 11659 2060
rect 11877 2055 12277 2060
rect 12859 2055 13259 2060
rect 13477 2055 13877 2060
rect 14459 2055 14859 2060
rect 15077 2055 15477 2060
rect 16059 2055 16459 2060
rect 16677 2055 17077 2060
rect 17659 2055 18059 2060
rect 18277 2055 18677 2060
rect 19259 2055 19659 2060
rect 19877 2055 20277 2060
rect 20859 2055 21259 2060
rect 21477 2055 21877 2060
rect 22459 2055 22859 2060
rect 23077 2055 23477 2060
rect 24059 2055 24459 2060
rect 24677 2055 25077 2060
rect 25659 2055 26059 2060
rect 26277 2055 26677 2060
rect 27259 2055 27659 2060
rect 27877 2055 28277 2060
rect 28859 2055 29259 2060
rect 29477 2055 29877 2060
rect 30459 2055 30859 2060
rect 31077 2055 31477 2060
rect 32059 2055 32459 2060
rect 32677 2055 33077 2060
rect 33659 2055 34059 2060
rect 34277 2055 34677 2060
rect 35259 2055 35659 2060
rect 35877 2055 36277 2060
rect 36859 2055 37259 2060
rect 37477 2055 37877 2060
rect 59 1237 480 1243
rect 59 1203 71 1237
rect 447 1203 480 1237
rect 59 1197 480 1203
rect 440 955 480 1197
rect 59 949 480 955
rect 59 915 71 949
rect 447 915 480 949
rect 59 909 480 915
rect -140 870 27 882
rect -140 736 -13 870
rect 21 736 27 870
rect -140 724 27 736
rect -140 460 0 724
rect 440 697 480 909
rect 660 1243 710 2055
rect 14900 2007 15040 2010
rect 1109 1995 1155 2007
rect 1109 1303 1115 1995
rect 1149 1303 1155 1995
rect 1109 1291 1155 1303
rect 1581 1995 1627 2007
rect 1581 1303 1587 1995
rect 1621 1303 1627 1995
rect 1581 1291 1627 1303
rect 2091 2000 2137 2007
rect 2199 2000 2245 2007
rect 2091 1995 2245 2000
rect 2091 1303 2097 1995
rect 2131 1990 2205 1995
rect 2131 1303 2205 1310
rect 2239 1303 2245 1995
rect 2091 1300 2245 1303
rect 2091 1291 2137 1300
rect 2199 1291 2245 1300
rect 2709 1995 2755 2007
rect 2709 1303 2715 1995
rect 2749 1303 2755 1995
rect 2709 1291 2755 1303
rect 3181 1995 3227 2007
rect 3181 1303 3187 1995
rect 3221 1303 3227 1995
rect 3181 1291 3227 1303
rect 3691 2000 3737 2007
rect 3799 2000 3845 2007
rect 3691 1995 3845 2000
rect 3691 1303 3697 1995
rect 3731 1990 3805 1995
rect 3731 1303 3805 1310
rect 3839 1303 3845 1995
rect 3691 1300 3845 1303
rect 3691 1291 3737 1300
rect 3799 1291 3845 1300
rect 4309 1995 4355 2007
rect 4309 1303 4315 1995
rect 4349 1303 4355 1995
rect 4309 1291 4355 1303
rect 4781 1995 4827 2007
rect 4781 1303 4787 1995
rect 4821 1303 4827 1995
rect 4781 1291 4827 1303
rect 5291 2000 5337 2007
rect 5399 2000 5445 2007
rect 5291 1995 5445 2000
rect 5291 1303 5297 1995
rect 5331 1990 5405 1995
rect 5331 1303 5405 1310
rect 5439 1303 5445 1995
rect 5291 1300 5445 1303
rect 5291 1291 5337 1300
rect 5399 1291 5445 1300
rect 5909 1995 5955 2007
rect 5909 1303 5915 1995
rect 5949 1303 5955 1995
rect 5909 1291 5955 1303
rect 6381 1995 6427 2007
rect 6381 1303 6387 1995
rect 6421 1303 6427 1995
rect 6381 1291 6427 1303
rect 6891 2000 6937 2007
rect 6999 2000 7045 2007
rect 6891 1995 7045 2000
rect 6891 1303 6897 1995
rect 6931 1990 7005 1995
rect 6931 1303 7005 1310
rect 7039 1303 7045 1995
rect 6891 1300 7045 1303
rect 6891 1291 6937 1300
rect 6999 1291 7045 1300
rect 7509 1995 7555 2007
rect 7509 1303 7515 1995
rect 7549 1303 7555 1995
rect 7509 1291 7555 1303
rect 7981 1995 8027 2007
rect 7981 1303 7987 1995
rect 8021 1303 8027 1995
rect 7981 1291 8027 1303
rect 8491 2000 8537 2007
rect 8599 2000 8645 2007
rect 8491 1995 8645 2000
rect 8491 1303 8497 1995
rect 8531 1990 8605 1995
rect 8531 1303 8605 1310
rect 8639 1303 8645 1995
rect 8491 1300 8645 1303
rect 8491 1291 8537 1300
rect 8599 1291 8645 1300
rect 9109 1995 9155 2007
rect 9109 1303 9115 1995
rect 9149 1303 9155 1995
rect 9109 1291 9155 1303
rect 9581 1995 9627 2007
rect 9581 1303 9587 1995
rect 9621 1303 9627 1995
rect 9581 1291 9627 1303
rect 10091 2000 10137 2007
rect 10199 2000 10245 2007
rect 10091 1995 10245 2000
rect 10091 1303 10097 1995
rect 10131 1990 10205 1995
rect 10131 1303 10205 1310
rect 10239 1303 10245 1995
rect 10091 1300 10245 1303
rect 10091 1291 10137 1300
rect 10199 1291 10245 1300
rect 10709 1995 10755 2007
rect 10709 1303 10715 1995
rect 10749 1303 10755 1995
rect 11181 1995 11227 2007
rect 11181 1960 11187 1995
rect 11020 1950 11187 1960
rect 11020 1330 11030 1950
rect 11150 1330 11187 1950
rect 11020 1320 11187 1330
rect 10709 1291 10755 1303
rect 11181 1303 11187 1320
rect 11221 1303 11227 1995
rect 11181 1291 11227 1303
rect 11691 2000 11737 2007
rect 11799 2000 11845 2007
rect 11691 1995 11845 2000
rect 11691 1303 11697 1995
rect 11731 1303 11805 1995
rect 11839 1303 11845 1995
rect 11691 1300 11845 1303
rect 11691 1291 11737 1300
rect 11799 1291 11845 1300
rect 12309 1995 12355 2007
rect 12309 1303 12315 1995
rect 12349 1960 12355 1995
rect 12781 1995 12827 2007
rect 12781 1960 12787 1995
rect 12349 1950 12787 1960
rect 12349 1330 12610 1950
rect 12730 1330 12787 1950
rect 12349 1320 12787 1330
rect 12349 1303 12355 1320
rect 12309 1291 12355 1303
rect 12781 1303 12787 1320
rect 12821 1303 12827 1995
rect 12781 1291 12827 1303
rect 13291 2000 13337 2007
rect 13399 2000 13445 2007
rect 13291 1995 13445 2000
rect 13291 1303 13297 1995
rect 13331 1303 13405 1995
rect 13439 1303 13445 1995
rect 13291 1300 13445 1303
rect 13291 1291 13337 1300
rect 13399 1291 13445 1300
rect 13909 1995 13955 2007
rect 13909 1303 13915 1995
rect 13949 1960 13955 1995
rect 14381 1995 14427 2007
rect 13949 1950 14120 1960
rect 13949 1330 13990 1950
rect 14110 1330 14120 1950
rect 13949 1303 14120 1330
rect 13909 1291 14120 1303
rect 14381 1303 14387 1995
rect 14421 1303 14427 1995
rect 14381 1291 14427 1303
rect 14891 1995 15045 2007
rect 14891 1303 14897 1995
rect 14931 1980 15005 1995
rect 14931 1303 15005 1320
rect 15039 1303 15045 1995
rect 14891 1291 15045 1303
rect 15509 1995 15555 2007
rect 15509 1303 15515 1995
rect 15549 1303 15555 1995
rect 15509 1291 15555 1303
rect 15981 1995 16027 2007
rect 15981 1303 15987 1995
rect 16021 1303 16027 1995
rect 15981 1291 16027 1303
rect 16491 2000 16537 2007
rect 16599 2000 16645 2007
rect 16491 1995 16645 2000
rect 16491 1303 16497 1995
rect 16531 1990 16605 1995
rect 16531 1303 16605 1310
rect 16639 1303 16645 1995
rect 16491 1300 16645 1303
rect 16491 1291 16537 1300
rect 16599 1291 16645 1300
rect 17109 1995 17155 2007
rect 17109 1303 17115 1995
rect 17149 1303 17155 1995
rect 17109 1291 17155 1303
rect 17581 1995 17627 2007
rect 17581 1303 17587 1995
rect 17621 1303 17627 1995
rect 17581 1291 17627 1303
rect 18091 2000 18137 2007
rect 18199 2000 18245 2007
rect 18091 1995 18245 2000
rect 18091 1303 18097 1995
rect 18131 1990 18205 1995
rect 18131 1303 18205 1310
rect 18239 1303 18245 1995
rect 18091 1300 18245 1303
rect 18091 1291 18137 1300
rect 18199 1291 18245 1300
rect 18709 1995 18755 2007
rect 18709 1303 18715 1995
rect 18749 1303 18755 1995
rect 18709 1291 18755 1303
rect 19181 1995 19227 2007
rect 19181 1303 19187 1995
rect 19221 1303 19227 1995
rect 19181 1291 19227 1303
rect 19691 2000 19737 2007
rect 19799 2000 19845 2007
rect 19691 1995 19845 2000
rect 19691 1303 19697 1995
rect 19731 1990 19805 1995
rect 19731 1303 19805 1310
rect 19839 1303 19845 1995
rect 19691 1300 19845 1303
rect 19691 1291 19737 1300
rect 19799 1291 19845 1300
rect 20309 1995 20355 2007
rect 20309 1303 20315 1995
rect 20349 1303 20355 1995
rect 20309 1291 20355 1303
rect 20781 1995 20827 2007
rect 20781 1303 20787 1995
rect 20821 1303 20827 1995
rect 20781 1291 20827 1303
rect 21291 2000 21337 2007
rect 21399 2000 21445 2007
rect 21291 1995 21445 2000
rect 21291 1303 21297 1995
rect 21331 1990 21405 1995
rect 21331 1303 21405 1310
rect 21439 1303 21445 1995
rect 21291 1300 21445 1303
rect 21291 1291 21337 1300
rect 21399 1291 21445 1300
rect 21909 1995 21955 2007
rect 21909 1303 21915 1995
rect 21949 1303 21955 1995
rect 21909 1291 21955 1303
rect 22381 1995 22427 2007
rect 22381 1303 22387 1995
rect 22421 1303 22427 1995
rect 22381 1291 22427 1303
rect 22891 2000 22937 2007
rect 22999 2000 23045 2007
rect 22891 1995 23045 2000
rect 22891 1303 22897 1995
rect 22931 1990 23005 1995
rect 22931 1303 23005 1310
rect 23039 1303 23045 1995
rect 22891 1300 23045 1303
rect 22891 1291 22937 1300
rect 22999 1291 23045 1300
rect 23509 1995 23555 2007
rect 23509 1303 23515 1995
rect 23549 1303 23555 1995
rect 23509 1291 23555 1303
rect 23981 1995 24027 2007
rect 23981 1303 23987 1995
rect 24021 1303 24027 1995
rect 23981 1291 24027 1303
rect 24491 2000 24537 2007
rect 24599 2000 24645 2007
rect 24491 1995 24645 2000
rect 24491 1303 24497 1995
rect 24531 1990 24605 1995
rect 24531 1303 24605 1310
rect 24639 1303 24645 1995
rect 24491 1300 24645 1303
rect 24491 1291 24537 1300
rect 24599 1291 24645 1300
rect 25109 1995 25155 2007
rect 25109 1303 25115 1995
rect 25149 1303 25155 1995
rect 25109 1291 25155 1303
rect 25581 1995 25627 2007
rect 25581 1303 25587 1995
rect 25621 1303 25627 1995
rect 25581 1291 25627 1303
rect 26091 2000 26137 2007
rect 26199 2000 26245 2007
rect 26091 1995 26245 2000
rect 26091 1303 26097 1995
rect 26131 1990 26205 1995
rect 26131 1303 26205 1310
rect 26239 1303 26245 1995
rect 26091 1300 26245 1303
rect 26091 1291 26137 1300
rect 26199 1291 26245 1300
rect 26709 1995 26755 2007
rect 26709 1303 26715 1995
rect 26749 1303 26755 1995
rect 26709 1291 26755 1303
rect 27181 1995 27227 2007
rect 27181 1303 27187 1995
rect 27221 1303 27227 1995
rect 27181 1291 27227 1303
rect 27691 2000 27737 2007
rect 27799 2000 27845 2007
rect 27691 1995 27845 2000
rect 27691 1303 27697 1995
rect 27731 1990 27805 1995
rect 27731 1303 27805 1310
rect 27839 1303 27845 1995
rect 27691 1300 27845 1303
rect 27691 1291 27737 1300
rect 27799 1291 27845 1300
rect 28309 1995 28355 2007
rect 28309 1303 28315 1995
rect 28349 1303 28355 1995
rect 28309 1291 28355 1303
rect 28781 1995 28827 2007
rect 28781 1303 28787 1995
rect 28821 1303 28827 1995
rect 28781 1291 28827 1303
rect 29291 2000 29337 2007
rect 29399 2000 29445 2007
rect 29291 1995 29445 2000
rect 29291 1303 29297 1995
rect 29331 1990 29405 1995
rect 29331 1303 29405 1310
rect 29439 1303 29445 1995
rect 29291 1300 29445 1303
rect 29291 1291 29337 1300
rect 29399 1291 29445 1300
rect 29909 1995 29955 2007
rect 29909 1303 29915 1995
rect 29949 1303 29955 1995
rect 29909 1291 29955 1303
rect 30381 1995 30427 2007
rect 30381 1303 30387 1995
rect 30421 1303 30427 1995
rect 30381 1291 30427 1303
rect 30891 2000 30937 2007
rect 30999 2000 31045 2007
rect 30891 1995 31045 2000
rect 30891 1303 30897 1995
rect 30931 1990 31005 1995
rect 30931 1303 31005 1310
rect 31039 1303 31045 1995
rect 30891 1300 31045 1303
rect 30891 1291 30937 1300
rect 30999 1291 31045 1300
rect 31509 1995 31555 2007
rect 31509 1303 31515 1995
rect 31549 1303 31555 1995
rect 31509 1291 31555 1303
rect 31981 1995 32027 2007
rect 31981 1303 31987 1995
rect 32021 1303 32027 1995
rect 31981 1291 32027 1303
rect 32491 2000 32537 2007
rect 32599 2000 32645 2007
rect 32491 1995 32645 2000
rect 32491 1303 32497 1995
rect 32531 1990 32605 1995
rect 32531 1303 32605 1310
rect 32639 1303 32645 1995
rect 32491 1300 32645 1303
rect 32491 1291 32537 1300
rect 32599 1291 32645 1300
rect 33109 1995 33155 2007
rect 33109 1303 33115 1995
rect 33149 1303 33155 1995
rect 33109 1291 33155 1303
rect 33581 1995 33627 2007
rect 33581 1303 33587 1995
rect 33621 1303 33627 1995
rect 33581 1291 33627 1303
rect 34091 2000 34137 2007
rect 34199 2000 34245 2007
rect 34091 1995 34245 2000
rect 34091 1303 34097 1995
rect 34131 1990 34205 1995
rect 34131 1303 34205 1310
rect 34239 1303 34245 1995
rect 34091 1300 34245 1303
rect 34091 1291 34137 1300
rect 34199 1291 34245 1300
rect 34709 1995 34755 2007
rect 34709 1303 34715 1995
rect 34749 1303 34755 1995
rect 34709 1291 34755 1303
rect 35181 1995 35227 2007
rect 35181 1303 35187 1995
rect 35221 1303 35227 1995
rect 35181 1291 35227 1303
rect 35691 2000 35737 2007
rect 35799 2000 35845 2007
rect 35691 1995 35845 2000
rect 35691 1303 35697 1995
rect 35731 1990 35805 1995
rect 35731 1303 35805 1310
rect 35839 1303 35845 1995
rect 35691 1300 35845 1303
rect 35691 1291 35737 1300
rect 35799 1291 35845 1300
rect 36309 1995 36355 2007
rect 36309 1303 36315 1995
rect 36349 1303 36355 1995
rect 36309 1291 36355 1303
rect 36781 1995 36827 2007
rect 36781 1303 36787 1995
rect 36821 1303 36827 1995
rect 36781 1291 36827 1303
rect 37291 2000 37337 2007
rect 37399 2000 37445 2007
rect 37291 1995 37445 2000
rect 37291 1303 37297 1995
rect 37331 1990 37405 1995
rect 37331 1303 37405 1310
rect 37439 1303 37445 1995
rect 37291 1300 37445 1303
rect 37291 1291 37337 1300
rect 37399 1291 37445 1300
rect 37909 1995 37955 2007
rect 37909 1303 37915 1995
rect 37949 1303 37955 1995
rect 37909 1291 37955 1303
rect 660 1237 1077 1243
rect 660 1203 689 1237
rect 1065 1203 1077 1237
rect 660 1197 1077 1203
rect 1659 1237 2059 1243
rect 1659 1203 1671 1237
rect 2047 1203 2059 1237
rect 1659 1197 2059 1203
rect 2277 1237 2677 1243
rect 2277 1203 2289 1237
rect 2665 1203 2677 1237
rect 2277 1197 2677 1203
rect 3259 1237 3659 1243
rect 3259 1203 3271 1237
rect 3647 1203 3659 1237
rect 3259 1197 3659 1203
rect 3877 1237 4277 1243
rect 3877 1203 3889 1237
rect 4265 1203 4277 1237
rect 3877 1197 4277 1203
rect 4859 1237 5259 1243
rect 4859 1203 4871 1237
rect 5247 1203 5259 1237
rect 4859 1197 5259 1203
rect 5477 1237 5877 1243
rect 5477 1203 5489 1237
rect 5865 1203 5877 1237
rect 5477 1197 5877 1203
rect 6459 1237 6859 1243
rect 6459 1203 6471 1237
rect 6847 1203 6859 1237
rect 6459 1197 6859 1203
rect 7077 1237 7477 1243
rect 7077 1203 7089 1237
rect 7465 1203 7477 1237
rect 7077 1197 7477 1203
rect 8059 1237 8459 1243
rect 8059 1203 8071 1237
rect 8447 1203 8459 1237
rect 8059 1197 8459 1203
rect 8677 1237 9077 1243
rect 8677 1203 8689 1237
rect 9065 1203 9077 1237
rect 8677 1197 9077 1203
rect 9659 1237 10059 1243
rect 9659 1203 9671 1237
rect 10047 1203 10059 1237
rect 9659 1197 10059 1203
rect 10277 1237 10677 1243
rect 11259 1240 11659 1243
rect 11877 1240 12277 1243
rect 12859 1240 13259 1243
rect 13477 1240 13877 1243
rect 13910 1240 14120 1291
rect 10277 1203 10289 1237
rect 10665 1203 10677 1237
rect 10277 1197 10677 1203
rect 11240 1237 11680 1240
rect 11240 1230 11271 1237
rect 11647 1230 11680 1237
rect 660 955 710 1197
rect 1680 1160 2040 1197
rect 2300 1160 2660 1197
rect 3280 1160 3640 1197
rect 3900 1160 4260 1197
rect 4880 1160 5240 1197
rect 5500 1160 5860 1197
rect 6480 1160 6840 1197
rect 7100 1160 7460 1197
rect 8080 1160 8440 1197
rect 8700 1160 9060 1197
rect 9680 1160 10040 1197
rect 10300 1160 10660 1197
rect 1400 1150 10660 1160
rect 1400 1030 1410 1150
rect 1530 1030 3010 1150
rect 3130 1030 4610 1150
rect 4730 1030 6210 1150
rect 6330 1030 7810 1150
rect 7930 1030 9410 1150
rect 9530 1030 10660 1150
rect 11240 1070 11250 1230
rect 11670 1070 11680 1230
rect 11860 1237 13280 1240
rect 11860 1203 11889 1237
rect 12265 1203 12871 1237
rect 13247 1203 13280 1237
rect 11860 1120 13280 1203
rect 13477 1237 14120 1240
rect 13477 1203 13489 1237
rect 13865 1203 14120 1237
rect 13477 1197 14120 1203
rect 14459 1240 14859 1243
rect 14900 1240 15040 1291
rect 15077 1240 15477 1243
rect 14459 1237 15480 1240
rect 14459 1203 14471 1237
rect 14847 1203 15089 1237
rect 15465 1203 15480 1237
rect 14459 1197 15480 1203
rect 16059 1237 16459 1243
rect 16059 1203 16071 1237
rect 16447 1203 16459 1237
rect 16059 1197 16459 1203
rect 16677 1237 17077 1243
rect 16677 1203 16689 1237
rect 17065 1203 17077 1237
rect 16677 1197 17077 1203
rect 17659 1237 18059 1243
rect 17659 1203 17671 1237
rect 18047 1203 18059 1237
rect 17659 1197 18059 1203
rect 18277 1237 18677 1243
rect 18277 1203 18289 1237
rect 18665 1203 18677 1237
rect 18277 1197 18677 1203
rect 19259 1237 19659 1243
rect 19259 1203 19271 1237
rect 19647 1203 19659 1237
rect 19259 1197 19659 1203
rect 19877 1237 20277 1243
rect 19877 1203 19889 1237
rect 20265 1203 20277 1237
rect 19877 1197 20277 1203
rect 20859 1237 21259 1243
rect 20859 1203 20871 1237
rect 21247 1203 21259 1237
rect 20859 1197 21259 1203
rect 21477 1237 21877 1243
rect 21477 1203 21489 1237
rect 21865 1203 21877 1237
rect 21477 1197 21877 1203
rect 22459 1237 22859 1243
rect 22459 1203 22471 1237
rect 22847 1203 22859 1237
rect 22459 1197 22859 1203
rect 23077 1237 23477 1243
rect 23077 1203 23089 1237
rect 23465 1203 23477 1237
rect 23077 1197 23477 1203
rect 24059 1237 24459 1243
rect 24059 1203 24071 1237
rect 24447 1203 24459 1237
rect 24059 1197 24459 1203
rect 24677 1237 25077 1243
rect 24677 1203 24689 1237
rect 25065 1203 25077 1237
rect 24677 1197 25077 1203
rect 25659 1237 26059 1243
rect 25659 1203 25671 1237
rect 26047 1203 26059 1237
rect 25659 1197 26059 1203
rect 26277 1237 26677 1243
rect 26277 1203 26289 1237
rect 26665 1203 26677 1237
rect 26277 1197 26677 1203
rect 27259 1237 27659 1243
rect 27259 1203 27271 1237
rect 27647 1203 27659 1237
rect 27259 1197 27659 1203
rect 27877 1237 28277 1243
rect 27877 1203 27889 1237
rect 28265 1203 28277 1237
rect 27877 1197 28277 1203
rect 28859 1237 29259 1243
rect 28859 1203 28871 1237
rect 29247 1203 29259 1237
rect 28859 1197 29259 1203
rect 29477 1237 29877 1243
rect 29477 1203 29489 1237
rect 29865 1203 29877 1237
rect 29477 1197 29877 1203
rect 30459 1237 30859 1243
rect 30459 1203 30471 1237
rect 30847 1203 30859 1237
rect 30459 1197 30859 1203
rect 31077 1237 31477 1243
rect 31077 1203 31089 1237
rect 31465 1203 31477 1237
rect 31077 1197 31477 1203
rect 32059 1237 32459 1243
rect 32059 1203 32071 1237
rect 32447 1203 32459 1237
rect 32059 1197 32459 1203
rect 32677 1237 33077 1243
rect 32677 1203 32689 1237
rect 33065 1203 33077 1237
rect 32677 1197 33077 1203
rect 33659 1237 34059 1243
rect 33659 1203 33671 1237
rect 34047 1203 34059 1237
rect 33659 1197 34059 1203
rect 34277 1237 34677 1243
rect 34277 1203 34289 1237
rect 34665 1203 34677 1237
rect 34277 1197 34677 1203
rect 35259 1237 35659 1243
rect 35259 1203 35271 1237
rect 35647 1203 35659 1237
rect 35259 1197 35659 1203
rect 35877 1237 36277 1243
rect 35877 1203 35889 1237
rect 36265 1203 36277 1237
rect 35877 1197 36277 1203
rect 36859 1237 37259 1243
rect 36859 1203 36871 1237
rect 37247 1230 37259 1237
rect 37477 1237 37877 1243
rect 37247 1203 37260 1230
rect 36859 1197 37260 1203
rect 37477 1203 37489 1237
rect 37865 1203 37877 1237
rect 37477 1197 37877 1203
rect 13480 1120 14120 1197
rect 14460 1150 15480 1197
rect 16080 1160 16440 1197
rect 16700 1160 17060 1197
rect 17680 1160 18040 1197
rect 18300 1160 18660 1197
rect 19280 1160 19640 1197
rect 19900 1160 20260 1197
rect 20880 1160 21240 1197
rect 21500 1160 21860 1197
rect 22480 1160 22840 1197
rect 23100 1160 23460 1197
rect 24080 1160 24440 1197
rect 24700 1160 25060 1197
rect 25680 1160 26040 1197
rect 26300 1160 26660 1197
rect 27280 1160 27640 1197
rect 27900 1160 28260 1197
rect 28880 1160 29240 1197
rect 29500 1160 29860 1197
rect 30480 1160 30840 1197
rect 31100 1160 31460 1197
rect 32080 1160 32440 1197
rect 32700 1160 33060 1197
rect 33680 1160 34040 1197
rect 34300 1160 34660 1197
rect 35280 1160 35640 1197
rect 35900 1160 36260 1197
rect 15590 1150 17060 1160
rect 11240 1060 11680 1070
rect 1400 1020 10660 1030
rect 15590 1030 15600 1150
rect 15700 1030 17060 1150
rect 15590 1020 17060 1030
rect 17190 1150 18660 1160
rect 17190 1030 17200 1150
rect 17300 1030 18660 1150
rect 17190 1020 18660 1030
rect 18790 1150 20260 1160
rect 18790 1030 18800 1150
rect 18900 1030 20260 1150
rect 18790 1020 20260 1030
rect 20390 1150 21860 1160
rect 20390 1030 20400 1150
rect 20500 1030 21860 1150
rect 20390 1020 21860 1030
rect 21990 1150 23460 1160
rect 21990 1030 22000 1150
rect 22100 1030 23460 1150
rect 21990 1020 23460 1030
rect 23590 1150 25060 1160
rect 23590 1030 23600 1150
rect 23700 1030 25060 1150
rect 23590 1020 25060 1030
rect 25660 1150 28260 1160
rect 25660 1030 26800 1150
rect 26900 1030 28260 1150
rect 25660 1020 28260 1030
rect 28391 1150 31460 1160
rect 28391 1030 28400 1150
rect 28500 1030 31460 1150
rect 28391 1020 31460 1030
rect 32060 1020 34660 1160
rect 35260 1020 36260 1160
rect 1680 955 2040 1020
rect 2300 955 2660 1020
rect 3280 955 3640 1020
rect 3900 955 4260 1020
rect 4880 955 5240 1020
rect 5500 955 5860 1020
rect 6480 955 6840 1020
rect 7100 955 7460 1020
rect 8080 955 8440 1020
rect 8700 955 9060 1020
rect 9680 955 10040 1020
rect 10300 955 10660 1020
rect 16080 975 16440 1020
rect 16700 975 17060 1020
rect 17680 975 18040 1020
rect 18300 975 18660 1020
rect 19280 975 19640 1020
rect 19900 975 20260 1020
rect 20880 975 21240 1020
rect 21500 975 21860 1020
rect 22480 975 22840 1020
rect 23100 975 23460 1020
rect 24080 975 24440 1020
rect 24700 975 25060 1020
rect 25680 975 26040 1020
rect 26300 975 26660 1020
rect 27280 975 27640 1020
rect 27900 975 28260 1020
rect 28880 975 29240 1020
rect 29500 975 29860 1020
rect 30480 975 30840 1020
rect 31100 975 31460 1020
rect 32080 975 32440 1020
rect 32700 975 33060 1020
rect 33680 975 34040 1020
rect 34300 975 34660 1020
rect 35280 975 35640 1020
rect 35900 975 36260 1020
rect 16059 970 16459 975
rect 660 949 1077 955
rect 660 915 689 949
rect 1065 915 1077 949
rect 660 909 1077 915
rect 1659 949 2059 955
rect 1659 915 1671 949
rect 2047 915 2059 949
rect 1659 909 2059 915
rect 2277 949 2677 955
rect 2277 915 2289 949
rect 2665 915 2677 949
rect 2277 909 2677 915
rect 3259 949 3659 955
rect 3259 915 3271 949
rect 3647 915 3659 949
rect 3259 909 3659 915
rect 3877 949 4277 955
rect 3877 915 3889 949
rect 4265 915 4277 949
rect 3877 909 4277 915
rect 4859 949 5259 955
rect 4859 915 4871 949
rect 5247 915 5259 949
rect 4859 909 5259 915
rect 5477 949 5877 955
rect 5477 915 5489 949
rect 5865 915 5877 949
rect 5477 909 5877 915
rect 6459 949 6859 955
rect 6459 915 6471 949
rect 6847 915 6859 949
rect 6459 909 6859 915
rect 7077 949 7477 955
rect 7077 915 7089 949
rect 7465 915 7477 949
rect 7077 909 7477 915
rect 8059 949 8459 955
rect 8059 915 8071 949
rect 8447 915 8459 949
rect 8059 909 8459 915
rect 8677 949 9077 955
rect 8677 915 8689 949
rect 9065 915 9077 949
rect 8677 909 9077 915
rect 9659 949 10059 955
rect 9659 915 9671 949
rect 10047 915 10059 949
rect 9659 909 10059 915
rect 10277 949 10677 955
rect 10277 915 10289 949
rect 10665 915 10677 949
rect 10277 909 10677 915
rect 11259 949 11659 955
rect 11259 915 11271 949
rect 11647 915 11659 949
rect 11259 909 11659 915
rect 11877 949 12277 955
rect 11877 915 11889 949
rect 12265 915 12277 949
rect 11877 909 12277 915
rect 12859 949 13259 955
rect 12859 915 12871 949
rect 13247 915 13259 949
rect 12859 909 13259 915
rect 13477 949 13877 955
rect 13477 915 13489 949
rect 13865 915 13877 949
rect 13477 909 13877 915
rect 14459 949 14859 955
rect 14459 915 14471 949
rect 14847 915 14859 949
rect 14459 909 14859 915
rect 15077 949 15477 955
rect 15077 915 15089 949
rect 15465 915 15477 949
rect 15077 909 15477 915
rect 16059 949 16460 970
rect 16059 915 16071 949
rect 16447 915 16460 949
rect 16059 910 16460 915
rect 16677 949 17077 975
rect 16677 915 16689 949
rect 17065 915 17077 949
rect 16059 909 16459 910
rect 16677 909 17077 915
rect 17659 970 18059 975
rect 17659 949 18060 970
rect 17659 915 17671 949
rect 18047 915 18060 949
rect 17659 910 18060 915
rect 18277 949 18677 975
rect 18277 915 18289 949
rect 18665 915 18677 949
rect 17659 909 18059 910
rect 18277 909 18677 915
rect 19259 970 19659 975
rect 19259 949 19660 970
rect 19259 915 19271 949
rect 19647 915 19660 949
rect 19259 910 19660 915
rect 19877 949 20277 975
rect 19877 915 19889 949
rect 20265 915 20277 949
rect 19259 909 19659 910
rect 19877 909 20277 915
rect 20859 970 21259 975
rect 20859 949 21260 970
rect 20859 915 20871 949
rect 21247 915 21260 949
rect 20859 910 21260 915
rect 21477 949 21877 975
rect 21477 915 21489 949
rect 21865 915 21877 949
rect 20859 909 21259 910
rect 21477 909 21877 915
rect 22459 970 22859 975
rect 22459 949 22860 970
rect 22459 915 22471 949
rect 22847 915 22860 949
rect 22459 910 22860 915
rect 23077 949 23477 975
rect 23077 915 23089 949
rect 23465 915 23477 949
rect 22459 909 22859 910
rect 23077 909 23477 915
rect 24059 970 24459 975
rect 24059 949 24460 970
rect 24059 915 24071 949
rect 24447 915 24460 949
rect 24059 910 24460 915
rect 24677 949 25077 975
rect 24677 915 24689 949
rect 25065 915 25077 949
rect 24059 909 24459 910
rect 24677 909 25077 915
rect 25659 970 26059 975
rect 25659 949 26060 970
rect 25659 915 25671 949
rect 26047 915 26060 949
rect 25659 910 26060 915
rect 26277 949 26677 975
rect 26277 915 26289 949
rect 26665 915 26677 949
rect 25659 909 26059 910
rect 26277 909 26677 915
rect 27259 970 27659 975
rect 27259 949 27660 970
rect 27259 915 27271 949
rect 27647 915 27660 949
rect 27259 910 27660 915
rect 27877 949 28277 975
rect 27877 915 27889 949
rect 28265 915 28277 949
rect 27259 909 27659 910
rect 27877 909 28277 915
rect 28859 970 29259 975
rect 28859 949 29260 970
rect 28859 915 28871 949
rect 29247 915 29260 949
rect 28859 910 29260 915
rect 29477 949 29877 975
rect 29477 915 29489 949
rect 29865 915 29877 949
rect 28859 909 29259 910
rect 29477 909 29877 915
rect 30459 970 30859 975
rect 30459 949 30860 970
rect 30459 915 30471 949
rect 30847 915 30860 949
rect 30459 910 30860 915
rect 31077 949 31477 975
rect 32060 970 32459 975
rect 32060 955 32460 970
rect 31077 915 31089 949
rect 31465 915 31477 949
rect 30459 909 30859 910
rect 31077 909 31477 915
rect 32059 949 32460 955
rect 32059 915 32071 949
rect 32447 915 32460 949
rect 32059 910 32460 915
rect 32677 949 33077 975
rect 32677 915 32689 949
rect 33065 915 33077 949
rect 32059 909 32459 910
rect 32677 909 33077 915
rect 33659 970 34059 975
rect 33659 949 34060 970
rect 33659 915 33671 949
rect 34047 915 34060 949
rect 33659 910 34060 915
rect 34277 949 34677 975
rect 34277 915 34289 949
rect 34665 915 34677 949
rect 33659 909 34059 910
rect 34277 909 34677 915
rect 35259 970 35659 975
rect 35259 949 35660 970
rect 35259 915 35271 949
rect 35647 915 35660 949
rect 35259 910 35660 915
rect 35877 949 36277 975
rect 36870 955 37260 1197
rect 37480 955 37870 1197
rect 35877 915 35889 949
rect 36265 915 36277 949
rect 35259 909 35659 910
rect 35877 909 36277 915
rect 36859 949 37260 955
rect 36859 915 36871 949
rect 37247 930 37260 949
rect 37477 949 37877 955
rect 37247 915 37259 930
rect 36859 909 37259 915
rect 37477 915 37489 949
rect 37865 915 37877 949
rect 37477 909 37877 915
rect 59 691 480 697
rect 59 657 71 691
rect 447 657 480 691
rect 59 651 480 657
rect 440 460 480 651
rect -140 429 480 460
rect 660 697 710 909
rect 1109 870 1155 882
rect 1581 870 1627 882
rect 2091 870 2137 882
rect 2199 870 2245 882
rect 2709 870 2755 882
rect 3181 870 3227 882
rect 3691 870 3737 882
rect 3799 870 3845 882
rect 4309 870 4355 882
rect 4781 870 4827 882
rect 5291 870 5337 882
rect 5399 870 5445 882
rect 5909 870 5955 882
rect 6381 870 6427 882
rect 6891 870 6937 882
rect 6999 870 7045 882
rect 7509 870 7555 882
rect 7981 870 8027 882
rect 8491 870 8537 882
rect 8599 870 8645 882
rect 9109 870 9155 882
rect 9581 870 9627 882
rect 10091 870 10137 882
rect 10199 870 10245 882
rect 10709 870 10755 882
rect 11181 870 11227 882
rect 11420 870 11500 909
rect 11691 870 11737 882
rect 11799 870 11845 882
rect 12040 870 12120 909
rect 12309 880 12355 882
rect 12309 870 12520 880
rect 12781 870 12827 882
rect 13020 870 13100 909
rect 13291 870 13337 882
rect 13399 870 13445 882
rect 13640 870 13720 909
rect 13909 870 13955 882
rect 14381 870 14427 882
rect 14620 870 14700 909
rect 14891 870 14937 882
rect 14999 870 15045 882
rect 15240 870 15320 909
rect 15509 870 15555 882
rect 15981 870 16027 882
rect 16491 870 16537 882
rect 16599 870 16645 882
rect 17109 870 17155 882
rect 17581 870 17627 882
rect 18091 870 18137 882
rect 18199 870 18245 882
rect 18709 870 18755 882
rect 19181 870 19227 882
rect 19691 870 19737 882
rect 19799 870 19845 882
rect 20309 870 20355 882
rect 20781 870 20827 882
rect 21291 870 21337 882
rect 21399 870 21445 882
rect 21909 870 21955 882
rect 22381 870 22427 882
rect 22891 870 22937 882
rect 22999 870 23045 882
rect 23509 870 23555 882
rect 23981 870 24027 882
rect 24491 870 24537 882
rect 24599 870 24645 882
rect 25109 870 25155 882
rect 25581 870 25627 882
rect 26091 870 26137 882
rect 26199 870 26245 882
rect 26709 870 26755 882
rect 27181 870 27227 882
rect 27691 870 27737 882
rect 27799 870 27845 882
rect 28309 870 28355 882
rect 28781 870 28827 882
rect 29291 870 29337 882
rect 29399 870 29445 882
rect 29909 870 29955 882
rect 30381 870 30427 882
rect 30891 870 30937 882
rect 30999 870 31045 882
rect 31509 870 31555 882
rect 31981 870 32027 882
rect 32491 870 32537 882
rect 32599 870 32645 882
rect 33109 870 33155 882
rect 33581 870 33627 882
rect 34091 870 34137 882
rect 34199 870 34245 882
rect 34709 870 34755 882
rect 35181 870 35227 882
rect 35691 870 35737 882
rect 35799 870 35845 882
rect 36309 870 36355 882
rect 36781 870 36827 882
rect 37291 870 37337 882
rect 37399 870 37445 882
rect 37909 870 37955 882
rect 1109 736 1115 870
rect 1149 736 1155 870
rect 1540 740 1587 870
rect 1109 724 1155 736
rect 1581 736 1587 740
rect 1621 740 2097 870
rect 1621 736 1627 740
rect 1581 724 1627 736
rect 2091 736 2097 740
rect 2131 740 2205 870
rect 2131 736 2137 740
rect 2091 724 2137 736
rect 2199 736 2205 740
rect 2239 740 2715 870
rect 2239 736 2245 740
rect 2199 724 2245 736
rect 2709 736 2715 740
rect 2749 740 3187 870
rect 2749 736 2755 740
rect 2709 724 2755 736
rect 3181 736 3187 740
rect 3221 740 3697 870
rect 3221 736 3227 740
rect 3181 724 3227 736
rect 3691 736 3697 740
rect 3731 740 3805 870
rect 3731 736 3737 740
rect 3691 724 3737 736
rect 3799 736 3805 740
rect 3839 740 4315 870
rect 3839 736 3845 740
rect 3799 724 3845 736
rect 4309 736 4315 740
rect 4349 740 4787 870
rect 4349 736 4355 740
rect 4309 724 4355 736
rect 4781 736 4787 740
rect 4821 740 5297 870
rect 4821 736 4827 740
rect 4781 724 4827 736
rect 5291 736 5297 740
rect 5331 740 5405 870
rect 5331 736 5337 740
rect 5291 724 5337 736
rect 5399 736 5405 740
rect 5439 740 5915 870
rect 5439 736 5445 740
rect 5399 724 5445 736
rect 5909 736 5915 740
rect 5949 740 6387 870
rect 5949 736 5955 740
rect 5909 724 5955 736
rect 6381 736 6387 740
rect 6421 740 6897 870
rect 6421 736 6427 740
rect 6381 724 6427 736
rect 6891 736 6897 740
rect 6931 740 7005 870
rect 6931 736 6937 740
rect 6891 724 6937 736
rect 6999 736 7005 740
rect 7039 740 7515 870
rect 7039 736 7045 740
rect 6999 724 7045 736
rect 7509 736 7515 740
rect 7549 740 7987 870
rect 7549 736 7555 740
rect 7509 724 7555 736
rect 7981 736 7987 740
rect 8021 740 8497 870
rect 8021 736 8027 740
rect 7981 724 8027 736
rect 8491 736 8497 740
rect 8531 740 8605 870
rect 8531 736 8537 740
rect 8491 724 8537 736
rect 8599 736 8605 740
rect 8639 740 9115 870
rect 8639 736 8645 740
rect 8599 724 8645 736
rect 9109 736 9115 740
rect 9149 740 9587 870
rect 9149 736 9155 740
rect 9109 724 9155 736
rect 9581 736 9587 740
rect 9621 740 10097 870
rect 9621 736 9627 740
rect 9581 724 9627 736
rect 10091 736 10097 740
rect 10131 740 10205 870
rect 10131 736 10137 740
rect 10091 724 10137 736
rect 10199 736 10205 740
rect 10239 740 10715 870
rect 10239 736 10245 740
rect 10199 724 10245 736
rect 10709 736 10715 740
rect 10749 740 11187 870
rect 10749 736 10755 740
rect 10709 724 10755 736
rect 11181 736 11187 740
rect 11221 740 11697 870
rect 11221 736 11227 740
rect 11181 724 11227 736
rect 11420 697 11500 740
rect 11691 736 11697 740
rect 11731 740 11805 870
rect 11731 736 11737 740
rect 11691 724 11737 736
rect 11799 736 11805 740
rect 11839 740 12315 870
rect 11839 736 11845 740
rect 11799 724 11845 736
rect 12040 697 12120 740
rect 12309 736 12315 740
rect 12349 750 12390 870
rect 12510 750 12787 870
rect 12349 740 12787 750
rect 12349 736 12355 740
rect 12309 724 12355 736
rect 12781 736 12787 740
rect 12821 740 13297 870
rect 12821 736 12827 740
rect 12781 724 12827 736
rect 13020 697 13100 740
rect 13291 736 13297 740
rect 13331 740 13405 870
rect 13331 736 13337 740
rect 13291 724 13337 736
rect 13399 736 13405 740
rect 13439 740 13915 870
rect 13439 736 13445 740
rect 13399 724 13445 736
rect 13640 697 13720 740
rect 13909 736 13915 740
rect 13949 740 14387 870
rect 13949 736 13955 740
rect 13909 724 13955 736
rect 14381 736 14387 740
rect 14421 740 14897 870
rect 14421 736 14427 740
rect 14381 724 14427 736
rect 14620 697 14700 740
rect 14891 736 14897 740
rect 14931 740 15005 870
rect 14931 736 14937 740
rect 14891 724 14937 736
rect 14999 736 15005 740
rect 15039 740 15515 870
rect 15039 736 15045 740
rect 14999 724 15045 736
rect 15240 697 15320 740
rect 15509 736 15515 740
rect 15549 740 15987 870
rect 15549 736 15555 740
rect 15509 724 15555 736
rect 15981 736 15987 740
rect 16021 740 16497 870
rect 16021 736 16027 740
rect 15981 724 16027 736
rect 16491 736 16497 740
rect 16531 740 16605 870
rect 16531 736 16537 740
rect 16491 724 16537 736
rect 16599 736 16605 740
rect 16639 740 17115 870
rect 16639 736 16645 740
rect 16599 724 16645 736
rect 17109 736 17115 740
rect 17149 740 17587 870
rect 17149 736 17155 740
rect 17109 724 17155 736
rect 17581 736 17587 740
rect 17621 740 18097 870
rect 17621 736 17627 740
rect 17581 724 17627 736
rect 18091 736 18097 740
rect 18131 740 18205 870
rect 18131 736 18137 740
rect 18091 724 18137 736
rect 18199 736 18205 740
rect 18239 740 18715 870
rect 18239 736 18245 740
rect 18199 724 18245 736
rect 18709 736 18715 740
rect 18749 740 19187 870
rect 18749 736 18755 740
rect 18709 724 18755 736
rect 19181 736 19187 740
rect 19221 740 19697 870
rect 19221 736 19227 740
rect 19181 724 19227 736
rect 19691 736 19697 740
rect 19731 740 19805 870
rect 19731 736 19737 740
rect 19691 724 19737 736
rect 19799 736 19805 740
rect 19839 740 20315 870
rect 19839 736 19845 740
rect 19799 724 19845 736
rect 20309 736 20315 740
rect 20349 740 20787 870
rect 20349 736 20355 740
rect 20309 724 20355 736
rect 20781 736 20787 740
rect 20821 740 21297 870
rect 20821 736 20827 740
rect 20781 724 20827 736
rect 21291 736 21297 740
rect 21331 740 21405 870
rect 21331 736 21337 740
rect 21291 724 21337 736
rect 21399 736 21405 740
rect 21439 740 21915 870
rect 21439 736 21445 740
rect 21399 724 21445 736
rect 21909 736 21915 740
rect 21949 740 22387 870
rect 21949 736 21955 740
rect 21909 724 21955 736
rect 22381 736 22387 740
rect 22421 740 22897 870
rect 22421 736 22427 740
rect 22381 724 22427 736
rect 22891 736 22897 740
rect 22931 740 23005 870
rect 22931 736 22937 740
rect 22891 724 22937 736
rect 22999 736 23005 740
rect 23039 740 23515 870
rect 23039 736 23045 740
rect 22999 724 23045 736
rect 23509 736 23515 740
rect 23549 740 23987 870
rect 23549 736 23555 740
rect 23509 724 23555 736
rect 23981 736 23987 740
rect 24021 740 24497 870
rect 24021 736 24027 740
rect 23981 724 24027 736
rect 24491 736 24497 740
rect 24531 740 24605 870
rect 24531 736 24537 740
rect 24491 724 24537 736
rect 24599 736 24605 740
rect 24639 740 25115 870
rect 24639 736 24645 740
rect 24599 724 24645 736
rect 25109 736 25115 740
rect 25149 740 25587 870
rect 25149 736 25155 740
rect 25109 724 25155 736
rect 25581 736 25587 740
rect 25621 740 26097 870
rect 25621 736 25627 740
rect 25581 724 25627 736
rect 26091 736 26097 740
rect 26131 740 26205 870
rect 26131 736 26137 740
rect 26091 724 26137 736
rect 26199 736 26205 740
rect 26239 740 26715 870
rect 26239 736 26245 740
rect 26199 724 26245 736
rect 26709 736 26715 740
rect 26749 740 27187 870
rect 26749 736 26755 740
rect 26709 724 26755 736
rect 27181 736 27187 740
rect 27221 740 27697 870
rect 27221 736 27227 740
rect 27181 724 27227 736
rect 27691 736 27697 740
rect 27731 740 27805 870
rect 27731 736 27737 740
rect 27691 724 27737 736
rect 27799 736 27805 740
rect 27839 740 28315 870
rect 27839 736 27845 740
rect 27799 724 27845 736
rect 28309 736 28315 740
rect 28349 740 28787 870
rect 28349 736 28355 740
rect 28309 724 28355 736
rect 28781 736 28787 740
rect 28821 740 29297 870
rect 28821 736 28827 740
rect 28781 724 28827 736
rect 29291 736 29297 740
rect 29331 740 29405 870
rect 29331 736 29337 740
rect 29291 724 29337 736
rect 29399 736 29405 740
rect 29439 740 29915 870
rect 29439 736 29445 740
rect 29399 724 29445 736
rect 29909 736 29915 740
rect 29949 740 30387 870
rect 29949 736 29955 740
rect 29909 724 29955 736
rect 30381 736 30387 740
rect 30421 740 30897 870
rect 30421 736 30427 740
rect 30381 724 30427 736
rect 30891 736 30897 740
rect 30931 740 31005 870
rect 30931 736 30937 740
rect 30891 724 30937 736
rect 30999 736 31005 740
rect 31039 740 31515 870
rect 31039 736 31045 740
rect 30999 724 31045 736
rect 31509 736 31515 740
rect 31549 740 31987 870
rect 31549 736 31555 740
rect 31509 724 31555 736
rect 31981 736 31987 740
rect 32021 740 32497 870
rect 32021 736 32027 740
rect 31981 724 32027 736
rect 32491 736 32497 740
rect 32531 740 32605 870
rect 32531 736 32537 740
rect 32491 724 32537 736
rect 32599 736 32605 740
rect 32639 740 33115 870
rect 32639 736 32645 740
rect 32599 724 32645 736
rect 33109 736 33115 740
rect 33149 740 33587 870
rect 33149 736 33155 740
rect 33109 724 33155 736
rect 33581 736 33587 740
rect 33621 740 34097 870
rect 33621 736 33627 740
rect 33581 724 33627 736
rect 34091 736 34097 740
rect 34131 740 34205 870
rect 34131 736 34137 740
rect 34091 724 34137 736
rect 34199 736 34205 740
rect 34239 740 34715 870
rect 34239 736 34245 740
rect 34199 724 34245 736
rect 34709 736 34715 740
rect 34749 740 35187 870
rect 34749 736 34755 740
rect 34709 724 34755 736
rect 35181 736 35187 740
rect 35221 740 35697 870
rect 35221 736 35227 740
rect 35181 724 35227 736
rect 35691 736 35697 740
rect 35731 740 35805 870
rect 35731 736 35737 740
rect 35691 724 35737 736
rect 35799 736 35805 740
rect 35839 740 36315 870
rect 35839 736 35845 740
rect 35799 724 35845 736
rect 36309 736 36315 740
rect 36349 740 36787 870
rect 36349 736 36355 740
rect 36309 724 36355 736
rect 36781 736 36787 740
rect 36821 740 37297 870
rect 36821 736 36827 740
rect 36781 724 36827 736
rect 37291 736 37297 740
rect 37331 740 37405 870
rect 37331 736 37337 740
rect 37291 724 37337 736
rect 37399 736 37405 740
rect 37439 740 37915 870
rect 37439 736 37445 740
rect 37399 724 37445 736
rect 37909 736 37915 740
rect 37949 736 37955 870
rect 37909 724 37955 736
rect 660 691 1077 697
rect 660 657 689 691
rect 1065 657 1077 691
rect 1659 691 2059 697
rect 660 651 1077 657
rect 1180 680 1320 690
rect 1659 680 1671 691
rect 660 460 710 651
rect 1180 560 1190 680
rect 1310 657 1671 680
rect 2047 680 2059 691
rect 2277 691 2677 697
rect 2277 680 2289 691
rect 2047 657 2289 680
rect 2665 680 2677 691
rect 3259 691 3659 697
rect 2780 680 2920 690
rect 3259 680 3271 691
rect 2665 657 2790 680
rect 1310 560 2790 657
rect 2910 657 3271 680
rect 3647 680 3659 691
rect 3877 691 4277 697
rect 3877 680 3889 691
rect 3647 657 3889 680
rect 4265 680 4277 691
rect 4859 691 5259 697
rect 4380 680 4520 690
rect 4859 680 4871 691
rect 4265 657 4390 680
rect 2910 560 4390 657
rect 4510 657 4871 680
rect 5247 680 5259 691
rect 5477 691 5877 697
rect 5477 680 5489 691
rect 5247 657 5489 680
rect 5865 680 5877 691
rect 6459 691 6859 697
rect 5980 680 6120 690
rect 6459 680 6471 691
rect 5865 657 5990 680
rect 4510 560 5990 657
rect 6110 657 6471 680
rect 6847 680 6859 691
rect 7077 691 7477 697
rect 7077 680 7089 691
rect 6847 657 7089 680
rect 7465 680 7477 691
rect 8059 691 8459 697
rect 7580 680 7720 690
rect 8059 680 8071 691
rect 7465 657 7590 680
rect 6110 560 7590 657
rect 7710 657 8071 680
rect 8447 680 8459 691
rect 8677 691 9077 697
rect 8677 680 8689 691
rect 8447 657 8689 680
rect 9065 680 9077 691
rect 9659 691 10059 697
rect 9180 680 9320 690
rect 9659 680 9671 691
rect 9065 657 9190 680
rect 7710 560 9190 657
rect 9310 657 9671 680
rect 10047 680 10059 691
rect 10277 691 10677 697
rect 10277 680 10289 691
rect 10047 657 10289 680
rect 10665 680 10677 691
rect 11259 691 11659 697
rect 10665 657 10720 680
rect 9310 560 10720 657
rect 11259 657 11271 691
rect 11647 657 11659 691
rect 11259 651 11659 657
rect 11877 691 12277 697
rect 11877 657 11889 691
rect 12265 657 12277 691
rect 11877 651 12277 657
rect 12859 691 13259 697
rect 12859 657 12871 691
rect 13247 657 13259 691
rect 12859 651 13259 657
rect 13477 691 13877 697
rect 13477 657 13489 691
rect 13865 657 13877 691
rect 13477 651 13877 657
rect 14459 691 14859 697
rect 14459 657 14471 691
rect 14847 657 14859 691
rect 14459 651 14859 657
rect 15077 691 15477 697
rect 15077 657 15089 691
rect 15465 657 15477 691
rect 16059 691 16459 697
rect 15077 651 15477 657
rect 15810 680 15930 690
rect 16059 680 16071 691
rect 15810 560 15820 680
rect 15920 657 16071 680
rect 16447 680 16459 691
rect 16677 691 17077 697
rect 16677 680 16689 691
rect 16447 657 16689 680
rect 17065 680 17077 691
rect 17659 691 18059 697
rect 17410 680 17530 690
rect 17659 680 17671 691
rect 17065 657 17120 680
rect 15920 560 17120 657
rect 17410 560 17420 680
rect 17520 657 17671 680
rect 18047 680 18059 691
rect 18277 691 18677 697
rect 18277 680 18289 691
rect 18047 657 18289 680
rect 18665 680 18677 691
rect 19259 691 19659 697
rect 19010 680 19130 690
rect 19259 680 19271 691
rect 18665 657 18720 680
rect 17520 560 18720 657
rect 19010 560 19020 680
rect 19120 657 19271 680
rect 19647 680 19659 691
rect 19877 691 20277 697
rect 19877 680 19889 691
rect 19647 657 19889 680
rect 20265 680 20277 691
rect 20859 691 21259 697
rect 20610 680 20730 690
rect 20859 680 20871 691
rect 20265 657 20320 680
rect 19120 560 20320 657
rect 20610 560 20620 680
rect 20720 657 20871 680
rect 21247 680 21259 691
rect 21477 691 21877 697
rect 21477 680 21489 691
rect 21247 657 21489 680
rect 21865 680 21877 691
rect 22459 691 22859 697
rect 22210 680 22330 690
rect 22459 680 22471 691
rect 21865 657 21920 680
rect 20720 560 21920 657
rect 22210 560 22220 680
rect 22320 657 22471 680
rect 22847 680 22859 691
rect 23077 691 23477 697
rect 23077 680 23089 691
rect 22847 657 23089 680
rect 23465 680 23477 691
rect 24059 691 24459 697
rect 23810 680 23930 690
rect 24059 680 24071 691
rect 23465 657 23520 680
rect 22320 560 23520 657
rect 23810 560 23820 680
rect 23920 657 24071 680
rect 24447 680 24459 691
rect 24677 691 25077 697
rect 24677 680 24689 691
rect 24447 657 24689 680
rect 25065 680 25077 691
rect 25659 691 26059 697
rect 25659 680 25671 691
rect 25065 657 25120 680
rect 23920 560 25120 657
rect 25620 657 25671 680
rect 26047 680 26059 691
rect 26277 691 26677 697
rect 26277 680 26289 691
rect 26047 657 26289 680
rect 26665 680 26677 691
rect 27259 691 27659 697
rect 27010 680 27130 690
rect 27259 680 27271 691
rect 26665 657 27020 680
rect 25620 560 27020 657
rect 27120 657 27271 680
rect 27647 680 27659 691
rect 27877 691 28277 697
rect 27877 680 27889 691
rect 27647 657 27889 680
rect 28265 680 28277 691
rect 28859 691 29259 697
rect 28859 690 28871 691
rect 28610 680 28871 690
rect 28265 657 28320 680
rect 27120 560 28320 657
rect 28610 560 28620 680
rect 28720 657 28871 680
rect 29247 690 29259 691
rect 29477 691 29877 697
rect 29477 690 29489 691
rect 29247 657 29489 690
rect 29865 690 29877 691
rect 30459 691 30859 697
rect 30459 690 30471 691
rect 29865 657 30471 690
rect 30847 690 30859 691
rect 31077 691 31477 697
rect 31077 690 31089 691
rect 30847 657 31089 690
rect 31465 690 31477 691
rect 32059 691 32459 697
rect 31465 657 31520 690
rect 28720 560 31520 657
rect 1180 550 1320 560
rect 2780 550 2920 560
rect 4380 550 4520 560
rect 5980 550 6120 560
rect 7580 550 7720 560
rect 9180 550 9320 560
rect 15810 550 15930 560
rect 17410 550 17530 560
rect 19010 550 19130 560
rect 20610 550 20730 560
rect 22210 550 22330 560
rect 23810 550 23930 560
rect 27010 550 27130 560
rect 28610 550 31520 560
rect 31810 680 31930 690
rect 32059 680 32071 691
rect 31810 560 31820 680
rect 31920 657 32071 680
rect 32447 680 32459 691
rect 32677 691 33077 697
rect 32677 680 32689 691
rect 32447 657 32689 680
rect 33065 680 33077 691
rect 33659 691 34059 697
rect 33659 680 33671 691
rect 33065 657 33671 680
rect 34047 680 34059 691
rect 34277 691 34677 697
rect 34277 680 34289 691
rect 34047 657 34289 680
rect 34665 680 34677 691
rect 35259 691 35659 697
rect 35259 680 35271 691
rect 34665 657 35271 680
rect 35647 680 35659 691
rect 35877 691 36277 697
rect 35877 680 35889 691
rect 35647 657 35889 680
rect 36265 657 36277 691
rect 36859 691 37259 697
rect 31920 651 36277 657
rect 36590 670 36730 680
rect 31920 560 36270 651
rect 31810 550 31930 560
rect 36590 550 36600 670
rect 36720 660 36730 670
rect 36859 660 36871 691
rect 36720 657 36871 660
rect 37247 657 37259 691
rect 36720 651 37259 657
rect 37477 691 37877 697
rect 37477 657 37489 691
rect 37865 660 37877 691
rect 37865 657 37980 660
rect 37477 651 37980 657
rect 36720 560 37252 651
rect 37480 650 37980 651
rect 37480 560 37850 650
rect 36720 550 36730 560
rect 36590 540 36730 550
rect 37840 530 37850 560
rect 37970 530 37980 650
rect 37840 520 37980 530
rect 660 435 38060 460
rect 660 429 38065 435
rect -140 395 -117 429
rect 1253 395 1483 429
rect 2853 395 3083 429
rect 4453 395 4683 429
rect 6053 395 6283 429
rect 7653 395 7883 429
rect 9253 395 9483 429
rect 10853 395 11083 429
rect 12453 395 12683 429
rect 14053 395 14283 429
rect 15653 395 15883 429
rect 17253 395 17483 429
rect 18853 395 19083 429
rect 20453 395 20683 429
rect 22053 395 22283 429
rect 23653 395 23883 429
rect 25253 395 25483 429
rect 26853 395 27083 429
rect 28453 395 28683 429
rect 30053 395 30283 429
rect 31653 395 31883 429
rect 33253 395 33483 429
rect 34853 395 35083 429
rect 36453 395 36683 429
rect 38053 395 38065 429
rect -140 295 480 395
rect -140 261 71 295
rect 447 261 480 295
rect -140 260 480 261
rect -140 207 0 260
rect 59 255 480 260
rect -140 195 27 207
rect -140 -497 -13 195
rect 21 -497 27 195
rect -140 -509 27 -497
rect -140 -918 0 -509
rect 440 -557 480 255
rect 660 389 38065 395
rect 660 295 38060 389
rect 660 261 689 295
rect 1065 261 1671 295
rect 2047 261 2289 295
rect 2665 261 3271 295
rect 3647 261 3889 295
rect 4265 261 4871 295
rect 5247 261 5489 295
rect 5865 261 6471 295
rect 6847 261 7089 295
rect 7465 261 8071 295
rect 8447 261 8689 295
rect 9065 261 9671 295
rect 10047 261 10289 295
rect 10665 261 11271 295
rect 11647 261 11889 295
rect 12265 261 12871 295
rect 13247 261 13489 295
rect 13865 261 14471 295
rect 14847 261 15089 295
rect 15465 261 16071 295
rect 16447 261 16689 295
rect 17065 261 17671 295
rect 18047 261 18289 295
rect 18665 261 19271 295
rect 19647 261 19889 295
rect 20265 261 20871 295
rect 21247 261 21489 295
rect 21865 261 22471 295
rect 22847 261 23089 295
rect 23465 261 24071 295
rect 24447 261 24689 295
rect 25065 261 25671 295
rect 26047 261 26289 295
rect 26665 261 27271 295
rect 27647 261 27889 295
rect 28265 261 28871 295
rect 29247 261 29489 295
rect 29865 261 30471 295
rect 30847 261 31089 295
rect 31465 261 32071 295
rect 32447 261 32689 295
rect 33065 261 33671 295
rect 34047 261 34289 295
rect 34665 261 35271 295
rect 35647 261 35889 295
rect 36265 261 36871 295
rect 37247 261 37489 295
rect 37865 261 38060 295
rect 660 260 38060 261
rect 660 255 1077 260
rect 1659 255 2059 260
rect 2277 255 2677 260
rect 3259 255 3659 260
rect 3877 255 4277 260
rect 4859 255 5259 260
rect 5477 255 5877 260
rect 6459 255 6859 260
rect 7077 255 7477 260
rect 8059 255 8459 260
rect 8677 255 9077 260
rect 9659 255 10059 260
rect 10277 255 10677 260
rect 11259 255 11659 260
rect 11877 255 12277 260
rect 12859 255 13259 260
rect 13477 255 13877 260
rect 14459 255 14859 260
rect 15077 255 15477 260
rect 16059 255 16459 260
rect 16677 255 17077 260
rect 17659 255 18059 260
rect 18277 255 18677 260
rect 19259 255 19659 260
rect 19877 255 20277 260
rect 20859 255 21259 260
rect 21477 255 21877 260
rect 22459 255 22859 260
rect 23077 255 23477 260
rect 24059 255 24459 260
rect 24677 255 25077 260
rect 25659 255 26059 260
rect 26277 255 26677 260
rect 27259 255 27659 260
rect 27877 255 28277 260
rect 28859 255 29259 260
rect 29477 255 29877 260
rect 30459 255 30859 260
rect 31077 255 31477 260
rect 32059 255 32459 260
rect 32677 255 33077 260
rect 33659 255 34059 260
rect 34277 255 34677 260
rect 35259 255 35659 260
rect 35877 255 36277 260
rect 59 -563 480 -557
rect 59 -597 71 -563
rect 447 -597 480 -563
rect 59 -603 480 -597
rect 440 -845 480 -603
rect 59 -851 480 -845
rect 59 -885 71 -851
rect 447 -885 480 -851
rect 59 -891 480 -885
rect -140 -930 27 -918
rect -140 -1064 -13 -930
rect 21 -1064 27 -930
rect -140 -1076 27 -1064
rect -140 -1340 0 -1076
rect 440 -1103 480 -891
rect 660 -557 710 255
rect 36660 207 36800 260
rect 36859 255 37259 260
rect 37300 207 37440 260
rect 37477 255 37877 260
rect 37920 207 38060 260
rect 1109 195 1155 207
rect 1109 -497 1115 195
rect 1149 -497 1155 195
rect 1109 -509 1155 -497
rect 1581 195 1627 207
rect 1581 -497 1587 195
rect 1621 -497 1627 195
rect 1581 -509 1627 -497
rect 2091 200 2137 207
rect 2199 200 2245 207
rect 2091 195 2245 200
rect 2091 -497 2097 195
rect 2131 190 2205 195
rect 2131 -497 2205 -490
rect 2239 -497 2245 195
rect 2091 -500 2245 -497
rect 2091 -509 2137 -500
rect 2199 -509 2245 -500
rect 2709 195 2755 207
rect 2709 -497 2715 195
rect 2749 -497 2755 195
rect 2709 -509 2755 -497
rect 3181 195 3227 207
rect 3181 -497 3187 195
rect 3221 -497 3227 195
rect 3181 -509 3227 -497
rect 3691 200 3737 207
rect 3799 200 3845 207
rect 3691 195 3845 200
rect 3691 -497 3697 195
rect 3731 190 3805 195
rect 3731 -497 3805 -490
rect 3839 -497 3845 195
rect 3691 -500 3845 -497
rect 3691 -509 3737 -500
rect 3799 -509 3845 -500
rect 4309 195 4355 207
rect 4309 -497 4315 195
rect 4349 -497 4355 195
rect 4309 -509 4355 -497
rect 4781 195 4827 207
rect 4781 -497 4787 195
rect 4821 -497 4827 195
rect 4781 -509 4827 -497
rect 5291 200 5337 207
rect 5399 200 5445 207
rect 5291 195 5445 200
rect 5291 -497 5297 195
rect 5331 190 5405 195
rect 5331 -497 5405 -490
rect 5439 -497 5445 195
rect 5291 -500 5445 -497
rect 5291 -509 5337 -500
rect 5399 -509 5445 -500
rect 5909 195 5955 207
rect 5909 -497 5915 195
rect 5949 -497 5955 195
rect 5909 -509 5955 -497
rect 6381 195 6427 207
rect 6381 -497 6387 195
rect 6421 -497 6427 195
rect 6381 -509 6427 -497
rect 6891 200 6937 207
rect 6999 200 7045 207
rect 6891 195 7045 200
rect 6891 -497 6897 195
rect 6931 190 7005 195
rect 6931 -497 7005 -490
rect 7039 -497 7045 195
rect 6891 -500 7045 -497
rect 6891 -509 6937 -500
rect 6999 -509 7045 -500
rect 7509 195 7555 207
rect 7509 -497 7515 195
rect 7549 -497 7555 195
rect 7509 -509 7555 -497
rect 7981 195 8027 207
rect 7981 -497 7987 195
rect 8021 -497 8027 195
rect 7981 -509 8027 -497
rect 8491 200 8537 207
rect 8599 200 8645 207
rect 8491 195 8645 200
rect 8491 -497 8497 195
rect 8531 190 8605 195
rect 8531 -497 8605 -490
rect 8639 -497 8645 195
rect 8491 -500 8645 -497
rect 8491 -509 8537 -500
rect 8599 -509 8645 -500
rect 9109 195 9155 207
rect 9109 -497 9115 195
rect 9149 -497 9155 195
rect 9109 -509 9155 -497
rect 9581 195 9627 207
rect 9581 -497 9587 195
rect 9621 -497 9627 195
rect 9581 -509 9627 -497
rect 10091 200 10137 207
rect 10199 200 10245 207
rect 10091 195 10245 200
rect 10091 -497 10097 195
rect 10131 190 10205 195
rect 10131 -497 10205 -490
rect 10239 -497 10245 195
rect 10091 -500 10245 -497
rect 10091 -509 10137 -500
rect 10199 -509 10245 -500
rect 10709 195 10755 207
rect 10709 -497 10715 195
rect 10749 -497 10755 195
rect 10709 -509 10755 -497
rect 11181 195 11227 207
rect 11181 -497 11187 195
rect 11221 -497 11227 195
rect 11181 -509 11227 -497
rect 11691 200 11737 207
rect 11799 200 11845 207
rect 11691 195 11845 200
rect 11691 -497 11697 195
rect 11731 190 11805 195
rect 11839 -497 11845 195
rect 11691 -509 11710 -497
rect 660 -563 1077 -557
rect 660 -597 689 -563
rect 1065 -597 1077 -563
rect 660 -603 1077 -597
rect 1659 -563 2059 -557
rect 1659 -597 1671 -563
rect 2047 -597 2059 -563
rect 1659 -603 2059 -597
rect 2277 -563 2677 -557
rect 2277 -597 2289 -563
rect 2665 -597 2677 -563
rect 2277 -603 2677 -597
rect 3259 -563 3659 -557
rect 3259 -597 3271 -563
rect 3647 -597 3659 -563
rect 3259 -603 3659 -597
rect 3877 -563 4277 -557
rect 3877 -597 3889 -563
rect 4265 -597 4277 -563
rect 3877 -603 4277 -597
rect 4859 -563 5259 -557
rect 4859 -597 4871 -563
rect 5247 -597 5259 -563
rect 4859 -603 5259 -597
rect 5477 -563 5877 -557
rect 5477 -597 5489 -563
rect 5865 -597 5877 -563
rect 5477 -603 5877 -597
rect 6459 -563 6859 -557
rect 6459 -597 6471 -563
rect 6847 -597 6859 -563
rect 6459 -603 6859 -597
rect 7077 -563 7477 -557
rect 7077 -597 7089 -563
rect 7465 -597 7477 -563
rect 7077 -603 7477 -597
rect 8059 -563 8459 -557
rect 8059 -597 8071 -563
rect 8447 -597 8459 -563
rect 8059 -603 8459 -597
rect 8677 -563 9077 -557
rect 8677 -597 8689 -563
rect 9065 -597 9077 -563
rect 8677 -603 9077 -597
rect 9659 -563 10059 -557
rect 9659 -597 9671 -563
rect 10047 -597 10059 -563
rect 9659 -603 10059 -597
rect 10277 -563 10677 -557
rect 10277 -597 10289 -563
rect 10665 -597 10677 -563
rect 10277 -603 10677 -597
rect 11259 -560 11659 -557
rect 11700 -560 11710 -509
rect 11259 -563 11710 -560
rect 11259 -570 11271 -563
rect 11647 -570 11710 -563
rect 11830 -509 11845 -497
rect 12309 195 12355 207
rect 12309 -497 12315 195
rect 12349 -497 12355 195
rect 12309 -509 12355 -497
rect 12781 195 12827 207
rect 12781 -497 12787 195
rect 12821 -497 12827 195
rect 12781 -509 12827 -497
rect 13291 200 13337 207
rect 13399 200 13445 207
rect 13291 195 13445 200
rect 13291 -497 13297 195
rect 13331 190 13405 195
rect 13331 -497 13405 -490
rect 13439 -497 13445 195
rect 13291 -500 13445 -497
rect 13291 -509 13337 -500
rect 13399 -509 13445 -500
rect 13909 195 13955 207
rect 13909 -497 13915 195
rect 13949 -497 13955 195
rect 14381 195 14427 207
rect 14381 -490 14387 195
rect 13909 -509 13955 -497
rect 14380 -497 14387 -490
rect 14421 -490 14427 195
rect 14891 200 14937 207
rect 14999 200 15045 207
rect 14891 195 15045 200
rect 14421 -497 14430 -490
rect 11830 -560 11840 -509
rect 11877 -560 12277 -557
rect 11830 -563 12280 -560
rect 11830 -570 11889 -563
rect 12265 -570 12280 -563
rect 11259 -603 11270 -570
rect 660 -845 710 -603
rect 1680 -640 2040 -603
rect 2300 -640 2660 -603
rect 3280 -640 3640 -603
rect 3900 -640 4260 -603
rect 4880 -640 5240 -603
rect 5500 -640 5860 -603
rect 6480 -640 6840 -603
rect 7100 -640 7460 -603
rect 8080 -640 8440 -603
rect 8700 -640 9060 -603
rect 9680 -640 10040 -603
rect 10300 -640 10660 -603
rect 1400 -650 10660 -640
rect 1400 -770 1410 -650
rect 1530 -770 3010 -650
rect 3130 -770 4610 -650
rect 4730 -770 6210 -650
rect 6330 -770 7810 -650
rect 7930 -770 9410 -650
rect 9530 -770 10660 -650
rect 11260 -730 11270 -603
rect 12270 -730 12280 -570
rect 12859 -563 13259 -557
rect 12859 -597 12871 -563
rect 13247 -597 13259 -563
rect 12859 -603 13259 -597
rect 13477 -563 13877 -557
rect 13477 -597 13489 -563
rect 13865 -597 13877 -563
rect 13477 -603 13877 -597
rect 14380 -560 14430 -497
rect 14891 -497 14897 195
rect 14931 190 15005 195
rect 15039 -497 15045 195
rect 14891 -509 14910 -497
rect 14459 -560 14859 -557
rect 14900 -560 14910 -509
rect 14380 -563 14910 -560
rect 14380 -570 14471 -563
rect 14847 -570 14910 -563
rect 15030 -509 15045 -497
rect 15509 195 15555 207
rect 15509 -497 15515 195
rect 15549 -490 15555 195
rect 15981 195 16027 207
rect 15549 -497 15560 -490
rect 15509 -509 15560 -497
rect 15981 -497 15987 195
rect 16021 -497 16027 195
rect 15981 -509 16027 -497
rect 16491 200 16537 207
rect 16599 200 16645 207
rect 16491 195 16645 200
rect 16491 -497 16497 195
rect 16531 190 16605 195
rect 16531 -497 16605 -490
rect 16639 -497 16645 195
rect 16491 -500 16645 -497
rect 16491 -509 16537 -500
rect 16599 -509 16645 -500
rect 17109 195 17155 207
rect 17109 -497 17115 195
rect 17149 -497 17155 195
rect 17109 -509 17155 -497
rect 17581 195 17627 207
rect 17581 -497 17587 195
rect 17621 -497 17627 195
rect 17581 -509 17627 -497
rect 18091 200 18137 207
rect 18199 200 18245 207
rect 18091 195 18245 200
rect 18091 -497 18097 195
rect 18131 190 18205 195
rect 18131 -497 18205 -490
rect 18239 -497 18245 195
rect 18091 -500 18245 -497
rect 18091 -509 18137 -500
rect 18199 -509 18245 -500
rect 18709 195 18755 207
rect 18709 -497 18715 195
rect 18749 -497 18755 195
rect 18709 -509 18755 -497
rect 19181 195 19227 207
rect 19181 -497 19187 195
rect 19221 -497 19227 195
rect 19181 -509 19227 -497
rect 19691 200 19737 207
rect 19799 200 19845 207
rect 19691 195 19845 200
rect 19691 -497 19697 195
rect 19731 190 19805 195
rect 19731 -497 19805 -490
rect 19839 -497 19845 195
rect 19691 -500 19845 -497
rect 19691 -509 19737 -500
rect 19799 -509 19845 -500
rect 20309 195 20355 207
rect 20309 -497 20315 195
rect 20349 -497 20355 195
rect 20309 -509 20355 -497
rect 20781 195 20827 207
rect 20781 -497 20787 195
rect 20821 -497 20827 195
rect 20781 -509 20827 -497
rect 21291 200 21337 207
rect 21399 200 21445 207
rect 21291 195 21445 200
rect 21291 -497 21297 195
rect 21331 190 21405 195
rect 21331 -497 21405 -490
rect 21439 -497 21445 195
rect 21291 -500 21445 -497
rect 21291 -509 21337 -500
rect 21399 -509 21445 -500
rect 21909 195 21955 207
rect 21909 -497 21915 195
rect 21949 -497 21955 195
rect 21909 -509 21955 -497
rect 22381 195 22427 207
rect 22381 -497 22387 195
rect 22421 -497 22427 195
rect 22381 -509 22427 -497
rect 22891 200 22937 207
rect 22999 200 23045 207
rect 22891 195 23045 200
rect 22891 -497 22897 195
rect 22931 190 23005 195
rect 22931 -497 23005 -490
rect 23039 -497 23045 195
rect 22891 -500 23045 -497
rect 22891 -509 22937 -500
rect 22999 -509 23045 -500
rect 23509 195 23555 207
rect 23509 -497 23515 195
rect 23549 -497 23555 195
rect 23509 -509 23555 -497
rect 23981 195 24027 207
rect 23981 -497 23987 195
rect 24021 -497 24027 195
rect 23981 -509 24027 -497
rect 24491 200 24537 207
rect 24599 200 24645 207
rect 24491 195 24645 200
rect 24491 -497 24497 195
rect 24531 190 24605 195
rect 24531 -497 24605 -490
rect 24639 -497 24645 195
rect 24491 -500 24645 -497
rect 24491 -509 24537 -500
rect 24599 -509 24645 -500
rect 25109 195 25155 207
rect 25109 -497 25115 195
rect 25149 -497 25155 195
rect 25109 -509 25155 -497
rect 25581 195 25627 207
rect 25581 -497 25587 195
rect 25621 -497 25627 195
rect 25581 -509 25627 -497
rect 26091 200 26137 207
rect 26199 200 26245 207
rect 26091 195 26245 200
rect 26091 -497 26097 195
rect 26131 190 26205 195
rect 26131 -497 26205 -490
rect 26239 -497 26245 195
rect 26091 -500 26245 -497
rect 26091 -509 26137 -500
rect 26199 -509 26245 -500
rect 26709 195 26755 207
rect 26709 -497 26715 195
rect 26749 -497 26755 195
rect 26709 -509 26755 -497
rect 27181 195 27227 207
rect 27181 -497 27187 195
rect 27221 -497 27227 195
rect 27181 -509 27227 -497
rect 27691 200 27737 207
rect 27799 200 27845 207
rect 27691 195 27845 200
rect 27691 -497 27697 195
rect 27731 190 27805 195
rect 27731 -497 27805 -490
rect 27839 -497 27845 195
rect 27691 -500 27845 -497
rect 27691 -509 27737 -500
rect 27799 -509 27845 -500
rect 28309 195 28355 207
rect 28309 -497 28315 195
rect 28349 -497 28355 195
rect 28309 -509 28355 -497
rect 28781 195 28827 207
rect 28781 -497 28787 195
rect 28821 -497 28827 195
rect 28781 -509 28827 -497
rect 29291 200 29337 207
rect 29399 200 29445 207
rect 29291 195 29445 200
rect 29291 -497 29297 195
rect 29331 190 29405 195
rect 29331 -497 29405 -490
rect 29439 -497 29445 195
rect 29291 -500 29445 -497
rect 29291 -509 29337 -500
rect 29399 -509 29445 -500
rect 29909 195 29955 207
rect 29909 -497 29915 195
rect 29949 -497 29955 195
rect 29909 -509 29955 -497
rect 30381 195 30427 207
rect 30381 -497 30387 195
rect 30421 -497 30427 195
rect 30381 -509 30427 -497
rect 30891 200 30937 207
rect 30999 200 31045 207
rect 30891 195 31045 200
rect 30891 -497 30897 195
rect 30931 190 31005 195
rect 30931 -497 31005 -490
rect 31039 -497 31045 195
rect 30891 -500 31045 -497
rect 30891 -509 30937 -500
rect 30999 -509 31045 -500
rect 31509 195 31555 207
rect 31509 -497 31515 195
rect 31549 -497 31555 195
rect 31509 -509 31555 -497
rect 31981 195 32027 207
rect 31981 -497 31987 195
rect 32021 -497 32027 195
rect 31981 -509 32027 -497
rect 32491 200 32537 207
rect 32599 200 32645 207
rect 32491 195 32645 200
rect 32491 -497 32497 195
rect 32531 190 32605 195
rect 32531 -497 32605 -490
rect 32639 -497 32645 195
rect 32491 -500 32645 -497
rect 32491 -509 32537 -500
rect 32599 -509 32645 -500
rect 33109 195 33155 207
rect 33109 -497 33115 195
rect 33149 -497 33155 195
rect 33109 -509 33155 -497
rect 33581 195 33627 207
rect 33581 -497 33587 195
rect 33621 -497 33627 195
rect 33581 -509 33627 -497
rect 34091 200 34137 207
rect 34199 200 34245 207
rect 34091 195 34245 200
rect 34091 -497 34097 195
rect 34131 190 34205 195
rect 34131 -497 34205 -490
rect 34239 -497 34245 195
rect 34091 -500 34245 -497
rect 34091 -509 34137 -500
rect 34199 -509 34245 -500
rect 34709 195 34755 207
rect 34709 -497 34715 195
rect 34749 -497 34755 195
rect 34709 -509 34755 -497
rect 35181 195 35227 207
rect 35181 -497 35187 195
rect 35221 -497 35227 195
rect 35181 -509 35227 -497
rect 35691 200 35737 207
rect 35799 200 35845 207
rect 35691 195 35845 200
rect 35691 -497 35697 195
rect 35731 190 35805 195
rect 35731 -497 35805 -490
rect 35839 -497 35845 195
rect 35691 -500 35845 -497
rect 35691 -509 35737 -500
rect 35799 -509 35845 -500
rect 36309 195 36355 207
rect 36309 -497 36315 195
rect 36349 -497 36355 195
rect 36309 -509 36355 -497
rect 36660 195 36827 207
rect 36660 -497 36787 195
rect 36821 -497 36827 195
rect 36660 -509 36827 -497
rect 37291 195 37445 207
rect 37291 -497 37297 195
rect 37331 -497 37405 195
rect 37439 -497 37445 195
rect 37291 -509 37445 -497
rect 37909 195 38060 207
rect 37909 -497 37915 195
rect 37949 -497 38060 195
rect 37909 -509 38060 -497
rect 15030 -560 15040 -509
rect 15077 -560 15477 -557
rect 15510 -560 15560 -509
rect 15030 -563 15560 -560
rect 15030 -570 15089 -563
rect 15465 -570 15560 -563
rect 12880 -640 13240 -603
rect 13500 -640 13860 -603
rect 11260 -740 12280 -730
rect 12380 -650 14300 -640
rect 1400 -780 10660 -770
rect 1680 -845 2040 -780
rect 2300 -845 2660 -780
rect 3280 -845 3640 -780
rect 3900 -845 4260 -780
rect 4880 -845 5240 -780
rect 5500 -845 5860 -780
rect 6480 -845 6840 -780
rect 7100 -845 7460 -780
rect 8080 -845 8440 -780
rect 8700 -845 9060 -780
rect 9680 -845 10040 -780
rect 10300 -845 10660 -780
rect 12380 -810 12390 -650
rect 12510 -780 14300 -650
rect 14380 -730 14470 -570
rect 15470 -730 15560 -570
rect 16059 -563 16459 -557
rect 16059 -597 16071 -563
rect 16447 -597 16459 -563
rect 16059 -603 16459 -597
rect 16677 -563 17077 -557
rect 16677 -597 16689 -563
rect 17065 -597 17077 -563
rect 16677 -603 17077 -597
rect 17659 -563 18059 -557
rect 17659 -597 17671 -563
rect 18047 -597 18059 -563
rect 17659 -603 18059 -597
rect 18277 -563 18677 -557
rect 18277 -597 18289 -563
rect 18665 -597 18677 -563
rect 18277 -603 18677 -597
rect 19259 -563 19659 -557
rect 19259 -597 19271 -563
rect 19647 -597 19659 -563
rect 19259 -603 19659 -597
rect 19877 -563 20277 -557
rect 19877 -597 19889 -563
rect 20265 -597 20277 -563
rect 19877 -603 20277 -597
rect 20859 -563 21259 -557
rect 20859 -597 20871 -563
rect 21247 -597 21259 -563
rect 20859 -603 21259 -597
rect 21477 -563 21877 -557
rect 21477 -597 21489 -563
rect 21865 -597 21877 -563
rect 21477 -603 21877 -597
rect 22459 -563 22859 -557
rect 22459 -597 22471 -563
rect 22847 -597 22859 -563
rect 22459 -603 22859 -597
rect 23077 -563 23477 -557
rect 23077 -597 23089 -563
rect 23465 -597 23477 -563
rect 23077 -603 23477 -597
rect 24059 -563 24459 -557
rect 24059 -597 24071 -563
rect 24447 -597 24459 -563
rect 24059 -603 24459 -597
rect 24677 -563 25077 -557
rect 24677 -597 24689 -563
rect 25065 -597 25077 -563
rect 24677 -603 25077 -597
rect 25659 -563 26059 -557
rect 25659 -597 25671 -563
rect 26047 -597 26059 -563
rect 25659 -603 26059 -597
rect 26277 -563 26677 -557
rect 26277 -597 26289 -563
rect 26665 -597 26677 -563
rect 26277 -603 26677 -597
rect 27259 -563 27659 -557
rect 27259 -597 27271 -563
rect 27647 -597 27659 -563
rect 27259 -603 27659 -597
rect 27877 -563 28277 -557
rect 27877 -597 27889 -563
rect 28265 -597 28277 -563
rect 27877 -603 28277 -597
rect 28859 -563 29259 -557
rect 28859 -597 28871 -563
rect 29247 -597 29259 -563
rect 28859 -603 29259 -597
rect 29477 -563 29877 -557
rect 29477 -597 29489 -563
rect 29865 -597 29877 -563
rect 29477 -603 29877 -597
rect 30459 -563 30859 -557
rect 30459 -597 30471 -563
rect 30847 -597 30859 -563
rect 30459 -603 30859 -597
rect 31077 -563 31477 -557
rect 31077 -597 31089 -563
rect 31465 -597 31477 -563
rect 31077 -603 31477 -597
rect 32059 -563 32459 -557
rect 32059 -597 32071 -563
rect 32447 -597 32459 -563
rect 32059 -603 32459 -597
rect 32677 -563 33077 -557
rect 32677 -597 32689 -563
rect 33065 -597 33077 -563
rect 32677 -603 33077 -597
rect 33659 -563 34059 -557
rect 33659 -597 33671 -563
rect 34047 -597 34059 -563
rect 33659 -603 34059 -597
rect 34277 -563 34677 -557
rect 34277 -597 34289 -563
rect 34665 -597 34677 -563
rect 34277 -603 34677 -597
rect 35259 -563 35659 -557
rect 35259 -597 35271 -563
rect 35647 -597 35659 -563
rect 35259 -603 35659 -597
rect 35877 -563 36277 -557
rect 35877 -597 35889 -563
rect 36265 -597 36277 -563
rect 35877 -603 36277 -597
rect 16080 -640 16440 -603
rect 16700 -640 17060 -603
rect 17680 -640 18040 -603
rect 18300 -640 18660 -603
rect 19280 -640 19640 -603
rect 19900 -640 20260 -603
rect 20880 -640 21240 -603
rect 21500 -640 21860 -603
rect 22480 -640 22840 -603
rect 23100 -640 23460 -603
rect 24080 -640 24440 -603
rect 24700 -640 25060 -603
rect 25680 -640 26040 -603
rect 26300 -640 26660 -603
rect 27280 -640 27640 -603
rect 27900 -640 28260 -603
rect 28880 -640 29240 -603
rect 29500 -640 29860 -603
rect 30480 -640 30840 -603
rect 31100 -640 31460 -603
rect 32080 -640 32440 -603
rect 32700 -640 33060 -603
rect 33680 -640 34040 -603
rect 34300 -640 34660 -603
rect 35280 -640 35640 -603
rect 35900 -640 36260 -603
rect 14380 -740 15560 -730
rect 15590 -650 17060 -640
rect 15590 -770 15600 -650
rect 15700 -770 17060 -650
rect 15590 -780 17060 -770
rect 17190 -650 18660 -640
rect 17190 -770 17200 -650
rect 17300 -770 18660 -650
rect 17190 -780 18660 -770
rect 18790 -650 20260 -640
rect 18790 -770 18800 -650
rect 18900 -770 20260 -650
rect 18790 -780 20260 -770
rect 20390 -650 21860 -640
rect 20390 -770 20400 -650
rect 20500 -770 21860 -650
rect 20390 -780 21860 -770
rect 21990 -650 23460 -640
rect 21990 -770 22000 -650
rect 22100 -770 23460 -650
rect 21990 -780 23460 -770
rect 23590 -650 25060 -640
rect 23590 -770 23600 -650
rect 23700 -770 25060 -650
rect 23590 -780 25060 -770
rect 25660 -650 28260 -640
rect 25660 -770 26800 -650
rect 26900 -770 28260 -650
rect 25660 -780 28260 -770
rect 28390 -650 31460 -640
rect 28390 -770 28400 -650
rect 28500 -770 31460 -650
rect 28390 -780 31460 -770
rect 32060 -780 36260 -640
rect 12510 -810 12520 -780
rect 660 -851 1077 -845
rect 660 -885 689 -851
rect 1065 -885 1077 -851
rect 660 -891 1077 -885
rect 1659 -851 2059 -845
rect 1659 -885 1671 -851
rect 2047 -885 2059 -851
rect 1659 -891 2059 -885
rect 2277 -851 2677 -845
rect 2277 -885 2289 -851
rect 2665 -885 2677 -851
rect 2277 -891 2677 -885
rect 3259 -851 3659 -845
rect 3259 -885 3271 -851
rect 3647 -885 3659 -851
rect 3259 -891 3659 -885
rect 3877 -851 4277 -845
rect 3877 -885 3889 -851
rect 4265 -885 4277 -851
rect 3877 -891 4277 -885
rect 4859 -851 5259 -845
rect 4859 -885 4871 -851
rect 5247 -885 5259 -851
rect 4859 -891 5259 -885
rect 5477 -851 5877 -845
rect 5477 -885 5489 -851
rect 5865 -885 5877 -851
rect 5477 -891 5877 -885
rect 6459 -851 6859 -845
rect 6459 -885 6471 -851
rect 6847 -885 6859 -851
rect 6459 -891 6859 -885
rect 7077 -851 7477 -845
rect 7077 -885 7089 -851
rect 7465 -885 7477 -851
rect 7077 -891 7477 -885
rect 8059 -851 8459 -845
rect 8059 -885 8071 -851
rect 8447 -885 8459 -851
rect 8059 -891 8459 -885
rect 8677 -851 9077 -845
rect 8677 -885 8689 -851
rect 9065 -885 9077 -851
rect 8677 -891 9077 -885
rect 9659 -851 10059 -845
rect 9659 -885 9671 -851
rect 10047 -885 10059 -851
rect 9659 -891 10059 -885
rect 10277 -851 10677 -845
rect 10277 -885 10289 -851
rect 10665 -885 10677 -851
rect 10277 -891 10677 -885
rect 11259 -851 11659 -845
rect 11259 -885 11271 -851
rect 11647 -885 11659 -851
rect 11259 -891 11659 -885
rect 11877 -851 12277 -845
rect 11877 -885 11889 -851
rect 12265 -885 12277 -851
rect 11877 -891 12277 -885
rect 59 -1109 480 -1103
rect 59 -1143 71 -1109
rect 447 -1143 480 -1109
rect 59 -1149 480 -1143
rect 440 -1340 480 -1149
rect -140 -1371 480 -1340
rect 660 -1103 710 -891
rect 1109 -930 1155 -918
rect 1581 -930 1627 -918
rect 2091 -930 2137 -918
rect 2199 -930 2245 -918
rect 2709 -930 2755 -918
rect 3181 -930 3227 -918
rect 3691 -930 3737 -918
rect 3799 -930 3845 -918
rect 4309 -930 4355 -918
rect 4781 -930 4827 -918
rect 5291 -930 5337 -918
rect 5399 -930 5445 -918
rect 5909 -930 5955 -918
rect 6381 -930 6427 -918
rect 6891 -930 6937 -918
rect 6999 -930 7045 -918
rect 7509 -930 7555 -918
rect 7981 -930 8027 -918
rect 8491 -930 8537 -918
rect 8599 -930 8645 -918
rect 9109 -930 9155 -918
rect 9581 -930 9627 -918
rect 10091 -930 10137 -918
rect 10199 -930 10245 -918
rect 10709 -930 10755 -918
rect 11181 -930 11227 -918
rect 11400 -930 11480 -891
rect 11691 -930 11737 -918
rect 11799 -930 11845 -918
rect 12020 -930 12100 -891
rect 12380 -910 12520 -810
rect 12880 -845 13240 -780
rect 13500 -845 13860 -780
rect 12859 -851 13259 -845
rect 12859 -885 12871 -851
rect 13247 -885 13259 -851
rect 12859 -891 13259 -885
rect 13477 -851 13877 -845
rect 13477 -885 13489 -851
rect 13865 -885 13877 -851
rect 13477 -891 13877 -885
rect 12310 -918 12520 -910
rect 12309 -930 12520 -918
rect 12781 -920 12827 -918
rect 1109 -1064 1115 -930
rect 1149 -1064 1155 -930
rect 1540 -1060 1587 -930
rect 1109 -1076 1155 -1064
rect 1581 -1064 1587 -1060
rect 1621 -1060 2097 -930
rect 1621 -1064 1627 -1060
rect 1581 -1076 1627 -1064
rect 2091 -1064 2097 -1060
rect 2131 -1060 2205 -930
rect 2131 -1064 2137 -1060
rect 2091 -1076 2137 -1064
rect 2199 -1064 2205 -1060
rect 2239 -1060 2715 -930
rect 2239 -1064 2245 -1060
rect 2199 -1076 2245 -1064
rect 2709 -1064 2715 -1060
rect 2749 -1060 3187 -930
rect 2749 -1064 2755 -1060
rect 2709 -1076 2755 -1064
rect 3181 -1064 3187 -1060
rect 3221 -1060 3697 -930
rect 3221 -1064 3227 -1060
rect 3181 -1076 3227 -1064
rect 3691 -1064 3697 -1060
rect 3731 -1060 3805 -930
rect 3731 -1064 3737 -1060
rect 3691 -1076 3737 -1064
rect 3799 -1064 3805 -1060
rect 3839 -1060 4315 -930
rect 3839 -1064 3845 -1060
rect 3799 -1076 3845 -1064
rect 4309 -1064 4315 -1060
rect 4349 -1060 4787 -930
rect 4349 -1064 4355 -1060
rect 4309 -1076 4355 -1064
rect 4781 -1064 4787 -1060
rect 4821 -1060 5297 -930
rect 4821 -1064 4827 -1060
rect 4781 -1076 4827 -1064
rect 5291 -1064 5297 -1060
rect 5331 -1060 5405 -930
rect 5331 -1064 5337 -1060
rect 5291 -1076 5337 -1064
rect 5399 -1064 5405 -1060
rect 5439 -1060 5915 -930
rect 5439 -1064 5445 -1060
rect 5399 -1076 5445 -1064
rect 5909 -1064 5915 -1060
rect 5949 -1060 6387 -930
rect 5949 -1064 5955 -1060
rect 5909 -1076 5955 -1064
rect 6381 -1064 6387 -1060
rect 6421 -1060 6897 -930
rect 6421 -1064 6427 -1060
rect 6381 -1076 6427 -1064
rect 6891 -1064 6897 -1060
rect 6931 -1060 7005 -930
rect 6931 -1064 6937 -1060
rect 6891 -1076 6937 -1064
rect 6999 -1064 7005 -1060
rect 7039 -1060 7515 -930
rect 7039 -1064 7045 -1060
rect 6999 -1076 7045 -1064
rect 7509 -1064 7515 -1060
rect 7549 -1060 7987 -930
rect 7549 -1064 7555 -1060
rect 7509 -1076 7555 -1064
rect 7981 -1064 7987 -1060
rect 8021 -1060 8497 -930
rect 8021 -1064 8027 -1060
rect 7981 -1076 8027 -1064
rect 8491 -1064 8497 -1060
rect 8531 -1060 8605 -930
rect 8531 -1064 8537 -1060
rect 8491 -1076 8537 -1064
rect 8599 -1064 8605 -1060
rect 8639 -1060 9115 -930
rect 8639 -1064 8645 -1060
rect 8599 -1076 8645 -1064
rect 9109 -1064 9115 -1060
rect 9149 -1060 9587 -930
rect 9149 -1064 9155 -1060
rect 9109 -1076 9155 -1064
rect 9581 -1064 9587 -1060
rect 9621 -1060 10097 -930
rect 9621 -1064 9627 -1060
rect 9581 -1076 9627 -1064
rect 10091 -1064 10097 -1060
rect 10131 -1060 10205 -930
rect 10131 -1064 10137 -1060
rect 10091 -1076 10137 -1064
rect 10199 -1064 10205 -1060
rect 10239 -1060 10715 -930
rect 10239 -1064 10245 -1060
rect 10199 -1076 10245 -1064
rect 10709 -1064 10715 -1060
rect 10749 -1060 11187 -930
rect 10749 -1064 10755 -1060
rect 10709 -1076 10755 -1064
rect 11181 -1064 11187 -1060
rect 11221 -1060 11697 -930
rect 11221 -1064 11227 -1060
rect 11181 -1076 11227 -1064
rect 11400 -1103 11480 -1060
rect 11691 -1064 11697 -1060
rect 11731 -1060 11805 -930
rect 11731 -1064 11737 -1060
rect 11691 -1076 11737 -1064
rect 11799 -1064 11805 -1060
rect 11839 -1060 12315 -930
rect 11839 -1064 11845 -1060
rect 11799 -1076 11845 -1064
rect 12020 -1103 12100 -1060
rect 12309 -1064 12315 -1060
rect 12349 -980 12520 -930
rect 12349 -1050 12390 -980
rect 12510 -1050 12520 -980
rect 12349 -1060 12520 -1050
rect 12620 -930 12827 -920
rect 12349 -1064 12355 -1060
rect 12309 -1076 12355 -1064
rect 12620 -1070 12630 -930
rect 12750 -1064 12787 -930
rect 12821 -1064 12827 -930
rect 12750 -1070 12827 -1064
rect 12620 -1076 12827 -1070
rect 13291 -930 13337 -918
rect 13291 -1064 13297 -930
rect 13331 -1064 13337 -930
rect 13291 -1076 13337 -1064
rect 13399 -930 13445 -918
rect 13399 -1064 13405 -930
rect 13439 -1064 13445 -930
rect 13399 -1076 13445 -1064
rect 13909 -920 13955 -918
rect 13909 -930 14100 -920
rect 13909 -1064 13915 -930
rect 13949 -1064 13970 -930
rect 13909 -1070 13970 -1064
rect 14090 -1070 14100 -930
rect 14160 -930 14300 -780
rect 16080 -825 16440 -780
rect 16700 -825 17060 -780
rect 17680 -825 18040 -780
rect 18300 -825 18660 -780
rect 19280 -825 19640 -780
rect 19900 -825 20260 -780
rect 20880 -825 21240 -780
rect 21500 -825 21860 -780
rect 22480 -825 22840 -780
rect 23100 -825 23460 -780
rect 24080 -825 24440 -780
rect 24700 -825 25060 -780
rect 25680 -825 26040 -780
rect 26300 -825 26660 -780
rect 27280 -825 27640 -780
rect 27900 -825 28260 -780
rect 28880 -825 29240 -780
rect 29500 -825 29860 -780
rect 30480 -825 30840 -780
rect 31100 -825 31460 -780
rect 32080 -825 32440 -780
rect 32700 -825 33060 -780
rect 33680 -825 34040 -780
rect 34300 -825 34660 -780
rect 35280 -825 35640 -780
rect 35900 -825 36260 -780
rect 16059 -830 16459 -825
rect 14459 -851 14859 -845
rect 14459 -885 14471 -851
rect 14847 -885 14859 -851
rect 14459 -891 14859 -885
rect 15077 -851 15477 -845
rect 15077 -885 15089 -851
rect 15465 -885 15477 -851
rect 15077 -891 15477 -885
rect 16059 -851 16460 -830
rect 16059 -885 16071 -851
rect 16447 -885 16460 -851
rect 16059 -890 16460 -885
rect 16677 -851 17077 -825
rect 16677 -885 16689 -851
rect 17065 -885 17077 -851
rect 16059 -891 16459 -890
rect 16677 -891 17077 -885
rect 17659 -830 18059 -825
rect 17659 -851 18060 -830
rect 17659 -885 17671 -851
rect 18047 -885 18060 -851
rect 17659 -890 18060 -885
rect 18277 -851 18677 -825
rect 18277 -885 18289 -851
rect 18665 -885 18677 -851
rect 17659 -891 18059 -890
rect 18277 -891 18677 -885
rect 19259 -830 19659 -825
rect 19259 -851 19660 -830
rect 19259 -885 19271 -851
rect 19647 -885 19660 -851
rect 19259 -890 19660 -885
rect 19877 -851 20277 -825
rect 19877 -885 19889 -851
rect 20265 -885 20277 -851
rect 19259 -891 19659 -890
rect 19877 -891 20277 -885
rect 20859 -830 21259 -825
rect 20859 -851 21260 -830
rect 20859 -885 20871 -851
rect 21247 -885 21260 -851
rect 20859 -890 21260 -885
rect 21477 -851 21877 -825
rect 21477 -885 21489 -851
rect 21865 -885 21877 -851
rect 20859 -891 21259 -890
rect 21477 -891 21877 -885
rect 22459 -830 22859 -825
rect 22459 -851 22860 -830
rect 22459 -885 22471 -851
rect 22847 -885 22860 -851
rect 22459 -890 22860 -885
rect 23077 -851 23477 -825
rect 23077 -885 23089 -851
rect 23465 -885 23477 -851
rect 22459 -891 22859 -890
rect 23077 -891 23477 -885
rect 24059 -830 24459 -825
rect 24059 -851 24460 -830
rect 24059 -885 24071 -851
rect 24447 -885 24460 -851
rect 24059 -890 24460 -885
rect 24677 -851 25077 -825
rect 24677 -885 24689 -851
rect 25065 -885 25077 -851
rect 24059 -891 24459 -890
rect 24677 -891 25077 -885
rect 25659 -830 26059 -825
rect 25659 -851 26060 -830
rect 25659 -885 25671 -851
rect 26047 -885 26060 -851
rect 25659 -890 26060 -885
rect 26277 -851 26677 -825
rect 26277 -885 26289 -851
rect 26665 -885 26677 -851
rect 25659 -891 26059 -890
rect 26277 -891 26677 -885
rect 27259 -830 27659 -825
rect 27259 -851 27660 -830
rect 27259 -885 27271 -851
rect 27647 -885 27660 -851
rect 27259 -890 27660 -885
rect 27877 -851 28277 -825
rect 27877 -885 27889 -851
rect 28265 -885 28277 -851
rect 27259 -891 27659 -890
rect 27877 -891 28277 -885
rect 28859 -830 29259 -825
rect 28859 -851 29260 -830
rect 28859 -885 28871 -851
rect 29247 -885 29260 -851
rect 28859 -890 29260 -885
rect 29477 -851 29877 -825
rect 29477 -885 29489 -851
rect 29865 -885 29877 -851
rect 28859 -891 29259 -890
rect 29477 -891 29877 -885
rect 30459 -830 30859 -825
rect 30459 -851 30860 -830
rect 30459 -885 30471 -851
rect 30847 -885 30860 -851
rect 30459 -890 30860 -885
rect 31077 -851 31477 -825
rect 32060 -830 32459 -825
rect 32060 -845 32460 -830
rect 31077 -885 31089 -851
rect 31465 -885 31477 -851
rect 30459 -891 30859 -890
rect 31077 -891 31477 -885
rect 32059 -851 32460 -845
rect 32059 -885 32071 -851
rect 32447 -885 32460 -851
rect 32059 -890 32460 -885
rect 32677 -851 33077 -825
rect 32677 -885 32689 -851
rect 33065 -885 33077 -851
rect 32059 -891 32459 -890
rect 32677 -891 33077 -885
rect 33659 -830 34059 -825
rect 33659 -851 34060 -830
rect 33659 -885 33671 -851
rect 34047 -885 34060 -851
rect 33659 -890 34060 -885
rect 34277 -851 34677 -825
rect 34277 -885 34289 -851
rect 34665 -885 34677 -851
rect 33659 -891 34059 -890
rect 34277 -891 34677 -885
rect 35259 -830 35659 -825
rect 35259 -851 35660 -830
rect 35259 -885 35271 -851
rect 35647 -885 35660 -851
rect 35259 -890 35660 -885
rect 35877 -851 36277 -825
rect 35877 -885 35889 -851
rect 36265 -885 36277 -851
rect 35259 -891 35659 -890
rect 35877 -891 36277 -885
rect 14381 -930 14427 -918
rect 14620 -930 14700 -891
rect 14891 -930 14937 -918
rect 14999 -930 15045 -918
rect 15220 -930 15300 -891
rect 36660 -918 36800 -509
rect 36859 -563 37259 -557
rect 36859 -597 36871 -563
rect 37247 -597 37259 -563
rect 36859 -603 37259 -597
rect 36859 -851 37259 -845
rect 36859 -885 36871 -851
rect 37247 -885 37259 -851
rect 36859 -891 37259 -885
rect 37300 -918 37440 -509
rect 37477 -563 37877 -557
rect 37477 -597 37489 -563
rect 37865 -597 37877 -563
rect 37477 -603 37877 -597
rect 37477 -851 37877 -845
rect 37477 -885 37489 -851
rect 37865 -885 37877 -851
rect 37477 -891 37877 -885
rect 37920 -918 38060 -509
rect 15509 -930 15555 -918
rect 15981 -930 16027 -918
rect 16491 -930 16537 -918
rect 16599 -930 16645 -918
rect 17109 -930 17155 -918
rect 17581 -930 17627 -918
rect 18091 -930 18137 -918
rect 18199 -930 18245 -918
rect 18709 -930 18755 -918
rect 19181 -930 19227 -918
rect 19691 -930 19737 -918
rect 19799 -930 19845 -918
rect 20309 -930 20355 -918
rect 20781 -930 20827 -918
rect 21291 -930 21337 -918
rect 21399 -930 21445 -918
rect 21909 -930 21955 -918
rect 22381 -930 22427 -918
rect 22891 -930 22937 -918
rect 22999 -930 23045 -918
rect 23509 -930 23555 -918
rect 23981 -930 24027 -918
rect 24491 -930 24537 -918
rect 24599 -930 24645 -918
rect 25109 -930 25155 -918
rect 25581 -930 25627 -918
rect 26091 -930 26137 -918
rect 26199 -930 26245 -918
rect 26709 -930 26755 -918
rect 27181 -930 27227 -918
rect 27691 -930 27737 -918
rect 27799 -930 27845 -918
rect 28309 -930 28355 -918
rect 28781 -930 28827 -918
rect 29291 -930 29337 -918
rect 29399 -930 29445 -918
rect 29909 -930 29955 -918
rect 30381 -930 30427 -918
rect 30891 -930 30937 -918
rect 30999 -930 31045 -918
rect 31509 -930 31555 -918
rect 31981 -930 32027 -918
rect 32491 -930 32537 -918
rect 32599 -930 32645 -918
rect 33109 -930 33155 -918
rect 33581 -930 33627 -918
rect 34091 -930 34137 -918
rect 34199 -930 34245 -918
rect 34709 -930 34755 -918
rect 35181 -930 35227 -918
rect 35691 -930 35737 -918
rect 35799 -930 35845 -918
rect 36309 -930 36355 -918
rect 36660 -930 36827 -918
rect 14160 -1060 14387 -930
rect 13909 -1076 14100 -1070
rect 14381 -1064 14387 -1060
rect 14421 -1060 14897 -930
rect 14421 -1064 14427 -1060
rect 14381 -1076 14427 -1064
rect 12620 -1080 12820 -1076
rect 13920 -1080 14100 -1076
rect 12870 -1103 13250 -1100
rect 14620 -1103 14700 -1060
rect 14891 -1064 14897 -1060
rect 14931 -1060 15005 -930
rect 14931 -1064 14937 -1060
rect 14891 -1076 14937 -1064
rect 14999 -1064 15005 -1060
rect 15039 -1060 15515 -930
rect 15039 -1064 15045 -1060
rect 14999 -1076 15045 -1064
rect 15220 -1103 15300 -1060
rect 15509 -1064 15515 -1060
rect 15549 -1060 15987 -930
rect 15549 -1064 15555 -1060
rect 15509 -1076 15555 -1064
rect 15981 -1064 15987 -1060
rect 16021 -1060 16497 -930
rect 16021 -1064 16027 -1060
rect 15981 -1076 16027 -1064
rect 16491 -1064 16497 -1060
rect 16531 -1060 16605 -930
rect 16531 -1064 16537 -1060
rect 16491 -1076 16537 -1064
rect 16599 -1064 16605 -1060
rect 16639 -1060 17115 -930
rect 16639 -1064 16645 -1060
rect 16599 -1076 16645 -1064
rect 17109 -1064 17115 -1060
rect 17149 -1060 17587 -930
rect 17149 -1064 17155 -1060
rect 17109 -1076 17155 -1064
rect 17581 -1064 17587 -1060
rect 17621 -1060 18097 -930
rect 17621 -1064 17627 -1060
rect 17581 -1076 17627 -1064
rect 18091 -1064 18097 -1060
rect 18131 -1060 18205 -930
rect 18131 -1064 18137 -1060
rect 18091 -1076 18137 -1064
rect 18199 -1064 18205 -1060
rect 18239 -1060 18715 -930
rect 18239 -1064 18245 -1060
rect 18199 -1076 18245 -1064
rect 18709 -1064 18715 -1060
rect 18749 -1060 19187 -930
rect 18749 -1064 18755 -1060
rect 18709 -1076 18755 -1064
rect 19181 -1064 19187 -1060
rect 19221 -1060 19697 -930
rect 19221 -1064 19227 -1060
rect 19181 -1076 19227 -1064
rect 19691 -1064 19697 -1060
rect 19731 -1060 19805 -930
rect 19731 -1064 19737 -1060
rect 19691 -1076 19737 -1064
rect 19799 -1064 19805 -1060
rect 19839 -1060 20315 -930
rect 19839 -1064 19845 -1060
rect 19799 -1076 19845 -1064
rect 20309 -1064 20315 -1060
rect 20349 -1060 20787 -930
rect 20349 -1064 20355 -1060
rect 20309 -1076 20355 -1064
rect 20781 -1064 20787 -1060
rect 20821 -1060 21297 -930
rect 20821 -1064 20827 -1060
rect 20781 -1076 20827 -1064
rect 21291 -1064 21297 -1060
rect 21331 -1060 21405 -930
rect 21331 -1064 21337 -1060
rect 21291 -1076 21337 -1064
rect 21399 -1064 21405 -1060
rect 21439 -1060 21915 -930
rect 21439 -1064 21445 -1060
rect 21399 -1076 21445 -1064
rect 21909 -1064 21915 -1060
rect 21949 -1060 22387 -930
rect 21949 -1064 21955 -1060
rect 21909 -1076 21955 -1064
rect 22381 -1064 22387 -1060
rect 22421 -1060 22897 -930
rect 22421 -1064 22427 -1060
rect 22381 -1076 22427 -1064
rect 22891 -1064 22897 -1060
rect 22931 -1060 23005 -930
rect 22931 -1064 22937 -1060
rect 22891 -1076 22937 -1064
rect 22999 -1064 23005 -1060
rect 23039 -1060 23515 -930
rect 23039 -1064 23045 -1060
rect 22999 -1076 23045 -1064
rect 23509 -1064 23515 -1060
rect 23549 -1060 23987 -930
rect 23549 -1064 23555 -1060
rect 23509 -1076 23555 -1064
rect 23981 -1064 23987 -1060
rect 24021 -1060 24497 -930
rect 24021 -1064 24027 -1060
rect 23981 -1076 24027 -1064
rect 24491 -1064 24497 -1060
rect 24531 -1060 24605 -930
rect 24531 -1064 24537 -1060
rect 24491 -1076 24537 -1064
rect 24599 -1064 24605 -1060
rect 24639 -1060 25115 -930
rect 24639 -1064 24645 -1060
rect 24599 -1076 24645 -1064
rect 25109 -1064 25115 -1060
rect 25149 -1060 25587 -930
rect 25149 -1064 25155 -1060
rect 25109 -1076 25155 -1064
rect 25581 -1064 25587 -1060
rect 25621 -1060 26097 -930
rect 25621 -1064 25627 -1060
rect 25581 -1076 25627 -1064
rect 26091 -1064 26097 -1060
rect 26131 -1060 26205 -930
rect 26131 -1064 26137 -1060
rect 26091 -1076 26137 -1064
rect 26199 -1064 26205 -1060
rect 26239 -1060 26715 -930
rect 26239 -1064 26245 -1060
rect 26199 -1076 26245 -1064
rect 26709 -1064 26715 -1060
rect 26749 -1060 27187 -930
rect 26749 -1064 26755 -1060
rect 26709 -1076 26755 -1064
rect 27181 -1064 27187 -1060
rect 27221 -1060 27697 -930
rect 27221 -1064 27227 -1060
rect 27181 -1076 27227 -1064
rect 27691 -1064 27697 -1060
rect 27731 -1060 27805 -930
rect 27731 -1064 27737 -1060
rect 27691 -1076 27737 -1064
rect 27799 -1064 27805 -1060
rect 27839 -1060 28315 -930
rect 27839 -1064 27845 -1060
rect 27799 -1076 27845 -1064
rect 28309 -1064 28315 -1060
rect 28349 -1060 28787 -930
rect 28349 -1064 28355 -1060
rect 28309 -1076 28355 -1064
rect 28781 -1064 28787 -1060
rect 28821 -1060 29297 -930
rect 28821 -1064 28827 -1060
rect 28781 -1076 28827 -1064
rect 29291 -1064 29297 -1060
rect 29331 -1060 29405 -930
rect 29331 -1064 29337 -1060
rect 29291 -1076 29337 -1064
rect 29399 -1064 29405 -1060
rect 29439 -1060 29915 -930
rect 29439 -1064 29445 -1060
rect 29399 -1076 29445 -1064
rect 29909 -1064 29915 -1060
rect 29949 -1060 30387 -930
rect 29949 -1064 29955 -1060
rect 29909 -1076 29955 -1064
rect 30381 -1064 30387 -1060
rect 30421 -1060 30897 -930
rect 30421 -1064 30427 -1060
rect 30381 -1076 30427 -1064
rect 30891 -1064 30897 -1060
rect 30931 -1060 31005 -930
rect 30931 -1064 30937 -1060
rect 30891 -1076 30937 -1064
rect 30999 -1064 31005 -1060
rect 31039 -1060 31515 -930
rect 31039 -1064 31045 -1060
rect 30999 -1076 31045 -1064
rect 31509 -1064 31515 -1060
rect 31549 -1060 31987 -930
rect 31549 -1064 31555 -1060
rect 31509 -1076 31555 -1064
rect 31981 -1064 31987 -1060
rect 32021 -1060 32497 -930
rect 32021 -1064 32027 -1060
rect 31981 -1076 32027 -1064
rect 32491 -1064 32497 -1060
rect 32531 -1060 32605 -930
rect 32531 -1064 32537 -1060
rect 32491 -1076 32537 -1064
rect 32599 -1064 32605 -1060
rect 32639 -1060 33115 -930
rect 32639 -1064 32645 -1060
rect 32599 -1076 32645 -1064
rect 33109 -1064 33115 -1060
rect 33149 -1060 33587 -930
rect 33149 -1064 33155 -1060
rect 33109 -1076 33155 -1064
rect 33581 -1064 33587 -1060
rect 33621 -1060 34097 -930
rect 33621 -1064 33627 -1060
rect 33581 -1076 33627 -1064
rect 34091 -1064 34097 -1060
rect 34131 -1060 34205 -930
rect 34131 -1064 34137 -1060
rect 34091 -1076 34137 -1064
rect 34199 -1064 34205 -1060
rect 34239 -1060 34715 -930
rect 34239 -1064 34245 -1060
rect 34199 -1076 34245 -1064
rect 34709 -1064 34715 -1060
rect 34749 -1060 35187 -930
rect 34749 -1064 34755 -1060
rect 34709 -1076 34755 -1064
rect 35181 -1064 35187 -1060
rect 35221 -1060 35697 -930
rect 35221 -1064 35227 -1060
rect 35181 -1076 35227 -1064
rect 35691 -1064 35697 -1060
rect 35731 -1060 35805 -930
rect 35731 -1064 35737 -1060
rect 35691 -1076 35737 -1064
rect 35799 -1064 35805 -1060
rect 35839 -1060 36315 -930
rect 35839 -1064 35845 -1060
rect 35799 -1076 35845 -1064
rect 36309 -1064 36315 -1060
rect 36349 -1060 36400 -930
rect 36349 -1064 36355 -1060
rect 36309 -1076 36355 -1064
rect 36660 -1064 36787 -930
rect 36821 -1064 36827 -930
rect 36660 -1076 36827 -1064
rect 37291 -930 37445 -918
rect 37291 -1064 37297 -930
rect 37331 -1064 37405 -930
rect 37439 -1064 37445 -930
rect 37291 -1076 37445 -1064
rect 37909 -930 38060 -918
rect 37909 -1064 37915 -930
rect 37949 -1064 38060 -930
rect 37909 -1076 38060 -1064
rect 660 -1109 1077 -1103
rect 660 -1143 689 -1109
rect 1065 -1143 1077 -1109
rect 1659 -1109 2059 -1103
rect 660 -1149 1077 -1143
rect 1180 -1120 1320 -1110
rect 1659 -1120 1671 -1109
rect 660 -1340 710 -1149
rect 1180 -1240 1190 -1120
rect 1310 -1143 1671 -1120
rect 2047 -1120 2059 -1109
rect 2277 -1109 2677 -1103
rect 2277 -1120 2289 -1109
rect 2047 -1143 2289 -1120
rect 2665 -1120 2677 -1109
rect 3259 -1109 3659 -1103
rect 2780 -1120 2920 -1110
rect 3259 -1120 3271 -1109
rect 2665 -1143 2790 -1120
rect 1310 -1240 2790 -1143
rect 2910 -1143 3271 -1120
rect 3647 -1120 3659 -1109
rect 3877 -1109 4277 -1103
rect 3877 -1120 3889 -1109
rect 3647 -1143 3889 -1120
rect 4265 -1120 4277 -1109
rect 4859 -1109 5259 -1103
rect 4380 -1120 4520 -1110
rect 4859 -1120 4871 -1109
rect 4265 -1143 4390 -1120
rect 2910 -1240 4390 -1143
rect 4510 -1143 4871 -1120
rect 5247 -1120 5259 -1109
rect 5477 -1109 5877 -1103
rect 5477 -1120 5489 -1109
rect 5247 -1143 5489 -1120
rect 5865 -1120 5877 -1109
rect 6459 -1109 6859 -1103
rect 5980 -1120 6120 -1110
rect 6459 -1120 6471 -1109
rect 5865 -1143 5990 -1120
rect 4510 -1240 5990 -1143
rect 6110 -1143 6471 -1120
rect 6847 -1120 6859 -1109
rect 7077 -1109 7477 -1103
rect 7077 -1120 7089 -1109
rect 6847 -1143 7089 -1120
rect 7465 -1120 7477 -1109
rect 8059 -1109 8459 -1103
rect 7580 -1120 7720 -1110
rect 8059 -1120 8071 -1109
rect 7465 -1143 7590 -1120
rect 6110 -1240 7590 -1143
rect 7710 -1143 8071 -1120
rect 8447 -1120 8459 -1109
rect 8677 -1109 9077 -1103
rect 8677 -1120 8689 -1109
rect 8447 -1143 8689 -1120
rect 9065 -1120 9077 -1109
rect 9659 -1109 10059 -1103
rect 9180 -1120 9320 -1110
rect 9659 -1120 9671 -1109
rect 9065 -1143 9190 -1120
rect 7710 -1240 9190 -1143
rect 9310 -1143 9671 -1120
rect 10047 -1120 10059 -1109
rect 10277 -1109 10677 -1103
rect 10277 -1120 10289 -1109
rect 10047 -1143 10289 -1120
rect 10665 -1120 10677 -1109
rect 11259 -1109 11659 -1103
rect 10665 -1143 10720 -1120
rect 9310 -1240 10720 -1143
rect 11259 -1143 11271 -1109
rect 11647 -1143 11659 -1109
rect 11259 -1149 11659 -1143
rect 11877 -1109 12277 -1103
rect 11877 -1143 11889 -1109
rect 12265 -1143 12277 -1109
rect 11877 -1149 12277 -1143
rect 12859 -1109 13259 -1103
rect 12859 -1143 12871 -1109
rect 13247 -1120 13259 -1109
rect 13477 -1109 13877 -1103
rect 13477 -1120 13489 -1109
rect 13247 -1143 13489 -1120
rect 13865 -1143 13877 -1109
rect 12859 -1149 12880 -1143
rect 1180 -1250 1320 -1240
rect 2780 -1250 2920 -1240
rect 4380 -1250 4520 -1240
rect 5980 -1250 6120 -1240
rect 7580 -1250 7720 -1240
rect 9180 -1250 9320 -1240
rect 12870 -1260 12880 -1149
rect 13240 -1149 13877 -1143
rect 14459 -1109 14859 -1103
rect 14459 -1143 14471 -1109
rect 14847 -1143 14859 -1109
rect 14459 -1149 14859 -1143
rect 15077 -1109 15477 -1103
rect 15077 -1143 15089 -1109
rect 15465 -1143 15477 -1109
rect 16059 -1109 16459 -1103
rect 15077 -1149 15477 -1143
rect 15810 -1120 15930 -1110
rect 16059 -1120 16071 -1109
rect 13240 -1260 13860 -1149
rect 15810 -1240 15820 -1120
rect 15920 -1143 16071 -1120
rect 16447 -1120 16459 -1109
rect 16677 -1109 17077 -1103
rect 16677 -1120 16689 -1109
rect 16447 -1143 16689 -1120
rect 17065 -1120 17077 -1109
rect 17659 -1109 18059 -1103
rect 17410 -1120 17530 -1110
rect 17659 -1120 17671 -1109
rect 17065 -1143 17120 -1120
rect 15920 -1240 17120 -1143
rect 17410 -1240 17420 -1120
rect 17520 -1143 17671 -1120
rect 18047 -1120 18059 -1109
rect 18277 -1109 18677 -1103
rect 18277 -1120 18289 -1109
rect 18047 -1143 18289 -1120
rect 18665 -1120 18677 -1109
rect 19259 -1109 19659 -1103
rect 19010 -1120 19130 -1110
rect 19259 -1120 19271 -1109
rect 18665 -1143 18720 -1120
rect 17520 -1240 18720 -1143
rect 19010 -1240 19020 -1120
rect 19120 -1143 19271 -1120
rect 19647 -1120 19659 -1109
rect 19877 -1109 20277 -1103
rect 19877 -1120 19889 -1109
rect 19647 -1143 19889 -1120
rect 20265 -1120 20277 -1109
rect 20859 -1109 21259 -1103
rect 20610 -1120 20730 -1110
rect 20859 -1120 20871 -1109
rect 20265 -1143 20320 -1120
rect 19120 -1240 20320 -1143
rect 20610 -1240 20620 -1120
rect 20720 -1143 20871 -1120
rect 21247 -1120 21259 -1109
rect 21477 -1109 21877 -1103
rect 21477 -1120 21489 -1109
rect 21247 -1143 21489 -1120
rect 21865 -1120 21877 -1109
rect 22459 -1109 22859 -1103
rect 22210 -1120 22330 -1110
rect 22459 -1120 22471 -1109
rect 21865 -1143 21920 -1120
rect 20720 -1240 21920 -1143
rect 22210 -1240 22220 -1120
rect 22320 -1143 22471 -1120
rect 22847 -1120 22859 -1109
rect 23077 -1109 23477 -1103
rect 23077 -1120 23089 -1109
rect 22847 -1143 23089 -1120
rect 23465 -1120 23477 -1109
rect 24059 -1109 24459 -1103
rect 23810 -1120 23930 -1110
rect 24059 -1120 24071 -1109
rect 23465 -1143 23520 -1120
rect 22320 -1240 23520 -1143
rect 23810 -1240 23820 -1120
rect 23920 -1143 24071 -1120
rect 24447 -1120 24459 -1109
rect 24677 -1109 25077 -1103
rect 24677 -1120 24689 -1109
rect 24447 -1143 24689 -1120
rect 25065 -1120 25077 -1109
rect 25659 -1109 26059 -1103
rect 25659 -1120 25671 -1109
rect 25065 -1143 25120 -1120
rect 23920 -1240 25120 -1143
rect 25620 -1143 25671 -1120
rect 26047 -1120 26059 -1109
rect 26277 -1109 26677 -1103
rect 26277 -1120 26289 -1109
rect 26047 -1143 26289 -1120
rect 26665 -1120 26677 -1109
rect 27259 -1109 27659 -1103
rect 27259 -1110 27271 -1109
rect 27010 -1120 27271 -1110
rect 26665 -1143 27020 -1120
rect 25620 -1240 27020 -1143
rect 27120 -1143 27271 -1120
rect 27647 -1110 27659 -1109
rect 27877 -1109 28277 -1103
rect 27877 -1110 27889 -1109
rect 27647 -1143 27889 -1110
rect 28265 -1143 28277 -1109
rect 28859 -1109 29259 -1103
rect 28859 -1110 28871 -1109
rect 27120 -1149 28277 -1143
rect 28610 -1120 28871 -1110
rect 27120 -1240 28270 -1149
rect 15810 -1250 15930 -1240
rect 17410 -1250 17530 -1240
rect 19010 -1250 19130 -1240
rect 20610 -1250 20730 -1240
rect 22210 -1250 22330 -1240
rect 23810 -1250 23930 -1240
rect 27010 -1250 28270 -1240
rect 28610 -1240 28620 -1120
rect 28720 -1143 28871 -1120
rect 29247 -1110 29259 -1109
rect 29477 -1109 29877 -1103
rect 29477 -1110 29489 -1109
rect 29247 -1143 29489 -1110
rect 29865 -1110 29877 -1109
rect 30459 -1109 30859 -1103
rect 30459 -1110 30471 -1109
rect 29865 -1143 30471 -1110
rect 30847 -1110 30859 -1109
rect 31077 -1109 31477 -1103
rect 31077 -1110 31089 -1109
rect 30847 -1143 31089 -1110
rect 31465 -1110 31477 -1109
rect 32059 -1109 32459 -1103
rect 31465 -1143 31520 -1110
rect 28720 -1240 31520 -1143
rect 28610 -1250 31520 -1240
rect 31590 -1120 31710 -1110
rect 32059 -1120 32071 -1109
rect 31590 -1240 31600 -1120
rect 31700 -1143 32071 -1120
rect 32447 -1120 32459 -1109
rect 32677 -1109 33077 -1103
rect 32677 -1120 32689 -1109
rect 32447 -1143 32689 -1120
rect 33065 -1120 33077 -1109
rect 33659 -1109 34059 -1103
rect 33659 -1120 33671 -1109
rect 33065 -1143 33671 -1120
rect 34047 -1120 34059 -1109
rect 34277 -1109 34677 -1103
rect 34277 -1120 34289 -1109
rect 34047 -1143 34289 -1120
rect 34665 -1120 34677 -1109
rect 35259 -1109 35659 -1103
rect 35259 -1120 35271 -1109
rect 34665 -1143 35271 -1120
rect 35647 -1120 35659 -1109
rect 35877 -1109 36277 -1103
rect 35877 -1120 35889 -1109
rect 35647 -1143 35889 -1120
rect 36265 -1143 36277 -1109
rect 31700 -1149 36277 -1143
rect 31700 -1240 36270 -1149
rect 31590 -1250 31710 -1240
rect 12870 -1290 13860 -1260
rect 36660 -1300 36800 -1076
rect 36859 -1109 37259 -1103
rect 36859 -1143 36871 -1109
rect 37247 -1143 37259 -1109
rect 36859 -1149 37259 -1143
rect 37300 -1300 37440 -1076
rect 37477 -1109 37877 -1103
rect 37477 -1143 37489 -1109
rect 37865 -1143 37877 -1109
rect 37477 -1149 37877 -1143
rect 37920 -1300 38060 -1076
rect 31760 -1340 38060 -1300
rect 660 -1365 38060 -1340
rect 660 -1371 38065 -1365
rect -140 -1405 -117 -1371
rect 1253 -1405 1483 -1371
rect 2853 -1405 3083 -1371
rect 4453 -1405 4683 -1371
rect 6053 -1405 6283 -1371
rect 7653 -1405 7883 -1371
rect 9253 -1405 9483 -1371
rect 10853 -1405 11083 -1371
rect 12453 -1405 12683 -1371
rect 14053 -1405 14283 -1371
rect 15653 -1405 15883 -1371
rect 17253 -1405 17483 -1371
rect 18853 -1405 19083 -1371
rect 20453 -1405 20683 -1371
rect 22053 -1405 22283 -1371
rect 23653 -1405 23883 -1371
rect 25253 -1405 25483 -1371
rect 26853 -1405 27083 -1371
rect 28453 -1405 28683 -1371
rect 30053 -1405 30283 -1371
rect 31653 -1405 31883 -1371
rect 33253 -1405 33483 -1371
rect 34853 -1405 35083 -1371
rect 36453 -1405 36683 -1371
rect 38053 -1405 38065 -1371
rect -140 -1505 480 -1405
rect -140 -1539 71 -1505
rect 447 -1539 480 -1505
rect -140 -1540 480 -1539
rect -140 -1593 0 -1540
rect 59 -1545 480 -1540
rect -140 -1605 27 -1593
rect -140 -2297 -13 -1605
rect 21 -2297 27 -1605
rect -140 -2309 27 -2297
rect -140 -2718 0 -2309
rect 440 -2357 480 -1545
rect 660 -1411 38065 -1405
rect 660 -1420 38060 -1411
rect 660 -1505 31780 -1420
rect 32060 -1470 33490 -1460
rect 32060 -1499 33360 -1470
rect 660 -1539 689 -1505
rect 1065 -1539 1671 -1505
rect 2047 -1539 2289 -1505
rect 2665 -1539 3271 -1505
rect 3647 -1539 3889 -1505
rect 4265 -1539 4871 -1505
rect 5247 -1539 5489 -1505
rect 5865 -1539 6471 -1505
rect 6847 -1539 7089 -1505
rect 7465 -1539 8071 -1505
rect 8447 -1539 8689 -1505
rect 9065 -1539 9671 -1505
rect 10047 -1539 10289 -1505
rect 10665 -1539 11271 -1505
rect 11647 -1539 11889 -1505
rect 12265 -1539 12871 -1505
rect 13247 -1539 13489 -1505
rect 13865 -1539 14471 -1505
rect 14847 -1539 15089 -1505
rect 15465 -1539 16071 -1505
rect 16447 -1539 16689 -1505
rect 17065 -1539 17671 -1505
rect 18047 -1539 18289 -1505
rect 18665 -1539 19271 -1505
rect 19647 -1539 19889 -1505
rect 20265 -1539 20871 -1505
rect 21247 -1539 21489 -1505
rect 21865 -1539 22471 -1505
rect 22847 -1539 23089 -1505
rect 23465 -1539 24071 -1505
rect 24447 -1539 24689 -1505
rect 25065 -1539 25671 -1505
rect 26047 -1539 26289 -1505
rect 26665 -1539 27271 -1505
rect 27647 -1539 27889 -1505
rect 28265 -1539 28871 -1505
rect 29247 -1539 29489 -1505
rect 29865 -1539 30471 -1505
rect 30847 -1539 31089 -1505
rect 31465 -1539 31780 -1505
rect 660 -1540 31780 -1539
rect 32059 -1505 33360 -1499
rect 32059 -1539 32071 -1505
rect 32447 -1539 32689 -1505
rect 33065 -1539 33360 -1505
rect 32059 -1540 33360 -1539
rect 660 -1545 1077 -1540
rect 1659 -1545 2059 -1540
rect 2277 -1545 2677 -1540
rect 3259 -1545 3659 -1540
rect 3877 -1545 4277 -1540
rect 4859 -1545 5259 -1540
rect 5477 -1545 5877 -1540
rect 6459 -1545 6859 -1540
rect 7077 -1545 7477 -1540
rect 8059 -1545 8459 -1540
rect 8677 -1545 9077 -1540
rect 9659 -1545 10059 -1540
rect 10277 -1545 10677 -1540
rect 11259 -1545 11659 -1540
rect 11877 -1545 12277 -1540
rect 12859 -1545 13259 -1540
rect 13477 -1545 13877 -1540
rect 14459 -1545 14859 -1540
rect 15077 -1545 15477 -1540
rect 16059 -1545 16459 -1540
rect 16677 -1545 17077 -1540
rect 17659 -1545 18059 -1540
rect 18277 -1545 18677 -1540
rect 19259 -1545 19659 -1540
rect 19877 -1545 20277 -1540
rect 20859 -1545 21259 -1540
rect 21477 -1545 21877 -1540
rect 22459 -1545 22859 -1540
rect 23077 -1545 23477 -1540
rect 24059 -1545 24459 -1540
rect 24677 -1545 25077 -1540
rect 25659 -1545 26059 -1540
rect 26277 -1545 26677 -1540
rect 27259 -1545 27659 -1540
rect 27877 -1545 28277 -1540
rect 28859 -1545 29259 -1540
rect 29477 -1545 29877 -1540
rect 30459 -1545 30859 -1540
rect 31077 -1545 31477 -1540
rect 32059 -1545 32459 -1540
rect 32677 -1545 33077 -1540
rect 59 -2363 480 -2357
rect 59 -2397 71 -2363
rect 447 -2397 480 -2363
rect 59 -2403 480 -2397
rect 440 -2645 480 -2403
rect 59 -2651 480 -2645
rect 59 -2685 71 -2651
rect 447 -2685 480 -2651
rect 59 -2691 480 -2685
rect -140 -2730 27 -2718
rect -140 -2864 -13 -2730
rect 21 -2864 27 -2730
rect -140 -2876 27 -2864
rect -140 -3140 0 -2876
rect 440 -2903 480 -2691
rect 660 -2357 710 -1545
rect 33350 -1590 33360 -1540
rect 33480 -1590 33490 -1470
rect 33660 -1470 35650 -1460
rect 33660 -1499 35020 -1470
rect 33659 -1505 35020 -1499
rect 33659 -1539 33671 -1505
rect 34047 -1539 34289 -1505
rect 34665 -1539 35020 -1505
rect 33659 -1540 35020 -1539
rect 33659 -1545 34059 -1540
rect 34277 -1545 34677 -1540
rect 1109 -1605 1155 -1593
rect 1109 -2297 1115 -1605
rect 1149 -2297 1155 -1605
rect 1109 -2309 1155 -2297
rect 1581 -1605 1627 -1593
rect 1581 -2297 1587 -1605
rect 1621 -2297 1627 -1605
rect 1581 -2309 1627 -2297
rect 2091 -1600 2137 -1593
rect 2199 -1600 2245 -1593
rect 2091 -1605 2245 -1600
rect 2091 -2297 2097 -1605
rect 2131 -1610 2205 -1605
rect 2131 -2297 2205 -2290
rect 2239 -2297 2245 -1605
rect 2091 -2300 2245 -2297
rect 2091 -2309 2137 -2300
rect 2199 -2309 2245 -2300
rect 2709 -1605 2755 -1593
rect 2709 -2297 2715 -1605
rect 2749 -2297 2755 -1605
rect 2709 -2309 2755 -2297
rect 3181 -1605 3227 -1593
rect 3181 -2297 3187 -1605
rect 3221 -2297 3227 -1605
rect 3181 -2309 3227 -2297
rect 3691 -1600 3737 -1593
rect 3799 -1600 3845 -1593
rect 3691 -1605 3845 -1600
rect 3691 -2297 3697 -1605
rect 3731 -1610 3805 -1605
rect 3731 -2297 3805 -2290
rect 3839 -2297 3845 -1605
rect 3691 -2300 3845 -2297
rect 3691 -2309 3737 -2300
rect 3799 -2309 3845 -2300
rect 4309 -1605 4355 -1593
rect 4309 -2297 4315 -1605
rect 4349 -2297 4355 -1605
rect 4309 -2309 4355 -2297
rect 4781 -1605 4827 -1593
rect 4781 -2297 4787 -1605
rect 4821 -2297 4827 -1605
rect 4781 -2309 4827 -2297
rect 5291 -1600 5337 -1593
rect 5399 -1600 5445 -1593
rect 5291 -1605 5445 -1600
rect 5291 -2297 5297 -1605
rect 5331 -1610 5405 -1605
rect 5331 -2297 5405 -2290
rect 5439 -2297 5445 -1605
rect 5291 -2300 5445 -2297
rect 5291 -2309 5337 -2300
rect 5399 -2309 5445 -2300
rect 5909 -1605 5955 -1593
rect 5909 -2297 5915 -1605
rect 5949 -2297 5955 -1605
rect 5909 -2309 5955 -2297
rect 6381 -1605 6427 -1593
rect 6381 -2297 6387 -1605
rect 6421 -2297 6427 -1605
rect 6381 -2309 6427 -2297
rect 6891 -1600 6937 -1593
rect 6999 -1600 7045 -1593
rect 6891 -1605 7045 -1600
rect 6891 -2297 6897 -1605
rect 6931 -1610 7005 -1605
rect 6931 -2297 7005 -2290
rect 7039 -2297 7045 -1605
rect 6891 -2300 7045 -2297
rect 6891 -2309 6937 -2300
rect 6999 -2309 7045 -2300
rect 7509 -1605 7555 -1593
rect 7509 -2297 7515 -1605
rect 7549 -2297 7555 -1605
rect 7509 -2309 7555 -2297
rect 7981 -1605 8027 -1593
rect 7981 -2297 7987 -1605
rect 8021 -2297 8027 -1605
rect 7981 -2309 8027 -2297
rect 8491 -1600 8537 -1593
rect 8599 -1600 8645 -1593
rect 8491 -1605 8645 -1600
rect 8491 -2297 8497 -1605
rect 8531 -1610 8605 -1605
rect 8531 -2297 8605 -2290
rect 8639 -2297 8645 -1605
rect 8491 -2300 8645 -2297
rect 8491 -2309 8537 -2300
rect 8599 -2309 8645 -2300
rect 9109 -1605 9155 -1593
rect 9109 -2297 9115 -1605
rect 9149 -2297 9155 -1605
rect 9109 -2309 9155 -2297
rect 9581 -1605 9627 -1593
rect 9581 -2297 9587 -1605
rect 9621 -2297 9627 -1605
rect 9581 -2309 9627 -2297
rect 10091 -1600 10137 -1593
rect 10199 -1600 10245 -1593
rect 10091 -1605 10245 -1600
rect 10091 -2297 10097 -1605
rect 10131 -1610 10205 -1605
rect 10131 -2297 10205 -2290
rect 10239 -2297 10245 -1605
rect 10091 -2300 10245 -2297
rect 10091 -2309 10137 -2300
rect 10199 -2309 10245 -2300
rect 10709 -1605 10755 -1593
rect 10709 -2297 10715 -1605
rect 10749 -2297 10755 -1605
rect 10709 -2309 10755 -2297
rect 11181 -1605 11227 -1593
rect 11181 -2297 11187 -1605
rect 11221 -2297 11227 -1605
rect 11181 -2309 11227 -2297
rect 11691 -1600 11737 -1593
rect 11799 -1600 11845 -1593
rect 11691 -1605 11845 -1600
rect 11691 -2297 11697 -1605
rect 11731 -1610 11805 -1605
rect 11731 -2297 11805 -2290
rect 11839 -2297 11845 -1605
rect 11691 -2300 11845 -2297
rect 11691 -2309 11737 -2300
rect 11799 -2309 11845 -2300
rect 12309 -1605 12355 -1593
rect 12309 -2297 12315 -1605
rect 12349 -2297 12355 -1605
rect 12309 -2309 12355 -2297
rect 12781 -1605 12827 -1593
rect 12781 -2297 12787 -1605
rect 12821 -2297 12827 -1605
rect 12781 -2309 12827 -2297
rect 13291 -1600 13337 -1593
rect 13399 -1600 13445 -1593
rect 13291 -1605 13445 -1600
rect 13291 -2297 13297 -1605
rect 13331 -1610 13405 -1605
rect 13331 -2297 13405 -2290
rect 13439 -2297 13445 -1605
rect 13291 -2300 13445 -2297
rect 13291 -2309 13337 -2300
rect 13399 -2309 13445 -2300
rect 13909 -1605 13955 -1593
rect 13909 -2297 13915 -1605
rect 13949 -2297 13955 -1605
rect 13909 -2309 13955 -2297
rect 14381 -1605 14427 -1593
rect 14381 -2297 14387 -1605
rect 14421 -2297 14427 -1605
rect 14381 -2309 14427 -2297
rect 14891 -1600 14937 -1593
rect 14999 -1600 15045 -1593
rect 14891 -1605 15045 -1600
rect 14891 -2297 14897 -1605
rect 14931 -1610 15005 -1605
rect 14931 -2297 15005 -2290
rect 15039 -2297 15045 -1605
rect 14891 -2300 15045 -2297
rect 14891 -2309 14937 -2300
rect 14999 -2309 15045 -2300
rect 15509 -1605 15555 -1593
rect 15509 -2297 15515 -1605
rect 15549 -2297 15555 -1605
rect 15509 -2309 15555 -2297
rect 15981 -1605 16027 -1593
rect 15981 -2297 15987 -1605
rect 16021 -2297 16027 -1605
rect 15981 -2309 16027 -2297
rect 16491 -1600 16537 -1593
rect 16599 -1600 16645 -1593
rect 16491 -1605 16645 -1600
rect 16491 -2297 16497 -1605
rect 16531 -1610 16605 -1605
rect 16531 -2297 16605 -2290
rect 16639 -2297 16645 -1605
rect 16491 -2300 16645 -2297
rect 16491 -2309 16537 -2300
rect 16599 -2309 16645 -2300
rect 17109 -1605 17155 -1593
rect 17109 -2297 17115 -1605
rect 17149 -2297 17155 -1605
rect 17109 -2309 17155 -2297
rect 17581 -1605 17627 -1593
rect 17581 -2297 17587 -1605
rect 17621 -2297 17627 -1605
rect 17581 -2309 17627 -2297
rect 18091 -1600 18137 -1593
rect 18199 -1600 18245 -1593
rect 18091 -1605 18245 -1600
rect 18091 -2297 18097 -1605
rect 18131 -1610 18205 -1605
rect 18131 -2297 18205 -2290
rect 18239 -2297 18245 -1605
rect 18091 -2300 18245 -2297
rect 18091 -2309 18137 -2300
rect 18199 -2309 18245 -2300
rect 18709 -1605 18755 -1593
rect 18709 -2297 18715 -1605
rect 18749 -2297 18755 -1605
rect 18709 -2309 18755 -2297
rect 19181 -1605 19227 -1593
rect 19181 -2297 19187 -1605
rect 19221 -2297 19227 -1605
rect 19181 -2309 19227 -2297
rect 19691 -1600 19737 -1593
rect 19799 -1600 19845 -1593
rect 19691 -1605 19845 -1600
rect 19691 -2297 19697 -1605
rect 19731 -1610 19805 -1605
rect 19731 -2297 19805 -2290
rect 19839 -2297 19845 -1605
rect 19691 -2300 19845 -2297
rect 19691 -2309 19737 -2300
rect 19799 -2309 19845 -2300
rect 20309 -1605 20355 -1593
rect 20309 -2297 20315 -1605
rect 20349 -2297 20355 -1605
rect 20309 -2309 20355 -2297
rect 20781 -1605 20827 -1593
rect 20781 -2297 20787 -1605
rect 20821 -2297 20827 -1605
rect 20781 -2309 20827 -2297
rect 21291 -1600 21337 -1593
rect 21399 -1600 21445 -1593
rect 21291 -1605 21445 -1600
rect 21291 -2297 21297 -1605
rect 21331 -1610 21405 -1605
rect 21331 -2297 21405 -2290
rect 21439 -2297 21445 -1605
rect 21291 -2300 21445 -2297
rect 21291 -2309 21337 -2300
rect 21399 -2309 21445 -2300
rect 21909 -1605 21955 -1593
rect 21909 -2297 21915 -1605
rect 21949 -2297 21955 -1605
rect 21909 -2309 21955 -2297
rect 22381 -1605 22427 -1593
rect 22381 -2297 22387 -1605
rect 22421 -2297 22427 -1605
rect 22381 -2309 22427 -2297
rect 22891 -1600 22937 -1593
rect 22999 -1600 23045 -1593
rect 22891 -1605 23045 -1600
rect 22891 -2297 22897 -1605
rect 22931 -1610 23005 -1605
rect 22931 -2297 23005 -2290
rect 23039 -2297 23045 -1605
rect 22891 -2300 23045 -2297
rect 22891 -2309 22937 -2300
rect 22999 -2309 23045 -2300
rect 23509 -1605 23555 -1593
rect 23509 -2297 23515 -1605
rect 23549 -2297 23555 -1605
rect 23509 -2309 23555 -2297
rect 23981 -1605 24027 -1593
rect 23981 -2297 23987 -1605
rect 24021 -2297 24027 -1605
rect 23981 -2309 24027 -2297
rect 24491 -1600 24537 -1593
rect 24599 -1600 24645 -1593
rect 24491 -1605 24645 -1600
rect 24491 -2297 24497 -1605
rect 24531 -1610 24605 -1605
rect 24531 -2297 24605 -2290
rect 24639 -2297 24645 -1605
rect 24491 -2300 24645 -2297
rect 24491 -2309 24537 -2300
rect 24599 -2309 24645 -2300
rect 25109 -1605 25155 -1593
rect 25109 -2297 25115 -1605
rect 25149 -2297 25155 -1605
rect 25109 -2309 25155 -2297
rect 25581 -1605 25627 -1593
rect 25581 -2297 25587 -1605
rect 25621 -2297 25627 -1605
rect 25581 -2309 25627 -2297
rect 26091 -1600 26137 -1593
rect 26199 -1600 26245 -1593
rect 26091 -1605 26245 -1600
rect 26091 -2297 26097 -1605
rect 26131 -1610 26205 -1605
rect 26131 -2297 26205 -2290
rect 26239 -2297 26245 -1605
rect 26091 -2300 26245 -2297
rect 26091 -2309 26137 -2300
rect 26199 -2309 26245 -2300
rect 26709 -1605 26755 -1593
rect 26709 -2297 26715 -1605
rect 26749 -2297 26755 -1605
rect 26709 -2309 26755 -2297
rect 27181 -1605 27227 -1593
rect 27181 -2297 27187 -1605
rect 27221 -2297 27227 -1605
rect 27181 -2309 27227 -2297
rect 27691 -1600 27737 -1593
rect 27799 -1600 27845 -1593
rect 27691 -1605 27845 -1600
rect 27691 -2297 27697 -1605
rect 27731 -1610 27805 -1605
rect 27731 -2297 27805 -2290
rect 27839 -2297 27845 -1605
rect 27691 -2300 27845 -2297
rect 27691 -2309 27737 -2300
rect 27799 -2309 27845 -2300
rect 28309 -1605 28355 -1593
rect 28309 -2297 28315 -1605
rect 28349 -2297 28355 -1605
rect 28309 -2309 28355 -2297
rect 28781 -1605 28827 -1593
rect 28781 -2297 28787 -1605
rect 28821 -2297 28827 -1605
rect 28781 -2309 28827 -2297
rect 29291 -1600 29337 -1593
rect 29399 -1600 29445 -1593
rect 29291 -1605 29445 -1600
rect 29291 -2297 29297 -1605
rect 29331 -1610 29405 -1605
rect 29331 -2297 29405 -2290
rect 29439 -2297 29445 -1605
rect 29291 -2300 29445 -2297
rect 29291 -2309 29337 -2300
rect 29399 -2309 29445 -2300
rect 29909 -1605 29955 -1593
rect 29909 -2297 29915 -1605
rect 29949 -2297 29955 -1605
rect 29909 -2309 29955 -2297
rect 30381 -1605 30427 -1593
rect 30381 -2297 30387 -1605
rect 30421 -2297 30427 -1605
rect 30381 -2309 30427 -2297
rect 30891 -1600 30937 -1593
rect 30999 -1600 31045 -1593
rect 30891 -1605 31045 -1600
rect 30891 -2297 30897 -1605
rect 30931 -1610 31005 -1605
rect 30931 -2297 31005 -2290
rect 31039 -2297 31045 -1605
rect 30891 -2300 31045 -2297
rect 30891 -2309 30937 -2300
rect 30999 -2309 31045 -2300
rect 31509 -1605 31555 -1593
rect 31509 -2297 31515 -1605
rect 31549 -2297 31555 -1605
rect 31509 -2309 31555 -2297
rect 31981 -1605 32027 -1593
rect 31981 -2297 31987 -1605
rect 32021 -2297 32027 -1605
rect 31981 -2309 32027 -2297
rect 32491 -1600 32537 -1593
rect 32599 -1600 32645 -1593
rect 32491 -1605 32645 -1600
rect 32491 -2297 32497 -1605
rect 32531 -1610 32605 -1605
rect 32531 -2297 32605 -2290
rect 32639 -2297 32645 -1605
rect 32491 -2300 32645 -2297
rect 32491 -2309 32537 -2300
rect 32599 -2309 32645 -2300
rect 33109 -1605 33155 -1593
rect 33350 -1600 33490 -1590
rect 35010 -1590 35020 -1540
rect 35140 -1499 35650 -1470
rect 35880 -1499 36270 -1420
rect 35140 -1505 35659 -1499
rect 35140 -1539 35271 -1505
rect 35647 -1539 35659 -1505
rect 35140 -1540 35659 -1539
rect 35140 -1570 35160 -1540
rect 35259 -1545 35659 -1540
rect 35877 -1505 36277 -1499
rect 35877 -1539 35889 -1505
rect 36265 -1539 36277 -1505
rect 35877 -1545 36277 -1539
rect 35140 -1590 35150 -1570
rect 33109 -2297 33115 -1605
rect 33149 -2297 33155 -1605
rect 33109 -2309 33155 -2297
rect 33581 -1605 33627 -1593
rect 33581 -2297 33587 -1605
rect 33621 -2297 33627 -1605
rect 33581 -2309 33627 -2297
rect 34091 -1600 34137 -1593
rect 34199 -1600 34245 -1593
rect 34091 -1605 34245 -1600
rect 34091 -2297 34097 -1605
rect 34131 -1610 34205 -1605
rect 34131 -2297 34205 -2290
rect 34239 -2297 34245 -1605
rect 34091 -2300 34245 -2297
rect 34091 -2309 34137 -2300
rect 34199 -2309 34245 -2300
rect 34709 -1605 34755 -1593
rect 35010 -1600 35150 -1590
rect 34709 -2297 34715 -1605
rect 34749 -2297 34755 -1605
rect 34709 -2309 34755 -2297
rect 35181 -1605 35227 -1593
rect 35181 -2297 35187 -1605
rect 35221 -2297 35227 -1605
rect 35181 -2309 35227 -2297
rect 35690 -1600 35760 -1590
rect 35750 -2310 35760 -1600
rect 35799 -1605 35845 -1593
rect 35799 -2297 35805 -1605
rect 35839 -1838 35845 -1605
rect 36018 -1838 36102 -1545
rect 36660 -1593 36800 -1420
rect 36859 -1505 37259 -1499
rect 36859 -1539 36871 -1505
rect 37247 -1539 37259 -1505
rect 36859 -1545 37259 -1539
rect 37300 -1593 37440 -1420
rect 37477 -1505 37877 -1499
rect 37477 -1539 37489 -1505
rect 37865 -1539 37877 -1505
rect 37477 -1545 37877 -1539
rect 37920 -1593 38060 -1420
rect 36309 -1605 36355 -1593
rect 36309 -1838 36315 -1605
rect 35839 -2016 36315 -1838
rect 35839 -2297 35845 -2016
rect 35799 -2309 35845 -2297
rect 35690 -2320 35760 -2310
rect 36018 -2357 36102 -2016
rect 36309 -2297 36315 -2016
rect 36349 -2297 36355 -1605
rect 36309 -2309 36355 -2297
rect 36660 -1605 36827 -1593
rect 36660 -2297 36787 -1605
rect 36821 -2297 36827 -1605
rect 36660 -2309 36827 -2297
rect 37291 -1605 37445 -1593
rect 37291 -2297 37297 -1605
rect 37331 -2297 37405 -1605
rect 37439 -2297 37445 -1605
rect 37291 -2309 37445 -2297
rect 37909 -1605 38060 -1593
rect 37909 -2297 37915 -1605
rect 37949 -2297 38060 -1605
rect 37909 -2309 38060 -2297
rect 660 -2363 1077 -2357
rect 660 -2397 689 -2363
rect 1065 -2397 1077 -2363
rect 660 -2403 1077 -2397
rect 1659 -2363 2059 -2357
rect 1659 -2397 1671 -2363
rect 2047 -2397 2059 -2363
rect 1659 -2403 2059 -2397
rect 2277 -2363 2677 -2357
rect 2277 -2397 2289 -2363
rect 2665 -2397 2677 -2363
rect 2277 -2403 2677 -2397
rect 3259 -2363 3659 -2357
rect 3259 -2397 3271 -2363
rect 3647 -2397 3659 -2363
rect 3259 -2403 3659 -2397
rect 3877 -2363 4277 -2357
rect 3877 -2397 3889 -2363
rect 4265 -2397 4277 -2363
rect 3877 -2403 4277 -2397
rect 4859 -2363 5259 -2357
rect 4859 -2397 4871 -2363
rect 5247 -2397 5259 -2363
rect 4859 -2403 5259 -2397
rect 5477 -2363 5877 -2357
rect 5477 -2397 5489 -2363
rect 5865 -2397 5877 -2363
rect 5477 -2403 5877 -2397
rect 6459 -2363 6859 -2357
rect 6459 -2397 6471 -2363
rect 6847 -2397 6859 -2363
rect 6459 -2403 6859 -2397
rect 7077 -2363 7477 -2357
rect 7077 -2397 7089 -2363
rect 7465 -2397 7477 -2363
rect 7077 -2403 7477 -2397
rect 8059 -2363 8459 -2357
rect 8059 -2397 8071 -2363
rect 8447 -2397 8459 -2363
rect 8059 -2403 8459 -2397
rect 8677 -2363 9077 -2357
rect 8677 -2397 8689 -2363
rect 9065 -2397 9077 -2363
rect 8677 -2403 9077 -2397
rect 9659 -2363 10059 -2357
rect 9659 -2397 9671 -2363
rect 10047 -2397 10059 -2363
rect 9659 -2403 10059 -2397
rect 10277 -2363 10677 -2357
rect 10277 -2397 10289 -2363
rect 10665 -2397 10677 -2363
rect 10277 -2403 10677 -2397
rect 11259 -2363 11659 -2357
rect 11259 -2397 11271 -2363
rect 11647 -2397 11659 -2363
rect 11259 -2403 11659 -2397
rect 11877 -2363 12277 -2357
rect 11877 -2397 11889 -2363
rect 12265 -2397 12277 -2363
rect 11877 -2403 12277 -2397
rect 12859 -2363 13259 -2357
rect 12859 -2397 12871 -2363
rect 13247 -2397 13259 -2363
rect 12859 -2403 13259 -2397
rect 13477 -2363 13877 -2357
rect 13477 -2397 13489 -2363
rect 13865 -2397 13877 -2363
rect 13477 -2403 13877 -2397
rect 14459 -2363 14859 -2357
rect 14459 -2397 14471 -2363
rect 14847 -2397 14859 -2363
rect 14459 -2403 14859 -2397
rect 15077 -2363 15477 -2357
rect 15077 -2397 15089 -2363
rect 15465 -2397 15477 -2363
rect 15077 -2403 15477 -2397
rect 16059 -2363 16459 -2357
rect 16059 -2397 16071 -2363
rect 16447 -2397 16459 -2363
rect 16059 -2403 16459 -2397
rect 16677 -2363 17077 -2357
rect 16677 -2397 16689 -2363
rect 17065 -2397 17077 -2363
rect 16677 -2403 17077 -2397
rect 17659 -2363 18059 -2357
rect 17659 -2397 17671 -2363
rect 18047 -2397 18059 -2363
rect 17659 -2403 18059 -2397
rect 18277 -2363 18677 -2357
rect 18277 -2397 18289 -2363
rect 18665 -2397 18677 -2363
rect 18277 -2403 18677 -2397
rect 19259 -2363 19659 -2357
rect 19259 -2397 19271 -2363
rect 19647 -2397 19659 -2363
rect 19259 -2403 19659 -2397
rect 19877 -2363 20277 -2357
rect 19877 -2397 19889 -2363
rect 20265 -2397 20277 -2363
rect 19877 -2403 20277 -2397
rect 20859 -2363 21259 -2357
rect 20859 -2397 20871 -2363
rect 21247 -2397 21259 -2363
rect 20859 -2403 21259 -2397
rect 21477 -2363 21877 -2357
rect 21477 -2397 21489 -2363
rect 21865 -2397 21877 -2363
rect 21477 -2403 21877 -2397
rect 22459 -2363 22859 -2357
rect 22459 -2397 22471 -2363
rect 22847 -2397 22859 -2363
rect 22459 -2403 22859 -2397
rect 23077 -2363 23477 -2357
rect 23077 -2397 23089 -2363
rect 23465 -2397 23477 -2363
rect 23077 -2403 23477 -2397
rect 24059 -2363 24459 -2357
rect 24059 -2397 24071 -2363
rect 24447 -2397 24459 -2363
rect 24059 -2403 24459 -2397
rect 24677 -2363 25077 -2357
rect 24677 -2397 24689 -2363
rect 25065 -2397 25077 -2363
rect 24677 -2403 25077 -2397
rect 25659 -2363 26059 -2357
rect 25659 -2397 25671 -2363
rect 26047 -2397 26059 -2363
rect 25659 -2403 26059 -2397
rect 26277 -2363 26677 -2357
rect 26277 -2397 26289 -2363
rect 26665 -2397 26677 -2363
rect 26277 -2403 26677 -2397
rect 27259 -2363 27659 -2357
rect 27259 -2397 27271 -2363
rect 27647 -2397 27659 -2363
rect 27259 -2403 27659 -2397
rect 27877 -2363 28277 -2357
rect 27877 -2397 27889 -2363
rect 28265 -2397 28277 -2363
rect 27877 -2403 28277 -2397
rect 28859 -2363 29259 -2357
rect 28859 -2397 28871 -2363
rect 29247 -2397 29259 -2363
rect 28859 -2403 29259 -2397
rect 29477 -2363 29877 -2357
rect 29477 -2397 29489 -2363
rect 29865 -2397 29877 -2363
rect 29477 -2403 29877 -2397
rect 30459 -2363 30859 -2357
rect 30459 -2397 30471 -2363
rect 30847 -2397 30859 -2363
rect 30459 -2403 30859 -2397
rect 31077 -2363 31477 -2357
rect 31077 -2397 31089 -2363
rect 31465 -2397 31477 -2363
rect 31077 -2403 31477 -2397
rect 32059 -2363 32459 -2357
rect 32059 -2397 32071 -2363
rect 32447 -2397 32459 -2363
rect 32059 -2403 32459 -2397
rect 32677 -2363 33077 -2357
rect 32677 -2397 32689 -2363
rect 33065 -2397 33077 -2363
rect 32677 -2403 33077 -2397
rect 33659 -2363 34059 -2357
rect 33659 -2397 33671 -2363
rect 34047 -2397 34059 -2363
rect 33659 -2403 34059 -2397
rect 34277 -2363 34677 -2357
rect 34277 -2397 34289 -2363
rect 34665 -2397 34677 -2363
rect 34277 -2403 34677 -2397
rect 35259 -2363 35659 -2357
rect 35259 -2397 35271 -2363
rect 35647 -2397 35659 -2363
rect 35259 -2403 35659 -2397
rect 35877 -2363 36277 -2357
rect 35877 -2397 35889 -2363
rect 36265 -2397 36277 -2363
rect 35877 -2403 36277 -2397
rect 660 -2645 710 -2403
rect 1680 -2440 2040 -2403
rect 2300 -2440 2660 -2403
rect 3280 -2440 3640 -2403
rect 3900 -2440 4260 -2403
rect 4880 -2440 5240 -2403
rect 5500 -2440 5860 -2403
rect 6480 -2440 6840 -2403
rect 7100 -2440 7460 -2403
rect 8080 -2440 8440 -2403
rect 8700 -2440 9060 -2403
rect 9680 -2440 10040 -2403
rect 10300 -2440 10660 -2403
rect 11280 -2440 11640 -2403
rect 11900 -2440 12260 -2403
rect 12880 -2440 13240 -2403
rect 13500 -2440 13860 -2403
rect 14480 -2440 14840 -2403
rect 15100 -2440 15460 -2403
rect 16080 -2440 16440 -2403
rect 16700 -2440 17060 -2403
rect 17680 -2440 18040 -2403
rect 18300 -2440 18660 -2403
rect 19280 -2440 19640 -2403
rect 19900 -2440 20260 -2403
rect 20880 -2440 21240 -2403
rect 21500 -2440 21860 -2403
rect 22480 -2440 22840 -2403
rect 23100 -2440 23460 -2403
rect 24080 -2440 24440 -2403
rect 24700 -2440 25060 -2403
rect 25680 -2440 26040 -2403
rect 26300 -2440 26660 -2403
rect 27280 -2440 27640 -2403
rect 27900 -2440 28260 -2403
rect 28880 -2440 29240 -2403
rect 29500 -2440 29860 -2403
rect 30480 -2440 30840 -2403
rect 31100 -2440 31460 -2403
rect 32080 -2440 32440 -2403
rect 32700 -2440 33060 -2403
rect 33680 -2440 34040 -2403
rect 34300 -2440 34660 -2403
rect 35280 -2440 35640 -2403
rect 1400 -2450 10660 -2440
rect 1400 -2570 1410 -2450
rect 1530 -2570 3010 -2450
rect 3130 -2570 4610 -2450
rect 4730 -2570 6210 -2450
rect 6330 -2570 7810 -2450
rect 7930 -2570 9410 -2450
rect 9530 -2570 10660 -2450
rect 1400 -2580 10660 -2570
rect 11260 -2580 12260 -2440
rect 12860 -2580 13860 -2440
rect 14460 -2580 15460 -2440
rect 15590 -2450 17060 -2440
rect 15590 -2570 15600 -2450
rect 15700 -2570 17060 -2450
rect 15590 -2580 17060 -2570
rect 17190 -2450 18660 -2440
rect 17190 -2570 17200 -2450
rect 17300 -2570 18660 -2450
rect 17190 -2580 18660 -2570
rect 18790 -2450 20260 -2440
rect 18790 -2570 18800 -2450
rect 18900 -2570 20260 -2450
rect 18790 -2580 20260 -2570
rect 20390 -2450 21860 -2440
rect 20390 -2570 20400 -2450
rect 20500 -2570 21860 -2450
rect 20390 -2580 21860 -2570
rect 21990 -2450 23460 -2440
rect 21990 -2570 22000 -2450
rect 22100 -2570 23460 -2450
rect 21990 -2580 23460 -2570
rect 23590 -2450 25060 -2440
rect 23590 -2570 23600 -2450
rect 23700 -2570 25060 -2450
rect 23590 -2580 25060 -2570
rect 25190 -2450 26660 -2440
rect 25190 -2570 25200 -2450
rect 25300 -2570 26660 -2450
rect 25190 -2580 26660 -2570
rect 26791 -2450 28260 -2440
rect 26791 -2570 26800 -2450
rect 26900 -2570 28260 -2450
rect 26791 -2580 28260 -2570
rect 28390 -2450 29860 -2440
rect 28390 -2570 28400 -2450
rect 28500 -2570 29860 -2450
rect 28390 -2580 29860 -2570
rect 29990 -2450 31460 -2440
rect 29990 -2570 30000 -2450
rect 30100 -2570 31460 -2450
rect 29990 -2580 31460 -2570
rect 32060 -2450 33310 -2440
rect 32060 -2570 33180 -2450
rect 33300 -2570 33310 -2450
rect 32060 -2580 33310 -2570
rect 33660 -2580 35640 -2440
rect 1680 -2645 2040 -2580
rect 2300 -2645 2660 -2580
rect 3280 -2645 3640 -2580
rect 3900 -2645 4260 -2580
rect 4880 -2645 5240 -2580
rect 5500 -2645 5860 -2580
rect 6480 -2645 6840 -2580
rect 7100 -2645 7460 -2580
rect 8080 -2645 8440 -2580
rect 8700 -2645 9060 -2580
rect 9680 -2645 10040 -2580
rect 10300 -2645 10660 -2580
rect 11280 -2625 11640 -2580
rect 11900 -2625 12260 -2580
rect 12880 -2625 13240 -2580
rect 13500 -2625 13860 -2580
rect 14480 -2625 14840 -2580
rect 15100 -2625 15460 -2580
rect 16080 -2625 16440 -2580
rect 16700 -2625 17060 -2580
rect 17680 -2625 18040 -2580
rect 18300 -2625 18660 -2580
rect 19280 -2625 19640 -2580
rect 19900 -2625 20260 -2580
rect 20880 -2625 21240 -2580
rect 21500 -2625 21860 -2580
rect 22480 -2625 22840 -2580
rect 23100 -2625 23460 -2580
rect 24080 -2625 24440 -2580
rect 24700 -2625 25060 -2580
rect 25680 -2625 26040 -2580
rect 26300 -2625 26660 -2580
rect 27280 -2625 27640 -2580
rect 27900 -2625 28260 -2580
rect 28880 -2625 29240 -2580
rect 29500 -2625 29860 -2580
rect 30480 -2625 30840 -2580
rect 31100 -2625 31460 -2580
rect 32080 -2625 32440 -2580
rect 32700 -2625 33060 -2580
rect 33680 -2625 34040 -2580
rect 34300 -2625 34660 -2580
rect 35280 -2625 35640 -2580
rect 11260 -2645 11659 -2625
rect 660 -2651 1077 -2645
rect 660 -2685 689 -2651
rect 1065 -2685 1077 -2651
rect 660 -2691 1077 -2685
rect 1659 -2651 2059 -2645
rect 1659 -2685 1671 -2651
rect 2047 -2685 2059 -2651
rect 1659 -2691 2059 -2685
rect 2277 -2651 2677 -2645
rect 2277 -2685 2289 -2651
rect 2665 -2685 2677 -2651
rect 2277 -2691 2677 -2685
rect 3259 -2651 3659 -2645
rect 3259 -2685 3271 -2651
rect 3647 -2685 3659 -2651
rect 3259 -2691 3659 -2685
rect 3877 -2651 4277 -2645
rect 3877 -2685 3889 -2651
rect 4265 -2685 4277 -2651
rect 3877 -2691 4277 -2685
rect 4859 -2651 5259 -2645
rect 4859 -2685 4871 -2651
rect 5247 -2685 5259 -2651
rect 4859 -2691 5259 -2685
rect 5477 -2651 5877 -2645
rect 5477 -2685 5489 -2651
rect 5865 -2685 5877 -2651
rect 5477 -2691 5877 -2685
rect 6459 -2651 6859 -2645
rect 6459 -2685 6471 -2651
rect 6847 -2685 6859 -2651
rect 6459 -2691 6859 -2685
rect 7077 -2651 7477 -2645
rect 7077 -2685 7089 -2651
rect 7465 -2685 7477 -2651
rect 7077 -2691 7477 -2685
rect 8059 -2651 8459 -2645
rect 8059 -2685 8071 -2651
rect 8447 -2685 8459 -2651
rect 8059 -2691 8459 -2685
rect 8677 -2651 9077 -2645
rect 8677 -2685 8689 -2651
rect 9065 -2685 9077 -2651
rect 8677 -2691 9077 -2685
rect 9659 -2651 10059 -2645
rect 9659 -2685 9671 -2651
rect 10047 -2685 10059 -2651
rect 9659 -2691 10059 -2685
rect 10277 -2651 10677 -2645
rect 10277 -2685 10289 -2651
rect 10665 -2685 10677 -2651
rect 10277 -2691 10677 -2685
rect 11259 -2651 11659 -2645
rect 11259 -2685 11271 -2651
rect 11647 -2685 11659 -2651
rect 11259 -2691 11659 -2685
rect 11877 -2651 12277 -2625
rect 12860 -2645 13259 -2625
rect 11877 -2685 11889 -2651
rect 12265 -2685 12277 -2651
rect 11877 -2691 12277 -2685
rect 12859 -2651 13259 -2645
rect 12859 -2685 12871 -2651
rect 13247 -2685 13259 -2651
rect 12859 -2691 13259 -2685
rect 13477 -2651 13877 -2625
rect 13477 -2685 13489 -2651
rect 13865 -2685 13877 -2651
rect 13477 -2691 13877 -2685
rect 14459 -2651 14859 -2625
rect 14459 -2685 14471 -2651
rect 14847 -2685 14859 -2651
rect 14459 -2691 14859 -2685
rect 15077 -2651 15477 -2625
rect 15077 -2685 15089 -2651
rect 15465 -2685 15477 -2651
rect 15077 -2691 15477 -2685
rect 16059 -2630 16459 -2625
rect 16059 -2651 16460 -2630
rect 16059 -2685 16071 -2651
rect 16447 -2685 16460 -2651
rect 16059 -2690 16460 -2685
rect 16677 -2651 17077 -2625
rect 16677 -2685 16689 -2651
rect 17065 -2685 17077 -2651
rect 16059 -2691 16459 -2690
rect 16677 -2691 17077 -2685
rect 17659 -2630 18059 -2625
rect 17659 -2651 18060 -2630
rect 17659 -2685 17671 -2651
rect 18047 -2685 18060 -2651
rect 17659 -2690 18060 -2685
rect 18277 -2651 18677 -2625
rect 18277 -2685 18289 -2651
rect 18665 -2685 18677 -2651
rect 17659 -2691 18059 -2690
rect 18277 -2691 18677 -2685
rect 19259 -2630 19659 -2625
rect 19259 -2651 19660 -2630
rect 19259 -2685 19271 -2651
rect 19647 -2685 19660 -2651
rect 19259 -2690 19660 -2685
rect 19877 -2651 20277 -2625
rect 19877 -2685 19889 -2651
rect 20265 -2685 20277 -2651
rect 19259 -2691 19659 -2690
rect 19877 -2691 20277 -2685
rect 20859 -2630 21259 -2625
rect 20859 -2651 21260 -2630
rect 20859 -2685 20871 -2651
rect 21247 -2685 21260 -2651
rect 20859 -2690 21260 -2685
rect 21477 -2651 21877 -2625
rect 21477 -2685 21489 -2651
rect 21865 -2685 21877 -2651
rect 20859 -2691 21259 -2690
rect 21477 -2691 21877 -2685
rect 22459 -2630 22859 -2625
rect 22459 -2651 22860 -2630
rect 22459 -2685 22471 -2651
rect 22847 -2685 22860 -2651
rect 22459 -2690 22860 -2685
rect 23077 -2651 23477 -2625
rect 23077 -2685 23089 -2651
rect 23465 -2685 23477 -2651
rect 22459 -2691 22859 -2690
rect 23077 -2691 23477 -2685
rect 24059 -2630 24459 -2625
rect 24059 -2651 24460 -2630
rect 24059 -2685 24071 -2651
rect 24447 -2685 24460 -2651
rect 24059 -2690 24460 -2685
rect 24677 -2651 25077 -2625
rect 24677 -2685 24689 -2651
rect 25065 -2685 25077 -2651
rect 24059 -2691 24459 -2690
rect 24677 -2691 25077 -2685
rect 25659 -2630 26059 -2625
rect 25659 -2651 26060 -2630
rect 25659 -2685 25671 -2651
rect 26047 -2685 26060 -2651
rect 25659 -2690 26060 -2685
rect 26277 -2651 26677 -2625
rect 26277 -2685 26289 -2651
rect 26665 -2685 26677 -2651
rect 25659 -2691 26059 -2690
rect 26277 -2691 26677 -2685
rect 27259 -2630 27659 -2625
rect 27259 -2651 27660 -2630
rect 27259 -2685 27271 -2651
rect 27647 -2685 27660 -2651
rect 27259 -2690 27660 -2685
rect 27877 -2651 28277 -2625
rect 27877 -2685 27889 -2651
rect 28265 -2685 28277 -2651
rect 27259 -2691 27659 -2690
rect 27877 -2691 28277 -2685
rect 28859 -2630 29259 -2625
rect 28859 -2651 29260 -2630
rect 28859 -2685 28871 -2651
rect 29247 -2685 29260 -2651
rect 28859 -2690 29260 -2685
rect 29477 -2651 29877 -2625
rect 29477 -2685 29489 -2651
rect 29865 -2685 29877 -2651
rect 28859 -2691 29259 -2690
rect 29477 -2691 29877 -2685
rect 30459 -2630 30859 -2625
rect 30459 -2651 30860 -2630
rect 30459 -2685 30471 -2651
rect 30847 -2685 30860 -2651
rect 30459 -2690 30860 -2685
rect 31077 -2651 31477 -2625
rect 32060 -2630 32459 -2625
rect 32060 -2645 32460 -2630
rect 31077 -2685 31089 -2651
rect 31465 -2685 31477 -2651
rect 30459 -2691 30859 -2690
rect 31077 -2691 31477 -2685
rect 32059 -2651 32460 -2645
rect 32059 -2685 32071 -2651
rect 32447 -2685 32460 -2651
rect 32059 -2690 32460 -2685
rect 32677 -2651 33077 -2625
rect 32677 -2685 32689 -2651
rect 33065 -2685 33077 -2651
rect 32059 -2691 32459 -2690
rect 32677 -2691 33077 -2685
rect 33659 -2630 34059 -2625
rect 33659 -2651 34060 -2630
rect 33659 -2685 33671 -2651
rect 34047 -2685 34060 -2651
rect 33659 -2690 34060 -2685
rect 34277 -2651 34677 -2625
rect 34277 -2685 34289 -2651
rect 34665 -2685 34677 -2651
rect 33659 -2691 34059 -2690
rect 34277 -2691 34677 -2685
rect 35259 -2630 35659 -2625
rect 35259 -2651 35660 -2630
rect 35259 -2685 35271 -2651
rect 35647 -2685 35660 -2651
rect 35259 -2690 35660 -2685
rect 35877 -2651 36277 -2645
rect 35877 -2685 35889 -2651
rect 36265 -2685 36277 -2651
rect 35259 -2691 35659 -2690
rect 35877 -2691 36277 -2685
rect 59 -2909 480 -2903
rect 59 -2943 71 -2909
rect 447 -2943 480 -2909
rect 59 -2949 480 -2943
rect 440 -3140 480 -2949
rect -140 -3171 480 -3140
rect 660 -2903 710 -2691
rect 1109 -2730 1155 -2718
rect 1581 -2730 1627 -2718
rect 2091 -2730 2137 -2718
rect 2199 -2730 2245 -2718
rect 2709 -2730 2755 -2718
rect 3181 -2730 3227 -2718
rect 3691 -2730 3737 -2718
rect 3799 -2730 3845 -2718
rect 4309 -2730 4355 -2718
rect 4781 -2730 4827 -2718
rect 5291 -2730 5337 -2718
rect 5399 -2730 5445 -2718
rect 5909 -2730 5955 -2718
rect 6381 -2730 6427 -2718
rect 6891 -2730 6937 -2718
rect 6999 -2730 7045 -2718
rect 7509 -2730 7555 -2718
rect 7981 -2730 8027 -2718
rect 8491 -2730 8537 -2718
rect 8599 -2730 8645 -2718
rect 9109 -2730 9155 -2718
rect 9581 -2730 9627 -2718
rect 10091 -2730 10137 -2718
rect 10199 -2730 10245 -2718
rect 10709 -2730 10755 -2718
rect 11181 -2730 11227 -2718
rect 11691 -2730 11737 -2718
rect 11799 -2730 11845 -2718
rect 12309 -2720 12355 -2718
rect 12309 -2730 12520 -2720
rect 12781 -2730 12827 -2718
rect 13291 -2730 13337 -2718
rect 13399 -2730 13445 -2718
rect 13909 -2730 13955 -2718
rect 14381 -2730 14427 -2718
rect 14891 -2730 14937 -2718
rect 14999 -2730 15045 -2718
rect 15509 -2730 15555 -2718
rect 15981 -2730 16027 -2718
rect 16491 -2730 16537 -2718
rect 16599 -2730 16645 -2718
rect 17109 -2730 17155 -2718
rect 17581 -2730 17627 -2718
rect 18091 -2730 18137 -2718
rect 18199 -2730 18245 -2718
rect 18709 -2730 18755 -2718
rect 19181 -2730 19227 -2718
rect 19691 -2730 19737 -2718
rect 19799 -2730 19845 -2718
rect 20309 -2730 20355 -2718
rect 20781 -2730 20827 -2718
rect 21291 -2730 21337 -2718
rect 21399 -2730 21445 -2718
rect 21909 -2730 21955 -2718
rect 22381 -2730 22427 -2718
rect 22891 -2730 22937 -2718
rect 22999 -2730 23045 -2718
rect 23509 -2730 23555 -2718
rect 23981 -2730 24027 -2718
rect 24491 -2730 24537 -2718
rect 24599 -2730 24645 -2718
rect 25109 -2730 25155 -2718
rect 25581 -2730 25627 -2718
rect 26091 -2730 26137 -2718
rect 26199 -2730 26245 -2718
rect 26709 -2730 26755 -2718
rect 27181 -2730 27227 -2718
rect 27691 -2730 27737 -2718
rect 27799 -2730 27845 -2718
rect 28309 -2730 28355 -2718
rect 28781 -2730 28827 -2718
rect 29291 -2730 29337 -2718
rect 29399 -2730 29445 -2718
rect 29909 -2730 29955 -2718
rect 30381 -2730 30427 -2718
rect 30891 -2730 30937 -2718
rect 30999 -2730 31045 -2718
rect 31509 -2730 31555 -2718
rect 31981 -2730 32027 -2718
rect 32491 -2730 32537 -2718
rect 32599 -2730 32645 -2718
rect 33109 -2730 33155 -2718
rect 33581 -2730 33627 -2718
rect 34091 -2730 34137 -2718
rect 34199 -2730 34245 -2718
rect 34709 -2730 34755 -2718
rect 35181 -2730 35227 -2718
rect 35691 -2730 35737 -2718
rect 35799 -2730 35845 -2718
rect 36026 -2730 36116 -2691
rect 36660 -2718 36800 -2309
rect 36859 -2363 37259 -2357
rect 36859 -2397 36871 -2363
rect 37247 -2397 37259 -2363
rect 36859 -2403 37259 -2397
rect 36859 -2651 37259 -2645
rect 36859 -2685 36871 -2651
rect 37247 -2685 37259 -2651
rect 36859 -2691 37259 -2685
rect 37300 -2718 37440 -2309
rect 37477 -2363 37877 -2357
rect 37477 -2397 37489 -2363
rect 37865 -2397 37877 -2363
rect 37477 -2403 37877 -2397
rect 37477 -2651 37877 -2645
rect 37477 -2685 37489 -2651
rect 37865 -2685 37877 -2651
rect 37477 -2691 37877 -2685
rect 37920 -2718 38060 -2309
rect 36309 -2730 36355 -2718
rect 36660 -2730 36827 -2718
rect 1109 -2864 1115 -2730
rect 1149 -2864 1155 -2730
rect 1540 -2860 1587 -2730
rect 1109 -2876 1155 -2864
rect 1581 -2864 1587 -2860
rect 1621 -2860 2097 -2730
rect 1621 -2864 1627 -2860
rect 1581 -2876 1627 -2864
rect 2091 -2864 2097 -2860
rect 2131 -2860 2205 -2730
rect 2131 -2864 2137 -2860
rect 2091 -2876 2137 -2864
rect 2199 -2864 2205 -2860
rect 2239 -2860 2715 -2730
rect 2239 -2864 2245 -2860
rect 2199 -2876 2245 -2864
rect 2709 -2864 2715 -2860
rect 2749 -2860 3187 -2730
rect 2749 -2864 2755 -2860
rect 2709 -2876 2755 -2864
rect 3181 -2864 3187 -2860
rect 3221 -2860 3697 -2730
rect 3221 -2864 3227 -2860
rect 3181 -2876 3227 -2864
rect 3691 -2864 3697 -2860
rect 3731 -2860 3805 -2730
rect 3731 -2864 3737 -2860
rect 3691 -2876 3737 -2864
rect 3799 -2864 3805 -2860
rect 3839 -2860 4315 -2730
rect 3839 -2864 3845 -2860
rect 3799 -2876 3845 -2864
rect 4309 -2864 4315 -2860
rect 4349 -2860 4787 -2730
rect 4349 -2864 4355 -2860
rect 4309 -2876 4355 -2864
rect 4781 -2864 4787 -2860
rect 4821 -2860 5297 -2730
rect 4821 -2864 4827 -2860
rect 4781 -2876 4827 -2864
rect 5291 -2864 5297 -2860
rect 5331 -2860 5405 -2730
rect 5331 -2864 5337 -2860
rect 5291 -2876 5337 -2864
rect 5399 -2864 5405 -2860
rect 5439 -2860 5915 -2730
rect 5439 -2864 5445 -2860
rect 5399 -2876 5445 -2864
rect 5909 -2864 5915 -2860
rect 5949 -2860 6387 -2730
rect 5949 -2864 5955 -2860
rect 5909 -2876 5955 -2864
rect 6381 -2864 6387 -2860
rect 6421 -2860 6897 -2730
rect 6421 -2864 6427 -2860
rect 6381 -2876 6427 -2864
rect 6891 -2864 6897 -2860
rect 6931 -2860 7005 -2730
rect 6931 -2864 6937 -2860
rect 6891 -2876 6937 -2864
rect 6999 -2864 7005 -2860
rect 7039 -2860 7515 -2730
rect 7039 -2864 7045 -2860
rect 6999 -2876 7045 -2864
rect 7509 -2864 7515 -2860
rect 7549 -2860 7987 -2730
rect 7549 -2864 7555 -2860
rect 7509 -2876 7555 -2864
rect 7981 -2864 7987 -2860
rect 8021 -2860 8497 -2730
rect 8021 -2864 8027 -2860
rect 7981 -2876 8027 -2864
rect 8491 -2864 8497 -2860
rect 8531 -2860 8605 -2730
rect 8531 -2864 8537 -2860
rect 8491 -2876 8537 -2864
rect 8599 -2864 8605 -2860
rect 8639 -2860 9115 -2730
rect 8639 -2864 8645 -2860
rect 8599 -2876 8645 -2864
rect 9109 -2864 9115 -2860
rect 9149 -2860 9587 -2730
rect 9149 -2864 9155 -2860
rect 9109 -2876 9155 -2864
rect 9581 -2864 9587 -2860
rect 9621 -2860 10097 -2730
rect 9621 -2864 9627 -2860
rect 9581 -2876 9627 -2864
rect 10091 -2864 10097 -2860
rect 10131 -2860 10205 -2730
rect 10131 -2864 10137 -2860
rect 10091 -2876 10137 -2864
rect 10199 -2864 10205 -2860
rect 10239 -2860 10715 -2730
rect 10239 -2864 10245 -2860
rect 10199 -2876 10245 -2864
rect 10709 -2864 10715 -2860
rect 10749 -2860 11187 -2730
rect 10749 -2864 10755 -2860
rect 10709 -2876 10755 -2864
rect 11181 -2864 11187 -2860
rect 11221 -2860 11697 -2730
rect 11221 -2864 11227 -2860
rect 11181 -2876 11227 -2864
rect 11691 -2864 11697 -2860
rect 11731 -2860 11805 -2730
rect 11731 -2864 11737 -2860
rect 11691 -2876 11737 -2864
rect 11799 -2864 11805 -2860
rect 11839 -2860 12315 -2730
rect 11839 -2864 11845 -2860
rect 11799 -2876 11845 -2864
rect 12309 -2864 12315 -2860
rect 12349 -2850 12390 -2730
rect 12510 -2850 12787 -2730
rect 12349 -2860 12787 -2850
rect 12349 -2864 12355 -2860
rect 12309 -2876 12355 -2864
rect 12781 -2864 12787 -2860
rect 12821 -2860 13297 -2730
rect 12821 -2864 12827 -2860
rect 12781 -2876 12827 -2864
rect 13291 -2864 13297 -2860
rect 13331 -2860 13405 -2730
rect 13331 -2864 13337 -2860
rect 13291 -2876 13337 -2864
rect 13399 -2864 13405 -2860
rect 13439 -2860 13915 -2730
rect 13439 -2864 13445 -2860
rect 13399 -2876 13445 -2864
rect 13909 -2864 13915 -2860
rect 13949 -2860 14387 -2730
rect 13949 -2864 13955 -2860
rect 13909 -2876 13955 -2864
rect 14381 -2864 14387 -2860
rect 14421 -2860 14897 -2730
rect 14421 -2864 14427 -2860
rect 14381 -2876 14427 -2864
rect 14891 -2864 14897 -2860
rect 14931 -2860 15005 -2730
rect 14931 -2864 14937 -2860
rect 14891 -2876 14937 -2864
rect 14999 -2864 15005 -2860
rect 15039 -2860 15515 -2730
rect 15039 -2864 15045 -2860
rect 14999 -2876 15045 -2864
rect 15509 -2864 15515 -2860
rect 15549 -2860 15987 -2730
rect 15549 -2864 15555 -2860
rect 15509 -2876 15555 -2864
rect 15981 -2864 15987 -2860
rect 16021 -2860 16497 -2730
rect 16021 -2864 16027 -2860
rect 15981 -2876 16027 -2864
rect 16491 -2864 16497 -2860
rect 16531 -2860 16605 -2730
rect 16531 -2864 16537 -2860
rect 16491 -2876 16537 -2864
rect 16599 -2864 16605 -2860
rect 16639 -2860 17115 -2730
rect 16639 -2864 16645 -2860
rect 16599 -2876 16645 -2864
rect 17109 -2864 17115 -2860
rect 17149 -2860 17587 -2730
rect 17149 -2864 17155 -2860
rect 17109 -2876 17155 -2864
rect 17581 -2864 17587 -2860
rect 17621 -2860 18097 -2730
rect 17621 -2864 17627 -2860
rect 17581 -2876 17627 -2864
rect 18091 -2864 18097 -2860
rect 18131 -2860 18205 -2730
rect 18131 -2864 18137 -2860
rect 18091 -2876 18137 -2864
rect 18199 -2864 18205 -2860
rect 18239 -2860 18715 -2730
rect 18239 -2864 18245 -2860
rect 18199 -2876 18245 -2864
rect 18709 -2864 18715 -2860
rect 18749 -2860 19187 -2730
rect 18749 -2864 18755 -2860
rect 18709 -2876 18755 -2864
rect 19181 -2864 19187 -2860
rect 19221 -2860 19697 -2730
rect 19221 -2864 19227 -2860
rect 19181 -2876 19227 -2864
rect 19691 -2864 19697 -2860
rect 19731 -2860 19805 -2730
rect 19731 -2864 19737 -2860
rect 19691 -2876 19737 -2864
rect 19799 -2864 19805 -2860
rect 19839 -2860 20315 -2730
rect 19839 -2864 19845 -2860
rect 19799 -2876 19845 -2864
rect 20309 -2864 20315 -2860
rect 20349 -2860 20787 -2730
rect 20349 -2864 20355 -2860
rect 20309 -2876 20355 -2864
rect 20781 -2864 20787 -2860
rect 20821 -2860 21297 -2730
rect 20821 -2864 20827 -2860
rect 20781 -2876 20827 -2864
rect 21291 -2864 21297 -2860
rect 21331 -2860 21405 -2730
rect 21331 -2864 21337 -2860
rect 21291 -2876 21337 -2864
rect 21399 -2864 21405 -2860
rect 21439 -2860 21915 -2730
rect 21439 -2864 21445 -2860
rect 21399 -2876 21445 -2864
rect 21909 -2864 21915 -2860
rect 21949 -2860 22387 -2730
rect 21949 -2864 21955 -2860
rect 21909 -2876 21955 -2864
rect 22381 -2864 22387 -2860
rect 22421 -2860 22897 -2730
rect 22421 -2864 22427 -2860
rect 22381 -2876 22427 -2864
rect 22891 -2864 22897 -2860
rect 22931 -2860 23005 -2730
rect 22931 -2864 22937 -2860
rect 22891 -2876 22937 -2864
rect 22999 -2864 23005 -2860
rect 23039 -2860 23515 -2730
rect 23039 -2864 23045 -2860
rect 22999 -2876 23045 -2864
rect 23509 -2864 23515 -2860
rect 23549 -2860 23987 -2730
rect 23549 -2864 23555 -2860
rect 23509 -2876 23555 -2864
rect 23981 -2864 23987 -2860
rect 24021 -2860 24497 -2730
rect 24021 -2864 24027 -2860
rect 23981 -2876 24027 -2864
rect 24491 -2864 24497 -2860
rect 24531 -2860 24605 -2730
rect 24531 -2864 24537 -2860
rect 24491 -2876 24537 -2864
rect 24599 -2864 24605 -2860
rect 24639 -2860 25115 -2730
rect 24639 -2864 24645 -2860
rect 24599 -2876 24645 -2864
rect 25109 -2864 25115 -2860
rect 25149 -2860 25587 -2730
rect 25149 -2864 25155 -2860
rect 25109 -2876 25155 -2864
rect 25581 -2864 25587 -2860
rect 25621 -2860 26097 -2730
rect 25621 -2864 25627 -2860
rect 25581 -2876 25627 -2864
rect 26091 -2864 26097 -2860
rect 26131 -2860 26205 -2730
rect 26131 -2864 26137 -2860
rect 26091 -2876 26137 -2864
rect 26199 -2864 26205 -2860
rect 26239 -2860 26715 -2730
rect 26239 -2864 26245 -2860
rect 26199 -2876 26245 -2864
rect 26709 -2864 26715 -2860
rect 26749 -2860 27187 -2730
rect 26749 -2864 26755 -2860
rect 26709 -2876 26755 -2864
rect 27181 -2864 27187 -2860
rect 27221 -2860 27697 -2730
rect 27221 -2864 27227 -2860
rect 27181 -2876 27227 -2864
rect 27691 -2864 27697 -2860
rect 27731 -2860 27805 -2730
rect 27731 -2864 27737 -2860
rect 27691 -2876 27737 -2864
rect 27799 -2864 27805 -2860
rect 27839 -2860 28315 -2730
rect 27839 -2864 27845 -2860
rect 27799 -2876 27845 -2864
rect 28309 -2864 28315 -2860
rect 28349 -2860 28787 -2730
rect 28349 -2864 28355 -2860
rect 28309 -2876 28355 -2864
rect 28781 -2864 28787 -2860
rect 28821 -2860 29297 -2730
rect 28821 -2864 28827 -2860
rect 28781 -2876 28827 -2864
rect 29291 -2864 29297 -2860
rect 29331 -2860 29405 -2730
rect 29331 -2864 29337 -2860
rect 29291 -2876 29337 -2864
rect 29399 -2864 29405 -2860
rect 29439 -2860 29915 -2730
rect 29439 -2864 29445 -2860
rect 29399 -2876 29445 -2864
rect 29909 -2864 29915 -2860
rect 29949 -2860 30387 -2730
rect 29949 -2864 29955 -2860
rect 29909 -2876 29955 -2864
rect 30381 -2864 30387 -2860
rect 30421 -2860 30897 -2730
rect 30421 -2864 30427 -2860
rect 30381 -2876 30427 -2864
rect 30891 -2864 30897 -2860
rect 30931 -2860 31005 -2730
rect 30931 -2864 30937 -2860
rect 30891 -2876 30937 -2864
rect 30999 -2864 31005 -2860
rect 31039 -2860 31515 -2730
rect 31039 -2864 31045 -2860
rect 30999 -2876 31045 -2864
rect 31509 -2864 31515 -2860
rect 31549 -2860 31987 -2730
rect 31549 -2864 31555 -2860
rect 31509 -2876 31555 -2864
rect 31981 -2864 31987 -2860
rect 32021 -2860 32497 -2730
rect 32021 -2864 32027 -2860
rect 31981 -2876 32027 -2864
rect 32491 -2864 32497 -2860
rect 32531 -2860 32605 -2730
rect 32531 -2864 32537 -2860
rect 32491 -2876 32537 -2864
rect 32599 -2864 32605 -2860
rect 32639 -2860 33115 -2730
rect 32639 -2864 32645 -2860
rect 32599 -2876 32645 -2864
rect 33109 -2864 33115 -2860
rect 33149 -2860 33587 -2730
rect 33149 -2864 33155 -2860
rect 33109 -2876 33155 -2864
rect 33581 -2864 33587 -2860
rect 33621 -2860 34097 -2730
rect 33621 -2864 33627 -2860
rect 33581 -2876 33627 -2864
rect 34091 -2864 34097 -2860
rect 34131 -2860 34205 -2730
rect 34131 -2864 34137 -2860
rect 34091 -2876 34137 -2864
rect 34199 -2864 34205 -2860
rect 34239 -2860 34715 -2730
rect 34239 -2864 34245 -2860
rect 34199 -2876 34245 -2864
rect 34709 -2864 34715 -2860
rect 34749 -2860 35187 -2730
rect 34749 -2864 34755 -2860
rect 34709 -2876 34755 -2864
rect 35181 -2864 35187 -2860
rect 35221 -2860 35697 -2730
rect 35221 -2864 35227 -2860
rect 35181 -2876 35227 -2864
rect 35691 -2864 35697 -2860
rect 35731 -2860 35805 -2730
rect 35731 -2864 35737 -2860
rect 35691 -2876 35737 -2864
rect 35799 -2864 35805 -2860
rect 35839 -2860 36315 -2730
rect 35839 -2864 35845 -2860
rect 35799 -2876 35845 -2864
rect 36026 -2903 36116 -2860
rect 36309 -2864 36315 -2860
rect 36349 -2860 36400 -2730
rect 36349 -2864 36355 -2860
rect 36309 -2876 36355 -2864
rect 36660 -2864 36787 -2730
rect 36821 -2864 36827 -2730
rect 36660 -2876 36827 -2864
rect 37291 -2730 37445 -2718
rect 37291 -2864 37297 -2730
rect 37331 -2864 37405 -2730
rect 37439 -2864 37445 -2730
rect 37291 -2876 37445 -2864
rect 37909 -2730 38060 -2718
rect 37909 -2864 37915 -2730
rect 37949 -2864 38060 -2730
rect 37909 -2876 38060 -2864
rect 660 -2909 1077 -2903
rect 660 -2943 689 -2909
rect 1065 -2943 1077 -2909
rect 1659 -2909 2059 -2903
rect 660 -2949 1077 -2943
rect 1180 -2920 1320 -2910
rect 1659 -2920 1671 -2909
rect 660 -3140 710 -2949
rect 1180 -3040 1190 -2920
rect 1310 -2943 1671 -2920
rect 2047 -2920 2059 -2909
rect 2277 -2909 2677 -2903
rect 2277 -2920 2289 -2909
rect 2047 -2943 2289 -2920
rect 2665 -2920 2677 -2909
rect 3259 -2909 3659 -2903
rect 2780 -2920 2920 -2910
rect 3259 -2920 3271 -2909
rect 2665 -2943 2790 -2920
rect 1310 -3040 2790 -2943
rect 2910 -2943 3271 -2920
rect 3647 -2920 3659 -2909
rect 3877 -2909 4277 -2903
rect 3877 -2920 3889 -2909
rect 3647 -2943 3889 -2920
rect 4265 -2920 4277 -2909
rect 4859 -2909 5259 -2903
rect 4380 -2920 4520 -2910
rect 4859 -2920 4871 -2909
rect 4265 -2943 4390 -2920
rect 2910 -3040 4390 -2943
rect 4510 -2943 4871 -2920
rect 5247 -2920 5259 -2909
rect 5477 -2909 5877 -2903
rect 5477 -2920 5489 -2909
rect 5247 -2943 5489 -2920
rect 5865 -2920 5877 -2909
rect 6459 -2909 6859 -2903
rect 5980 -2920 6120 -2910
rect 6459 -2920 6471 -2909
rect 5865 -2943 5990 -2920
rect 4510 -3040 5990 -2943
rect 6110 -2943 6471 -2920
rect 6847 -2920 6859 -2909
rect 7077 -2909 7477 -2903
rect 7077 -2920 7089 -2909
rect 6847 -2943 7089 -2920
rect 7465 -2920 7477 -2909
rect 8059 -2909 8459 -2903
rect 7580 -2920 7720 -2910
rect 8059 -2920 8071 -2909
rect 7465 -2943 7590 -2920
rect 6110 -3040 7590 -2943
rect 7710 -2943 8071 -2920
rect 8447 -2920 8459 -2909
rect 8677 -2909 9077 -2903
rect 8677 -2920 8689 -2909
rect 8447 -2943 8689 -2920
rect 9065 -2920 9077 -2909
rect 9659 -2909 10059 -2903
rect 9180 -2920 9320 -2910
rect 9659 -2920 9671 -2909
rect 9065 -2943 9190 -2920
rect 7710 -3040 9190 -2943
rect 9310 -2943 9671 -2920
rect 10047 -2920 10059 -2909
rect 10277 -2909 10677 -2903
rect 10277 -2920 10289 -2909
rect 10047 -2943 10289 -2920
rect 10665 -2920 10677 -2909
rect 11259 -2909 11659 -2903
rect 11000 -2920 11140 -2910
rect 11259 -2920 11271 -2909
rect 10665 -2943 10720 -2920
rect 9310 -3040 10720 -2943
rect 11000 -3040 11010 -2920
rect 11130 -2943 11271 -2920
rect 11647 -2920 11659 -2909
rect 11877 -2909 12277 -2903
rect 11877 -2920 11889 -2909
rect 11647 -2943 11889 -2920
rect 12265 -2920 12277 -2909
rect 12859 -2909 13259 -2903
rect 12859 -2920 12871 -2909
rect 12265 -2943 12320 -2920
rect 11130 -3040 12320 -2943
rect 12820 -2943 12871 -2920
rect 13247 -2920 13259 -2909
rect 13477 -2909 13877 -2903
rect 13477 -2920 13489 -2909
rect 13247 -2943 13489 -2920
rect 13865 -2920 13877 -2909
rect 14459 -2909 14859 -2903
rect 14459 -2910 14471 -2909
rect 14200 -2920 14340 -2910
rect 13865 -2943 14210 -2920
rect 12820 -3040 14210 -2943
rect 14330 -3040 14340 -2920
rect 1180 -3050 1320 -3040
rect 2780 -3050 2920 -3040
rect 4380 -3050 4520 -3040
rect 5980 -3050 6120 -3040
rect 7580 -3050 7720 -3040
rect 9180 -3050 9320 -3040
rect 11000 -3050 11140 -3040
rect 14200 -3050 14340 -3040
rect 14420 -2920 14471 -2910
rect 14847 -2920 14859 -2909
rect 15077 -2909 15477 -2903
rect 15077 -2920 15089 -2909
rect 14420 -3040 14430 -2920
rect 14847 -2943 15089 -2920
rect 15465 -2920 15477 -2909
rect 16059 -2909 16459 -2903
rect 15810 -2920 15930 -2910
rect 16059 -2920 16071 -2909
rect 15465 -2943 15520 -2920
rect 14550 -3040 15520 -2943
rect 15810 -3040 15820 -2920
rect 15920 -2943 16071 -2920
rect 16447 -2920 16459 -2909
rect 16677 -2909 17077 -2903
rect 16677 -2920 16689 -2909
rect 16447 -2943 16689 -2920
rect 17065 -2920 17077 -2909
rect 17659 -2909 18059 -2903
rect 17410 -2920 17530 -2910
rect 17659 -2920 17671 -2909
rect 17065 -2943 17120 -2920
rect 15920 -3040 17120 -2943
rect 17410 -3040 17420 -2920
rect 17520 -2943 17671 -2920
rect 18047 -2920 18059 -2909
rect 18277 -2909 18677 -2903
rect 18277 -2920 18289 -2909
rect 18047 -2943 18289 -2920
rect 18665 -2920 18677 -2909
rect 19259 -2909 19659 -2903
rect 19010 -2920 19130 -2910
rect 19259 -2920 19271 -2909
rect 18665 -2943 18720 -2920
rect 17520 -3040 18720 -2943
rect 19010 -3040 19020 -2920
rect 19120 -2943 19271 -2920
rect 19647 -2920 19659 -2909
rect 19877 -2909 20277 -2903
rect 19877 -2920 19889 -2909
rect 19647 -2943 19889 -2920
rect 20265 -2920 20277 -2909
rect 20859 -2909 21259 -2903
rect 20610 -2920 20730 -2910
rect 20859 -2920 20871 -2909
rect 20265 -2943 20320 -2920
rect 19120 -3040 20320 -2943
rect 20610 -3040 20620 -2920
rect 20720 -2943 20871 -2920
rect 21247 -2920 21259 -2909
rect 21477 -2909 21877 -2903
rect 21477 -2920 21489 -2909
rect 21247 -2943 21489 -2920
rect 21865 -2920 21877 -2909
rect 22459 -2909 22859 -2903
rect 22210 -2920 22330 -2910
rect 22459 -2920 22471 -2909
rect 21865 -2943 21920 -2920
rect 20720 -3040 21920 -2943
rect 22210 -3040 22220 -2920
rect 22320 -2943 22471 -2920
rect 22847 -2920 22859 -2909
rect 23077 -2909 23477 -2903
rect 23077 -2920 23089 -2909
rect 22847 -2943 23089 -2920
rect 23465 -2920 23477 -2909
rect 24059 -2909 24459 -2903
rect 23810 -2920 23930 -2910
rect 24059 -2920 24071 -2909
rect 23465 -2943 23520 -2920
rect 22320 -3040 23520 -2943
rect 23810 -3040 23820 -2920
rect 23920 -2943 24071 -2920
rect 24447 -2920 24459 -2909
rect 24677 -2909 25077 -2903
rect 24677 -2920 24689 -2909
rect 24447 -2943 24689 -2920
rect 25065 -2920 25077 -2909
rect 25659 -2909 26059 -2903
rect 25410 -2920 25530 -2910
rect 25659 -2920 25671 -2909
rect 25065 -2943 25120 -2920
rect 23920 -3040 25120 -2943
rect 25410 -3040 25420 -2920
rect 25520 -2943 25671 -2920
rect 26047 -2920 26059 -2909
rect 26277 -2909 26677 -2903
rect 26277 -2920 26289 -2909
rect 26047 -2943 26289 -2920
rect 26665 -2920 26677 -2909
rect 27259 -2909 27659 -2903
rect 27011 -2920 27130 -2910
rect 27259 -2920 27271 -2909
rect 26665 -2943 26720 -2920
rect 25520 -3040 26720 -2943
rect 27011 -3040 27020 -2920
rect 27120 -2943 27271 -2920
rect 27647 -2920 27659 -2909
rect 27877 -2909 28277 -2903
rect 27877 -2920 27889 -2909
rect 27647 -2943 27889 -2920
rect 28265 -2920 28277 -2909
rect 28859 -2909 29259 -2903
rect 28859 -2910 28871 -2909
rect 28610 -2920 28871 -2910
rect 28265 -2943 28320 -2920
rect 27120 -3040 28320 -2943
rect 28610 -3040 28620 -2920
rect 28720 -2943 28871 -2920
rect 29247 -2910 29259 -2909
rect 29477 -2909 29877 -2903
rect 29477 -2910 29489 -2909
rect 29247 -2943 29489 -2910
rect 29865 -2910 29877 -2909
rect 30459 -2909 30859 -2903
rect 29865 -2943 29880 -2910
rect 28720 -3040 29880 -2943
rect 14420 -3050 14560 -3040
rect 15810 -3050 15930 -3040
rect 17410 -3050 17530 -3040
rect 19010 -3050 19130 -3040
rect 20610 -3050 20730 -3040
rect 22210 -3050 22330 -3040
rect 23810 -3050 23930 -3040
rect 25410 -3050 25530 -3040
rect 27011 -3050 27130 -3040
rect 28610 -3050 29880 -3040
rect 30210 -2920 30330 -2910
rect 30459 -2920 30471 -2909
rect 30210 -3040 30220 -2920
rect 30320 -2943 30471 -2920
rect 30847 -2920 30859 -2909
rect 31077 -2909 31477 -2903
rect 31077 -2920 31089 -2909
rect 30847 -2943 31089 -2920
rect 31465 -2920 31477 -2909
rect 32059 -2909 32459 -2903
rect 31465 -2943 31480 -2920
rect 30320 -3040 31480 -2943
rect 32059 -2943 32071 -2909
rect 32447 -2920 32459 -2909
rect 32677 -2909 33077 -2903
rect 32677 -2920 32689 -2909
rect 32447 -2943 32689 -2920
rect 33065 -2920 33077 -2909
rect 33659 -2909 34059 -2903
rect 33659 -2920 33671 -2909
rect 33065 -2943 33671 -2920
rect 34047 -2920 34059 -2909
rect 34277 -2909 34677 -2903
rect 34277 -2920 34289 -2909
rect 34047 -2943 34289 -2920
rect 34665 -2920 34677 -2909
rect 35259 -2909 35659 -2903
rect 35259 -2920 35271 -2909
rect 34665 -2943 35271 -2920
rect 35647 -2920 35659 -2909
rect 35877 -2909 36277 -2903
rect 35647 -2943 35840 -2920
rect 32059 -2949 35840 -2943
rect 35877 -2943 35889 -2909
rect 36265 -2943 36277 -2909
rect 36390 -2910 36510 -2900
rect 36390 -2920 36400 -2910
rect 35877 -2949 36277 -2943
rect 32060 -2980 35840 -2949
rect 36320 -2980 36400 -2920
rect 32060 -3030 36400 -2980
rect 36500 -3030 36510 -2910
rect 32060 -3040 36510 -3030
rect 30210 -3050 30330 -3040
rect 36660 -3100 36800 -2876
rect 36859 -2909 37259 -2903
rect 36859 -2943 36871 -2909
rect 37247 -2943 37259 -2909
rect 36859 -2949 37259 -2943
rect 37300 -3100 37440 -2876
rect 37477 -2909 37877 -2903
rect 37477 -2943 37489 -2909
rect 37865 -2943 37877 -2909
rect 37477 -2949 37877 -2943
rect 37920 -3100 38060 -2876
rect 31720 -3140 38100 -3100
rect 660 -3171 38100 -3140
rect -140 -3205 -117 -3171
rect 1253 -3205 1483 -3171
rect 2853 -3205 3083 -3171
rect 4453 -3205 4683 -3171
rect 6053 -3205 6283 -3171
rect 7653 -3205 7883 -3171
rect 9253 -3205 9483 -3171
rect 10853 -3205 11083 -3171
rect 12453 -3205 12683 -3171
rect 14053 -3205 14283 -3171
rect 15653 -3205 15883 -3171
rect 17253 -3205 17483 -3171
rect 18853 -3205 19083 -3171
rect 20453 -3205 20683 -3171
rect 22053 -3205 22283 -3171
rect 23653 -3205 23883 -3171
rect 25253 -3205 25483 -3171
rect 26853 -3205 27083 -3171
rect 28453 -3205 28683 -3171
rect 30053 -3205 30283 -3171
rect 31653 -3205 31883 -3171
rect 33253 -3205 33483 -3171
rect 34853 -3205 35083 -3171
rect 36453 -3205 36683 -3171
rect 38053 -3205 38100 -3171
rect -140 -3305 480 -3205
rect -140 -3339 71 -3305
rect 447 -3339 480 -3305
rect -140 -3340 480 -3339
rect -140 -3393 0 -3340
rect 59 -3345 480 -3340
rect -140 -3405 27 -3393
rect -140 -4097 -13 -3405
rect 21 -4097 27 -3405
rect -140 -4109 27 -4097
rect -140 -4518 0 -4109
rect 440 -4157 480 -3345
rect 660 -3220 38100 -3205
rect 660 -3240 31960 -3220
rect 660 -3305 12520 -3240
rect 660 -3339 689 -3305
rect 1065 -3339 1671 -3305
rect 2047 -3339 2289 -3305
rect 2665 -3339 3271 -3305
rect 3647 -3339 3889 -3305
rect 4265 -3339 4871 -3305
rect 5247 -3339 5489 -3305
rect 5865 -3339 6471 -3305
rect 6847 -3339 7089 -3305
rect 7465 -3339 8071 -3305
rect 8447 -3339 8689 -3305
rect 9065 -3339 9671 -3305
rect 10047 -3339 10289 -3305
rect 10665 -3339 11271 -3305
rect 11647 -3339 11889 -3305
rect 12265 -3339 12520 -3305
rect 660 -3340 12520 -3339
rect 12600 -3290 13260 -3280
rect 660 -3345 1077 -3340
rect 1659 -3345 2059 -3340
rect 2277 -3345 2677 -3340
rect 3259 -3345 3659 -3340
rect 3877 -3345 4277 -3340
rect 4859 -3345 5259 -3340
rect 5477 -3345 5877 -3340
rect 6459 -3345 6859 -3340
rect 7077 -3345 7477 -3340
rect 8059 -3345 8459 -3340
rect 8677 -3345 9077 -3340
rect 9659 -3345 10059 -3340
rect 10277 -3345 10677 -3340
rect 11259 -3345 11659 -3340
rect 11877 -3345 12277 -3340
rect 59 -4163 480 -4157
rect 59 -4197 71 -4163
rect 447 -4197 480 -4163
rect 59 -4203 480 -4197
rect 440 -4445 480 -4203
rect 59 -4451 480 -4445
rect 59 -4485 71 -4451
rect 447 -4485 480 -4451
rect 59 -4491 480 -4485
rect -140 -4530 27 -4518
rect -140 -4664 -13 -4530
rect 21 -4664 27 -4530
rect -140 -4676 27 -4664
rect -140 -4680 0 -4676
rect 440 -4703 480 -4491
rect 660 -4157 710 -3345
rect 12600 -3390 12610 -3290
rect 12730 -3305 13260 -3290
rect 12730 -3339 12871 -3305
rect 13247 -3339 13260 -3305
rect 12730 -3340 13260 -3339
rect 13380 -3305 14120 -3240
rect 13380 -3339 13489 -3305
rect 13865 -3339 14120 -3305
rect 13380 -3340 14120 -3339
rect 14200 -3290 14860 -3280
rect 12730 -3390 12740 -3340
rect 12859 -3345 13259 -3340
rect 13477 -3345 13877 -3340
rect 1109 -3405 1155 -3393
rect 1109 -4097 1115 -3405
rect 1149 -4097 1155 -3405
rect 1109 -4109 1155 -4097
rect 1581 -3405 1627 -3393
rect 1581 -4097 1587 -3405
rect 1621 -4097 1627 -3405
rect 1581 -4109 1627 -4097
rect 2091 -3400 2137 -3393
rect 2199 -3400 2245 -3393
rect 2091 -3405 2245 -3400
rect 2091 -4097 2097 -3405
rect 2131 -3410 2205 -3405
rect 2131 -4097 2205 -4090
rect 2239 -4097 2245 -3405
rect 2091 -4100 2245 -4097
rect 2091 -4109 2137 -4100
rect 2199 -4109 2245 -4100
rect 2709 -3405 2755 -3393
rect 2709 -4097 2715 -3405
rect 2749 -4097 2755 -3405
rect 2709 -4109 2755 -4097
rect 3181 -3405 3227 -3393
rect 3181 -4097 3187 -3405
rect 3221 -4097 3227 -3405
rect 3181 -4109 3227 -4097
rect 3691 -3400 3737 -3393
rect 3799 -3400 3845 -3393
rect 3691 -3405 3845 -3400
rect 3691 -4097 3697 -3405
rect 3731 -3410 3805 -3405
rect 3731 -4097 3805 -4090
rect 3839 -4097 3845 -3405
rect 3691 -4100 3845 -4097
rect 3691 -4109 3737 -4100
rect 3799 -4109 3845 -4100
rect 4309 -3405 4355 -3393
rect 4309 -4097 4315 -3405
rect 4349 -4097 4355 -3405
rect 4309 -4109 4355 -4097
rect 4781 -3405 4827 -3393
rect 4781 -4097 4787 -3405
rect 4821 -4097 4827 -3405
rect 4781 -4109 4827 -4097
rect 5291 -3400 5337 -3393
rect 5399 -3400 5445 -3393
rect 5291 -3405 5445 -3400
rect 5291 -4097 5297 -3405
rect 5331 -3410 5405 -3405
rect 5331 -4097 5405 -4090
rect 5439 -4097 5445 -3405
rect 5291 -4100 5445 -4097
rect 5291 -4109 5337 -4100
rect 5399 -4109 5445 -4100
rect 5909 -3405 5955 -3393
rect 5909 -4097 5915 -3405
rect 5949 -4097 5955 -3405
rect 5909 -4109 5955 -4097
rect 6381 -3405 6427 -3393
rect 6381 -4097 6387 -3405
rect 6421 -4097 6427 -3405
rect 6381 -4109 6427 -4097
rect 6891 -3400 6937 -3393
rect 6999 -3400 7045 -3393
rect 6891 -3405 7045 -3400
rect 6891 -4097 6897 -3405
rect 6931 -3410 7005 -3405
rect 6931 -4097 7005 -4090
rect 7039 -4097 7045 -3405
rect 6891 -4100 7045 -4097
rect 6891 -4109 6937 -4100
rect 6999 -4109 7045 -4100
rect 7509 -3405 7555 -3393
rect 7509 -4097 7515 -3405
rect 7549 -4097 7555 -3405
rect 7509 -4109 7555 -4097
rect 7981 -3405 8027 -3393
rect 7981 -4097 7987 -3405
rect 8021 -4097 8027 -3405
rect 7981 -4109 8027 -4097
rect 8491 -3400 8537 -3393
rect 8599 -3400 8645 -3393
rect 8491 -3405 8645 -3400
rect 8491 -4097 8497 -3405
rect 8531 -3410 8605 -3405
rect 8531 -4097 8605 -4090
rect 8639 -4097 8645 -3405
rect 8491 -4100 8645 -4097
rect 8491 -4109 8537 -4100
rect 8599 -4109 8645 -4100
rect 9109 -3405 9155 -3393
rect 9109 -4097 9115 -3405
rect 9149 -4097 9155 -3405
rect 9109 -4109 9155 -4097
rect 9581 -3405 9627 -3393
rect 9581 -4097 9587 -3405
rect 9621 -4097 9627 -3405
rect 9581 -4109 9627 -4097
rect 10091 -3400 10137 -3393
rect 10199 -3400 10245 -3393
rect 10091 -3405 10245 -3400
rect 10091 -4097 10097 -3405
rect 10131 -3410 10205 -3405
rect 10131 -4097 10205 -4090
rect 10239 -4097 10245 -3405
rect 10091 -4100 10245 -4097
rect 10091 -4109 10137 -4100
rect 10199 -4109 10245 -4100
rect 10709 -3405 10755 -3393
rect 10709 -4097 10715 -3405
rect 10749 -4097 10755 -3405
rect 10709 -4109 10755 -4097
rect 11181 -3405 11227 -3393
rect 11181 -4097 11187 -3405
rect 11221 -4097 11227 -3405
rect 11181 -4109 11227 -4097
rect 11691 -3400 11737 -3393
rect 11799 -3400 11845 -3393
rect 11691 -3405 11845 -3400
rect 11691 -4097 11697 -3405
rect 11731 -3410 11805 -3405
rect 11731 -4097 11805 -4090
rect 11839 -4097 11845 -3405
rect 11691 -4100 11845 -4097
rect 11691 -4109 11737 -4100
rect 11799 -4109 11845 -4100
rect 12309 -3405 12355 -3393
rect 12600 -3400 12740 -3390
rect 12309 -4097 12315 -3405
rect 12349 -4097 12355 -3405
rect 12309 -4109 12355 -4097
rect 12781 -3405 12827 -3393
rect 12781 -4097 12787 -3405
rect 12821 -4097 12827 -3405
rect 12781 -4109 12827 -4097
rect 13291 -3400 13337 -3393
rect 13399 -3400 13445 -3393
rect 13291 -3405 13445 -3400
rect 13291 -4097 13297 -3405
rect 13331 -3410 13405 -3405
rect 13331 -4097 13405 -4090
rect 13439 -4097 13445 -3405
rect 13291 -4100 13445 -4097
rect 13291 -4109 13337 -4100
rect 13399 -4109 13445 -4100
rect 13909 -3405 13955 -3393
rect 13909 -4097 13915 -3405
rect 13949 -4097 13955 -3405
rect 14200 -3410 14210 -3290
rect 14330 -3305 14860 -3290
rect 14330 -3339 14471 -3305
rect 14847 -3339 14860 -3305
rect 14330 -3340 14860 -3339
rect 14980 -3305 31960 -3240
rect 32060 -3280 36270 -3270
rect 32060 -3299 33400 -3280
rect 14980 -3339 15089 -3305
rect 15465 -3339 16071 -3305
rect 16447 -3339 16689 -3305
rect 17065 -3339 17671 -3305
rect 18047 -3339 18289 -3305
rect 18665 -3339 19271 -3305
rect 19647 -3339 19889 -3305
rect 20265 -3339 20871 -3305
rect 21247 -3339 21489 -3305
rect 21865 -3339 22471 -3305
rect 22847 -3339 23089 -3305
rect 23465 -3339 24071 -3305
rect 24447 -3339 24689 -3305
rect 25065 -3339 25671 -3305
rect 26047 -3339 26289 -3305
rect 26665 -3339 27271 -3305
rect 27647 -3339 27889 -3305
rect 28265 -3339 28871 -3305
rect 29247 -3339 29489 -3305
rect 29865 -3339 30471 -3305
rect 30847 -3339 31089 -3305
rect 31465 -3339 31960 -3305
rect 14980 -3340 31960 -3339
rect 32059 -3305 33400 -3299
rect 32059 -3339 32071 -3305
rect 32447 -3339 32689 -3305
rect 33065 -3339 33400 -3305
rect 32059 -3340 33400 -3339
rect 14330 -3410 14340 -3340
rect 14459 -3345 14859 -3340
rect 15077 -3345 15477 -3340
rect 16059 -3345 16459 -3340
rect 16677 -3345 17077 -3340
rect 17659 -3345 18059 -3340
rect 18277 -3345 18677 -3340
rect 19259 -3345 19659 -3340
rect 19877 -3345 20277 -3340
rect 20859 -3345 21259 -3340
rect 21477 -3345 21877 -3340
rect 22459 -3345 22859 -3340
rect 23077 -3345 23477 -3340
rect 24059 -3345 24459 -3340
rect 24677 -3345 25077 -3340
rect 25659 -3345 26059 -3340
rect 26277 -3345 26677 -3340
rect 27259 -3345 27659 -3340
rect 27877 -3345 28277 -3340
rect 28859 -3345 29259 -3340
rect 29477 -3345 29877 -3340
rect 30459 -3345 30859 -3340
rect 31077 -3345 31477 -3340
rect 32059 -3345 32459 -3340
rect 32677 -3345 33077 -3340
rect 14200 -3420 14340 -3410
rect 14381 -3405 14427 -3393
rect 13909 -4109 13955 -4097
rect 14381 -4097 14387 -3405
rect 14421 -4097 14427 -3405
rect 14381 -4109 14427 -4097
rect 14891 -3400 14937 -3393
rect 14999 -3400 15045 -3393
rect 14891 -3405 15045 -3400
rect 14891 -4097 14897 -3405
rect 14931 -3410 15005 -3405
rect 14931 -4097 15005 -4090
rect 15039 -4097 15045 -3405
rect 14891 -4100 15045 -4097
rect 14891 -4109 14937 -4100
rect 14999 -4109 15045 -4100
rect 15509 -3405 15555 -3393
rect 15509 -4097 15515 -3405
rect 15549 -4097 15555 -3405
rect 15509 -4109 15555 -4097
rect 15981 -3405 16027 -3393
rect 15981 -4097 15987 -3405
rect 16021 -4097 16027 -3405
rect 15981 -4109 16027 -4097
rect 16491 -3400 16537 -3393
rect 16599 -3400 16645 -3393
rect 16491 -3405 16645 -3400
rect 16491 -4097 16497 -3405
rect 16531 -3410 16605 -3405
rect 16531 -4097 16605 -4090
rect 16639 -4097 16645 -3405
rect 16491 -4100 16645 -4097
rect 16491 -4109 16537 -4100
rect 16599 -4109 16645 -4100
rect 17109 -3405 17155 -3393
rect 17109 -4097 17115 -3405
rect 17149 -4097 17155 -3405
rect 17109 -4109 17155 -4097
rect 17581 -3405 17627 -3393
rect 17581 -4097 17587 -3405
rect 17621 -4097 17627 -3405
rect 17581 -4109 17627 -4097
rect 18091 -3400 18137 -3393
rect 18199 -3400 18245 -3393
rect 18091 -3405 18245 -3400
rect 18091 -4097 18097 -3405
rect 18131 -3410 18205 -3405
rect 18131 -4097 18205 -4090
rect 18239 -4097 18245 -3405
rect 18091 -4100 18245 -4097
rect 18091 -4109 18137 -4100
rect 18199 -4109 18245 -4100
rect 18709 -3405 18755 -3393
rect 18709 -4097 18715 -3405
rect 18749 -4097 18755 -3405
rect 18709 -4109 18755 -4097
rect 19181 -3405 19227 -3393
rect 19181 -4097 19187 -3405
rect 19221 -4097 19227 -3405
rect 19181 -4109 19227 -4097
rect 19691 -3400 19737 -3393
rect 19799 -3400 19845 -3393
rect 19691 -3405 19845 -3400
rect 19691 -4097 19697 -3405
rect 19731 -3410 19805 -3405
rect 19731 -4097 19805 -4090
rect 19839 -4097 19845 -3405
rect 19691 -4100 19845 -4097
rect 19691 -4109 19737 -4100
rect 19799 -4109 19845 -4100
rect 20309 -3405 20355 -3393
rect 20309 -4097 20315 -3405
rect 20349 -4097 20355 -3405
rect 20309 -4109 20355 -4097
rect 20781 -3405 20827 -3393
rect 20781 -4097 20787 -3405
rect 20821 -4097 20827 -3405
rect 20781 -4109 20827 -4097
rect 21291 -3400 21337 -3393
rect 21399 -3400 21445 -3393
rect 21291 -3405 21445 -3400
rect 21291 -4097 21297 -3405
rect 21331 -3410 21405 -3405
rect 21331 -4097 21405 -4090
rect 21439 -4097 21445 -3405
rect 21291 -4100 21445 -4097
rect 21291 -4109 21337 -4100
rect 21399 -4109 21445 -4100
rect 21909 -3405 21955 -3393
rect 21909 -4097 21915 -3405
rect 21949 -4097 21955 -3405
rect 21909 -4109 21955 -4097
rect 22381 -3405 22427 -3393
rect 22381 -4097 22387 -3405
rect 22421 -4097 22427 -3405
rect 22381 -4109 22427 -4097
rect 22891 -3400 22937 -3393
rect 22999 -3400 23045 -3393
rect 22891 -3405 23045 -3400
rect 22891 -4097 22897 -3405
rect 22931 -3410 23005 -3405
rect 22931 -4097 23005 -4090
rect 23039 -4097 23045 -3405
rect 22891 -4100 23045 -4097
rect 22891 -4109 22937 -4100
rect 22999 -4109 23045 -4100
rect 23509 -3405 23555 -3393
rect 23509 -4097 23515 -3405
rect 23549 -4097 23555 -3405
rect 23509 -4109 23555 -4097
rect 23981 -3405 24027 -3393
rect 23981 -4097 23987 -3405
rect 24021 -4097 24027 -3405
rect 23981 -4109 24027 -4097
rect 24491 -3400 24537 -3393
rect 24599 -3400 24645 -3393
rect 24491 -3405 24645 -3400
rect 24491 -4097 24497 -3405
rect 24531 -3410 24605 -3405
rect 24531 -4097 24605 -4090
rect 24639 -4097 24645 -3405
rect 24491 -4100 24645 -4097
rect 24491 -4109 24537 -4100
rect 24599 -4109 24645 -4100
rect 25109 -3405 25155 -3393
rect 25109 -4097 25115 -3405
rect 25149 -4097 25155 -3405
rect 25109 -4109 25155 -4097
rect 25581 -3405 25627 -3393
rect 25581 -4097 25587 -3405
rect 25621 -4097 25627 -3405
rect 25581 -4109 25627 -4097
rect 26091 -3400 26137 -3393
rect 26199 -3400 26245 -3393
rect 26091 -3405 26245 -3400
rect 26091 -4097 26097 -3405
rect 26131 -3410 26205 -3405
rect 26131 -4097 26205 -4090
rect 26239 -4097 26245 -3405
rect 26091 -4100 26245 -4097
rect 26091 -4109 26137 -4100
rect 26199 -4109 26245 -4100
rect 26709 -3405 26755 -3393
rect 26709 -4097 26715 -3405
rect 26749 -4097 26755 -3405
rect 26709 -4109 26755 -4097
rect 27181 -3405 27227 -3393
rect 27181 -4097 27187 -3405
rect 27221 -4097 27227 -3405
rect 27181 -4109 27227 -4097
rect 27691 -3400 27737 -3393
rect 27799 -3400 27845 -3393
rect 27691 -3405 27845 -3400
rect 27691 -4097 27697 -3405
rect 27731 -3410 27805 -3405
rect 27731 -4097 27805 -4090
rect 27839 -4097 27845 -3405
rect 27691 -4100 27845 -4097
rect 27691 -4109 27737 -4100
rect 27799 -4109 27845 -4100
rect 28309 -3405 28355 -3393
rect 28309 -4097 28315 -3405
rect 28349 -4097 28355 -3405
rect 28309 -4109 28355 -4097
rect 28781 -3405 28827 -3393
rect 28781 -4097 28787 -3405
rect 28821 -4097 28827 -3405
rect 28781 -4109 28827 -4097
rect 29291 -3400 29337 -3393
rect 29399 -3400 29445 -3393
rect 29291 -3405 29445 -3400
rect 29291 -4097 29297 -3405
rect 29331 -3410 29405 -3405
rect 29331 -4097 29405 -4090
rect 29439 -4097 29445 -3405
rect 29291 -4100 29445 -4097
rect 29291 -4109 29337 -4100
rect 29399 -4109 29445 -4100
rect 29909 -3405 29955 -3393
rect 29909 -4097 29915 -3405
rect 29949 -4097 29955 -3405
rect 29909 -4109 29955 -4097
rect 30381 -3405 30427 -3393
rect 30381 -4097 30387 -3405
rect 30421 -4097 30427 -3405
rect 30381 -4109 30427 -4097
rect 30891 -3400 30937 -3393
rect 30999 -3400 31045 -3393
rect 30891 -3405 31045 -3400
rect 30891 -4097 30897 -3405
rect 30931 -3410 31005 -3405
rect 30931 -4097 31005 -4090
rect 31039 -4097 31045 -3405
rect 30891 -4100 31045 -4097
rect 30891 -4109 30937 -4100
rect 30999 -4109 31045 -4100
rect 31509 -3405 31555 -3393
rect 31509 -4097 31515 -3405
rect 31549 -4097 31555 -3405
rect 31509 -4109 31555 -4097
rect 31981 -3405 32027 -3393
rect 31981 -4097 31987 -3405
rect 32021 -4097 32027 -3405
rect 31981 -4109 32027 -4097
rect 32491 -3400 32537 -3393
rect 32599 -3400 32645 -3393
rect 32491 -3405 32645 -3400
rect 32491 -4097 32497 -3405
rect 32531 -3410 32605 -3405
rect 32531 -4097 32605 -4090
rect 32639 -4097 32645 -3405
rect 32491 -4100 32645 -4097
rect 32491 -4109 32537 -4100
rect 32599 -4109 32645 -4100
rect 33109 -3405 33155 -3393
rect 33109 -4097 33115 -3405
rect 33149 -4097 33155 -3405
rect 33390 -3400 33400 -3340
rect 33530 -3299 36270 -3280
rect 33530 -3305 36277 -3299
rect 33530 -3339 33671 -3305
rect 34047 -3339 34289 -3305
rect 34665 -3339 35271 -3305
rect 35647 -3339 35889 -3305
rect 36265 -3339 36277 -3305
rect 33530 -3340 36277 -3339
rect 36530 -3305 38100 -3220
rect 36530 -3339 36871 -3305
rect 37247 -3339 37489 -3305
rect 37865 -3339 38100 -3305
rect 36530 -3340 38100 -3339
rect 33659 -3345 34059 -3340
rect 34277 -3345 34677 -3340
rect 35259 -3345 35659 -3340
rect 35877 -3345 36277 -3340
rect 36660 -3393 36800 -3340
rect 36859 -3345 37259 -3340
rect 37300 -3393 37440 -3340
rect 37477 -3345 37877 -3340
rect 37920 -3393 38060 -3340
rect 33390 -3410 33530 -3400
rect 33581 -3405 33627 -3393
rect 33109 -4109 33155 -4097
rect 33581 -4097 33587 -3405
rect 33621 -4097 33627 -3405
rect 33581 -4109 33627 -4097
rect 34091 -3400 34137 -3393
rect 34199 -3400 34245 -3393
rect 34091 -3405 34245 -3400
rect 34091 -4097 34097 -3405
rect 34131 -3410 34205 -3405
rect 34131 -4097 34205 -4090
rect 34239 -4097 34245 -3405
rect 34091 -4100 34245 -4097
rect 34091 -4109 34137 -4100
rect 34199 -4109 34245 -4100
rect 34709 -3405 34755 -3393
rect 34709 -4097 34715 -3405
rect 34749 -4097 34755 -3405
rect 34709 -4109 34755 -4097
rect 35181 -3405 35227 -3393
rect 35181 -4097 35187 -3405
rect 35221 -4097 35227 -3405
rect 35181 -4109 35227 -4097
rect 35691 -3400 35737 -3393
rect 35799 -3400 35845 -3393
rect 35691 -3405 35845 -3400
rect 35691 -4097 35697 -3405
rect 35731 -3410 35805 -3405
rect 35731 -4097 35805 -4090
rect 35839 -4097 35845 -3405
rect 35691 -4100 35845 -4097
rect 35691 -4109 35737 -4100
rect 35799 -4109 35845 -4100
rect 36309 -3405 36355 -3393
rect 36309 -4097 36315 -3405
rect 36349 -4097 36355 -3405
rect 36309 -4109 36355 -4097
rect 36660 -3405 36827 -3393
rect 36660 -4097 36787 -3405
rect 36821 -4097 36827 -3405
rect 36660 -4109 36827 -4097
rect 37291 -3405 37445 -3393
rect 37291 -4097 37297 -3405
rect 37331 -4097 37405 -3405
rect 37439 -4097 37445 -3405
rect 37291 -4109 37445 -4097
rect 37909 -3405 38060 -3393
rect 37909 -4097 37915 -3405
rect 37949 -4097 38060 -3405
rect 37909 -4109 38060 -4097
rect 660 -4163 1077 -4157
rect 660 -4197 689 -4163
rect 1065 -4197 1077 -4163
rect 660 -4203 1077 -4197
rect 1659 -4163 2059 -4157
rect 1659 -4197 1671 -4163
rect 2047 -4197 2059 -4163
rect 1659 -4203 2059 -4197
rect 2277 -4163 2677 -4157
rect 2277 -4197 2289 -4163
rect 2665 -4197 2677 -4163
rect 2277 -4203 2677 -4197
rect 3259 -4163 3659 -4157
rect 3259 -4197 3271 -4163
rect 3647 -4197 3659 -4163
rect 3259 -4203 3659 -4197
rect 3877 -4163 4277 -4157
rect 3877 -4197 3889 -4163
rect 4265 -4197 4277 -4163
rect 3877 -4203 4277 -4197
rect 4859 -4163 5259 -4157
rect 4859 -4197 4871 -4163
rect 5247 -4197 5259 -4163
rect 4859 -4203 5259 -4197
rect 5477 -4163 5877 -4157
rect 5477 -4197 5489 -4163
rect 5865 -4197 5877 -4163
rect 5477 -4203 5877 -4197
rect 6459 -4163 6859 -4157
rect 6459 -4197 6471 -4163
rect 6847 -4197 6859 -4163
rect 6459 -4203 6859 -4197
rect 7077 -4163 7477 -4157
rect 7077 -4197 7089 -4163
rect 7465 -4197 7477 -4163
rect 7077 -4203 7477 -4197
rect 8059 -4163 8459 -4157
rect 8059 -4197 8071 -4163
rect 8447 -4197 8459 -4163
rect 8059 -4203 8459 -4197
rect 8677 -4163 9077 -4157
rect 8677 -4197 8689 -4163
rect 9065 -4197 9077 -4163
rect 8677 -4203 9077 -4197
rect 9659 -4163 10059 -4157
rect 9659 -4197 9671 -4163
rect 10047 -4197 10059 -4163
rect 9659 -4203 10059 -4197
rect 10277 -4163 10677 -4157
rect 10277 -4197 10289 -4163
rect 10665 -4197 10677 -4163
rect 10277 -4203 10677 -4197
rect 11259 -4163 11659 -4157
rect 11259 -4197 11271 -4163
rect 11647 -4197 11659 -4163
rect 11259 -4203 11659 -4197
rect 11877 -4163 12277 -4157
rect 11877 -4197 11889 -4163
rect 12265 -4197 12277 -4163
rect 12859 -4163 13259 -4157
rect 12859 -4180 12871 -4163
rect 11877 -4203 12277 -4197
rect 12840 -4197 12871 -4180
rect 13247 -4180 13259 -4163
rect 13477 -4163 13877 -4157
rect 13477 -4180 13489 -4163
rect 13247 -4197 13489 -4180
rect 13865 -4180 13877 -4163
rect 14459 -4163 14859 -4157
rect 14459 -4180 14471 -4163
rect 13865 -4197 13880 -4180
rect 660 -4445 710 -4203
rect 1680 -4240 2040 -4203
rect 2300 -4240 2660 -4203
rect 3280 -4240 3640 -4203
rect 3900 -4240 4260 -4203
rect 4880 -4240 5240 -4203
rect 5500 -4240 5860 -4203
rect 6480 -4240 6840 -4203
rect 7100 -4240 7460 -4203
rect 8080 -4240 8440 -4203
rect 8700 -4240 9060 -4203
rect 9680 -4240 10040 -4203
rect 10300 -4240 10660 -4203
rect 11280 -4240 11640 -4203
rect 11900 -4240 12260 -4203
rect 1400 -4250 10660 -4240
rect 1400 -4370 1410 -4250
rect 1530 -4370 3010 -4250
rect 3130 -4370 4610 -4250
rect 4730 -4370 6210 -4250
rect 6330 -4370 7810 -4250
rect 7930 -4370 9410 -4250
rect 9530 -4370 10660 -4250
rect 1400 -4380 10660 -4370
rect 11260 -4380 12260 -4240
rect 12840 -4260 13880 -4197
rect 14440 -4197 14471 -4180
rect 14847 -4180 14859 -4163
rect 15077 -4163 15477 -4157
rect 15077 -4180 15089 -4163
rect 14847 -4197 15089 -4180
rect 15465 -4180 15477 -4163
rect 16059 -4163 16459 -4157
rect 15465 -4197 15480 -4180
rect 14440 -4260 15480 -4197
rect 16059 -4197 16071 -4163
rect 16447 -4197 16459 -4163
rect 16059 -4203 16459 -4197
rect 16677 -4163 17077 -4157
rect 16677 -4197 16689 -4163
rect 17065 -4197 17077 -4163
rect 16677 -4203 17077 -4197
rect 17659 -4163 18059 -4157
rect 17659 -4197 17671 -4163
rect 18047 -4197 18059 -4163
rect 17659 -4203 18059 -4197
rect 18277 -4163 18677 -4157
rect 18277 -4197 18289 -4163
rect 18665 -4197 18677 -4163
rect 18277 -4203 18677 -4197
rect 19259 -4163 19659 -4157
rect 19259 -4197 19271 -4163
rect 19647 -4197 19659 -4163
rect 19259 -4203 19659 -4197
rect 19877 -4163 20277 -4157
rect 19877 -4197 19889 -4163
rect 20265 -4197 20277 -4163
rect 19877 -4203 20277 -4197
rect 20859 -4163 21259 -4157
rect 20859 -4197 20871 -4163
rect 21247 -4197 21259 -4163
rect 20859 -4203 21259 -4197
rect 21477 -4163 21877 -4157
rect 21477 -4197 21489 -4163
rect 21865 -4197 21877 -4163
rect 21477 -4203 21877 -4197
rect 22459 -4163 22859 -4157
rect 22459 -4197 22471 -4163
rect 22847 -4197 22859 -4163
rect 22459 -4203 22859 -4197
rect 23077 -4163 23477 -4157
rect 23077 -4197 23089 -4163
rect 23465 -4197 23477 -4163
rect 23077 -4203 23477 -4197
rect 24059 -4163 24459 -4157
rect 24059 -4197 24071 -4163
rect 24447 -4197 24459 -4163
rect 24059 -4203 24459 -4197
rect 24677 -4163 25077 -4157
rect 24677 -4197 24689 -4163
rect 25065 -4197 25077 -4163
rect 24677 -4203 25077 -4197
rect 25659 -4163 26059 -4157
rect 25659 -4197 25671 -4163
rect 26047 -4197 26059 -4163
rect 25659 -4203 26059 -4197
rect 26277 -4163 26677 -4157
rect 26277 -4197 26289 -4163
rect 26665 -4197 26677 -4163
rect 26277 -4203 26677 -4197
rect 27259 -4163 27659 -4157
rect 27259 -4197 27271 -4163
rect 27647 -4197 27659 -4163
rect 27259 -4203 27659 -4197
rect 27877 -4163 28277 -4157
rect 27877 -4197 27889 -4163
rect 28265 -4197 28277 -4163
rect 27877 -4203 28277 -4197
rect 28859 -4163 29259 -4157
rect 28859 -4197 28871 -4163
rect 29247 -4197 29259 -4163
rect 28859 -4203 29259 -4197
rect 29477 -4163 29877 -4157
rect 29477 -4197 29489 -4163
rect 29865 -4197 29877 -4163
rect 29477 -4203 29877 -4197
rect 30459 -4163 30859 -4157
rect 30459 -4197 30471 -4163
rect 30847 -4197 30859 -4163
rect 30459 -4203 30859 -4197
rect 31077 -4163 31477 -4157
rect 31077 -4197 31089 -4163
rect 31465 -4197 31477 -4163
rect 31077 -4203 31477 -4197
rect 32059 -4163 32459 -4157
rect 32059 -4197 32071 -4163
rect 32447 -4197 32459 -4163
rect 32059 -4203 32459 -4197
rect 32677 -4163 33077 -4157
rect 32677 -4197 32689 -4163
rect 33065 -4197 33077 -4163
rect 32677 -4203 33077 -4197
rect 33659 -4163 34059 -4157
rect 33659 -4197 33671 -4163
rect 34047 -4197 34059 -4163
rect 33659 -4203 34059 -4197
rect 34277 -4163 34677 -4157
rect 34277 -4197 34289 -4163
rect 34665 -4197 34677 -4163
rect 34277 -4203 34677 -4197
rect 35259 -4163 35659 -4157
rect 35259 -4197 35271 -4163
rect 35647 -4197 35659 -4163
rect 35259 -4203 35659 -4197
rect 35877 -4163 36277 -4157
rect 35877 -4197 35889 -4163
rect 36265 -4197 36277 -4163
rect 35877 -4203 36277 -4197
rect 16080 -4240 16440 -4203
rect 16700 -4240 17060 -4203
rect 17680 -4240 18040 -4203
rect 18300 -4240 18660 -4203
rect 19280 -4240 19640 -4203
rect 19900 -4240 20260 -4203
rect 20880 -4240 21240 -4203
rect 21500 -4240 21860 -4203
rect 22480 -4240 22840 -4203
rect 23100 -4240 23460 -4203
rect 24080 -4240 24440 -4203
rect 24700 -4240 25060 -4203
rect 25680 -4240 26040 -4203
rect 26300 -4240 26660 -4203
rect 27280 -4240 27640 -4203
rect 27900 -4240 28260 -4203
rect 28880 -4240 29240 -4203
rect 29500 -4240 29860 -4203
rect 30480 -4240 30840 -4203
rect 31100 -4240 31460 -4203
rect 32080 -4240 32440 -4203
rect 32700 -4240 33060 -4203
rect 33680 -4240 34040 -4203
rect 34300 -4240 34660 -4203
rect 35280 -4240 35640 -4203
rect 35900 -4240 36260 -4203
rect 15590 -4250 17060 -4240
rect 15590 -4370 15600 -4250
rect 15700 -4370 17060 -4250
rect 1680 -4445 2040 -4380
rect 2300 -4445 2660 -4380
rect 3280 -4445 3640 -4380
rect 3900 -4445 4260 -4380
rect 4880 -4445 5240 -4380
rect 5500 -4445 5860 -4380
rect 6480 -4445 6840 -4380
rect 7100 -4445 7460 -4380
rect 8080 -4445 8440 -4380
rect 8700 -4445 9060 -4380
rect 9680 -4445 10040 -4380
rect 10300 -4445 10660 -4380
rect 11280 -4425 11640 -4380
rect 11900 -4425 12260 -4380
rect 11260 -4430 11659 -4425
rect 11260 -4445 11660 -4430
rect 660 -4451 1077 -4445
rect 660 -4485 689 -4451
rect 1065 -4485 1077 -4451
rect 660 -4491 1077 -4485
rect 1659 -4451 2059 -4445
rect 1659 -4485 1671 -4451
rect 2047 -4485 2059 -4451
rect 1659 -4491 2059 -4485
rect 2277 -4451 2677 -4445
rect 2277 -4485 2289 -4451
rect 2665 -4485 2677 -4451
rect 2277 -4491 2677 -4485
rect 3259 -4451 3659 -4445
rect 3259 -4485 3271 -4451
rect 3647 -4485 3659 -4451
rect 3259 -4491 3659 -4485
rect 3877 -4451 4277 -4445
rect 3877 -4485 3889 -4451
rect 4265 -4485 4277 -4451
rect 3877 -4491 4277 -4485
rect 4859 -4451 5259 -4445
rect 4859 -4485 4871 -4451
rect 5247 -4485 5259 -4451
rect 4859 -4491 5259 -4485
rect 5477 -4451 5877 -4445
rect 5477 -4485 5489 -4451
rect 5865 -4485 5877 -4451
rect 5477 -4491 5877 -4485
rect 6459 -4451 6859 -4445
rect 6459 -4485 6471 -4451
rect 6847 -4485 6859 -4451
rect 6459 -4491 6859 -4485
rect 7077 -4451 7477 -4445
rect 7077 -4485 7089 -4451
rect 7465 -4485 7477 -4451
rect 7077 -4491 7477 -4485
rect 8059 -4451 8459 -4445
rect 8059 -4485 8071 -4451
rect 8447 -4485 8459 -4451
rect 8059 -4491 8459 -4485
rect 8677 -4451 9077 -4445
rect 8677 -4485 8689 -4451
rect 9065 -4485 9077 -4451
rect 8677 -4491 9077 -4485
rect 9659 -4451 10059 -4445
rect 9659 -4485 9671 -4451
rect 10047 -4485 10059 -4451
rect 9659 -4491 10059 -4485
rect 10277 -4451 10677 -4445
rect 10277 -4485 10289 -4451
rect 10665 -4485 10677 -4451
rect 10277 -4491 10677 -4485
rect 11259 -4451 11660 -4445
rect 11259 -4485 11271 -4451
rect 11647 -4485 11660 -4451
rect 11259 -4490 11660 -4485
rect 11877 -4451 12277 -4425
rect 11877 -4485 11889 -4451
rect 12265 -4485 12277 -4451
rect 12850 -4451 13880 -4370
rect 12850 -4460 12871 -4451
rect 11259 -4491 11659 -4490
rect 11877 -4491 12277 -4485
rect 12859 -4485 12871 -4460
rect 13247 -4460 13489 -4451
rect 13247 -4485 13259 -4460
rect 12859 -4491 13259 -4485
rect 13477 -4485 13489 -4460
rect 13865 -4460 13880 -4451
rect 14450 -4451 15480 -4370
rect 15590 -4380 17060 -4370
rect 17190 -4250 18660 -4240
rect 17190 -4370 17200 -4250
rect 17300 -4370 18660 -4250
rect 17190 -4380 18660 -4370
rect 18790 -4250 20260 -4240
rect 18790 -4370 18800 -4250
rect 18900 -4370 20260 -4250
rect 18790 -4380 20260 -4370
rect 20390 -4250 21860 -4240
rect 20390 -4370 20400 -4250
rect 20500 -4370 21860 -4250
rect 20390 -4380 21860 -4370
rect 21990 -4250 23460 -4240
rect 21990 -4370 22000 -4250
rect 22100 -4370 23460 -4250
rect 21990 -4380 23460 -4370
rect 23590 -4250 25060 -4240
rect 23590 -4370 23600 -4250
rect 23700 -4370 25060 -4250
rect 23590 -4380 25060 -4370
rect 25190 -4250 26660 -4240
rect 25190 -4370 25200 -4250
rect 25300 -4370 26660 -4250
rect 25190 -4380 26660 -4370
rect 26791 -4250 28260 -4240
rect 26791 -4370 26800 -4250
rect 26900 -4370 28260 -4250
rect 26791 -4380 28260 -4370
rect 28391 -4250 29860 -4240
rect 28391 -4370 28400 -4250
rect 28500 -4370 29860 -4250
rect 28391 -4380 29860 -4370
rect 29990 -4250 31460 -4240
rect 29990 -4370 30000 -4250
rect 30100 -4370 31460 -4250
rect 29990 -4380 31460 -4370
rect 32060 -4250 36260 -4240
rect 32060 -4370 33180 -4250
rect 33300 -4370 36260 -4250
rect 36660 -4320 36800 -4109
rect 36859 -4163 37259 -4157
rect 36859 -4197 36871 -4163
rect 37247 -4197 37259 -4163
rect 36859 -4203 37259 -4197
rect 37300 -4320 37440 -4109
rect 37477 -4163 37877 -4157
rect 37477 -4197 37489 -4163
rect 37865 -4197 37877 -4163
rect 37477 -4203 37877 -4197
rect 37920 -4320 38060 -4109
rect 32060 -4380 36260 -4370
rect 16080 -4425 16440 -4380
rect 16700 -4425 17060 -4380
rect 17680 -4425 18040 -4380
rect 18300 -4425 18660 -4380
rect 19280 -4425 19640 -4380
rect 19900 -4425 20260 -4380
rect 20880 -4425 21240 -4380
rect 21500 -4425 21860 -4380
rect 22480 -4425 22840 -4380
rect 23100 -4425 23460 -4380
rect 24080 -4425 24440 -4380
rect 24700 -4425 25060 -4380
rect 25680 -4425 26040 -4380
rect 26300 -4425 26660 -4380
rect 27280 -4425 27640 -4380
rect 27900 -4425 28260 -4380
rect 28880 -4425 29240 -4380
rect 29500 -4425 29860 -4380
rect 30480 -4425 30840 -4380
rect 31100 -4425 31460 -4380
rect 32080 -4425 32440 -4380
rect 32700 -4425 33060 -4380
rect 33680 -4425 34040 -4380
rect 34300 -4425 34660 -4380
rect 35280 -4425 35640 -4380
rect 35900 -4425 36260 -4380
rect 14450 -4460 14471 -4451
rect 13865 -4485 13877 -4460
rect 13477 -4491 13877 -4485
rect 14459 -4485 14471 -4460
rect 14847 -4460 15089 -4451
rect 14847 -4485 14859 -4460
rect 14459 -4491 14859 -4485
rect 15077 -4485 15089 -4460
rect 15465 -4460 15480 -4451
rect 16059 -4430 16459 -4425
rect 16059 -4451 16460 -4430
rect 15465 -4485 15477 -4460
rect 15077 -4491 15477 -4485
rect 16059 -4485 16071 -4451
rect 16447 -4485 16460 -4451
rect 16059 -4490 16460 -4485
rect 16677 -4451 17077 -4425
rect 16677 -4485 16689 -4451
rect 17065 -4485 17077 -4451
rect 16059 -4491 16459 -4490
rect 16677 -4491 17077 -4485
rect 17659 -4430 18059 -4425
rect 17659 -4451 18060 -4430
rect 17659 -4485 17671 -4451
rect 18047 -4485 18060 -4451
rect 17659 -4490 18060 -4485
rect 18277 -4451 18677 -4425
rect 18277 -4485 18289 -4451
rect 18665 -4485 18677 -4451
rect 17659 -4491 18059 -4490
rect 18277 -4491 18677 -4485
rect 19259 -4430 19659 -4425
rect 19259 -4451 19660 -4430
rect 19259 -4485 19271 -4451
rect 19647 -4485 19660 -4451
rect 19259 -4490 19660 -4485
rect 19877 -4451 20277 -4425
rect 19877 -4485 19889 -4451
rect 20265 -4485 20277 -4451
rect 19259 -4491 19659 -4490
rect 19877 -4491 20277 -4485
rect 20859 -4430 21259 -4425
rect 20859 -4451 21260 -4430
rect 20859 -4485 20871 -4451
rect 21247 -4485 21260 -4451
rect 20859 -4490 21260 -4485
rect 21477 -4451 21877 -4425
rect 21477 -4485 21489 -4451
rect 21865 -4485 21877 -4451
rect 20859 -4491 21259 -4490
rect 21477 -4491 21877 -4485
rect 22459 -4430 22859 -4425
rect 22459 -4451 22860 -4430
rect 22459 -4485 22471 -4451
rect 22847 -4485 22860 -4451
rect 22459 -4490 22860 -4485
rect 23077 -4451 23477 -4425
rect 23077 -4485 23089 -4451
rect 23465 -4485 23477 -4451
rect 22459 -4491 22859 -4490
rect 23077 -4491 23477 -4485
rect 24059 -4430 24459 -4425
rect 24059 -4451 24460 -4430
rect 24059 -4485 24071 -4451
rect 24447 -4485 24460 -4451
rect 24059 -4490 24460 -4485
rect 24677 -4451 25077 -4425
rect 24677 -4485 24689 -4451
rect 25065 -4485 25077 -4451
rect 24059 -4491 24459 -4490
rect 24677 -4491 25077 -4485
rect 25659 -4430 26059 -4425
rect 25659 -4451 26060 -4430
rect 25659 -4485 25671 -4451
rect 26047 -4485 26060 -4451
rect 25659 -4490 26060 -4485
rect 26277 -4451 26677 -4425
rect 26277 -4485 26289 -4451
rect 26665 -4485 26677 -4451
rect 25659 -4491 26059 -4490
rect 26277 -4491 26677 -4485
rect 27259 -4430 27659 -4425
rect 27259 -4451 27660 -4430
rect 27259 -4485 27271 -4451
rect 27647 -4485 27660 -4451
rect 27259 -4490 27660 -4485
rect 27877 -4451 28277 -4425
rect 27877 -4485 27889 -4451
rect 28265 -4485 28277 -4451
rect 27259 -4491 27659 -4490
rect 27877 -4491 28277 -4485
rect 28859 -4430 29259 -4425
rect 28859 -4451 29260 -4430
rect 28859 -4485 28871 -4451
rect 29247 -4485 29260 -4451
rect 28859 -4490 29260 -4485
rect 29477 -4451 29877 -4425
rect 29477 -4485 29489 -4451
rect 29865 -4485 29877 -4451
rect 28859 -4491 29259 -4490
rect 29477 -4491 29877 -4485
rect 30459 -4430 30859 -4425
rect 30459 -4451 30860 -4430
rect 30459 -4485 30471 -4451
rect 30847 -4485 30860 -4451
rect 30459 -4490 30860 -4485
rect 31077 -4451 31477 -4425
rect 32060 -4430 32459 -4425
rect 32060 -4445 32460 -4430
rect 31077 -4485 31089 -4451
rect 31465 -4485 31477 -4451
rect 30459 -4491 30859 -4490
rect 31077 -4491 31477 -4485
rect 32059 -4451 32460 -4445
rect 32059 -4485 32071 -4451
rect 32447 -4485 32460 -4451
rect 32059 -4490 32460 -4485
rect 32677 -4451 33077 -4425
rect 32677 -4485 32689 -4451
rect 33065 -4485 33077 -4451
rect 32059 -4491 32459 -4490
rect 32677 -4491 33077 -4485
rect 33659 -4430 34059 -4425
rect 33659 -4451 34060 -4430
rect 33659 -4485 33671 -4451
rect 34047 -4485 34060 -4451
rect 33659 -4490 34060 -4485
rect 34277 -4451 34677 -4425
rect 34277 -4485 34289 -4451
rect 34665 -4485 34677 -4451
rect 33659 -4491 34059 -4490
rect 34277 -4491 34677 -4485
rect 35259 -4430 35659 -4425
rect 35259 -4451 35660 -4430
rect 35259 -4485 35271 -4451
rect 35647 -4485 35660 -4451
rect 35259 -4490 35660 -4485
rect 35877 -4451 36277 -4425
rect 35877 -4485 35889 -4451
rect 36265 -4485 36277 -4451
rect 35259 -4491 35659 -4490
rect 35877 -4491 36277 -4485
rect 36859 -4451 37259 -4445
rect 36859 -4485 36871 -4451
rect 37247 -4485 37259 -4451
rect 36859 -4491 37259 -4485
rect 37477 -4451 37877 -4445
rect 37477 -4485 37489 -4451
rect 37865 -4485 37877 -4451
rect 37477 -4491 37877 -4485
rect 59 -4709 480 -4703
rect 59 -4743 71 -4709
rect 447 -4743 480 -4709
rect 59 -4749 480 -4743
rect 440 -4780 480 -4749
rect 660 -4703 710 -4491
rect 1109 -4530 1155 -4518
rect 1581 -4530 1627 -4518
rect 2091 -4530 2137 -4518
rect 2199 -4530 2245 -4518
rect 2709 -4530 2755 -4518
rect 3181 -4530 3227 -4518
rect 3691 -4530 3737 -4518
rect 3799 -4530 3845 -4518
rect 4309 -4530 4355 -4518
rect 4781 -4530 4827 -4518
rect 5291 -4530 5337 -4518
rect 5399 -4530 5445 -4518
rect 5909 -4530 5955 -4518
rect 6381 -4530 6427 -4518
rect 6891 -4530 6937 -4518
rect 6999 -4530 7045 -4518
rect 7509 -4530 7555 -4518
rect 7981 -4530 8027 -4518
rect 8491 -4530 8537 -4518
rect 8599 -4530 8645 -4518
rect 9109 -4530 9155 -4518
rect 9581 -4530 9627 -4518
rect 10091 -4530 10137 -4518
rect 10199 -4530 10245 -4518
rect 10709 -4530 10755 -4518
rect 11181 -4530 11227 -4518
rect 11691 -4530 11737 -4518
rect 11799 -4530 11845 -4518
rect 12309 -4520 12355 -4518
rect 12309 -4530 12520 -4520
rect 12781 -4530 12827 -4518
rect 13291 -4530 13337 -4518
rect 13399 -4530 13445 -4518
rect 13909 -4530 13955 -4518
rect 14381 -4530 14427 -4518
rect 14891 -4530 14937 -4518
rect 14999 -4530 15045 -4518
rect 15509 -4530 15555 -4518
rect 15981 -4530 16027 -4518
rect 16491 -4530 16537 -4518
rect 16599 -4530 16645 -4518
rect 17109 -4530 17155 -4518
rect 17581 -4530 17627 -4518
rect 18091 -4530 18137 -4518
rect 18199 -4530 18245 -4518
rect 18709 -4530 18755 -4518
rect 19181 -4530 19227 -4518
rect 19691 -4530 19737 -4518
rect 19799 -4530 19845 -4518
rect 20309 -4530 20355 -4518
rect 20781 -4530 20827 -4518
rect 21291 -4530 21337 -4518
rect 21399 -4530 21445 -4518
rect 21909 -4530 21955 -4518
rect 22381 -4530 22427 -4518
rect 22891 -4530 22937 -4518
rect 22999 -4530 23045 -4518
rect 23509 -4530 23555 -4518
rect 23981 -4530 24027 -4518
rect 24491 -4530 24537 -4518
rect 24599 -4530 24645 -4518
rect 25109 -4530 25155 -4518
rect 25581 -4530 25627 -4518
rect 26091 -4530 26137 -4518
rect 26199 -4530 26245 -4518
rect 26709 -4530 26755 -4518
rect 27181 -4530 27227 -4518
rect 27691 -4530 27737 -4518
rect 27799 -4530 27845 -4518
rect 28309 -4530 28355 -4518
rect 28781 -4530 28827 -4518
rect 29291 -4530 29337 -4518
rect 29399 -4530 29445 -4518
rect 29909 -4530 29955 -4518
rect 30381 -4530 30427 -4518
rect 30891 -4530 30937 -4518
rect 30999 -4530 31045 -4518
rect 31509 -4530 31555 -4518
rect 31981 -4530 32027 -4518
rect 32491 -4530 32537 -4518
rect 32599 -4530 32645 -4518
rect 33109 -4530 33155 -4518
rect 33581 -4530 33627 -4518
rect 34091 -4530 34137 -4518
rect 34199 -4530 34245 -4518
rect 34709 -4530 34755 -4518
rect 35181 -4530 35227 -4518
rect 35691 -4530 35737 -4518
rect 35799 -4530 35845 -4518
rect 36309 -4530 36355 -4518
rect 36781 -4530 36827 -4518
rect 1109 -4664 1115 -4530
rect 1149 -4664 1155 -4530
rect 1540 -4660 1587 -4530
rect 1109 -4676 1155 -4664
rect 1581 -4664 1587 -4660
rect 1621 -4660 2097 -4530
rect 1621 -4664 1627 -4660
rect 1581 -4676 1627 -4664
rect 2091 -4664 2097 -4660
rect 2131 -4660 2205 -4530
rect 2131 -4664 2137 -4660
rect 2091 -4676 2137 -4664
rect 2199 -4664 2205 -4660
rect 2239 -4660 2715 -4530
rect 2239 -4664 2245 -4660
rect 2199 -4676 2245 -4664
rect 2709 -4664 2715 -4660
rect 2749 -4660 3187 -4530
rect 2749 -4664 2755 -4660
rect 2709 -4676 2755 -4664
rect 3181 -4664 3187 -4660
rect 3221 -4660 3697 -4530
rect 3221 -4664 3227 -4660
rect 3181 -4676 3227 -4664
rect 3691 -4664 3697 -4660
rect 3731 -4660 3805 -4530
rect 3731 -4664 3737 -4660
rect 3691 -4676 3737 -4664
rect 3799 -4664 3805 -4660
rect 3839 -4660 4315 -4530
rect 3839 -4664 3845 -4660
rect 3799 -4676 3845 -4664
rect 4309 -4664 4315 -4660
rect 4349 -4660 4787 -4530
rect 4349 -4664 4355 -4660
rect 4309 -4676 4355 -4664
rect 4781 -4664 4787 -4660
rect 4821 -4660 5297 -4530
rect 4821 -4664 4827 -4660
rect 4781 -4676 4827 -4664
rect 5291 -4664 5297 -4660
rect 5331 -4660 5405 -4530
rect 5331 -4664 5337 -4660
rect 5291 -4676 5337 -4664
rect 5399 -4664 5405 -4660
rect 5439 -4660 5915 -4530
rect 5439 -4664 5445 -4660
rect 5399 -4676 5445 -4664
rect 5909 -4664 5915 -4660
rect 5949 -4660 6387 -4530
rect 5949 -4664 5955 -4660
rect 5909 -4676 5955 -4664
rect 6381 -4664 6387 -4660
rect 6421 -4660 6897 -4530
rect 6421 -4664 6427 -4660
rect 6381 -4676 6427 -4664
rect 6891 -4664 6897 -4660
rect 6931 -4660 7005 -4530
rect 6931 -4664 6937 -4660
rect 6891 -4676 6937 -4664
rect 6999 -4664 7005 -4660
rect 7039 -4660 7515 -4530
rect 7039 -4664 7045 -4660
rect 6999 -4676 7045 -4664
rect 7509 -4664 7515 -4660
rect 7549 -4660 7987 -4530
rect 7549 -4664 7555 -4660
rect 7509 -4676 7555 -4664
rect 7981 -4664 7987 -4660
rect 8021 -4660 8497 -4530
rect 8021 -4664 8027 -4660
rect 7981 -4676 8027 -4664
rect 8491 -4664 8497 -4660
rect 8531 -4660 8605 -4530
rect 8531 -4664 8537 -4660
rect 8491 -4676 8537 -4664
rect 8599 -4664 8605 -4660
rect 8639 -4660 9115 -4530
rect 8639 -4664 8645 -4660
rect 8599 -4676 8645 -4664
rect 9109 -4664 9115 -4660
rect 9149 -4660 9587 -4530
rect 9149 -4664 9155 -4660
rect 9109 -4676 9155 -4664
rect 9581 -4664 9587 -4660
rect 9621 -4660 10097 -4530
rect 9621 -4664 9627 -4660
rect 9581 -4676 9627 -4664
rect 10091 -4664 10097 -4660
rect 10131 -4660 10205 -4530
rect 10131 -4664 10137 -4660
rect 10091 -4676 10137 -4664
rect 10199 -4664 10205 -4660
rect 10239 -4660 10715 -4530
rect 10239 -4664 10245 -4660
rect 10199 -4676 10245 -4664
rect 10709 -4664 10715 -4660
rect 10749 -4660 11187 -4530
rect 10749 -4664 10755 -4660
rect 10709 -4676 10755 -4664
rect 11181 -4664 11187 -4660
rect 11221 -4660 11697 -4530
rect 11221 -4664 11227 -4660
rect 11181 -4676 11227 -4664
rect 11691 -4664 11697 -4660
rect 11731 -4660 11805 -4530
rect 11731 -4664 11737 -4660
rect 11691 -4676 11737 -4664
rect 11799 -4664 11805 -4660
rect 11839 -4660 12315 -4530
rect 11839 -4664 11845 -4660
rect 11799 -4676 11845 -4664
rect 12309 -4664 12315 -4660
rect 12349 -4650 12390 -4530
rect 12510 -4650 12787 -4530
rect 12349 -4660 12787 -4650
rect 12349 -4664 12355 -4660
rect 12309 -4676 12355 -4664
rect 12781 -4664 12787 -4660
rect 12821 -4660 13297 -4530
rect 12821 -4664 12827 -4660
rect 12781 -4676 12827 -4664
rect 13291 -4664 13297 -4660
rect 13331 -4660 13405 -4530
rect 13331 -4664 13337 -4660
rect 13291 -4676 13337 -4664
rect 13399 -4664 13405 -4660
rect 13439 -4660 13915 -4530
rect 13439 -4664 13445 -4660
rect 13399 -4676 13445 -4664
rect 13909 -4664 13915 -4660
rect 13949 -4660 14387 -4530
rect 13949 -4664 13955 -4660
rect 13909 -4676 13955 -4664
rect 14381 -4664 14387 -4660
rect 14421 -4660 14897 -4530
rect 14421 -4664 14427 -4660
rect 14381 -4676 14427 -4664
rect 14891 -4664 14897 -4660
rect 14931 -4660 15005 -4530
rect 14931 -4664 14937 -4660
rect 14891 -4676 14937 -4664
rect 14999 -4664 15005 -4660
rect 15039 -4660 15515 -4530
rect 15039 -4664 15045 -4660
rect 14999 -4676 15045 -4664
rect 15509 -4664 15515 -4660
rect 15549 -4660 15987 -4530
rect 15549 -4664 15555 -4660
rect 15509 -4676 15555 -4664
rect 15981 -4664 15987 -4660
rect 16021 -4660 16497 -4530
rect 16021 -4664 16027 -4660
rect 15981 -4676 16027 -4664
rect 16491 -4664 16497 -4660
rect 16531 -4660 16605 -4530
rect 16531 -4664 16537 -4660
rect 16491 -4676 16537 -4664
rect 16599 -4664 16605 -4660
rect 16639 -4660 17115 -4530
rect 16639 -4664 16645 -4660
rect 16599 -4676 16645 -4664
rect 17109 -4664 17115 -4660
rect 17149 -4660 17587 -4530
rect 17149 -4664 17155 -4660
rect 17109 -4676 17155 -4664
rect 17581 -4664 17587 -4660
rect 17621 -4660 18097 -4530
rect 17621 -4664 17627 -4660
rect 17581 -4676 17627 -4664
rect 18091 -4664 18097 -4660
rect 18131 -4660 18205 -4530
rect 18131 -4664 18137 -4660
rect 18091 -4676 18137 -4664
rect 18199 -4664 18205 -4660
rect 18239 -4660 18715 -4530
rect 18239 -4664 18245 -4660
rect 18199 -4676 18245 -4664
rect 18709 -4664 18715 -4660
rect 18749 -4660 19187 -4530
rect 18749 -4664 18755 -4660
rect 18709 -4676 18755 -4664
rect 19181 -4664 19187 -4660
rect 19221 -4660 19697 -4530
rect 19221 -4664 19227 -4660
rect 19181 -4676 19227 -4664
rect 19691 -4664 19697 -4660
rect 19731 -4660 19805 -4530
rect 19731 -4664 19737 -4660
rect 19691 -4676 19737 -4664
rect 19799 -4664 19805 -4660
rect 19839 -4660 20315 -4530
rect 19839 -4664 19845 -4660
rect 19799 -4676 19845 -4664
rect 20309 -4664 20315 -4660
rect 20349 -4660 20787 -4530
rect 20349 -4664 20355 -4660
rect 20309 -4676 20355 -4664
rect 20781 -4664 20787 -4660
rect 20821 -4660 21297 -4530
rect 20821 -4664 20827 -4660
rect 20781 -4676 20827 -4664
rect 21291 -4664 21297 -4660
rect 21331 -4660 21405 -4530
rect 21331 -4664 21337 -4660
rect 21291 -4676 21337 -4664
rect 21399 -4664 21405 -4660
rect 21439 -4660 21915 -4530
rect 21439 -4664 21445 -4660
rect 21399 -4676 21445 -4664
rect 21909 -4664 21915 -4660
rect 21949 -4660 22387 -4530
rect 21949 -4664 21955 -4660
rect 21909 -4676 21955 -4664
rect 22381 -4664 22387 -4660
rect 22421 -4660 22897 -4530
rect 22421 -4664 22427 -4660
rect 22381 -4676 22427 -4664
rect 22891 -4664 22897 -4660
rect 22931 -4660 23005 -4530
rect 22931 -4664 22937 -4660
rect 22891 -4676 22937 -4664
rect 22999 -4664 23005 -4660
rect 23039 -4660 23515 -4530
rect 23039 -4664 23045 -4660
rect 22999 -4676 23045 -4664
rect 23509 -4664 23515 -4660
rect 23549 -4660 23987 -4530
rect 23549 -4664 23555 -4660
rect 23509 -4676 23555 -4664
rect 23981 -4664 23987 -4660
rect 24021 -4660 24497 -4530
rect 24021 -4664 24027 -4660
rect 23981 -4676 24027 -4664
rect 24491 -4664 24497 -4660
rect 24531 -4660 24605 -4530
rect 24531 -4664 24537 -4660
rect 24491 -4676 24537 -4664
rect 24599 -4664 24605 -4660
rect 24639 -4660 25115 -4530
rect 24639 -4664 24645 -4660
rect 24599 -4676 24645 -4664
rect 25109 -4664 25115 -4660
rect 25149 -4660 25587 -4530
rect 25149 -4664 25155 -4660
rect 25109 -4676 25155 -4664
rect 25581 -4664 25587 -4660
rect 25621 -4660 26097 -4530
rect 25621 -4664 25627 -4660
rect 25581 -4676 25627 -4664
rect 26091 -4664 26097 -4660
rect 26131 -4660 26205 -4530
rect 26131 -4664 26137 -4660
rect 26091 -4676 26137 -4664
rect 26199 -4664 26205 -4660
rect 26239 -4660 26715 -4530
rect 26239 -4664 26245 -4660
rect 26199 -4676 26245 -4664
rect 26709 -4664 26715 -4660
rect 26749 -4660 27187 -4530
rect 26749 -4664 26755 -4660
rect 26709 -4676 26755 -4664
rect 27181 -4664 27187 -4660
rect 27221 -4660 27697 -4530
rect 27221 -4664 27227 -4660
rect 27181 -4676 27227 -4664
rect 27691 -4664 27697 -4660
rect 27731 -4660 27805 -4530
rect 27731 -4664 27737 -4660
rect 27691 -4676 27737 -4664
rect 27799 -4664 27805 -4660
rect 27839 -4660 28315 -4530
rect 27839 -4664 27845 -4660
rect 27799 -4676 27845 -4664
rect 28309 -4664 28315 -4660
rect 28349 -4660 28787 -4530
rect 28349 -4664 28355 -4660
rect 28309 -4676 28355 -4664
rect 28781 -4664 28787 -4660
rect 28821 -4660 29297 -4530
rect 28821 -4664 28827 -4660
rect 28781 -4676 28827 -4664
rect 29291 -4664 29297 -4660
rect 29331 -4660 29405 -4530
rect 29331 -4664 29337 -4660
rect 29291 -4676 29337 -4664
rect 29399 -4664 29405 -4660
rect 29439 -4660 29915 -4530
rect 29439 -4664 29445 -4660
rect 29399 -4676 29445 -4664
rect 29909 -4664 29915 -4660
rect 29949 -4660 30387 -4530
rect 29949 -4664 29955 -4660
rect 29909 -4676 29955 -4664
rect 30381 -4664 30387 -4660
rect 30421 -4660 30897 -4530
rect 30421 -4664 30427 -4660
rect 30381 -4676 30427 -4664
rect 30891 -4664 30897 -4660
rect 30931 -4660 31005 -4530
rect 30931 -4664 30937 -4660
rect 30891 -4676 30937 -4664
rect 30999 -4664 31005 -4660
rect 31039 -4660 31515 -4530
rect 31039 -4664 31045 -4660
rect 30999 -4676 31045 -4664
rect 31509 -4664 31515 -4660
rect 31549 -4660 31987 -4530
rect 31549 -4664 31555 -4660
rect 31509 -4676 31555 -4664
rect 31981 -4664 31987 -4660
rect 32021 -4660 32497 -4530
rect 32021 -4664 32027 -4660
rect 31981 -4676 32027 -4664
rect 32491 -4664 32497 -4660
rect 32531 -4660 32605 -4530
rect 32531 -4664 32537 -4660
rect 32491 -4676 32537 -4664
rect 32599 -4664 32605 -4660
rect 32639 -4660 33115 -4530
rect 32639 -4664 32645 -4660
rect 32599 -4676 32645 -4664
rect 33109 -4664 33115 -4660
rect 33149 -4660 33587 -4530
rect 33149 -4664 33155 -4660
rect 33109 -4676 33155 -4664
rect 33581 -4664 33587 -4660
rect 33621 -4660 34097 -4530
rect 33621 -4664 33627 -4660
rect 33581 -4676 33627 -4664
rect 34091 -4664 34097 -4660
rect 34131 -4660 34205 -4530
rect 34131 -4664 34137 -4660
rect 34091 -4676 34137 -4664
rect 34199 -4664 34205 -4660
rect 34239 -4660 34715 -4530
rect 34239 -4664 34245 -4660
rect 34199 -4676 34245 -4664
rect 34709 -4664 34715 -4660
rect 34749 -4660 35187 -4530
rect 34749 -4664 34755 -4660
rect 34709 -4676 34755 -4664
rect 35181 -4664 35187 -4660
rect 35221 -4660 35697 -4530
rect 35221 -4664 35227 -4660
rect 35181 -4676 35227 -4664
rect 35691 -4664 35697 -4660
rect 35731 -4660 35805 -4530
rect 35731 -4664 35737 -4660
rect 35691 -4676 35737 -4664
rect 35799 -4664 35805 -4660
rect 35839 -4660 36315 -4530
rect 35839 -4664 35845 -4660
rect 35799 -4676 35845 -4664
rect 36309 -4664 36315 -4660
rect 36349 -4660 36400 -4530
rect 36349 -4664 36355 -4660
rect 36309 -4676 36355 -4664
rect 36781 -4664 36787 -4530
rect 36821 -4664 36827 -4530
rect 36781 -4676 36827 -4664
rect 37291 -4530 37337 -4518
rect 37291 -4664 37297 -4530
rect 37331 -4664 37337 -4530
rect 37291 -4676 37337 -4664
rect 37399 -4530 37445 -4518
rect 37399 -4664 37405 -4530
rect 37439 -4664 37445 -4530
rect 37399 -4676 37445 -4664
rect 37909 -4530 37955 -4518
rect 37909 -4664 37915 -4530
rect 37949 -4664 37955 -4530
rect 37909 -4676 37955 -4664
rect 660 -4709 1077 -4703
rect 660 -4743 689 -4709
rect 1065 -4743 1077 -4709
rect 1659 -4709 2059 -4703
rect 660 -4749 1077 -4743
rect 1180 -4720 1320 -4710
rect 1659 -4720 1671 -4709
rect 660 -4780 710 -4749
rect 440 -4800 710 -4780
rect 1180 -4840 1190 -4720
rect 1310 -4743 1671 -4720
rect 2047 -4720 2059 -4709
rect 2277 -4709 2677 -4703
rect 2277 -4720 2289 -4709
rect 2047 -4743 2289 -4720
rect 2665 -4720 2677 -4709
rect 3259 -4709 3659 -4703
rect 2780 -4720 2920 -4710
rect 3259 -4720 3271 -4709
rect 2665 -4743 2790 -4720
rect 1310 -4840 2790 -4743
rect 2910 -4743 3271 -4720
rect 3647 -4720 3659 -4709
rect 3877 -4709 4277 -4703
rect 3877 -4720 3889 -4709
rect 3647 -4743 3889 -4720
rect 4265 -4720 4277 -4709
rect 4859 -4709 5259 -4703
rect 4380 -4720 4520 -4710
rect 4859 -4720 4871 -4709
rect 4265 -4743 4390 -4720
rect 2910 -4840 4390 -4743
rect 4510 -4743 4871 -4720
rect 5247 -4720 5259 -4709
rect 5477 -4709 5877 -4703
rect 5477 -4720 5489 -4709
rect 5247 -4743 5489 -4720
rect 5865 -4720 5877 -4709
rect 6459 -4709 6859 -4703
rect 5980 -4720 6120 -4710
rect 6459 -4720 6471 -4709
rect 5865 -4743 5990 -4720
rect 4510 -4840 5990 -4743
rect 6110 -4743 6471 -4720
rect 6847 -4720 6859 -4709
rect 7077 -4709 7477 -4703
rect 7077 -4720 7089 -4709
rect 6847 -4743 7089 -4720
rect 7465 -4720 7477 -4709
rect 8059 -4709 8459 -4703
rect 7580 -4720 7720 -4710
rect 8059 -4720 8071 -4709
rect 7465 -4743 7590 -4720
rect 6110 -4840 7590 -4743
rect 7710 -4743 8071 -4720
rect 8447 -4720 8459 -4709
rect 8677 -4709 9077 -4703
rect 8677 -4720 8689 -4709
rect 8447 -4743 8689 -4720
rect 9065 -4720 9077 -4709
rect 9659 -4709 10059 -4703
rect 9180 -4720 9320 -4710
rect 9659 -4720 9671 -4709
rect 9065 -4743 9190 -4720
rect 7710 -4840 9190 -4743
rect 9310 -4743 9671 -4720
rect 10047 -4720 10059 -4709
rect 10277 -4709 10677 -4703
rect 10277 -4720 10289 -4709
rect 10047 -4743 10289 -4720
rect 10665 -4720 10677 -4709
rect 11259 -4709 11659 -4703
rect 11259 -4720 11271 -4709
rect 10665 -4743 10720 -4720
rect 9310 -4840 10720 -4743
rect 11220 -4743 11271 -4720
rect 11647 -4720 11659 -4709
rect 11877 -4709 12277 -4703
rect 11877 -4720 11889 -4709
rect 11647 -4743 11889 -4720
rect 12265 -4720 12277 -4709
rect 12859 -4709 13259 -4703
rect 12265 -4743 12350 -4720
rect 11220 -4810 12350 -4743
rect 11220 -4840 11710 -4810
rect 1180 -4850 1320 -4840
rect 2780 -4850 2920 -4840
rect 4380 -4850 4520 -4840
rect 5980 -4850 6120 -4840
rect 7580 -4850 7720 -4840
rect 9180 -4850 9320 -4840
rect 11700 -4930 11710 -4840
rect 11830 -4840 12350 -4810
rect 12600 -4730 12740 -4720
rect 11830 -4930 11840 -4840
rect 12600 -4850 12610 -4730
rect 12730 -4740 12740 -4730
rect 12859 -4740 12871 -4709
rect 12730 -4743 12871 -4740
rect 13247 -4740 13259 -4709
rect 13477 -4709 13877 -4703
rect 13477 -4720 13489 -4709
rect 13247 -4743 13260 -4740
rect 12730 -4840 13260 -4743
rect 13470 -4743 13489 -4720
rect 13865 -4720 13877 -4709
rect 14459 -4709 14859 -4703
rect 13865 -4743 13890 -4720
rect 13470 -4790 13890 -4743
rect 13470 -4840 13630 -4790
rect 12730 -4850 12740 -4840
rect 12600 -4860 12740 -4850
rect 13620 -4910 13630 -4840
rect 13750 -4840 13890 -4790
rect 14200 -4730 14340 -4720
rect 13750 -4910 13760 -4840
rect 14200 -4850 14210 -4730
rect 14330 -4740 14340 -4730
rect 14459 -4740 14471 -4709
rect 14330 -4743 14471 -4740
rect 14847 -4740 14859 -4709
rect 15077 -4709 15477 -4703
rect 15077 -4720 15089 -4709
rect 14847 -4743 14860 -4740
rect 14330 -4840 14860 -4743
rect 15070 -4743 15089 -4720
rect 15465 -4720 15477 -4709
rect 16059 -4709 16459 -4703
rect 15810 -4720 15930 -4710
rect 16059 -4720 16071 -4709
rect 15465 -4743 15490 -4720
rect 15070 -4790 15490 -4743
rect 15070 -4840 15230 -4790
rect 14330 -4850 14340 -4840
rect 14200 -4860 14340 -4850
rect 13620 -4920 13760 -4910
rect 15220 -4910 15230 -4840
rect 15350 -4840 15490 -4790
rect 15810 -4840 15820 -4720
rect 15920 -4743 16071 -4720
rect 16447 -4720 16459 -4709
rect 16677 -4709 17077 -4703
rect 16677 -4720 16689 -4709
rect 16447 -4743 16689 -4720
rect 17065 -4720 17077 -4709
rect 17659 -4709 18059 -4703
rect 17410 -4720 17530 -4710
rect 17659 -4720 17671 -4709
rect 17065 -4743 17120 -4720
rect 15920 -4840 17120 -4743
rect 17410 -4840 17420 -4720
rect 17520 -4743 17671 -4720
rect 18047 -4720 18059 -4709
rect 18277 -4709 18677 -4703
rect 18277 -4720 18289 -4709
rect 18047 -4743 18289 -4720
rect 18665 -4720 18677 -4709
rect 19259 -4709 19659 -4703
rect 19010 -4720 19130 -4710
rect 19259 -4720 19271 -4709
rect 18665 -4743 18720 -4720
rect 17520 -4840 18720 -4743
rect 19010 -4840 19020 -4720
rect 19120 -4743 19271 -4720
rect 19647 -4720 19659 -4709
rect 19877 -4709 20277 -4703
rect 19877 -4720 19889 -4709
rect 19647 -4743 19889 -4720
rect 20265 -4720 20277 -4709
rect 20859 -4709 21259 -4703
rect 20610 -4720 20730 -4710
rect 20859 -4720 20871 -4709
rect 20265 -4743 20320 -4720
rect 19120 -4840 20320 -4743
rect 20610 -4840 20620 -4720
rect 20720 -4743 20871 -4720
rect 21247 -4720 21259 -4709
rect 21477 -4709 21877 -4703
rect 21477 -4720 21489 -4709
rect 21247 -4743 21489 -4720
rect 21865 -4720 21877 -4709
rect 22459 -4709 22859 -4703
rect 22210 -4720 22330 -4710
rect 22459 -4720 22471 -4709
rect 21865 -4743 21920 -4720
rect 20720 -4840 21920 -4743
rect 22210 -4840 22220 -4720
rect 22320 -4743 22471 -4720
rect 22847 -4720 22859 -4709
rect 23077 -4709 23477 -4703
rect 23077 -4720 23089 -4709
rect 22847 -4743 23089 -4720
rect 23465 -4720 23477 -4709
rect 24059 -4709 24459 -4703
rect 23810 -4720 23930 -4710
rect 24059 -4720 24071 -4709
rect 23465 -4743 23520 -4720
rect 22320 -4840 23520 -4743
rect 23810 -4840 23820 -4720
rect 23920 -4743 24071 -4720
rect 24447 -4720 24459 -4709
rect 24677 -4709 25077 -4703
rect 24677 -4720 24689 -4709
rect 24447 -4743 24689 -4720
rect 25065 -4720 25077 -4709
rect 25659 -4709 26059 -4703
rect 25410 -4720 25530 -4710
rect 25659 -4720 25671 -4709
rect 25065 -4743 25120 -4720
rect 23920 -4840 25120 -4743
rect 25410 -4840 25420 -4720
rect 25520 -4743 25671 -4720
rect 26047 -4720 26059 -4709
rect 26277 -4709 26677 -4703
rect 26277 -4720 26289 -4709
rect 26047 -4743 26289 -4720
rect 26665 -4720 26677 -4709
rect 27259 -4709 27659 -4703
rect 27011 -4720 27130 -4710
rect 27259 -4720 27271 -4709
rect 26665 -4743 26720 -4720
rect 25520 -4840 26720 -4743
rect 27011 -4840 27020 -4720
rect 27120 -4743 27271 -4720
rect 27647 -4720 27659 -4709
rect 27877 -4709 28277 -4703
rect 27877 -4720 27889 -4709
rect 27647 -4743 27889 -4720
rect 28265 -4720 28277 -4709
rect 28859 -4709 29259 -4703
rect 28611 -4720 28730 -4710
rect 28859 -4720 28871 -4709
rect 28265 -4743 28320 -4720
rect 27120 -4840 28320 -4743
rect 28611 -4840 28620 -4720
rect 28720 -4743 28871 -4720
rect 29247 -4720 29259 -4709
rect 29477 -4709 29877 -4703
rect 29477 -4720 29489 -4709
rect 29247 -4743 29489 -4720
rect 29865 -4720 29877 -4709
rect 30459 -4709 30859 -4703
rect 30211 -4720 30330 -4710
rect 30459 -4720 30471 -4709
rect 29865 -4743 29920 -4720
rect 28720 -4840 29920 -4743
rect 30211 -4840 30220 -4720
rect 30320 -4743 30471 -4720
rect 30847 -4720 30859 -4709
rect 31077 -4709 31477 -4703
rect 31077 -4720 31089 -4709
rect 30847 -4743 31089 -4720
rect 31465 -4720 31477 -4709
rect 32059 -4709 32459 -4703
rect 31465 -4743 31520 -4720
rect 30320 -4840 31520 -4743
rect 32059 -4743 32071 -4709
rect 32447 -4720 32459 -4709
rect 32677 -4709 33077 -4703
rect 32677 -4720 32689 -4709
rect 32447 -4743 32689 -4720
rect 33065 -4720 33077 -4709
rect 33659 -4709 34059 -4703
rect 33659 -4720 33671 -4709
rect 33065 -4743 33671 -4720
rect 34047 -4720 34059 -4709
rect 34277 -4709 34677 -4703
rect 34277 -4720 34289 -4709
rect 34047 -4743 34289 -4720
rect 34665 -4720 34677 -4709
rect 35259 -4709 35659 -4703
rect 35259 -4720 35271 -4709
rect 34665 -4743 35271 -4720
rect 35647 -4720 35659 -4709
rect 35877 -4709 36277 -4703
rect 35877 -4720 35889 -4709
rect 35647 -4743 35889 -4720
rect 36265 -4720 36277 -4709
rect 36390 -4710 36510 -4700
rect 36390 -4720 36400 -4710
rect 36265 -4743 36400 -4720
rect 32059 -4749 36400 -4743
rect 32060 -4830 36400 -4749
rect 36500 -4830 36510 -4710
rect 36859 -4709 37259 -4703
rect 36859 -4743 36871 -4709
rect 37247 -4743 37259 -4709
rect 36859 -4749 37259 -4743
rect 37477 -4709 37877 -4703
rect 37477 -4743 37489 -4709
rect 37865 -4743 37877 -4709
rect 37477 -4749 37877 -4743
rect 32060 -4840 36510 -4830
rect 15350 -4910 15360 -4840
rect 15810 -4850 15930 -4840
rect 17410 -4850 17530 -4840
rect 19010 -4850 19130 -4840
rect 20610 -4850 20730 -4840
rect 22210 -4850 22330 -4840
rect 23810 -4850 23930 -4840
rect 25410 -4850 25530 -4840
rect 27011 -4850 27130 -4840
rect 28611 -4850 28730 -4840
rect 30211 -4850 30330 -4840
rect 15220 -4920 15360 -4910
rect 11700 -4940 11840 -4930
rect 11700 -5830 11840 -5820
rect 11700 -5950 11710 -5830
rect 11830 -5840 11840 -5830
rect 13300 -5830 13440 -5820
rect 13300 -5840 13310 -5830
rect 11830 -5940 13310 -5840
rect 11830 -5950 11840 -5940
rect 11700 -5960 11840 -5950
rect 13300 -5950 13310 -5940
rect 13430 -5950 13440 -5830
rect 13300 -5960 13440 -5950
rect 11700 -6050 11840 -6040
rect 11700 -6170 11710 -6050
rect 11830 -6060 11840 -6050
rect 13620 -6050 13760 -6040
rect 13620 -6060 13630 -6050
rect 11830 -6160 13630 -6060
rect 11830 -6170 11840 -6160
rect 11700 -6180 11840 -6170
rect 13620 -6170 13630 -6160
rect 13750 -6170 13760 -6050
rect 13620 -6180 13760 -6170
rect 14220 -6050 14360 -6040
rect 14220 -6170 14230 -6050
rect 14350 -6060 14360 -6050
rect 15220 -6050 15360 -6040
rect 15220 -6060 15230 -6050
rect 14350 -6160 15230 -6060
rect 14350 -6170 14360 -6160
rect 14220 -6180 14360 -6170
rect 15220 -6170 15230 -6160
rect 15350 -6170 15360 -6050
rect 15220 -6180 15360 -6170
rect 12620 -6270 12760 -6260
rect 12620 -6390 12630 -6270
rect 12750 -6280 12760 -6270
rect 16500 -6270 16640 -6260
rect 16500 -6280 16510 -6270
rect 12750 -6380 16510 -6280
rect 12750 -6390 12760 -6380
rect 12620 -6400 12760 -6390
rect 16500 -6390 16510 -6380
rect 16630 -6390 16640 -6270
rect 16500 -6400 16640 -6390
rect 12400 -6490 12540 -6480
rect 12400 -6610 12410 -6490
rect 12530 -6500 12540 -6490
rect 14900 -6490 15040 -6480
rect 14900 -6500 14910 -6490
rect 12530 -6600 14910 -6500
rect 12530 -6610 12540 -6600
rect 12400 -6620 12540 -6610
rect 14900 -6610 14910 -6600
rect 15030 -6610 15040 -6490
rect 14900 -6620 15040 -6610
rect 12940 -6830 13120 -6820
rect 12940 -6900 12950 -6830
rect 440 -6990 12950 -6900
rect 13110 -6990 13120 -6830
rect 440 -8090 720 -6990
rect 12940 -7000 13120 -6990
rect 7800 -7870 7940 -7860
rect 7800 -7990 7810 -7870
rect 7930 -7880 7940 -7870
rect 14900 -7880 15050 -7870
rect 7930 -7990 14910 -7880
rect 7800 -8000 14910 -7990
rect 15040 -8000 15050 -7880
rect 14900 -8010 15050 -8000
rect 440 -8164 490 -8090
rect 57 -8170 490 -8164
rect 57 -8204 69 -8170
rect 445 -8204 490 -8170
rect 57 -8210 490 -8204
rect -30 -8257 16 -8245
rect -30 -8375 -24 -8257
rect 10 -8375 16 -8257
rect -30 -8387 16 -8375
rect 440 -8422 490 -8210
rect 670 -8164 720 -8090
rect 1200 -8070 1340 -8060
rect 670 -8170 1093 -8164
rect 670 -8204 705 -8170
rect 1081 -8204 1093 -8170
rect 1200 -8190 1210 -8070
rect 1330 -8080 1340 -8070
rect 2800 -8070 2940 -8060
rect 2800 -8080 2810 -8070
rect 1330 -8170 2810 -8080
rect 1330 -8180 1669 -8170
rect 1330 -8190 1340 -8180
rect 1200 -8200 1340 -8190
rect 670 -8210 1093 -8204
rect 1657 -8204 1669 -8180
rect 2045 -8180 2305 -8170
rect 2045 -8204 2057 -8180
rect 1657 -8210 2057 -8204
rect 2293 -8204 2305 -8180
rect 2681 -8180 2810 -8170
rect 2681 -8204 2693 -8180
rect 2800 -8190 2810 -8180
rect 2930 -8080 2940 -8070
rect 4400 -8070 4540 -8060
rect 4400 -8080 4410 -8070
rect 2930 -8170 4410 -8080
rect 2930 -8180 3269 -8170
rect 2930 -8190 2940 -8180
rect 2800 -8200 2940 -8190
rect 2293 -8210 2693 -8204
rect 3257 -8204 3269 -8180
rect 3645 -8180 3905 -8170
rect 3645 -8204 3657 -8180
rect 3257 -8210 3657 -8204
rect 3893 -8204 3905 -8180
rect 4281 -8180 4410 -8170
rect 4281 -8204 4293 -8180
rect 4400 -8190 4410 -8180
rect 4530 -8080 4540 -8070
rect 6000 -8070 6140 -8060
rect 6000 -8080 6010 -8070
rect 4530 -8170 6010 -8080
rect 4530 -8180 4869 -8170
rect 4530 -8190 4540 -8180
rect 4400 -8200 4540 -8190
rect 3893 -8210 4293 -8204
rect 4857 -8204 4869 -8180
rect 5245 -8180 5505 -8170
rect 5245 -8204 5257 -8180
rect 4857 -8210 5257 -8204
rect 5493 -8204 5505 -8180
rect 5881 -8180 6010 -8170
rect 5881 -8204 5893 -8180
rect 6000 -8190 6010 -8180
rect 6130 -8080 6140 -8070
rect 7600 -8070 7740 -8060
rect 7600 -8080 7610 -8070
rect 6130 -8170 7610 -8080
rect 6130 -8180 6469 -8170
rect 6130 -8190 6140 -8180
rect 6000 -8200 6140 -8190
rect 5493 -8210 5893 -8204
rect 6457 -8204 6469 -8180
rect 6845 -8180 7105 -8170
rect 6845 -8204 6857 -8180
rect 6457 -8210 6857 -8204
rect 7093 -8204 7105 -8180
rect 7481 -8180 7610 -8170
rect 7481 -8204 7493 -8180
rect 7600 -8190 7610 -8180
rect 7730 -8080 7740 -8070
rect 9200 -8070 9340 -8060
rect 9200 -8080 9210 -8070
rect 7730 -8170 9210 -8080
rect 7730 -8180 8069 -8170
rect 7730 -8190 7740 -8180
rect 7600 -8200 7740 -8190
rect 7093 -8210 7493 -8204
rect 8057 -8204 8069 -8180
rect 8445 -8180 8705 -8170
rect 8445 -8204 8457 -8180
rect 8057 -8210 8457 -8204
rect 8693 -8204 8705 -8180
rect 9081 -8180 9210 -8170
rect 9081 -8204 9093 -8180
rect 9200 -8190 9210 -8180
rect 9330 -8080 9340 -8070
rect 15820 -8070 15960 -8060
rect 9330 -8170 10700 -8080
rect 11270 -8110 15480 -8100
rect 11270 -8164 11710 -8110
rect 9330 -8180 9669 -8170
rect 9330 -8190 9340 -8180
rect 9200 -8200 9340 -8190
rect 8693 -8210 9093 -8204
rect 9657 -8204 9669 -8180
rect 10045 -8180 10305 -8170
rect 10045 -8204 10057 -8180
rect 9657 -8210 10057 -8204
rect 10293 -8204 10305 -8180
rect 10681 -8180 10700 -8170
rect 11257 -8170 11710 -8164
rect 10681 -8204 10693 -8180
rect 10293 -8210 10693 -8204
rect 11257 -8204 11269 -8170
rect 11645 -8200 11710 -8170
rect 11645 -8204 11657 -8200
rect 11257 -8210 11657 -8204
rect 57 -8428 490 -8422
rect 57 -8462 69 -8428
rect 445 -8462 490 -8428
rect 57 -8468 490 -8462
rect 440 -8690 490 -8468
rect 57 -8696 490 -8690
rect 57 -8730 69 -8696
rect 445 -8730 490 -8696
rect 57 -8736 490 -8730
rect -30 -8796 16 -8784
rect -30 -9488 -24 -8796
rect 10 -9488 16 -8796
rect -30 -9500 16 -9488
rect 440 -9548 490 -8736
rect 670 -8422 720 -8210
rect 11690 -8230 11710 -8200
rect 11840 -8164 15480 -8110
rect 11840 -8170 15493 -8164
rect 11840 -8200 11905 -8170
rect 11840 -8230 11860 -8200
rect 11893 -8204 11905 -8200
rect 12281 -8200 12869 -8170
rect 12281 -8204 12293 -8200
rect 11893 -8210 12293 -8204
rect 12857 -8204 12869 -8200
rect 13245 -8200 13505 -8170
rect 13245 -8204 13257 -8200
rect 12857 -8210 13257 -8204
rect 11690 -8240 11860 -8230
rect 13290 -8240 13460 -8200
rect 13493 -8204 13505 -8200
rect 13881 -8200 14469 -8170
rect 13881 -8204 13893 -8200
rect 13493 -8210 13893 -8204
rect 14457 -8204 14469 -8200
rect 14845 -8200 15105 -8170
rect 14845 -8204 14857 -8200
rect 14457 -8210 14857 -8204
rect 14890 -8240 15060 -8200
rect 15093 -8204 15105 -8200
rect 15481 -8204 15493 -8170
rect 15820 -8190 15830 -8070
rect 15950 -8100 15960 -8070
rect 17420 -8070 17560 -8060
rect 15950 -8164 17090 -8100
rect 15950 -8170 17093 -8164
rect 15950 -8190 16069 -8170
rect 15820 -8200 16069 -8190
rect 15093 -8210 15493 -8204
rect 16057 -8204 16069 -8200
rect 16445 -8200 16705 -8170
rect 16445 -8204 16457 -8200
rect 16057 -8210 16457 -8204
rect 16693 -8204 16705 -8200
rect 17081 -8204 17093 -8170
rect 17420 -8190 17430 -8070
rect 17550 -8100 17560 -8070
rect 19020 -8070 19160 -8060
rect 17550 -8164 18690 -8100
rect 17550 -8170 18693 -8164
rect 17550 -8190 17669 -8170
rect 17420 -8200 17669 -8190
rect 16693 -8210 17093 -8204
rect 17657 -8204 17669 -8200
rect 18045 -8200 18305 -8170
rect 18045 -8204 18057 -8200
rect 17657 -8210 18057 -8204
rect 18293 -8204 18305 -8200
rect 18681 -8204 18693 -8170
rect 19020 -8190 19030 -8070
rect 19150 -8100 19160 -8070
rect 20620 -8070 20760 -8060
rect 19150 -8164 20290 -8100
rect 19150 -8170 20293 -8164
rect 19150 -8190 19269 -8170
rect 19020 -8200 19269 -8190
rect 18293 -8210 18693 -8204
rect 19257 -8204 19269 -8200
rect 19645 -8200 19905 -8170
rect 19645 -8204 19657 -8200
rect 19257 -8210 19657 -8204
rect 19893 -8204 19905 -8200
rect 20281 -8204 20293 -8170
rect 20620 -8190 20630 -8070
rect 20750 -8100 20760 -8070
rect 22220 -8070 22360 -8060
rect 20750 -8164 21890 -8100
rect 20750 -8170 21893 -8164
rect 20750 -8190 20869 -8170
rect 20620 -8200 20869 -8190
rect 19893 -8210 20293 -8204
rect 20857 -8204 20869 -8200
rect 21245 -8200 21505 -8170
rect 21245 -8204 21257 -8200
rect 20857 -8210 21257 -8204
rect 21493 -8204 21505 -8200
rect 21881 -8204 21893 -8170
rect 22220 -8190 22230 -8070
rect 22350 -8100 22360 -8070
rect 23820 -8070 23960 -8060
rect 22350 -8164 23490 -8100
rect 22350 -8170 23493 -8164
rect 22350 -8190 22469 -8170
rect 22220 -8200 22469 -8190
rect 21493 -8210 21893 -8204
rect 22457 -8204 22469 -8200
rect 22845 -8200 23105 -8170
rect 22845 -8204 22857 -8200
rect 22457 -8210 22857 -8204
rect 23093 -8204 23105 -8200
rect 23481 -8204 23493 -8170
rect 23820 -8190 23830 -8070
rect 23950 -8100 23960 -8070
rect 25420 -8070 25560 -8060
rect 23950 -8164 25090 -8100
rect 23950 -8170 25093 -8164
rect 23950 -8190 24069 -8170
rect 23820 -8200 24069 -8190
rect 23093 -8210 23493 -8204
rect 24057 -8204 24069 -8200
rect 24445 -8200 24705 -8170
rect 24445 -8204 24457 -8200
rect 24057 -8210 24457 -8204
rect 24693 -8204 24705 -8200
rect 25081 -8204 25093 -8170
rect 25420 -8190 25430 -8070
rect 25550 -8100 25560 -8070
rect 27020 -8070 27160 -8060
rect 25550 -8164 26680 -8100
rect 25550 -8170 26693 -8164
rect 25550 -8190 25669 -8170
rect 25420 -8200 25669 -8190
rect 24693 -8210 25093 -8204
rect 25657 -8204 25669 -8200
rect 26045 -8200 26305 -8170
rect 26045 -8204 26057 -8200
rect 25657 -8210 26057 -8204
rect 26293 -8204 26305 -8200
rect 26681 -8204 26693 -8170
rect 27020 -8190 27030 -8070
rect 27150 -8100 27160 -8070
rect 28620 -8070 28760 -8060
rect 27150 -8164 28290 -8100
rect 27150 -8170 28293 -8164
rect 27150 -8190 27269 -8170
rect 27020 -8200 27269 -8190
rect 26293 -8210 26693 -8204
rect 27257 -8204 27269 -8200
rect 27645 -8200 27905 -8170
rect 27645 -8204 27657 -8200
rect 27257 -8210 27657 -8204
rect 27893 -8204 27905 -8200
rect 28281 -8204 28293 -8170
rect 28620 -8190 28630 -8070
rect 28750 -8100 28760 -8070
rect 30220 -8070 30360 -8060
rect 28750 -8164 29890 -8100
rect 28750 -8170 29893 -8164
rect 28750 -8190 28869 -8170
rect 28620 -8200 28869 -8190
rect 27893 -8210 28293 -8204
rect 28857 -8204 28869 -8200
rect 29245 -8200 29505 -8170
rect 29245 -8204 29257 -8200
rect 28857 -8210 29257 -8204
rect 29493 -8204 29505 -8200
rect 29881 -8204 29893 -8170
rect 30220 -8190 30230 -8070
rect 30350 -8100 30360 -8070
rect 31820 -8070 31960 -8060
rect 30350 -8164 31490 -8100
rect 30350 -8170 31493 -8164
rect 30350 -8190 30469 -8170
rect 30220 -8200 30469 -8190
rect 29493 -8210 29893 -8204
rect 30457 -8204 30469 -8200
rect 30845 -8200 31105 -8170
rect 30845 -8204 30857 -8200
rect 30457 -8210 30857 -8204
rect 31093 -8204 31105 -8200
rect 31481 -8204 31493 -8170
rect 31820 -8190 31830 -8070
rect 31950 -8100 31960 -8070
rect 34800 -8070 34940 -8060
rect 34800 -8100 34810 -8070
rect 31950 -8170 34810 -8100
rect 31950 -8190 32069 -8170
rect 31820 -8200 32069 -8190
rect 31093 -8210 31493 -8204
rect 32057 -8204 32069 -8200
rect 32445 -8200 32705 -8170
rect 32445 -8204 32457 -8200
rect 32057 -8210 32457 -8204
rect 32693 -8204 32705 -8200
rect 33081 -8200 33669 -8170
rect 33081 -8204 33093 -8200
rect 32693 -8210 33093 -8204
rect 33657 -8204 33669 -8200
rect 34045 -8200 34305 -8170
rect 34045 -8204 34057 -8200
rect 33657 -8210 34057 -8204
rect 34293 -8204 34305 -8200
rect 34681 -8190 34810 -8170
rect 34930 -8100 34940 -8070
rect 34930 -8164 36280 -8100
rect 34930 -8170 36293 -8164
rect 34930 -8190 35269 -8170
rect 34681 -8200 35269 -8190
rect 34681 -8204 34693 -8200
rect 34293 -8210 34693 -8204
rect 35257 -8204 35269 -8200
rect 35645 -8200 35905 -8170
rect 35645 -8204 35657 -8200
rect 35257 -8210 35657 -8204
rect 35893 -8204 35905 -8200
rect 36281 -8204 36293 -8170
rect 35893 -8210 36293 -8204
rect 36857 -8170 37257 -8164
rect 36857 -8204 36869 -8170
rect 37245 -8204 37257 -8170
rect 36857 -8210 37257 -8204
rect 37493 -8170 37893 -8164
rect 37493 -8204 37505 -8170
rect 37881 -8204 37893 -8170
rect 37493 -8210 37893 -8204
rect 11180 -8245 15570 -8240
rect 1134 -8257 1180 -8245
rect 1134 -8375 1140 -8257
rect 1174 -8375 1180 -8257
rect 1570 -8257 1616 -8245
rect 1570 -8260 1576 -8257
rect 1134 -8387 1180 -8375
rect 1560 -8375 1576 -8260
rect 1610 -8260 1616 -8257
rect 2098 -8257 2144 -8245
rect 2098 -8260 2104 -8257
rect 1610 -8375 2104 -8260
rect 2138 -8260 2144 -8257
rect 2206 -8257 2252 -8245
rect 2206 -8260 2212 -8257
rect 2138 -8375 2212 -8260
rect 2246 -8260 2252 -8257
rect 2734 -8257 2780 -8245
rect 2734 -8260 2740 -8257
rect 2246 -8375 2740 -8260
rect 2774 -8260 2780 -8257
rect 3170 -8257 3216 -8245
rect 3170 -8260 3176 -8257
rect 2774 -8375 3176 -8260
rect 3210 -8260 3216 -8257
rect 3698 -8257 3744 -8245
rect 3698 -8260 3704 -8257
rect 3210 -8375 3704 -8260
rect 3738 -8260 3744 -8257
rect 3806 -8257 3852 -8245
rect 3806 -8260 3812 -8257
rect 3738 -8375 3812 -8260
rect 3846 -8260 3852 -8257
rect 4334 -8257 4380 -8245
rect 4334 -8260 4340 -8257
rect 3846 -8375 4340 -8260
rect 4374 -8260 4380 -8257
rect 4770 -8257 4816 -8245
rect 4770 -8260 4776 -8257
rect 4374 -8375 4776 -8260
rect 4810 -8260 4816 -8257
rect 5298 -8257 5344 -8245
rect 5298 -8260 5304 -8257
rect 4810 -8375 5304 -8260
rect 5338 -8260 5344 -8257
rect 5406 -8257 5452 -8245
rect 5406 -8260 5412 -8257
rect 5338 -8375 5412 -8260
rect 5446 -8260 5452 -8257
rect 5934 -8257 5980 -8245
rect 5934 -8260 5940 -8257
rect 5446 -8375 5940 -8260
rect 5974 -8260 5980 -8257
rect 6370 -8257 6416 -8245
rect 6370 -8260 6376 -8257
rect 5974 -8375 6376 -8260
rect 6410 -8260 6416 -8257
rect 6898 -8257 6944 -8245
rect 6898 -8260 6904 -8257
rect 6410 -8375 6904 -8260
rect 6938 -8260 6944 -8257
rect 7006 -8257 7052 -8245
rect 7006 -8260 7012 -8257
rect 6938 -8375 7012 -8260
rect 7046 -8260 7052 -8257
rect 7534 -8257 7580 -8245
rect 7534 -8260 7540 -8257
rect 7046 -8375 7540 -8260
rect 7574 -8260 7580 -8257
rect 7970 -8257 8016 -8245
rect 7970 -8260 7976 -8257
rect 7574 -8375 7976 -8260
rect 8010 -8260 8016 -8257
rect 8498 -8257 8544 -8245
rect 8498 -8260 8504 -8257
rect 8010 -8375 8504 -8260
rect 8538 -8260 8544 -8257
rect 8606 -8257 8652 -8245
rect 8606 -8260 8612 -8257
rect 8538 -8375 8612 -8260
rect 8646 -8260 8652 -8257
rect 9134 -8257 9180 -8245
rect 9134 -8260 9140 -8257
rect 8646 -8375 9140 -8260
rect 9174 -8260 9180 -8257
rect 9570 -8257 9616 -8245
rect 9570 -8260 9576 -8257
rect 9174 -8375 9576 -8260
rect 9610 -8260 9616 -8257
rect 10098 -8257 10144 -8245
rect 10098 -8260 10104 -8257
rect 9610 -8375 10104 -8260
rect 10138 -8260 10144 -8257
rect 10206 -8257 10252 -8245
rect 10206 -8260 10212 -8257
rect 10138 -8375 10212 -8260
rect 10246 -8260 10252 -8257
rect 10734 -8250 10780 -8245
rect 10734 -8257 10940 -8250
rect 10734 -8260 10740 -8257
rect 10246 -8375 10740 -8260
rect 10774 -8260 10940 -8257
rect 10774 -8375 10810 -8260
rect 1560 -8380 10810 -8375
rect 10930 -8380 10940 -8260
rect 1570 -8387 1616 -8380
rect 2098 -8387 2144 -8380
rect 2206 -8387 2252 -8380
rect 2734 -8387 2780 -8380
rect 3170 -8387 3216 -8380
rect 3698 -8387 3744 -8380
rect 3806 -8387 3852 -8380
rect 4334 -8387 4380 -8380
rect 4770 -8387 4816 -8380
rect 5298 -8387 5344 -8380
rect 5406 -8387 5452 -8380
rect 5934 -8387 5980 -8380
rect 6370 -8387 6416 -8380
rect 6898 -8387 6944 -8380
rect 7006 -8387 7052 -8380
rect 7534 -8387 7580 -8380
rect 7970 -8387 8016 -8380
rect 8498 -8387 8544 -8380
rect 8606 -8387 8652 -8380
rect 9134 -8387 9180 -8380
rect 9570 -8387 9616 -8380
rect 10098 -8387 10144 -8380
rect 10206 -8387 10252 -8380
rect 10734 -8387 10940 -8380
rect 11170 -8257 15580 -8245
rect 11170 -8375 11176 -8257
rect 11210 -8375 11704 -8257
rect 11738 -8375 11812 -8257
rect 11846 -8375 12340 -8257
rect 12374 -8375 12776 -8257
rect 12810 -8375 13304 -8257
rect 13338 -8375 13412 -8257
rect 13446 -8375 13940 -8257
rect 13974 -8375 14376 -8257
rect 14410 -8375 14904 -8257
rect 14938 -8375 15012 -8257
rect 15046 -8375 15540 -8257
rect 15574 -8375 15580 -8257
rect 11170 -8387 15580 -8375
rect 15970 -8257 16016 -8245
rect 15970 -8375 15976 -8257
rect 16010 -8260 16016 -8257
rect 16498 -8250 16544 -8245
rect 16606 -8250 16652 -8245
rect 16498 -8257 16652 -8250
rect 16498 -8260 16504 -8257
rect 16538 -8260 16612 -8257
rect 16646 -8260 16652 -8257
rect 17134 -8257 17180 -8245
rect 17134 -8260 17140 -8257
rect 16010 -8375 16504 -8260
rect 16646 -8375 17140 -8260
rect 17174 -8260 17180 -8257
rect 17570 -8257 17616 -8245
rect 17570 -8260 17576 -8257
rect 17174 -8375 17576 -8260
rect 17610 -8260 17616 -8257
rect 18098 -8257 18144 -8245
rect 18098 -8260 18104 -8257
rect 17610 -8375 18104 -8260
rect 18138 -8260 18144 -8257
rect 18206 -8257 18252 -8245
rect 18206 -8260 18212 -8257
rect 18138 -8375 18212 -8260
rect 18246 -8260 18252 -8257
rect 18734 -8257 18780 -8245
rect 18734 -8260 18740 -8257
rect 18246 -8375 18740 -8260
rect 18774 -8260 18780 -8257
rect 19170 -8257 19216 -8245
rect 19170 -8260 19176 -8257
rect 18774 -8375 19176 -8260
rect 19210 -8260 19216 -8257
rect 19698 -8257 19744 -8245
rect 19698 -8260 19704 -8257
rect 19210 -8375 19704 -8260
rect 19738 -8260 19744 -8257
rect 19806 -8257 19852 -8245
rect 19806 -8260 19812 -8257
rect 19738 -8375 19812 -8260
rect 19846 -8260 19852 -8257
rect 20334 -8257 20380 -8245
rect 20334 -8260 20340 -8257
rect 19846 -8375 20340 -8260
rect 20374 -8260 20380 -8257
rect 20770 -8257 20816 -8245
rect 20770 -8260 20776 -8257
rect 20374 -8375 20776 -8260
rect 20810 -8260 20816 -8257
rect 21298 -8257 21344 -8245
rect 21298 -8260 21304 -8257
rect 20810 -8375 21304 -8260
rect 21338 -8260 21344 -8257
rect 21406 -8257 21452 -8245
rect 21406 -8260 21412 -8257
rect 21338 -8375 21412 -8260
rect 21446 -8260 21452 -8257
rect 21934 -8257 21980 -8245
rect 21934 -8260 21940 -8257
rect 21446 -8375 21940 -8260
rect 21974 -8260 21980 -8257
rect 22370 -8257 22416 -8245
rect 22370 -8260 22376 -8257
rect 21974 -8375 22376 -8260
rect 22410 -8260 22416 -8257
rect 22898 -8257 22944 -8245
rect 22898 -8260 22904 -8257
rect 22410 -8375 22904 -8260
rect 22938 -8260 22944 -8257
rect 23006 -8257 23052 -8245
rect 23006 -8260 23012 -8257
rect 22938 -8375 23012 -8260
rect 23046 -8260 23052 -8257
rect 23534 -8257 23580 -8245
rect 23534 -8260 23540 -8257
rect 23046 -8375 23540 -8260
rect 23574 -8260 23580 -8257
rect 23970 -8257 24016 -8245
rect 23970 -8260 23976 -8257
rect 23574 -8375 23976 -8260
rect 24010 -8260 24016 -8257
rect 24498 -8257 24544 -8245
rect 24498 -8260 24504 -8257
rect 24010 -8375 24504 -8260
rect 24538 -8260 24544 -8257
rect 24606 -8257 24652 -8245
rect 24606 -8260 24612 -8257
rect 24538 -8375 24612 -8260
rect 24646 -8260 24652 -8257
rect 25134 -8257 25180 -8245
rect 25134 -8260 25140 -8257
rect 24646 -8375 25140 -8260
rect 25174 -8260 25180 -8257
rect 25570 -8257 25616 -8245
rect 25570 -8260 25576 -8257
rect 25174 -8375 25576 -8260
rect 25610 -8260 25616 -8257
rect 26098 -8257 26144 -8245
rect 26098 -8260 26104 -8257
rect 25610 -8375 26104 -8260
rect 26138 -8260 26144 -8257
rect 26206 -8257 26252 -8245
rect 26206 -8260 26212 -8257
rect 26138 -8375 26212 -8260
rect 26246 -8260 26252 -8257
rect 26734 -8257 26780 -8245
rect 26734 -8260 26740 -8257
rect 26246 -8375 26740 -8260
rect 26774 -8260 26780 -8257
rect 27170 -8257 27216 -8245
rect 27170 -8260 27176 -8257
rect 26774 -8375 27176 -8260
rect 27210 -8260 27216 -8257
rect 27698 -8257 27744 -8245
rect 27698 -8260 27704 -8257
rect 27210 -8375 27704 -8260
rect 27738 -8260 27744 -8257
rect 27806 -8257 27852 -8245
rect 27806 -8260 27812 -8257
rect 27738 -8375 27812 -8260
rect 27846 -8260 27852 -8257
rect 28334 -8257 28380 -8245
rect 28334 -8260 28340 -8257
rect 27846 -8375 28340 -8260
rect 28374 -8260 28380 -8257
rect 28770 -8257 28816 -8245
rect 28770 -8260 28776 -8257
rect 28374 -8375 28776 -8260
rect 28810 -8260 28816 -8257
rect 29298 -8257 29344 -8245
rect 29298 -8260 29304 -8257
rect 28810 -8375 29304 -8260
rect 29338 -8260 29344 -8257
rect 29406 -8257 29452 -8245
rect 29406 -8260 29412 -8257
rect 29338 -8375 29412 -8260
rect 29446 -8260 29452 -8257
rect 29934 -8257 29980 -8245
rect 29934 -8260 29940 -8257
rect 29446 -8375 29940 -8260
rect 29974 -8260 29980 -8257
rect 30370 -8257 30416 -8237
rect 30370 -8260 30376 -8257
rect 29974 -8375 30376 -8260
rect 30410 -8260 30416 -8257
rect 30898 -8257 30944 -8237
rect 30898 -8260 30904 -8257
rect 30410 -8375 30904 -8260
rect 30938 -8260 30944 -8257
rect 31006 -8257 31052 -8237
rect 31006 -8260 31012 -8257
rect 30938 -8375 31012 -8260
rect 31046 -8260 31052 -8257
rect 31534 -8257 31580 -8245
rect 31534 -8260 31540 -8257
rect 31046 -8375 31540 -8260
rect 31574 -8260 31580 -8257
rect 31970 -8257 32016 -8245
rect 31970 -8260 31976 -8257
rect 31574 -8375 31976 -8260
rect 32010 -8260 32016 -8257
rect 32498 -8257 32544 -8245
rect 32498 -8260 32504 -8257
rect 32010 -8375 32504 -8260
rect 32538 -8260 32544 -8257
rect 32606 -8257 32652 -8245
rect 32606 -8260 32612 -8257
rect 32538 -8375 32612 -8260
rect 32646 -8260 32652 -8257
rect 33134 -8257 33180 -8245
rect 33134 -8260 33140 -8257
rect 32646 -8375 33140 -8260
rect 33174 -8260 33180 -8257
rect 33570 -8257 33616 -8245
rect 33570 -8260 33576 -8257
rect 33174 -8375 33576 -8260
rect 33610 -8260 33616 -8257
rect 34098 -8257 34144 -8245
rect 34098 -8260 34104 -8257
rect 33610 -8375 34104 -8260
rect 34138 -8260 34144 -8257
rect 34206 -8257 34252 -8245
rect 34206 -8260 34212 -8257
rect 34138 -8375 34212 -8260
rect 34246 -8260 34252 -8257
rect 34734 -8257 34780 -8245
rect 34734 -8260 34740 -8257
rect 34246 -8375 34740 -8260
rect 34774 -8260 34780 -8257
rect 35170 -8257 35216 -8245
rect 35170 -8260 35176 -8257
rect 34774 -8375 35176 -8260
rect 35210 -8260 35216 -8257
rect 35698 -8257 35744 -8245
rect 35698 -8260 35704 -8257
rect 35210 -8375 35704 -8260
rect 35738 -8260 35744 -8257
rect 35806 -8257 35852 -8245
rect 35806 -8260 35812 -8257
rect 35738 -8375 35812 -8260
rect 35846 -8260 35852 -8257
rect 36334 -8257 36380 -8245
rect 36334 -8260 36340 -8257
rect 35846 -8375 36340 -8260
rect 36374 -8375 36380 -8257
rect 15970 -8380 16510 -8375
rect 16640 -8380 36380 -8375
rect 15970 -8387 16016 -8380
rect 16498 -8387 16652 -8380
rect 17134 -8387 17180 -8380
rect 17570 -8387 17616 -8380
rect 18098 -8387 18144 -8380
rect 18206 -8387 18252 -8380
rect 18734 -8387 18780 -8380
rect 19170 -8387 19216 -8380
rect 19698 -8387 19744 -8380
rect 19806 -8387 19852 -8380
rect 20334 -8387 20380 -8380
rect 20770 -8387 20816 -8380
rect 21298 -8387 21344 -8380
rect 21406 -8387 21452 -8380
rect 21934 -8387 21980 -8380
rect 22370 -8387 22416 -8380
rect 22898 -8387 22944 -8380
rect 23006 -8387 23052 -8380
rect 23534 -8387 23580 -8380
rect 23970 -8387 24016 -8380
rect 24498 -8387 24544 -8380
rect 24606 -8387 24652 -8380
rect 25134 -8387 25180 -8380
rect 25570 -8387 25616 -8380
rect 26098 -8387 26144 -8380
rect 26206 -8387 26252 -8380
rect 26734 -8387 26780 -8380
rect 27170 -8387 27216 -8380
rect 27698 -8387 27744 -8380
rect 27806 -8387 27852 -8380
rect 28334 -8387 28380 -8380
rect 28770 -8387 28816 -8380
rect 29298 -8387 29344 -8380
rect 29406 -8387 29452 -8380
rect 29934 -8387 29980 -8380
rect 10750 -8390 10940 -8387
rect 11180 -8390 15570 -8387
rect 16500 -8390 16650 -8387
rect 30370 -8395 30416 -8380
rect 30898 -8395 30944 -8380
rect 31006 -8395 31052 -8380
rect 31534 -8387 31580 -8380
rect 31970 -8387 32016 -8380
rect 32498 -8387 32544 -8380
rect 32606 -8387 32652 -8380
rect 33134 -8387 33180 -8380
rect 33570 -8387 33616 -8380
rect 34098 -8387 34144 -8380
rect 34206 -8387 34252 -8380
rect 34734 -8387 34780 -8380
rect 35170 -8387 35216 -8380
rect 35698 -8387 35744 -8380
rect 35806 -8387 35852 -8380
rect 36334 -8387 36380 -8380
rect 36770 -8257 36816 -8245
rect 36770 -8375 36776 -8257
rect 36810 -8375 36816 -8257
rect 36770 -8387 36816 -8375
rect 37298 -8257 37344 -8245
rect 37298 -8375 37304 -8257
rect 37338 -8375 37344 -8257
rect 37298 -8387 37344 -8375
rect 37406 -8257 37452 -8245
rect 37406 -8375 37412 -8257
rect 37446 -8375 37452 -8257
rect 37406 -8387 37452 -8375
rect 37934 -8257 37980 -8245
rect 37934 -8375 37940 -8257
rect 37974 -8375 37980 -8257
rect 37934 -8387 37980 -8375
rect 670 -8428 1093 -8422
rect 670 -8462 705 -8428
rect 1081 -8462 1093 -8428
rect 670 -8468 1093 -8462
rect 1657 -8428 2057 -8422
rect 1657 -8462 1669 -8428
rect 2045 -8430 2057 -8428
rect 2293 -8428 2693 -8422
rect 2293 -8430 2305 -8428
rect 2045 -8462 2060 -8430
rect 1657 -8468 2060 -8462
rect 670 -8690 720 -8468
rect 1420 -8510 1560 -8500
rect 1420 -8630 1430 -8510
rect 1550 -8520 1560 -8510
rect 1660 -8520 2060 -8468
rect 2290 -8462 2305 -8430
rect 2681 -8462 2693 -8428
rect 2290 -8468 2693 -8462
rect 3257 -8428 3657 -8422
rect 3257 -8462 3269 -8428
rect 3645 -8430 3657 -8428
rect 3893 -8428 4293 -8422
rect 3893 -8430 3905 -8428
rect 3645 -8462 3660 -8430
rect 3257 -8468 3660 -8462
rect 2290 -8520 2690 -8468
rect 3020 -8510 3160 -8500
rect 3020 -8520 3030 -8510
rect 1550 -8620 3030 -8520
rect 1550 -8630 1560 -8620
rect 1420 -8640 1560 -8630
rect 1660 -8640 2690 -8620
rect 3020 -8630 3030 -8620
rect 3150 -8520 3160 -8510
rect 3260 -8520 3660 -8468
rect 3890 -8462 3905 -8430
rect 4281 -8462 4293 -8428
rect 3890 -8468 4293 -8462
rect 4857 -8428 5257 -8422
rect 4857 -8462 4869 -8428
rect 5245 -8430 5257 -8428
rect 5493 -8428 5893 -8422
rect 5493 -8430 5505 -8428
rect 5245 -8462 5260 -8430
rect 4857 -8468 5260 -8462
rect 3890 -8520 4290 -8468
rect 4620 -8510 4760 -8500
rect 4620 -8520 4630 -8510
rect 3150 -8620 4630 -8520
rect 3150 -8630 3160 -8620
rect 3020 -8640 3160 -8630
rect 3260 -8640 4290 -8620
rect 4620 -8630 4630 -8620
rect 4750 -8520 4760 -8510
rect 4860 -8520 5260 -8468
rect 5490 -8462 5505 -8430
rect 5881 -8462 5893 -8428
rect 5490 -8468 5893 -8462
rect 6457 -8428 6857 -8422
rect 6457 -8462 6469 -8428
rect 6845 -8430 6857 -8428
rect 7093 -8428 7493 -8422
rect 7093 -8430 7105 -8428
rect 6845 -8462 6860 -8430
rect 6457 -8468 6860 -8462
rect 5490 -8520 5890 -8468
rect 6220 -8510 6360 -8500
rect 6220 -8520 6230 -8510
rect 4750 -8620 6230 -8520
rect 4750 -8630 4760 -8620
rect 4620 -8640 4760 -8630
rect 4860 -8640 5890 -8620
rect 6220 -8630 6230 -8620
rect 6350 -8520 6360 -8510
rect 6460 -8520 6860 -8468
rect 7090 -8462 7105 -8430
rect 7481 -8462 7493 -8428
rect 7090 -8468 7493 -8462
rect 8057 -8428 8457 -8422
rect 8057 -8462 8069 -8428
rect 8445 -8430 8457 -8428
rect 8693 -8428 9093 -8422
rect 8693 -8430 8705 -8428
rect 8445 -8462 8460 -8430
rect 8057 -8468 8460 -8462
rect 7090 -8520 7490 -8468
rect 7820 -8510 7960 -8500
rect 7820 -8520 7830 -8510
rect 6350 -8620 7830 -8520
rect 6350 -8630 6360 -8620
rect 6220 -8640 6360 -8630
rect 6460 -8640 7490 -8620
rect 7820 -8630 7830 -8620
rect 7950 -8520 7960 -8510
rect 8060 -8520 8460 -8468
rect 8690 -8462 8705 -8430
rect 9081 -8462 9093 -8428
rect 8690 -8468 9093 -8462
rect 9657 -8428 10057 -8422
rect 9657 -8462 9669 -8428
rect 10045 -8430 10057 -8428
rect 10293 -8428 10693 -8422
rect 10293 -8430 10305 -8428
rect 10045 -8462 10060 -8430
rect 9657 -8468 10060 -8462
rect 8690 -8520 9090 -8468
rect 9420 -8510 9560 -8500
rect 9420 -8520 9430 -8510
rect 7950 -8620 9430 -8520
rect 7950 -8630 7960 -8620
rect 7820 -8640 7960 -8630
rect 8060 -8640 9090 -8620
rect 9420 -8630 9430 -8620
rect 9550 -8520 9560 -8510
rect 9660 -8520 10060 -8468
rect 10290 -8462 10305 -8430
rect 10681 -8462 10693 -8428
rect 10290 -8468 10693 -8462
rect 11257 -8428 11657 -8422
rect 11257 -8462 11269 -8428
rect 11645 -8430 11657 -8428
rect 11893 -8428 12293 -8422
rect 11893 -8430 11905 -8428
rect 11645 -8462 11905 -8430
rect 12281 -8430 12293 -8428
rect 12857 -8428 13257 -8422
rect 12857 -8430 12869 -8428
rect 12281 -8462 12869 -8430
rect 13245 -8430 13257 -8428
rect 13493 -8428 13893 -8422
rect 13493 -8430 13505 -8428
rect 13245 -8462 13505 -8430
rect 13881 -8430 13893 -8428
rect 14457 -8428 14857 -8422
rect 14457 -8430 14469 -8428
rect 13881 -8462 14469 -8430
rect 14845 -8430 14857 -8428
rect 15093 -8428 15493 -8422
rect 15093 -8430 15105 -8428
rect 14845 -8462 15105 -8430
rect 15481 -8462 15493 -8428
rect 11257 -8468 15493 -8462
rect 16057 -8428 16457 -8422
rect 16057 -8462 16069 -8428
rect 16445 -8462 16457 -8428
rect 16057 -8468 16457 -8462
rect 16693 -8428 17093 -8422
rect 16693 -8462 16705 -8428
rect 17081 -8462 17093 -8428
rect 16693 -8468 17093 -8462
rect 17657 -8428 18057 -8422
rect 17657 -8462 17669 -8428
rect 18045 -8462 18057 -8428
rect 17657 -8468 18057 -8462
rect 18293 -8428 18693 -8422
rect 18293 -8462 18305 -8428
rect 18681 -8462 18693 -8428
rect 18293 -8468 18693 -8462
rect 19257 -8428 19657 -8422
rect 19257 -8462 19269 -8428
rect 19645 -8462 19657 -8428
rect 19257 -8468 19657 -8462
rect 19893 -8428 20293 -8422
rect 19893 -8462 19905 -8428
rect 20281 -8462 20293 -8428
rect 19893 -8468 20293 -8462
rect 20857 -8428 21257 -8422
rect 20857 -8462 20869 -8428
rect 21245 -8462 21257 -8428
rect 20857 -8468 21257 -8462
rect 21493 -8428 21893 -8422
rect 21493 -8462 21505 -8428
rect 21881 -8462 21893 -8428
rect 21493 -8468 21893 -8462
rect 22457 -8428 22857 -8422
rect 22457 -8462 22469 -8428
rect 22845 -8462 22857 -8428
rect 22457 -8468 22857 -8462
rect 23093 -8428 23493 -8422
rect 23093 -8462 23105 -8428
rect 23481 -8462 23493 -8428
rect 23093 -8468 23493 -8462
rect 24057 -8428 24457 -8422
rect 24057 -8462 24069 -8428
rect 24445 -8462 24457 -8428
rect 24057 -8468 24457 -8462
rect 24693 -8428 25093 -8422
rect 24693 -8462 24705 -8428
rect 25081 -8462 25093 -8428
rect 24693 -8468 25093 -8462
rect 25657 -8428 26057 -8422
rect 25657 -8462 25669 -8428
rect 26045 -8462 26057 -8428
rect 25657 -8468 26057 -8462
rect 26293 -8428 26693 -8422
rect 26293 -8462 26305 -8428
rect 26681 -8462 26693 -8428
rect 26293 -8468 26693 -8462
rect 27257 -8428 27657 -8422
rect 27257 -8462 27269 -8428
rect 27645 -8462 27657 -8428
rect 27257 -8468 27657 -8462
rect 27893 -8428 28293 -8422
rect 27893 -8462 27905 -8428
rect 28281 -8462 28293 -8428
rect 27893 -8468 28293 -8462
rect 28857 -8428 29257 -8422
rect 28857 -8462 28869 -8428
rect 29245 -8462 29257 -8428
rect 28857 -8468 29257 -8462
rect 29493 -8428 29893 -8422
rect 29493 -8462 29505 -8428
rect 29881 -8462 29893 -8428
rect 29493 -8468 29893 -8462
rect 30457 -8428 30857 -8422
rect 30457 -8462 30469 -8428
rect 30845 -8462 30857 -8428
rect 30457 -8468 30857 -8462
rect 31093 -8428 31493 -8422
rect 31093 -8462 31105 -8428
rect 31481 -8462 31493 -8428
rect 31093 -8468 31493 -8462
rect 32057 -8428 32457 -8422
rect 32057 -8462 32069 -8428
rect 32445 -8462 32457 -8428
rect 32057 -8468 32457 -8462
rect 32693 -8428 33093 -8422
rect 32693 -8462 32705 -8428
rect 33081 -8462 33093 -8428
rect 32693 -8468 33093 -8462
rect 33657 -8428 34057 -8422
rect 33657 -8462 33669 -8428
rect 34045 -8462 34057 -8428
rect 33657 -8468 34057 -8462
rect 34293 -8428 34693 -8422
rect 34293 -8462 34305 -8428
rect 34681 -8462 34693 -8428
rect 34293 -8468 34693 -8462
rect 35257 -8428 35657 -8422
rect 35257 -8462 35269 -8428
rect 35645 -8462 35657 -8428
rect 35257 -8468 35657 -8462
rect 35893 -8428 36293 -8422
rect 35893 -8462 35905 -8428
rect 36281 -8462 36293 -8428
rect 35893 -8468 36293 -8462
rect 36857 -8428 37257 -8422
rect 36857 -8462 36869 -8428
rect 37245 -8462 37257 -8428
rect 36857 -8468 37257 -8462
rect 37493 -8428 37893 -8422
rect 37493 -8462 37505 -8428
rect 37881 -8462 37893 -8428
rect 37493 -8468 37893 -8462
rect 10290 -8520 10690 -8468
rect 11260 -8490 15490 -8468
rect 9550 -8620 10690 -8520
rect 9550 -8630 9560 -8620
rect 9420 -8640 9560 -8630
rect 9660 -8640 10690 -8620
rect 1660 -8690 2060 -8640
rect 670 -8696 1093 -8690
rect 670 -8730 705 -8696
rect 1081 -8730 1093 -8696
rect 670 -8736 1093 -8730
rect 1657 -8696 2060 -8690
rect 1657 -8730 1669 -8696
rect 2045 -8730 2060 -8696
rect 2290 -8690 2690 -8640
rect 3260 -8690 3660 -8640
rect 2290 -8696 2693 -8690
rect 2290 -8730 2305 -8696
rect 2681 -8730 2693 -8696
rect 1657 -8736 2057 -8730
rect 2293 -8736 2693 -8730
rect 3257 -8696 3660 -8690
rect 3257 -8730 3269 -8696
rect 3645 -8730 3660 -8696
rect 3890 -8690 4290 -8640
rect 4860 -8690 5260 -8640
rect 3890 -8696 4293 -8690
rect 3890 -8730 3905 -8696
rect 4281 -8730 4293 -8696
rect 3257 -8736 3657 -8730
rect 3893 -8736 4293 -8730
rect 4857 -8696 5260 -8690
rect 4857 -8730 4869 -8696
rect 5245 -8730 5260 -8696
rect 5490 -8690 5890 -8640
rect 6460 -8690 6860 -8640
rect 5490 -8696 5893 -8690
rect 5490 -8730 5505 -8696
rect 5881 -8730 5893 -8696
rect 4857 -8736 5257 -8730
rect 5493 -8736 5893 -8730
rect 6457 -8696 6860 -8690
rect 6457 -8730 6469 -8696
rect 6845 -8730 6860 -8696
rect 7090 -8690 7490 -8640
rect 8060 -8690 8460 -8640
rect 7090 -8696 7493 -8690
rect 7090 -8730 7105 -8696
rect 7481 -8730 7493 -8696
rect 6457 -8736 6857 -8730
rect 7093 -8736 7493 -8730
rect 8057 -8696 8460 -8690
rect 8057 -8730 8069 -8696
rect 8445 -8730 8460 -8696
rect 8690 -8690 9090 -8640
rect 9660 -8690 10060 -8640
rect 8690 -8696 9093 -8690
rect 8690 -8730 8705 -8696
rect 9081 -8730 9093 -8696
rect 8057 -8736 8457 -8730
rect 8693 -8736 9093 -8730
rect 9657 -8696 10060 -8690
rect 9657 -8730 9669 -8696
rect 10045 -8730 10060 -8696
rect 10290 -8690 10690 -8640
rect 11420 -8650 11480 -8490
rect 12070 -8650 12130 -8490
rect 11260 -8690 12290 -8650
rect 10290 -8696 10693 -8690
rect 10290 -8730 10305 -8696
rect 10681 -8730 10693 -8696
rect 9657 -8736 10057 -8730
rect 10293 -8736 10693 -8730
rect 11257 -8696 12293 -8690
rect 11257 -8730 11269 -8696
rect 11645 -8730 11905 -8696
rect 12281 -8730 12293 -8696
rect 11257 -8736 11657 -8730
rect 11893 -8736 12293 -8730
rect 57 -9554 490 -9548
rect 57 -9580 69 -9554
rect 0 -9588 69 -9580
rect 445 -9588 490 -9554
rect 0 -9688 490 -9588
rect 670 -9548 720 -8736
rect 1134 -8796 1180 -8784
rect 1134 -9488 1140 -8796
rect 1174 -9488 1180 -8796
rect 1134 -9500 1180 -9488
rect 1570 -8796 1616 -8784
rect 1570 -9488 1576 -8796
rect 1610 -9488 1616 -8796
rect 1570 -9500 1616 -9488
rect 2098 -8796 2144 -8784
rect 2098 -9488 2104 -8796
rect 2138 -8800 2144 -8796
rect 2206 -8796 2252 -8784
rect 2206 -8800 2212 -8796
rect 2138 -8810 2212 -8800
rect 2138 -9480 2212 -9470
rect 2138 -9488 2144 -9480
rect 2098 -9500 2144 -9488
rect 2206 -9488 2212 -9480
rect 2246 -9488 2252 -8796
rect 2206 -9500 2252 -9488
rect 2734 -8796 2780 -8784
rect 2734 -9488 2740 -8796
rect 2774 -9488 2780 -8796
rect 2734 -9500 2780 -9488
rect 3170 -8796 3216 -8784
rect 3170 -9488 3176 -8796
rect 3210 -9488 3216 -8796
rect 3170 -9500 3216 -9488
rect 3698 -8796 3744 -8784
rect 3698 -9488 3704 -8796
rect 3738 -8800 3744 -8796
rect 3806 -8796 3852 -8784
rect 3806 -8800 3812 -8796
rect 3738 -8810 3812 -8800
rect 3738 -9480 3812 -9470
rect 3738 -9488 3744 -9480
rect 3698 -9500 3744 -9488
rect 3806 -9488 3812 -9480
rect 3846 -9488 3852 -8796
rect 3806 -9500 3852 -9488
rect 4334 -8796 4380 -8784
rect 4334 -9488 4340 -8796
rect 4374 -9488 4380 -8796
rect 4334 -9500 4380 -9488
rect 4770 -8796 4816 -8784
rect 4770 -9488 4776 -8796
rect 4810 -9488 4816 -8796
rect 4770 -9500 4816 -9488
rect 5298 -8796 5344 -8784
rect 5298 -9488 5304 -8796
rect 5338 -8800 5344 -8796
rect 5406 -8796 5452 -8784
rect 5406 -8800 5412 -8796
rect 5338 -8810 5412 -8800
rect 5338 -9480 5412 -9470
rect 5338 -9488 5344 -9480
rect 5298 -9500 5344 -9488
rect 5406 -9488 5412 -9480
rect 5446 -9488 5452 -8796
rect 5406 -9500 5452 -9488
rect 5934 -8796 5980 -8784
rect 5934 -9488 5940 -8796
rect 5974 -9488 5980 -8796
rect 5934 -9500 5980 -9488
rect 6370 -8796 6416 -8784
rect 6370 -9488 6376 -8796
rect 6410 -9488 6416 -8796
rect 6370 -9500 6416 -9488
rect 6898 -8796 6944 -8784
rect 6898 -9488 6904 -8796
rect 6938 -8800 6944 -8796
rect 7006 -8796 7052 -8784
rect 7006 -8800 7012 -8796
rect 6938 -8810 7012 -8800
rect 6938 -9480 7012 -9470
rect 6938 -9488 6944 -9480
rect 6898 -9500 6944 -9488
rect 7006 -9488 7012 -9480
rect 7046 -9488 7052 -8796
rect 7006 -9500 7052 -9488
rect 7534 -8796 7580 -8784
rect 7534 -9488 7540 -8796
rect 7574 -9488 7580 -8796
rect 7534 -9500 7580 -9488
rect 7970 -8796 8016 -8784
rect 7970 -9488 7976 -8796
rect 8010 -9488 8016 -8796
rect 7970 -9500 8016 -9488
rect 8498 -8796 8544 -8784
rect 8498 -9488 8504 -8796
rect 8538 -8800 8544 -8796
rect 8606 -8796 8652 -8784
rect 8606 -8800 8612 -8796
rect 8538 -8810 8612 -8800
rect 8538 -9480 8612 -9470
rect 8538 -9488 8544 -9480
rect 8498 -9500 8544 -9488
rect 8606 -9488 8612 -9480
rect 8646 -9488 8652 -8796
rect 8606 -9500 8652 -9488
rect 9134 -8796 9180 -8784
rect 9134 -9488 9140 -8796
rect 9174 -9488 9180 -8796
rect 9134 -9500 9180 -9488
rect 9570 -8796 9616 -8784
rect 9570 -9488 9576 -8796
rect 9610 -9488 9616 -8796
rect 9570 -9500 9616 -9488
rect 10098 -8796 10144 -8784
rect 10098 -9488 10104 -8796
rect 10138 -8800 10144 -8796
rect 10206 -8796 10252 -8784
rect 10206 -8800 10212 -8796
rect 10138 -8810 10212 -8800
rect 10138 -9480 10212 -9470
rect 10138 -9488 10144 -9480
rect 10098 -9500 10144 -9488
rect 10206 -9488 10212 -9480
rect 10246 -9488 10252 -8796
rect 10206 -9500 10252 -9488
rect 10734 -8796 10780 -8784
rect 10734 -9488 10740 -8796
rect 10774 -9488 10780 -8796
rect 10734 -9500 10780 -9488
rect 11170 -8796 11216 -8784
rect 11170 -9488 11176 -8796
rect 11210 -9488 11216 -8796
rect 11170 -9500 11216 -9488
rect 11698 -8796 11744 -8784
rect 11698 -9488 11704 -8796
rect 11738 -8800 11744 -8796
rect 11806 -8796 11852 -8784
rect 11806 -8800 11812 -8796
rect 11738 -8810 11812 -8800
rect 11738 -9480 11812 -9470
rect 11738 -9488 11744 -9480
rect 11698 -9500 11744 -9488
rect 11806 -9488 11812 -9480
rect 11846 -9488 11852 -8796
rect 11806 -9500 11852 -9488
rect 12334 -8796 12380 -8784
rect 12334 -9488 12340 -8796
rect 12374 -9488 12380 -8796
rect 12334 -9500 12380 -9488
rect 670 -9554 1093 -9548
rect 670 -9588 705 -9554
rect 1081 -9580 1093 -9554
rect 1657 -9554 2057 -9548
rect 1657 -9580 1669 -9554
rect 1081 -9588 1669 -9580
rect 2045 -9580 2057 -9554
rect 2293 -9554 2693 -9548
rect 2293 -9580 2305 -9554
rect 2045 -9588 2305 -9580
rect 2681 -9580 2693 -9554
rect 3257 -9554 3657 -9548
rect 3257 -9580 3269 -9554
rect 2681 -9588 3269 -9580
rect 3645 -9580 3657 -9554
rect 3893 -9554 4293 -9548
rect 3893 -9580 3905 -9554
rect 3645 -9588 3905 -9580
rect 4281 -9580 4293 -9554
rect 4857 -9554 5257 -9548
rect 4857 -9580 4869 -9554
rect 4281 -9588 4869 -9580
rect 5245 -9580 5257 -9554
rect 5493 -9554 5893 -9548
rect 5493 -9580 5505 -9554
rect 5245 -9588 5505 -9580
rect 5881 -9580 5893 -9554
rect 6457 -9554 6857 -9548
rect 6457 -9580 6469 -9554
rect 5881 -9588 6469 -9580
rect 6845 -9580 6857 -9554
rect 7093 -9554 7493 -9548
rect 7093 -9580 7105 -9554
rect 6845 -9588 7105 -9580
rect 7481 -9580 7493 -9554
rect 8057 -9554 8457 -9548
rect 8057 -9580 8069 -9554
rect 7481 -9588 8069 -9580
rect 8445 -9580 8457 -9554
rect 8693 -9554 9093 -9548
rect 8693 -9580 8705 -9554
rect 8445 -9588 8705 -9580
rect 9081 -9580 9093 -9554
rect 9657 -9554 10057 -9548
rect 9657 -9580 9669 -9554
rect 9081 -9588 9669 -9580
rect 10045 -9580 10057 -9554
rect 10293 -9554 10693 -9548
rect 10293 -9580 10305 -9554
rect 10045 -9588 10305 -9580
rect 10681 -9580 10693 -9554
rect 11257 -9554 11657 -9548
rect 11257 -9580 11269 -9554
rect 10681 -9588 11269 -9580
rect 11645 -9580 11657 -9554
rect 11893 -9554 12293 -9548
rect 11893 -9580 11905 -9554
rect 11645 -9588 11905 -9580
rect 12281 -9580 12293 -9554
rect 12480 -9550 12680 -8490
rect 15600 -8520 15740 -8510
rect 12860 -8690 15490 -8630
rect 15600 -8640 15610 -8520
rect 15730 -8530 15740 -8520
rect 16060 -8530 16450 -8468
rect 16700 -8530 17090 -8468
rect 15730 -8630 17090 -8530
rect 15730 -8640 15740 -8630
rect 15600 -8650 15740 -8640
rect 16060 -8690 16450 -8630
rect 16700 -8690 17090 -8630
rect 17200 -8520 17340 -8510
rect 17200 -8640 17210 -8520
rect 17330 -8530 17340 -8520
rect 17660 -8530 18050 -8468
rect 18300 -8530 18690 -8468
rect 17330 -8630 18690 -8530
rect 17330 -8640 17340 -8630
rect 17200 -8650 17340 -8640
rect 17660 -8690 18050 -8630
rect 18300 -8690 18690 -8630
rect 18800 -8520 18940 -8510
rect 18800 -8640 18810 -8520
rect 18930 -8530 18940 -8520
rect 19260 -8530 19650 -8468
rect 19900 -8530 20290 -8468
rect 18930 -8630 20290 -8530
rect 18930 -8640 18940 -8630
rect 18800 -8650 18940 -8640
rect 19260 -8690 19650 -8630
rect 19900 -8690 20290 -8630
rect 20400 -8520 20540 -8510
rect 20400 -8640 20410 -8520
rect 20530 -8530 20540 -8520
rect 20860 -8530 21250 -8468
rect 21500 -8530 21890 -8468
rect 20530 -8630 21890 -8530
rect 20530 -8640 20540 -8630
rect 20400 -8650 20540 -8640
rect 20860 -8690 21250 -8630
rect 21500 -8690 21890 -8630
rect 22000 -8520 22140 -8510
rect 22000 -8640 22010 -8520
rect 22130 -8530 22140 -8520
rect 22460 -8530 22850 -8468
rect 23100 -8530 23490 -8468
rect 22130 -8630 23490 -8530
rect 22130 -8640 22140 -8630
rect 22000 -8650 22140 -8640
rect 22460 -8690 22850 -8630
rect 23100 -8690 23490 -8630
rect 23600 -8520 23740 -8510
rect 23600 -8640 23610 -8520
rect 23730 -8530 23740 -8520
rect 24060 -8530 24450 -8468
rect 24700 -8530 25090 -8468
rect 23730 -8630 25090 -8530
rect 23730 -8640 23740 -8630
rect 23600 -8650 23740 -8640
rect 24060 -8690 24450 -8630
rect 24700 -8690 25090 -8630
rect 25200 -8520 25340 -8510
rect 25200 -8640 25210 -8520
rect 25330 -8530 25340 -8520
rect 25660 -8530 26050 -8468
rect 26300 -8530 26690 -8468
rect 25330 -8630 26690 -8530
rect 25330 -8640 25340 -8630
rect 25200 -8650 25340 -8640
rect 25660 -8690 26050 -8630
rect 26300 -8690 26690 -8630
rect 26800 -8520 26940 -8510
rect 26800 -8640 26810 -8520
rect 26930 -8530 26940 -8520
rect 27260 -8530 27650 -8468
rect 27900 -8530 28290 -8468
rect 26930 -8630 28290 -8530
rect 26930 -8640 26940 -8630
rect 26800 -8650 26940 -8640
rect 27260 -8690 27650 -8630
rect 27900 -8690 28290 -8630
rect 28400 -8520 28540 -8510
rect 28400 -8640 28410 -8520
rect 28530 -8530 28540 -8520
rect 28860 -8530 29250 -8468
rect 29500 -8530 29890 -8468
rect 28530 -8630 29890 -8530
rect 28530 -8640 28540 -8630
rect 28400 -8650 28540 -8640
rect 28860 -8690 29250 -8630
rect 29500 -8690 29890 -8630
rect 30000 -8520 30140 -8510
rect 30000 -8640 30010 -8520
rect 30130 -8530 30140 -8520
rect 30460 -8530 30850 -8468
rect 31100 -8530 31490 -8468
rect 30130 -8630 31490 -8530
rect 30130 -8640 30140 -8630
rect 30000 -8650 30140 -8640
rect 30460 -8690 30850 -8630
rect 31100 -8690 31490 -8630
rect 32060 -8530 32450 -8468
rect 32700 -8530 33090 -8468
rect 33660 -8530 34050 -8468
rect 34300 -8530 34690 -8468
rect 35260 -8530 35650 -8468
rect 35900 -8530 36290 -8468
rect 32060 -8630 36290 -8530
rect 32060 -8690 32450 -8630
rect 32700 -8690 33090 -8630
rect 33660 -8690 34050 -8630
rect 34300 -8690 34690 -8630
rect 35260 -8690 35650 -8630
rect 35900 -8690 36290 -8630
rect 12857 -8696 15493 -8690
rect 12857 -8730 12869 -8696
rect 13245 -8730 13505 -8696
rect 13881 -8730 14469 -8696
rect 14845 -8730 15105 -8696
rect 15481 -8730 15493 -8696
rect 12857 -8736 13257 -8730
rect 13310 -8784 13440 -8730
rect 13493 -8736 13893 -8730
rect 14457 -8736 14857 -8730
rect 14910 -8784 15040 -8730
rect 15093 -8736 15493 -8730
rect 16057 -8696 16457 -8690
rect 16057 -8730 16069 -8696
rect 16445 -8730 16457 -8696
rect 16057 -8736 16457 -8730
rect 16693 -8696 17093 -8690
rect 16693 -8730 16705 -8696
rect 17081 -8730 17093 -8696
rect 16693 -8736 17093 -8730
rect 17657 -8696 18057 -8690
rect 17657 -8730 17669 -8696
rect 18045 -8730 18057 -8696
rect 17657 -8736 18057 -8730
rect 18293 -8696 18693 -8690
rect 18293 -8730 18305 -8696
rect 18681 -8730 18693 -8696
rect 18293 -8736 18693 -8730
rect 19257 -8696 19657 -8690
rect 19257 -8730 19269 -8696
rect 19645 -8730 19657 -8696
rect 19257 -8736 19657 -8730
rect 19893 -8696 20293 -8690
rect 19893 -8730 19905 -8696
rect 20281 -8730 20293 -8696
rect 19893 -8736 20293 -8730
rect 20857 -8696 21257 -8690
rect 20857 -8730 20869 -8696
rect 21245 -8730 21257 -8696
rect 20857 -8736 21257 -8730
rect 21493 -8696 21893 -8690
rect 21493 -8730 21505 -8696
rect 21881 -8730 21893 -8696
rect 21493 -8736 21893 -8730
rect 22457 -8696 22857 -8690
rect 22457 -8730 22469 -8696
rect 22845 -8730 22857 -8696
rect 22457 -8736 22857 -8730
rect 23093 -8696 23493 -8690
rect 23093 -8730 23105 -8696
rect 23481 -8730 23493 -8696
rect 23093 -8736 23493 -8730
rect 24057 -8696 24457 -8690
rect 24057 -8730 24069 -8696
rect 24445 -8730 24457 -8696
rect 24057 -8736 24457 -8730
rect 24693 -8696 25093 -8690
rect 24693 -8730 24705 -8696
rect 25081 -8730 25093 -8696
rect 24693 -8736 25093 -8730
rect 25657 -8696 26057 -8690
rect 25657 -8730 25669 -8696
rect 26045 -8730 26057 -8696
rect 25657 -8736 26057 -8730
rect 26293 -8696 26693 -8690
rect 26293 -8730 26305 -8696
rect 26681 -8730 26693 -8696
rect 26293 -8736 26693 -8730
rect 27257 -8696 27657 -8690
rect 27257 -8730 27269 -8696
rect 27645 -8730 27657 -8696
rect 27257 -8736 27657 -8730
rect 27893 -8696 28293 -8690
rect 27893 -8730 27905 -8696
rect 28281 -8730 28293 -8696
rect 27893 -8736 28293 -8730
rect 28857 -8696 29257 -8690
rect 28857 -8730 28869 -8696
rect 29245 -8730 29257 -8696
rect 28857 -8736 29257 -8730
rect 29493 -8696 29893 -8690
rect 29493 -8730 29505 -8696
rect 29881 -8730 29893 -8696
rect 29493 -8736 29893 -8730
rect 30457 -8696 30857 -8690
rect 30457 -8730 30469 -8696
rect 30845 -8730 30857 -8696
rect 30457 -8736 30857 -8730
rect 31093 -8696 31493 -8690
rect 31093 -8730 31105 -8696
rect 31481 -8730 31493 -8696
rect 31093 -8736 31493 -8730
rect 32057 -8696 32457 -8690
rect 32057 -8730 32069 -8696
rect 32445 -8730 32457 -8696
rect 32057 -8736 32457 -8730
rect 32693 -8696 33093 -8690
rect 32693 -8730 32705 -8696
rect 33081 -8730 33093 -8696
rect 32693 -8736 33093 -8730
rect 33657 -8696 34057 -8690
rect 33657 -8730 33669 -8696
rect 34045 -8730 34057 -8696
rect 33657 -8736 34057 -8730
rect 34293 -8696 34693 -8690
rect 34293 -8730 34305 -8696
rect 34681 -8730 34693 -8696
rect 34293 -8736 34693 -8730
rect 35257 -8696 35657 -8690
rect 35257 -8730 35269 -8696
rect 35645 -8730 35657 -8696
rect 35257 -8736 35657 -8730
rect 35893 -8696 36293 -8690
rect 35893 -8730 35905 -8696
rect 36281 -8730 36293 -8696
rect 35893 -8736 36293 -8730
rect 36857 -8696 37257 -8690
rect 36857 -8730 36869 -8696
rect 37245 -8730 37257 -8696
rect 36857 -8736 37257 -8730
rect 37493 -8696 37893 -8690
rect 37493 -8730 37505 -8696
rect 37881 -8730 37893 -8696
rect 37493 -8736 37893 -8730
rect 12770 -8796 12816 -8784
rect 12770 -9488 12776 -8796
rect 12810 -9488 12816 -8796
rect 12770 -9500 12816 -9488
rect 13298 -8796 13452 -8784
rect 13298 -9488 13304 -8796
rect 13338 -8810 13412 -8796
rect 13338 -9480 13412 -9470
rect 13338 -9488 13344 -9480
rect 13298 -9500 13344 -9488
rect 13406 -9488 13412 -9480
rect 13446 -9488 13452 -8796
rect 13406 -9500 13452 -9488
rect 13934 -8796 13980 -8784
rect 13934 -9488 13940 -8796
rect 13974 -9488 13980 -8796
rect 13934 -9500 13980 -9488
rect 14370 -8796 14416 -8784
rect 14370 -9488 14376 -8796
rect 14410 -9488 14416 -8796
rect 14370 -9500 14416 -9488
rect 14898 -8796 15052 -8784
rect 14898 -9488 14904 -8796
rect 14938 -9480 15012 -8796
rect 14938 -9488 14944 -9480
rect 14898 -9500 14944 -9488
rect 15006 -9488 15012 -9480
rect 15046 -9488 15052 -8796
rect 15006 -9500 15052 -9488
rect 15534 -8796 15580 -8784
rect 15534 -9488 15540 -8796
rect 15574 -9488 15580 -8796
rect 15534 -9500 15580 -9488
rect 15970 -8796 16016 -8784
rect 15970 -9488 15976 -8796
rect 16010 -9488 16016 -8796
rect 15970 -9500 16016 -9488
rect 16498 -8790 16544 -8784
rect 16606 -8790 16652 -8784
rect 16498 -8796 16652 -8790
rect 16498 -9488 16504 -8796
rect 16538 -8800 16612 -8796
rect 16538 -9488 16612 -9480
rect 16646 -9488 16652 -8796
rect 16498 -9490 16652 -9488
rect 16498 -9500 16544 -9490
rect 16606 -9500 16652 -9490
rect 17134 -8796 17180 -8784
rect 17134 -9488 17140 -8796
rect 17174 -9488 17180 -8796
rect 17134 -9500 17180 -9488
rect 17570 -8796 17616 -8784
rect 17570 -9488 17576 -8796
rect 17610 -9488 17616 -8796
rect 17570 -9500 17616 -9488
rect 18098 -8790 18144 -8784
rect 18206 -8790 18252 -8784
rect 18098 -8796 18252 -8790
rect 18098 -9488 18104 -8796
rect 18138 -8800 18212 -8796
rect 18138 -9488 18212 -9480
rect 18246 -9488 18252 -8796
rect 18098 -9490 18252 -9488
rect 18098 -9500 18144 -9490
rect 18206 -9500 18252 -9490
rect 18734 -8796 18780 -8784
rect 18734 -9488 18740 -8796
rect 18774 -9488 18780 -8796
rect 18734 -9500 18780 -9488
rect 19170 -8796 19216 -8784
rect 19170 -9488 19176 -8796
rect 19210 -9488 19216 -8796
rect 19170 -9500 19216 -9488
rect 19698 -8790 19744 -8784
rect 19806 -8790 19852 -8784
rect 19698 -8796 19852 -8790
rect 19698 -9488 19704 -8796
rect 19738 -8800 19812 -8796
rect 19738 -9488 19812 -9480
rect 19846 -9488 19852 -8796
rect 19698 -9490 19852 -9488
rect 19698 -9500 19744 -9490
rect 19806 -9500 19852 -9490
rect 20334 -8796 20380 -8784
rect 20334 -9488 20340 -8796
rect 20374 -9488 20380 -8796
rect 20334 -9500 20380 -9488
rect 20770 -8796 20816 -8784
rect 20770 -9488 20776 -8796
rect 20810 -9488 20816 -8796
rect 20770 -9500 20816 -9488
rect 21298 -8790 21344 -8784
rect 21406 -8790 21452 -8784
rect 21298 -8796 21452 -8790
rect 21298 -9488 21304 -8796
rect 21338 -8800 21412 -8796
rect 21338 -9488 21412 -9480
rect 21446 -9488 21452 -8796
rect 21298 -9490 21452 -9488
rect 21298 -9500 21344 -9490
rect 21406 -9500 21452 -9490
rect 21934 -8796 21980 -8784
rect 21934 -9488 21940 -8796
rect 21974 -9488 21980 -8796
rect 21934 -9500 21980 -9488
rect 22370 -8796 22416 -8784
rect 22370 -9488 22376 -8796
rect 22410 -9488 22416 -8796
rect 22370 -9500 22416 -9488
rect 22898 -8790 22944 -8784
rect 23006 -8790 23052 -8784
rect 22898 -8796 23052 -8790
rect 22898 -9488 22904 -8796
rect 22938 -8800 23012 -8796
rect 22938 -9488 23012 -9480
rect 23046 -9488 23052 -8796
rect 22898 -9490 23052 -9488
rect 22898 -9500 22944 -9490
rect 23006 -9500 23052 -9490
rect 23534 -8796 23580 -8784
rect 23534 -9488 23540 -8796
rect 23574 -9488 23580 -8796
rect 23534 -9500 23580 -9488
rect 23970 -8796 24016 -8784
rect 23970 -9488 23976 -8796
rect 24010 -9488 24016 -8796
rect 23970 -9500 24016 -9488
rect 24498 -8790 24544 -8784
rect 24606 -8790 24652 -8784
rect 24498 -8796 24652 -8790
rect 24498 -9488 24504 -8796
rect 24538 -8800 24612 -8796
rect 24538 -9488 24612 -9480
rect 24646 -9488 24652 -8796
rect 24498 -9490 24652 -9488
rect 24498 -9500 24544 -9490
rect 24606 -9500 24652 -9490
rect 25134 -8796 25180 -8784
rect 25134 -9488 25140 -8796
rect 25174 -9488 25180 -8796
rect 25134 -9500 25180 -9488
rect 25570 -8796 25616 -8784
rect 25570 -9488 25576 -8796
rect 25610 -9488 25616 -8796
rect 25570 -9500 25616 -9488
rect 26098 -8790 26144 -8784
rect 26206 -8790 26252 -8784
rect 26098 -8796 26252 -8790
rect 26098 -9488 26104 -8796
rect 26138 -8800 26212 -8796
rect 26138 -9488 26212 -9480
rect 26246 -9488 26252 -8796
rect 26098 -9490 26252 -9488
rect 26098 -9500 26144 -9490
rect 26206 -9500 26252 -9490
rect 26734 -8796 26780 -8784
rect 26734 -9488 26740 -8796
rect 26774 -9488 26780 -8796
rect 26734 -9500 26780 -9488
rect 27170 -8796 27216 -8784
rect 27170 -9488 27176 -8796
rect 27210 -9488 27216 -8796
rect 27170 -9500 27216 -9488
rect 27698 -8790 27744 -8784
rect 27806 -8790 27852 -8784
rect 27698 -8796 27852 -8790
rect 27698 -9488 27704 -8796
rect 27738 -8800 27812 -8796
rect 27738 -9488 27812 -9480
rect 27846 -9488 27852 -8796
rect 27698 -9490 27852 -9488
rect 27698 -9500 27744 -9490
rect 27806 -9500 27852 -9490
rect 28334 -8796 28380 -8784
rect 28334 -9488 28340 -8796
rect 28374 -9488 28380 -8796
rect 28334 -9500 28380 -9488
rect 28770 -8796 28816 -8784
rect 28770 -9488 28776 -8796
rect 28810 -9488 28816 -8796
rect 28770 -9500 28816 -9488
rect 29298 -8790 29344 -8784
rect 29406 -8790 29452 -8784
rect 29298 -8796 29452 -8790
rect 29298 -9488 29304 -8796
rect 29338 -8800 29412 -8796
rect 29338 -9488 29412 -9480
rect 29446 -9488 29452 -8796
rect 29298 -9490 29452 -9488
rect 29298 -9500 29344 -9490
rect 29406 -9500 29452 -9490
rect 29934 -8796 29980 -8784
rect 29934 -9488 29940 -8796
rect 29974 -9488 29980 -8796
rect 29934 -9500 29980 -9488
rect 30370 -8796 30416 -8784
rect 30370 -9488 30376 -8796
rect 30410 -9488 30416 -8796
rect 30370 -9500 30416 -9488
rect 30898 -8790 30944 -8784
rect 31006 -8790 31052 -8784
rect 30898 -8796 31052 -8790
rect 30898 -9488 30904 -8796
rect 30938 -8800 31012 -8796
rect 30938 -9488 31012 -9480
rect 31046 -9488 31052 -8796
rect 30898 -9490 31052 -9488
rect 30898 -9500 30944 -9490
rect 31006 -9500 31052 -9490
rect 31534 -8796 31580 -8784
rect 31534 -9488 31540 -8796
rect 31574 -9488 31580 -8796
rect 31534 -9500 31580 -9488
rect 31970 -8796 32016 -8784
rect 31970 -9488 31976 -8796
rect 32010 -9488 32016 -8796
rect 31970 -9500 32016 -9488
rect 32498 -8790 32544 -8784
rect 32606 -8790 32652 -8784
rect 32498 -8796 32652 -8790
rect 32498 -9488 32504 -8796
rect 32538 -8800 32612 -8796
rect 32538 -9488 32544 -9360
rect 32498 -9500 32544 -9488
rect 32606 -9488 32612 -9360
rect 32646 -9488 32652 -8796
rect 32606 -9500 32652 -9488
rect 33134 -8796 33180 -8784
rect 33134 -9488 33140 -8796
rect 33174 -9488 33180 -8796
rect 33134 -9500 33180 -9488
rect 33570 -8796 33616 -8784
rect 33570 -9488 33576 -8796
rect 33610 -9488 33616 -8796
rect 33570 -9500 33616 -9488
rect 34098 -8790 34144 -8784
rect 34206 -8790 34252 -8784
rect 34098 -8796 34252 -8790
rect 34098 -9488 34104 -8796
rect 34138 -8800 34212 -8796
rect 34138 -9488 34144 -9360
rect 34098 -9500 34144 -9488
rect 34206 -9488 34212 -9360
rect 34246 -9488 34252 -8796
rect 34206 -9500 34252 -9488
rect 34734 -8796 34780 -8784
rect 34734 -9488 34740 -8796
rect 34774 -9488 34780 -8796
rect 34734 -9500 34780 -9488
rect 35170 -8796 35216 -8784
rect 35170 -9488 35176 -8796
rect 35210 -9488 35216 -8796
rect 35170 -9500 35216 -9488
rect 35698 -8790 35744 -8784
rect 35806 -8790 35852 -8784
rect 35698 -8796 35852 -8790
rect 35698 -9488 35704 -8796
rect 35738 -8800 35812 -8796
rect 35738 -9488 35744 -9360
rect 35698 -9500 35744 -9488
rect 35806 -9488 35812 -9360
rect 35846 -9488 35852 -8796
rect 35806 -9500 35852 -9488
rect 36334 -8796 36380 -8784
rect 36334 -9488 36340 -8796
rect 36374 -9488 36380 -8796
rect 36334 -9500 36380 -9488
rect 36770 -8796 36816 -8784
rect 36770 -9488 36776 -8796
rect 36810 -9488 36816 -8796
rect 36770 -9500 36816 -9488
rect 37298 -8796 37344 -8784
rect 37298 -9488 37304 -8796
rect 37338 -9488 37344 -8796
rect 37298 -9500 37344 -9488
rect 37406 -8796 37452 -8784
rect 37406 -9488 37412 -8796
rect 37446 -9488 37452 -8796
rect 37406 -9500 37452 -9488
rect 37934 -8796 37980 -8784
rect 37934 -9488 37940 -8796
rect 37974 -9488 37980 -8796
rect 37934 -9500 37980 -9488
rect 33400 -9510 33540 -9500
rect 12857 -9550 13257 -9548
rect 13493 -9550 13893 -9548
rect 14457 -9550 14857 -9548
rect 15093 -9550 15493 -9548
rect 12480 -9554 15493 -9550
rect 12281 -9588 12420 -9580
rect 670 -9688 12420 -9588
rect 12480 -9588 12869 -9554
rect 13245 -9588 13505 -9554
rect 13881 -9588 14469 -9554
rect 14845 -9588 15105 -9554
rect 15481 -9588 15493 -9554
rect 16057 -9554 16457 -9548
rect 16057 -9580 16069 -9554
rect 12480 -9594 15493 -9588
rect 15700 -9588 16069 -9580
rect 16445 -9580 16457 -9554
rect 16693 -9554 17093 -9548
rect 16693 -9580 16705 -9554
rect 16445 -9588 16705 -9580
rect 17081 -9580 17093 -9554
rect 17657 -9554 18057 -9548
rect 17657 -9580 17669 -9554
rect 17081 -9588 17669 -9580
rect 18045 -9580 18057 -9554
rect 18293 -9554 18693 -9548
rect 18293 -9580 18305 -9554
rect 18045 -9588 18305 -9580
rect 18681 -9580 18693 -9554
rect 19257 -9554 19657 -9548
rect 19257 -9580 19269 -9554
rect 18681 -9588 19269 -9580
rect 19645 -9580 19657 -9554
rect 19893 -9554 20293 -9548
rect 19893 -9580 19905 -9554
rect 19645 -9588 19905 -9580
rect 20281 -9580 20293 -9554
rect 20857 -9554 21257 -9548
rect 20857 -9580 20869 -9554
rect 20281 -9588 20869 -9580
rect 21245 -9580 21257 -9554
rect 21493 -9554 21893 -9548
rect 21493 -9580 21505 -9554
rect 21245 -9588 21505 -9580
rect 21881 -9580 21893 -9554
rect 22457 -9554 22857 -9548
rect 22457 -9580 22469 -9554
rect 21881 -9588 22469 -9580
rect 22845 -9580 22857 -9554
rect 23093 -9554 23493 -9548
rect 23093 -9580 23105 -9554
rect 22845 -9588 23105 -9580
rect 23481 -9580 23493 -9554
rect 24057 -9554 24457 -9548
rect 24057 -9580 24069 -9554
rect 23481 -9588 24069 -9580
rect 24445 -9580 24457 -9554
rect 24693 -9554 25093 -9548
rect 24693 -9580 24705 -9554
rect 24445 -9588 24705 -9580
rect 25081 -9580 25093 -9554
rect 25657 -9554 26057 -9548
rect 25657 -9580 25669 -9554
rect 25081 -9588 25669 -9580
rect 26045 -9580 26057 -9554
rect 26293 -9554 26693 -9548
rect 26293 -9580 26305 -9554
rect 26045 -9588 26305 -9580
rect 26681 -9580 26693 -9554
rect 27257 -9554 27657 -9548
rect 27257 -9580 27269 -9554
rect 26681 -9588 27269 -9580
rect 27645 -9580 27657 -9554
rect 27893 -9554 28293 -9548
rect 27893 -9580 27905 -9554
rect 27645 -9588 27905 -9580
rect 28281 -9580 28293 -9554
rect 28857 -9554 29257 -9548
rect 28857 -9580 28869 -9554
rect 28281 -9588 28869 -9580
rect 29245 -9580 29257 -9554
rect 29493 -9554 29893 -9548
rect 29493 -9580 29505 -9554
rect 29245 -9588 29505 -9580
rect 29881 -9580 29893 -9554
rect 30457 -9554 30857 -9548
rect 30457 -9580 30469 -9554
rect 29881 -9588 30469 -9580
rect 30845 -9580 30857 -9554
rect 31093 -9554 31493 -9548
rect 31093 -9580 31105 -9554
rect 30845 -9588 31105 -9580
rect 31481 -9580 31493 -9554
rect 32057 -9550 32457 -9548
rect 32693 -9550 33093 -9548
rect 33400 -9550 33410 -9510
rect 32057 -9554 33410 -9550
rect 31481 -9588 31760 -9580
rect 12480 -9620 15490 -9594
rect 0 -9722 13 -9688
rect 1137 -9722 1613 -9688
rect 2737 -9722 3213 -9688
rect 4337 -9722 4813 -9688
rect 5937 -9722 6413 -9688
rect 7537 -9722 8013 -9688
rect 9137 -9722 9613 -9688
rect 10737 -9722 11213 -9688
rect 12337 -9700 12420 -9688
rect 12801 -9688 13949 -9682
rect 12801 -9700 12813 -9688
rect 12337 -9722 12813 -9700
rect 13937 -9700 13949 -9688
rect 14401 -9688 15549 -9682
rect 14401 -9700 14413 -9688
rect 13937 -9722 14413 -9700
rect 15537 -9700 15549 -9688
rect 15700 -9688 31760 -9588
rect 32057 -9588 32069 -9554
rect 32445 -9588 32705 -9554
rect 33081 -9588 33410 -9554
rect 32057 -9594 33410 -9588
rect 32060 -9630 33410 -9594
rect 33530 -9550 33540 -9510
rect 33657 -9550 34057 -9548
rect 34293 -9550 34693 -9548
rect 35257 -9550 35657 -9548
rect 35893 -9550 36293 -9548
rect 33530 -9554 36293 -9550
rect 33530 -9588 33669 -9554
rect 34045 -9588 34305 -9554
rect 34681 -9588 35269 -9554
rect 35645 -9588 35905 -9554
rect 36281 -9588 36293 -9554
rect 33530 -9594 36293 -9588
rect 36857 -9554 37257 -9548
rect 36857 -9588 36869 -9554
rect 37245 -9588 37257 -9554
rect 36857 -9594 37257 -9588
rect 37493 -9554 37893 -9548
rect 37493 -9588 37505 -9554
rect 37881 -9588 37893 -9554
rect 37493 -9594 37893 -9588
rect 33530 -9630 36290 -9594
rect 32060 -9640 36290 -9630
rect 15700 -9700 16013 -9688
rect 15537 -9722 16013 -9700
rect 17137 -9722 17613 -9688
rect 18737 -9722 19213 -9688
rect 20337 -9722 20813 -9688
rect 21937 -9722 22413 -9688
rect 23537 -9722 24013 -9688
rect 25137 -9722 25613 -9688
rect 26737 -9722 27213 -9688
rect 28337 -9722 28813 -9688
rect 29937 -9722 30413 -9688
rect 31537 -9700 31760 -9688
rect 32001 -9688 33149 -9682
rect 32001 -9700 32013 -9688
rect 31537 -9722 32013 -9700
rect 33137 -9700 33149 -9688
rect 33601 -9688 34749 -9682
rect 33601 -9700 33613 -9688
rect 33137 -9722 33613 -9700
rect 34737 -9700 34749 -9688
rect 35201 -9688 36349 -9682
rect 35201 -9700 35213 -9688
rect 34737 -9722 35213 -9700
rect 36337 -9700 36349 -9688
rect 36801 -9688 37949 -9682
rect 36801 -9700 36813 -9688
rect 36337 -9722 36813 -9700
rect 37937 -9722 37949 -9688
rect 0 -9820 490 -9722
rect 440 -9964 490 -9820
rect 57 -9970 490 -9964
rect 57 -10004 69 -9970
rect 445 -10004 490 -9970
rect 57 -10010 490 -10004
rect -30 -10057 16 -10045
rect -30 -10175 -24 -10057
rect 10 -10175 16 -10057
rect -30 -10187 16 -10175
rect 440 -10222 490 -10010
rect 670 -9728 37949 -9722
rect 670 -9820 37940 -9728
rect 670 -9964 720 -9820
rect 1200 -9870 1340 -9860
rect 670 -9970 1093 -9964
rect 670 -10004 705 -9970
rect 1081 -10004 1093 -9970
rect 1200 -9990 1210 -9870
rect 1330 -9880 1340 -9870
rect 2800 -9870 2940 -9860
rect 2800 -9880 2810 -9870
rect 1330 -9970 2810 -9880
rect 1330 -9980 1669 -9970
rect 1330 -9990 1340 -9980
rect 1200 -10000 1340 -9990
rect 670 -10010 1093 -10004
rect 1657 -10004 1669 -9980
rect 2045 -9980 2305 -9970
rect 2045 -10004 2057 -9980
rect 1657 -10010 2057 -10004
rect 2293 -10004 2305 -9980
rect 2681 -9980 2810 -9970
rect 2681 -10004 2693 -9980
rect 2800 -9990 2810 -9980
rect 2930 -9880 2940 -9870
rect 4400 -9870 4540 -9860
rect 4400 -9880 4410 -9870
rect 2930 -9970 4410 -9880
rect 2930 -9980 3269 -9970
rect 2930 -9990 2940 -9980
rect 2800 -10000 2940 -9990
rect 2293 -10010 2693 -10004
rect 3257 -10004 3269 -9980
rect 3645 -9980 3905 -9970
rect 3645 -10004 3657 -9980
rect 3257 -10010 3657 -10004
rect 3893 -10004 3905 -9980
rect 4281 -9980 4410 -9970
rect 4281 -10004 4293 -9980
rect 4400 -9990 4410 -9980
rect 4530 -9880 4540 -9870
rect 6000 -9870 6140 -9860
rect 6000 -9880 6010 -9870
rect 4530 -9970 6010 -9880
rect 4530 -9980 4869 -9970
rect 4530 -9990 4540 -9980
rect 4400 -10000 4540 -9990
rect 3893 -10010 4293 -10004
rect 4857 -10004 4869 -9980
rect 5245 -9980 5505 -9970
rect 5245 -10004 5257 -9980
rect 4857 -10010 5257 -10004
rect 5493 -10004 5505 -9980
rect 5881 -9980 6010 -9970
rect 5881 -10004 5893 -9980
rect 6000 -9990 6010 -9980
rect 6130 -9880 6140 -9870
rect 7600 -9870 7740 -9860
rect 7600 -9880 7610 -9870
rect 6130 -9970 7610 -9880
rect 6130 -9980 6469 -9970
rect 6130 -9990 6140 -9980
rect 6000 -10000 6140 -9990
rect 5493 -10010 5893 -10004
rect 6457 -10004 6469 -9980
rect 6845 -9980 7105 -9970
rect 6845 -10004 6857 -9980
rect 6457 -10010 6857 -10004
rect 7093 -10004 7105 -9980
rect 7481 -9980 7610 -9970
rect 7481 -10004 7493 -9980
rect 7600 -9990 7610 -9980
rect 7730 -9880 7740 -9870
rect 9200 -9870 9340 -9860
rect 9200 -9880 9210 -9870
rect 7730 -9970 9210 -9880
rect 7730 -9980 8069 -9970
rect 7730 -9990 7740 -9980
rect 7600 -10000 7740 -9990
rect 7093 -10010 7493 -10004
rect 8057 -10004 8069 -9980
rect 8445 -9980 8705 -9970
rect 8445 -10004 8457 -9980
rect 8057 -10010 8457 -10004
rect 8693 -10004 8705 -9980
rect 9081 -9980 9210 -9970
rect 9081 -10004 9093 -9980
rect 9200 -9990 9210 -9980
rect 9330 -9880 9340 -9870
rect 15820 -9870 15960 -9860
rect 9330 -9970 10700 -9880
rect 9330 -9980 9669 -9970
rect 9330 -9990 9340 -9980
rect 9200 -10000 9340 -9990
rect 8693 -10010 9093 -10004
rect 9657 -10004 9669 -9980
rect 10045 -9980 10305 -9970
rect 10045 -10004 10057 -9980
rect 9657 -10010 10057 -10004
rect 10293 -10004 10305 -9980
rect 10681 -9980 10700 -9970
rect 11257 -9970 11657 -9964
rect 10681 -10004 10693 -9980
rect 10293 -10010 10693 -10004
rect 11257 -10004 11269 -9970
rect 11645 -10004 11657 -9970
rect 11257 -10010 11657 -10004
rect 11893 -9970 12293 -9964
rect 11893 -10004 11905 -9970
rect 12281 -10004 12293 -9970
rect 11893 -10010 12293 -10004
rect 12857 -9970 13257 -9964
rect 12857 -10004 12869 -9970
rect 13245 -10004 13257 -9970
rect 12857 -10010 13257 -10004
rect 13493 -9970 13893 -9964
rect 13493 -10004 13505 -9970
rect 13881 -10004 13893 -9970
rect 13493 -10010 13893 -10004
rect 14457 -9970 14857 -9964
rect 14457 -10004 14469 -9970
rect 14845 -10004 14857 -9970
rect 14457 -10010 14857 -10004
rect 15093 -9970 15493 -9964
rect 15093 -10004 15105 -9970
rect 15481 -10004 15493 -9970
rect 15820 -9990 15830 -9870
rect 15950 -9900 15960 -9870
rect 17420 -9870 17560 -9860
rect 15950 -9964 17090 -9900
rect 15950 -9970 17093 -9964
rect 15950 -9990 16069 -9970
rect 15820 -10000 16069 -9990
rect 15093 -10010 15493 -10004
rect 16057 -10004 16069 -10000
rect 16445 -10000 16705 -9970
rect 16445 -10004 16457 -10000
rect 16057 -10010 16457 -10004
rect 16693 -10004 16705 -10000
rect 17081 -10004 17093 -9970
rect 17420 -9990 17430 -9870
rect 17550 -9900 17560 -9870
rect 19020 -9870 19160 -9860
rect 17550 -9964 18690 -9900
rect 17550 -9970 18693 -9964
rect 17550 -9990 17669 -9970
rect 17420 -10000 17669 -9990
rect 16693 -10010 17093 -10004
rect 17657 -10004 17669 -10000
rect 18045 -10000 18305 -9970
rect 18045 -10004 18057 -10000
rect 17657 -10010 18057 -10004
rect 18293 -10004 18305 -10000
rect 18681 -10004 18693 -9970
rect 19020 -9990 19030 -9870
rect 19150 -9900 19160 -9870
rect 20620 -9870 20760 -9860
rect 19150 -9964 20290 -9900
rect 19150 -9970 20293 -9964
rect 19150 -9990 19269 -9970
rect 19020 -10000 19269 -9990
rect 18293 -10010 18693 -10004
rect 19257 -10004 19269 -10000
rect 19645 -10000 19905 -9970
rect 19645 -10004 19657 -10000
rect 19257 -10010 19657 -10004
rect 19893 -10004 19905 -10000
rect 20281 -10004 20293 -9970
rect 20620 -9990 20630 -9870
rect 20750 -9900 20760 -9870
rect 22220 -9870 22360 -9860
rect 20750 -9964 21890 -9900
rect 20750 -9970 21893 -9964
rect 20750 -9990 20869 -9970
rect 20620 -10000 20869 -9990
rect 19893 -10010 20293 -10004
rect 20857 -10004 20869 -10000
rect 21245 -10000 21505 -9970
rect 21245 -10004 21257 -10000
rect 20857 -10010 21257 -10004
rect 21493 -10004 21505 -10000
rect 21881 -10004 21893 -9970
rect 22220 -9990 22230 -9870
rect 22350 -9900 22360 -9870
rect 23820 -9870 23960 -9860
rect 22350 -9964 23490 -9900
rect 22350 -9970 23493 -9964
rect 22350 -9990 22469 -9970
rect 22220 -10000 22469 -9990
rect 21493 -10010 21893 -10004
rect 22457 -10004 22469 -10000
rect 22845 -10000 23105 -9970
rect 22845 -10004 22857 -10000
rect 22457 -10010 22857 -10004
rect 23093 -10004 23105 -10000
rect 23481 -10004 23493 -9970
rect 23820 -9990 23830 -9870
rect 23950 -9900 23960 -9870
rect 25420 -9870 25560 -9860
rect 23950 -9964 25090 -9900
rect 23950 -9970 25093 -9964
rect 23950 -9990 24069 -9970
rect 23820 -10000 24069 -9990
rect 23093 -10010 23493 -10004
rect 24057 -10004 24069 -10000
rect 24445 -10000 24705 -9970
rect 24445 -10004 24457 -10000
rect 24057 -10010 24457 -10004
rect 24693 -10004 24705 -10000
rect 25081 -10004 25093 -9970
rect 25420 -9990 25430 -9870
rect 25550 -9900 25560 -9870
rect 27020 -9870 27160 -9860
rect 25550 -9964 26680 -9900
rect 25550 -9970 26693 -9964
rect 25550 -9990 25669 -9970
rect 25420 -10000 25669 -9990
rect 24693 -10010 25093 -10004
rect 25657 -10004 25669 -10000
rect 26045 -10000 26305 -9970
rect 26045 -10004 26057 -10000
rect 25657 -10010 26057 -10004
rect 26293 -10004 26305 -10000
rect 26681 -10004 26693 -9970
rect 27020 -9990 27030 -9870
rect 27150 -9900 27160 -9870
rect 28620 -9870 28760 -9860
rect 27150 -9964 28290 -9900
rect 27150 -9970 28293 -9964
rect 27150 -9990 27269 -9970
rect 27020 -10000 27269 -9990
rect 26293 -10010 26693 -10004
rect 27257 -10004 27269 -10000
rect 27645 -10000 27905 -9970
rect 27645 -10004 27657 -10000
rect 27257 -10010 27657 -10004
rect 27893 -10004 27905 -10000
rect 28281 -10004 28293 -9970
rect 28620 -9990 28630 -9870
rect 28750 -9900 28760 -9870
rect 30220 -9870 30360 -9860
rect 28750 -9964 29890 -9900
rect 28750 -9970 29893 -9964
rect 28750 -9990 28869 -9970
rect 28620 -10000 28869 -9990
rect 27893 -10010 28293 -10004
rect 28857 -10004 28869 -10000
rect 29245 -10000 29505 -9970
rect 29245 -10004 29257 -10000
rect 28857 -10010 29257 -10004
rect 29493 -10004 29505 -10000
rect 29881 -10004 29893 -9970
rect 30220 -9990 30230 -9870
rect 30350 -9900 30360 -9870
rect 31820 -9870 31960 -9860
rect 30350 -9964 31490 -9900
rect 30350 -9970 31493 -9964
rect 30350 -9990 30469 -9970
rect 30220 -10000 30469 -9990
rect 29493 -10010 29893 -10004
rect 30457 -10004 30469 -10000
rect 30845 -10000 31105 -9970
rect 30845 -10004 30857 -10000
rect 30457 -10010 30857 -10004
rect 31093 -10004 31105 -10000
rect 31481 -10004 31493 -9970
rect 31820 -9990 31830 -9870
rect 31950 -9900 31960 -9870
rect 34800 -9870 34940 -9860
rect 34800 -9900 34810 -9870
rect 31950 -9970 34810 -9900
rect 31950 -9990 32069 -9970
rect 31820 -10000 32069 -9990
rect 31093 -10010 31493 -10004
rect 32057 -10004 32069 -10000
rect 32445 -10000 32705 -9970
rect 32445 -10004 32457 -10000
rect 32057 -10010 32457 -10004
rect 32693 -10004 32705 -10000
rect 33081 -10000 33669 -9970
rect 33081 -10004 33093 -10000
rect 32693 -10010 33093 -10004
rect 33657 -10004 33669 -10000
rect 34045 -10000 34305 -9970
rect 34045 -10004 34057 -10000
rect 33657 -10010 34057 -10004
rect 34293 -10004 34305 -10000
rect 34681 -9990 34810 -9970
rect 34930 -9900 34940 -9870
rect 34930 -9964 36280 -9900
rect 34930 -9970 36293 -9964
rect 34930 -9990 35269 -9970
rect 34681 -10000 35269 -9990
rect 34681 -10004 34693 -10000
rect 34293 -10010 34693 -10004
rect 35257 -10004 35269 -10000
rect 35645 -10000 35905 -9970
rect 35645 -10004 35657 -10000
rect 35257 -10010 35657 -10004
rect 35893 -10004 35905 -10000
rect 36281 -10004 36293 -9970
rect 35893 -10010 36293 -10004
rect 36857 -9970 37257 -9964
rect 36857 -10004 36869 -9970
rect 37245 -10004 37257 -9970
rect 36857 -10010 37257 -10004
rect 37493 -9970 37893 -9964
rect 37493 -10004 37505 -9970
rect 37881 -10004 37893 -9970
rect 37493 -10010 37893 -10004
rect 57 -10228 490 -10222
rect 57 -10262 69 -10228
rect 445 -10262 490 -10228
rect 57 -10268 490 -10262
rect 440 -10490 490 -10268
rect 57 -10496 490 -10490
rect 57 -10530 69 -10496
rect 445 -10530 490 -10496
rect 57 -10536 490 -10530
rect -30 -10596 16 -10584
rect -30 -11288 -24 -10596
rect 10 -11288 16 -10596
rect -30 -11300 16 -11288
rect 440 -11348 490 -10536
rect 670 -10222 720 -10010
rect 1134 -10057 1180 -10045
rect 1134 -10175 1140 -10057
rect 1174 -10175 1180 -10057
rect 1570 -10057 1616 -10045
rect 1570 -10060 1576 -10057
rect 1134 -10187 1180 -10175
rect 1560 -10175 1576 -10060
rect 1610 -10060 1616 -10057
rect 2098 -10057 2144 -10045
rect 2098 -10060 2104 -10057
rect 1610 -10175 2104 -10060
rect 2138 -10060 2144 -10057
rect 2206 -10057 2252 -10045
rect 2206 -10060 2212 -10057
rect 2138 -10175 2212 -10060
rect 2246 -10060 2252 -10057
rect 2734 -10057 2780 -10045
rect 2734 -10060 2740 -10057
rect 2246 -10175 2740 -10060
rect 2774 -10060 2780 -10057
rect 3170 -10057 3216 -10045
rect 3170 -10060 3176 -10057
rect 2774 -10175 3176 -10060
rect 3210 -10060 3216 -10057
rect 3698 -10057 3744 -10045
rect 3698 -10060 3704 -10057
rect 3210 -10175 3704 -10060
rect 3738 -10060 3744 -10057
rect 3806 -10057 3852 -10045
rect 3806 -10060 3812 -10057
rect 3738 -10175 3812 -10060
rect 3846 -10060 3852 -10057
rect 4334 -10057 4380 -10045
rect 4334 -10060 4340 -10057
rect 3846 -10175 4340 -10060
rect 4374 -10060 4380 -10057
rect 4770 -10057 4816 -10045
rect 4770 -10060 4776 -10057
rect 4374 -10175 4776 -10060
rect 4810 -10060 4816 -10057
rect 5298 -10057 5344 -10045
rect 5298 -10060 5304 -10057
rect 4810 -10175 5304 -10060
rect 5338 -10060 5344 -10057
rect 5406 -10057 5452 -10045
rect 5406 -10060 5412 -10057
rect 5338 -10175 5412 -10060
rect 5446 -10060 5452 -10057
rect 5934 -10057 5980 -10045
rect 5934 -10060 5940 -10057
rect 5446 -10175 5940 -10060
rect 5974 -10060 5980 -10057
rect 6370 -10057 6416 -10045
rect 6370 -10060 6376 -10057
rect 5974 -10175 6376 -10060
rect 6410 -10060 6416 -10057
rect 6898 -10057 6944 -10045
rect 6898 -10060 6904 -10057
rect 6410 -10175 6904 -10060
rect 6938 -10060 6944 -10057
rect 7006 -10057 7052 -10045
rect 7006 -10060 7012 -10057
rect 6938 -10175 7012 -10060
rect 7046 -10060 7052 -10057
rect 7534 -10057 7580 -10045
rect 7534 -10060 7540 -10057
rect 7046 -10175 7540 -10060
rect 7574 -10060 7580 -10057
rect 7970 -10057 8016 -10045
rect 7970 -10060 7976 -10057
rect 7574 -10175 7976 -10060
rect 8010 -10060 8016 -10057
rect 8498 -10057 8544 -10045
rect 8498 -10060 8504 -10057
rect 8010 -10175 8504 -10060
rect 8538 -10060 8544 -10057
rect 8606 -10057 8652 -10045
rect 8606 -10060 8612 -10057
rect 8538 -10175 8612 -10060
rect 8646 -10060 8652 -10057
rect 9134 -10057 9180 -10045
rect 9134 -10060 9140 -10057
rect 8646 -10175 9140 -10060
rect 9174 -10060 9180 -10057
rect 9570 -10057 9616 -10045
rect 9570 -10060 9576 -10057
rect 9174 -10175 9576 -10060
rect 9610 -10060 9616 -10057
rect 10098 -10057 10144 -10045
rect 10098 -10060 10104 -10057
rect 9610 -10175 10104 -10060
rect 10138 -10060 10144 -10057
rect 10206 -10057 10252 -10045
rect 10206 -10060 10212 -10057
rect 10138 -10175 10212 -10060
rect 10246 -10060 10252 -10057
rect 10734 -10050 10780 -10045
rect 10734 -10057 10940 -10050
rect 10734 -10060 10740 -10057
rect 10246 -10175 10740 -10060
rect 10774 -10060 10940 -10057
rect 11170 -10057 11216 -10045
rect 11170 -10060 11176 -10057
rect 10774 -10175 10810 -10060
rect 1560 -10180 10810 -10175
rect 10930 -10175 11176 -10060
rect 11210 -10060 11216 -10057
rect 11400 -10060 11520 -10010
rect 11698 -10057 11744 -10045
rect 11698 -10060 11704 -10057
rect 11210 -10175 11704 -10060
rect 11738 -10060 11744 -10057
rect 11806 -10057 11852 -10045
rect 11806 -10060 11812 -10057
rect 11738 -10175 11812 -10060
rect 11846 -10060 11852 -10057
rect 12040 -10060 12160 -10010
rect 12334 -10057 12380 -10045
rect 12334 -10060 12340 -10057
rect 11846 -10175 12340 -10060
rect 12374 -10060 12380 -10057
rect 12770 -10057 12816 -10045
rect 12770 -10060 12776 -10057
rect 12374 -10175 12776 -10060
rect 12810 -10060 12816 -10057
rect 13000 -10060 13120 -10010
rect 13298 -10057 13344 -10045
rect 13298 -10060 13304 -10057
rect 12810 -10175 13304 -10060
rect 13338 -10060 13344 -10057
rect 13406 -10057 13452 -10045
rect 13406 -10060 13412 -10057
rect 13338 -10175 13412 -10060
rect 13446 -10060 13452 -10057
rect 13640 -10060 13760 -10010
rect 13934 -10057 13980 -10045
rect 13934 -10060 13940 -10057
rect 13446 -10175 13940 -10060
rect 13974 -10060 13980 -10057
rect 14370 -10057 14416 -10045
rect 14370 -10060 14376 -10057
rect 13974 -10175 14376 -10060
rect 14410 -10060 14416 -10057
rect 14600 -10060 14720 -10010
rect 14898 -10057 14944 -10045
rect 14898 -10060 14904 -10057
rect 14410 -10175 14904 -10060
rect 14938 -10060 14944 -10057
rect 15006 -10057 15052 -10045
rect 15006 -10060 15012 -10057
rect 14938 -10175 15012 -10060
rect 15046 -10060 15052 -10057
rect 15240 -10060 15360 -10010
rect 15534 -10057 15580 -10045
rect 15534 -10060 15540 -10057
rect 15046 -10175 15540 -10060
rect 15574 -10060 15580 -10057
rect 15970 -10057 16016 -10045
rect 15970 -10060 15976 -10057
rect 15574 -10175 15976 -10060
rect 16010 -10060 16016 -10057
rect 16498 -10057 16544 -10045
rect 16498 -10060 16504 -10057
rect 16010 -10175 16504 -10060
rect 16538 -10060 16544 -10057
rect 16606 -10057 16652 -10045
rect 16606 -10060 16612 -10057
rect 16538 -10175 16612 -10060
rect 16646 -10060 16652 -10057
rect 17134 -10057 17180 -10045
rect 17134 -10060 17140 -10057
rect 16646 -10175 17140 -10060
rect 17174 -10060 17180 -10057
rect 17570 -10057 17616 -10045
rect 17570 -10060 17576 -10057
rect 17174 -10175 17576 -10060
rect 17610 -10060 17616 -10057
rect 18098 -10057 18144 -10045
rect 18098 -10060 18104 -10057
rect 17610 -10175 18104 -10060
rect 18138 -10060 18144 -10057
rect 18206 -10057 18252 -10045
rect 18206 -10060 18212 -10057
rect 18138 -10175 18212 -10060
rect 18246 -10060 18252 -10057
rect 18734 -10057 18780 -10045
rect 18734 -10060 18740 -10057
rect 18246 -10175 18740 -10060
rect 18774 -10060 18780 -10057
rect 19170 -10057 19216 -10045
rect 19170 -10060 19176 -10057
rect 18774 -10175 19176 -10060
rect 19210 -10060 19216 -10057
rect 19698 -10057 19744 -10045
rect 19698 -10060 19704 -10057
rect 19210 -10175 19704 -10060
rect 19738 -10060 19744 -10057
rect 19806 -10057 19852 -10045
rect 19806 -10060 19812 -10057
rect 19738 -10175 19812 -10060
rect 19846 -10060 19852 -10057
rect 20334 -10057 20380 -10045
rect 20334 -10060 20340 -10057
rect 19846 -10175 20340 -10060
rect 20374 -10060 20380 -10057
rect 20770 -10057 20816 -10045
rect 20770 -10060 20776 -10057
rect 20374 -10175 20776 -10060
rect 20810 -10060 20816 -10057
rect 21298 -10057 21344 -10045
rect 21298 -10060 21304 -10057
rect 20810 -10175 21304 -10060
rect 21338 -10060 21344 -10057
rect 21406 -10057 21452 -10045
rect 21406 -10060 21412 -10057
rect 21338 -10175 21412 -10060
rect 21446 -10060 21452 -10057
rect 21934 -10057 21980 -10045
rect 21934 -10060 21940 -10057
rect 21446 -10175 21940 -10060
rect 21974 -10060 21980 -10057
rect 22370 -10057 22416 -10045
rect 22370 -10060 22376 -10057
rect 21974 -10175 22376 -10060
rect 22410 -10060 22416 -10057
rect 22898 -10057 22944 -10045
rect 22898 -10060 22904 -10057
rect 22410 -10175 22904 -10060
rect 22938 -10060 22944 -10057
rect 23006 -10057 23052 -10045
rect 23006 -10060 23012 -10057
rect 22938 -10175 23012 -10060
rect 23046 -10060 23052 -10057
rect 23534 -10057 23580 -10045
rect 23534 -10060 23540 -10057
rect 23046 -10175 23540 -10060
rect 23574 -10060 23580 -10057
rect 23970 -10057 24016 -10045
rect 23970 -10060 23976 -10057
rect 23574 -10175 23976 -10060
rect 24010 -10060 24016 -10057
rect 24498 -10057 24544 -10045
rect 24498 -10060 24504 -10057
rect 24010 -10175 24504 -10060
rect 24538 -10060 24544 -10057
rect 24606 -10057 24652 -10045
rect 24606 -10060 24612 -10057
rect 24538 -10175 24612 -10060
rect 24646 -10060 24652 -10057
rect 25134 -10057 25180 -10045
rect 25134 -10060 25140 -10057
rect 24646 -10175 25140 -10060
rect 25174 -10060 25180 -10057
rect 25570 -10057 25616 -10045
rect 25570 -10060 25576 -10057
rect 25174 -10175 25576 -10060
rect 25610 -10060 25616 -10057
rect 26098 -10057 26144 -10045
rect 26098 -10060 26104 -10057
rect 25610 -10175 26104 -10060
rect 26138 -10060 26144 -10057
rect 26206 -10057 26252 -10045
rect 26206 -10060 26212 -10057
rect 26138 -10175 26212 -10060
rect 26246 -10060 26252 -10057
rect 26734 -10057 26780 -10045
rect 26734 -10060 26740 -10057
rect 26246 -10175 26740 -10060
rect 26774 -10060 26780 -10057
rect 27170 -10057 27216 -10045
rect 27170 -10060 27176 -10057
rect 26774 -10175 27176 -10060
rect 27210 -10060 27216 -10057
rect 27698 -10057 27744 -10045
rect 27698 -10060 27704 -10057
rect 27210 -10175 27704 -10060
rect 27738 -10060 27744 -10057
rect 27806 -10057 27852 -10045
rect 27806 -10060 27812 -10057
rect 27738 -10175 27812 -10060
rect 27846 -10060 27852 -10057
rect 28334 -10057 28380 -10045
rect 28334 -10060 28340 -10057
rect 27846 -10175 28340 -10060
rect 28374 -10060 28380 -10057
rect 28770 -10057 28816 -10045
rect 28770 -10060 28776 -10057
rect 28374 -10175 28776 -10060
rect 28810 -10060 28816 -10057
rect 29298 -10057 29344 -10045
rect 29298 -10060 29304 -10057
rect 28810 -10175 29304 -10060
rect 29338 -10060 29344 -10057
rect 29406 -10057 29452 -10045
rect 29406 -10060 29412 -10057
rect 29338 -10175 29412 -10060
rect 29446 -10060 29452 -10057
rect 29934 -10057 29980 -10045
rect 29934 -10060 29940 -10057
rect 29446 -10175 29940 -10060
rect 29974 -10060 29980 -10057
rect 30370 -10057 30416 -10037
rect 30370 -10060 30376 -10057
rect 29974 -10175 30376 -10060
rect 30410 -10060 30416 -10057
rect 30898 -10057 30944 -10037
rect 30898 -10060 30904 -10057
rect 30410 -10175 30904 -10060
rect 30938 -10060 30944 -10057
rect 31006 -10057 31052 -10037
rect 31006 -10060 31012 -10057
rect 30938 -10175 31012 -10060
rect 31046 -10060 31052 -10057
rect 31534 -10057 31580 -10045
rect 31534 -10060 31540 -10057
rect 31046 -10175 31540 -10060
rect 31574 -10060 31580 -10057
rect 31970 -10057 32016 -10045
rect 31970 -10060 31976 -10057
rect 31574 -10175 31976 -10060
rect 32010 -10060 32016 -10057
rect 32498 -10057 32544 -10045
rect 32498 -10060 32504 -10057
rect 32010 -10175 32504 -10060
rect 32538 -10060 32544 -10057
rect 32606 -10057 32652 -10045
rect 32606 -10060 32612 -10057
rect 32538 -10175 32612 -10060
rect 32646 -10060 32652 -10057
rect 33134 -10057 33180 -10045
rect 33134 -10060 33140 -10057
rect 32646 -10175 33140 -10060
rect 33174 -10060 33180 -10057
rect 33570 -10057 33616 -10045
rect 33570 -10060 33576 -10057
rect 33174 -10175 33576 -10060
rect 33610 -10060 33616 -10057
rect 34098 -10057 34144 -10045
rect 34098 -10060 34104 -10057
rect 33610 -10175 34104 -10060
rect 34138 -10060 34144 -10057
rect 34206 -10057 34252 -10045
rect 34206 -10060 34212 -10057
rect 34138 -10175 34212 -10060
rect 34246 -10060 34252 -10057
rect 34734 -10057 34780 -10045
rect 34734 -10060 34740 -10057
rect 34246 -10175 34740 -10060
rect 34774 -10060 34780 -10057
rect 35170 -10057 35216 -10045
rect 35170 -10060 35176 -10057
rect 34774 -10175 35176 -10060
rect 35210 -10060 35216 -10057
rect 35698 -10057 35744 -10045
rect 35698 -10060 35704 -10057
rect 35210 -10175 35704 -10060
rect 35738 -10060 35744 -10057
rect 35806 -10057 35852 -10045
rect 35806 -10060 35812 -10057
rect 35738 -10175 35812 -10060
rect 35846 -10060 35852 -10057
rect 36334 -10057 36380 -10045
rect 36334 -10060 36340 -10057
rect 35846 -10175 36340 -10060
rect 36374 -10175 36380 -10057
rect 10930 -10180 36380 -10175
rect 1570 -10187 1616 -10180
rect 2098 -10187 2144 -10180
rect 2206 -10187 2252 -10180
rect 2734 -10187 2780 -10180
rect 3170 -10187 3216 -10180
rect 3698 -10187 3744 -10180
rect 3806 -10187 3852 -10180
rect 4334 -10187 4380 -10180
rect 4770 -10187 4816 -10180
rect 5298 -10187 5344 -10180
rect 5406 -10187 5452 -10180
rect 5934 -10187 5980 -10180
rect 6370 -10187 6416 -10180
rect 6898 -10187 6944 -10180
rect 7006 -10187 7052 -10180
rect 7534 -10187 7580 -10180
rect 7970 -10187 8016 -10180
rect 8498 -10187 8544 -10180
rect 8606 -10187 8652 -10180
rect 9134 -10187 9180 -10180
rect 9570 -10187 9616 -10180
rect 10098 -10187 10144 -10180
rect 10206 -10187 10252 -10180
rect 10734 -10187 10940 -10180
rect 11170 -10187 11216 -10180
rect 10750 -10190 10940 -10187
rect 11400 -10222 11520 -10180
rect 11698 -10187 11744 -10180
rect 11806 -10187 11852 -10180
rect 12040 -10222 12160 -10180
rect 12334 -10187 12380 -10180
rect 12770 -10187 12816 -10180
rect 13000 -10222 13120 -10180
rect 13298 -10187 13344 -10180
rect 13406 -10187 13452 -10180
rect 13640 -10222 13760 -10180
rect 13934 -10187 13980 -10180
rect 14370 -10187 14416 -10180
rect 14600 -10222 14720 -10180
rect 14898 -10187 14944 -10180
rect 15006 -10187 15052 -10180
rect 15240 -10222 15360 -10180
rect 15534 -10187 15580 -10180
rect 15970 -10187 16016 -10180
rect 16498 -10187 16544 -10180
rect 16606 -10187 16652 -10180
rect 17134 -10187 17180 -10180
rect 17570 -10187 17616 -10180
rect 18098 -10187 18144 -10180
rect 18206 -10187 18252 -10180
rect 18734 -10187 18780 -10180
rect 19170 -10187 19216 -10180
rect 19698 -10187 19744 -10180
rect 19806 -10187 19852 -10180
rect 20334 -10187 20380 -10180
rect 20770 -10187 20816 -10180
rect 21298 -10187 21344 -10180
rect 21406 -10187 21452 -10180
rect 21934 -10187 21980 -10180
rect 22370 -10187 22416 -10180
rect 22898 -10187 22944 -10180
rect 23006 -10187 23052 -10180
rect 23534 -10187 23580 -10180
rect 23970 -10187 24016 -10180
rect 24498 -10187 24544 -10180
rect 24606 -10187 24652 -10180
rect 25134 -10187 25180 -10180
rect 25570 -10187 25616 -10180
rect 26098 -10187 26144 -10180
rect 26206 -10187 26252 -10180
rect 26734 -10187 26780 -10180
rect 27170 -10187 27216 -10180
rect 27698 -10187 27744 -10180
rect 27806 -10187 27852 -10180
rect 28334 -10187 28380 -10180
rect 28770 -10187 28816 -10180
rect 29298 -10187 29344 -10180
rect 29406 -10187 29452 -10180
rect 29934 -10187 29980 -10180
rect 30370 -10195 30416 -10180
rect 30898 -10195 30944 -10180
rect 31006 -10195 31052 -10180
rect 31534 -10187 31580 -10180
rect 31970 -10187 32016 -10180
rect 32498 -10187 32544 -10180
rect 32606 -10187 32652 -10180
rect 33134 -10187 33180 -10180
rect 33570 -10187 33616 -10180
rect 34098 -10187 34144 -10180
rect 34206 -10187 34252 -10180
rect 34734 -10187 34780 -10180
rect 35170 -10187 35216 -10180
rect 35698 -10187 35744 -10180
rect 35806 -10187 35852 -10180
rect 36334 -10187 36380 -10180
rect 36770 -10057 36816 -10045
rect 36770 -10175 36776 -10057
rect 36810 -10175 36816 -10057
rect 36770 -10187 36816 -10175
rect 37298 -10057 37344 -10045
rect 37298 -10175 37304 -10057
rect 37338 -10175 37344 -10057
rect 37298 -10187 37344 -10175
rect 37406 -10057 37452 -10045
rect 37406 -10175 37412 -10057
rect 37446 -10175 37452 -10057
rect 37406 -10187 37452 -10175
rect 37934 -10057 37980 -10045
rect 37934 -10175 37940 -10057
rect 37974 -10175 37980 -10057
rect 37934 -10187 37980 -10175
rect 670 -10228 1093 -10222
rect 670 -10262 705 -10228
rect 1081 -10262 1093 -10228
rect 670 -10268 1093 -10262
rect 1657 -10228 2057 -10222
rect 1657 -10262 1669 -10228
rect 2045 -10230 2057 -10228
rect 2293 -10228 2693 -10222
rect 2293 -10230 2305 -10228
rect 2045 -10262 2060 -10230
rect 1657 -10268 2060 -10262
rect 670 -10490 720 -10268
rect 1420 -10310 1560 -10300
rect 1420 -10430 1430 -10310
rect 1550 -10320 1560 -10310
rect 1660 -10320 2060 -10268
rect 2290 -10262 2305 -10230
rect 2681 -10262 2693 -10228
rect 2290 -10268 2693 -10262
rect 3257 -10228 3657 -10222
rect 3257 -10262 3269 -10228
rect 3645 -10230 3657 -10228
rect 3893 -10228 4293 -10222
rect 3893 -10230 3905 -10228
rect 3645 -10262 3660 -10230
rect 3257 -10268 3660 -10262
rect 2290 -10320 2690 -10268
rect 3020 -10310 3160 -10300
rect 3020 -10320 3030 -10310
rect 1550 -10420 3030 -10320
rect 1550 -10430 1560 -10420
rect 1420 -10440 1560 -10430
rect 1660 -10440 2690 -10420
rect 3020 -10430 3030 -10420
rect 3150 -10320 3160 -10310
rect 3260 -10320 3660 -10268
rect 3890 -10262 3905 -10230
rect 4281 -10262 4293 -10228
rect 3890 -10268 4293 -10262
rect 4857 -10228 5257 -10222
rect 4857 -10262 4869 -10228
rect 5245 -10230 5257 -10228
rect 5493 -10228 5893 -10222
rect 5493 -10230 5505 -10228
rect 5245 -10262 5260 -10230
rect 4857 -10268 5260 -10262
rect 3890 -10320 4290 -10268
rect 4620 -10310 4760 -10300
rect 4620 -10320 4630 -10310
rect 3150 -10420 4630 -10320
rect 3150 -10430 3160 -10420
rect 3020 -10440 3160 -10430
rect 3260 -10440 4290 -10420
rect 4620 -10430 4630 -10420
rect 4750 -10320 4760 -10310
rect 4860 -10320 5260 -10268
rect 5490 -10262 5505 -10230
rect 5881 -10262 5893 -10228
rect 5490 -10268 5893 -10262
rect 6457 -10228 6857 -10222
rect 6457 -10262 6469 -10228
rect 6845 -10230 6857 -10228
rect 7093 -10228 7493 -10222
rect 7093 -10230 7105 -10228
rect 6845 -10262 6860 -10230
rect 6457 -10268 6860 -10262
rect 5490 -10320 5890 -10268
rect 6220 -10310 6360 -10300
rect 6220 -10320 6230 -10310
rect 4750 -10420 6230 -10320
rect 4750 -10430 4760 -10420
rect 4620 -10440 4760 -10430
rect 4860 -10440 5890 -10420
rect 6220 -10430 6230 -10420
rect 6350 -10320 6360 -10310
rect 6460 -10320 6860 -10268
rect 7090 -10262 7105 -10230
rect 7481 -10262 7493 -10228
rect 7090 -10268 7493 -10262
rect 8057 -10228 8457 -10222
rect 8057 -10262 8069 -10228
rect 8445 -10230 8457 -10228
rect 8693 -10228 9093 -10222
rect 8693 -10230 8705 -10228
rect 8445 -10262 8460 -10230
rect 8057 -10268 8460 -10262
rect 7090 -10320 7490 -10268
rect 7820 -10310 7960 -10300
rect 7820 -10320 7830 -10310
rect 6350 -10420 7830 -10320
rect 6350 -10430 6360 -10420
rect 6220 -10440 6360 -10430
rect 6460 -10440 7490 -10420
rect 7820 -10430 7830 -10420
rect 7950 -10320 7960 -10310
rect 8060 -10320 8460 -10268
rect 8690 -10262 8705 -10230
rect 9081 -10262 9093 -10228
rect 8690 -10268 9093 -10262
rect 9657 -10228 10057 -10222
rect 9657 -10262 9669 -10228
rect 10045 -10230 10057 -10228
rect 10293 -10228 10693 -10222
rect 10293 -10230 10305 -10228
rect 10045 -10262 10060 -10230
rect 9657 -10268 10060 -10262
rect 8690 -10320 9090 -10268
rect 9420 -10310 9560 -10300
rect 9420 -10320 9430 -10310
rect 7950 -10420 9430 -10320
rect 7950 -10430 7960 -10420
rect 7820 -10440 7960 -10430
rect 8060 -10440 9090 -10420
rect 9420 -10430 9430 -10420
rect 9550 -10320 9560 -10310
rect 9660 -10320 10060 -10268
rect 10290 -10262 10305 -10230
rect 10681 -10262 10693 -10228
rect 10290 -10268 10693 -10262
rect 11257 -10228 11657 -10222
rect 11257 -10262 11269 -10228
rect 11645 -10262 11657 -10228
rect 11257 -10268 11657 -10262
rect 11893 -10228 12293 -10222
rect 11893 -10262 11905 -10228
rect 12281 -10262 12293 -10228
rect 11893 -10268 12293 -10262
rect 12857 -10228 13257 -10222
rect 12857 -10262 12869 -10228
rect 13245 -10262 13257 -10228
rect 12857 -10268 13257 -10262
rect 13493 -10228 13893 -10222
rect 13493 -10262 13505 -10228
rect 13881 -10262 13893 -10228
rect 13493 -10268 13893 -10262
rect 14457 -10228 14857 -10222
rect 14457 -10262 14469 -10228
rect 14845 -10262 14857 -10228
rect 14457 -10268 14857 -10262
rect 15093 -10228 15493 -10222
rect 15093 -10262 15105 -10228
rect 15481 -10262 15493 -10228
rect 15093 -10268 15493 -10262
rect 16057 -10228 16457 -10222
rect 16057 -10262 16069 -10228
rect 16445 -10262 16457 -10228
rect 16057 -10268 16457 -10262
rect 16693 -10228 17093 -10222
rect 16693 -10262 16705 -10228
rect 17081 -10262 17093 -10228
rect 16693 -10268 17093 -10262
rect 17657 -10228 18057 -10222
rect 17657 -10262 17669 -10228
rect 18045 -10262 18057 -10228
rect 17657 -10268 18057 -10262
rect 18293 -10228 18693 -10222
rect 18293 -10262 18305 -10228
rect 18681 -10262 18693 -10228
rect 18293 -10268 18693 -10262
rect 19257 -10228 19657 -10222
rect 19257 -10262 19269 -10228
rect 19645 -10262 19657 -10228
rect 19257 -10268 19657 -10262
rect 19893 -10228 20293 -10222
rect 19893 -10262 19905 -10228
rect 20281 -10262 20293 -10228
rect 19893 -10268 20293 -10262
rect 20857 -10228 21257 -10222
rect 20857 -10262 20869 -10228
rect 21245 -10262 21257 -10228
rect 20857 -10268 21257 -10262
rect 21493 -10228 21893 -10222
rect 21493 -10262 21505 -10228
rect 21881 -10262 21893 -10228
rect 21493 -10268 21893 -10262
rect 22457 -10228 22857 -10222
rect 22457 -10262 22469 -10228
rect 22845 -10262 22857 -10228
rect 22457 -10268 22857 -10262
rect 23093 -10228 23493 -10222
rect 23093 -10262 23105 -10228
rect 23481 -10262 23493 -10228
rect 23093 -10268 23493 -10262
rect 24057 -10228 24457 -10222
rect 24057 -10262 24069 -10228
rect 24445 -10262 24457 -10228
rect 24057 -10268 24457 -10262
rect 24693 -10228 25093 -10222
rect 24693 -10262 24705 -10228
rect 25081 -10262 25093 -10228
rect 24693 -10268 25093 -10262
rect 25657 -10228 26057 -10222
rect 25657 -10262 25669 -10228
rect 26045 -10262 26057 -10228
rect 25657 -10268 26057 -10262
rect 26293 -10228 26693 -10222
rect 26293 -10262 26305 -10228
rect 26681 -10262 26693 -10228
rect 26293 -10268 26693 -10262
rect 27257 -10228 27657 -10222
rect 27257 -10262 27269 -10228
rect 27645 -10262 27657 -10228
rect 27257 -10268 27657 -10262
rect 27893 -10228 28293 -10222
rect 27893 -10262 27905 -10228
rect 28281 -10262 28293 -10228
rect 27893 -10268 28293 -10262
rect 28857 -10228 29257 -10222
rect 28857 -10262 28869 -10228
rect 29245 -10262 29257 -10228
rect 28857 -10268 29257 -10262
rect 29493 -10228 29893 -10222
rect 29493 -10262 29505 -10228
rect 29881 -10262 29893 -10228
rect 29493 -10268 29893 -10262
rect 30457 -10228 30857 -10222
rect 30457 -10262 30469 -10228
rect 30845 -10262 30857 -10228
rect 30457 -10268 30857 -10262
rect 31093 -10228 31493 -10222
rect 31093 -10262 31105 -10228
rect 31481 -10262 31493 -10228
rect 31093 -10268 31493 -10262
rect 32057 -10228 32457 -10222
rect 32057 -10262 32069 -10228
rect 32445 -10262 32457 -10228
rect 32057 -10268 32457 -10262
rect 32693 -10228 33093 -10222
rect 32693 -10262 32705 -10228
rect 33081 -10262 33093 -10228
rect 32693 -10268 33093 -10262
rect 33657 -10228 34057 -10222
rect 33657 -10262 33669 -10228
rect 34045 -10262 34057 -10228
rect 33657 -10268 34057 -10262
rect 34293 -10228 34693 -10222
rect 34293 -10262 34305 -10228
rect 34681 -10262 34693 -10228
rect 34293 -10268 34693 -10262
rect 35257 -10228 35657 -10222
rect 35257 -10262 35269 -10228
rect 35645 -10262 35657 -10228
rect 35257 -10268 35657 -10262
rect 35893 -10228 36293 -10222
rect 35893 -10262 35905 -10228
rect 36281 -10262 36293 -10228
rect 35893 -10268 36293 -10262
rect 36857 -10228 37257 -10222
rect 36857 -10262 36869 -10228
rect 37245 -10262 37257 -10228
rect 36857 -10268 37257 -10262
rect 37493 -10228 37893 -10222
rect 37493 -10262 37505 -10228
rect 37881 -10262 37893 -10228
rect 37493 -10268 37893 -10262
rect 10290 -10320 10690 -10268
rect 9550 -10420 10690 -10320
rect 15600 -10320 15740 -10310
rect 9550 -10430 9560 -10420
rect 9420 -10440 9560 -10430
rect 9660 -10440 10690 -10420
rect 1660 -10490 2060 -10440
rect 670 -10496 1093 -10490
rect 670 -10530 705 -10496
rect 1081 -10530 1093 -10496
rect 670 -10536 1093 -10530
rect 1657 -10496 2060 -10490
rect 1657 -10530 1669 -10496
rect 2045 -10530 2060 -10496
rect 2290 -10490 2690 -10440
rect 3260 -10490 3660 -10440
rect 2290 -10496 2693 -10490
rect 2290 -10530 2305 -10496
rect 2681 -10530 2693 -10496
rect 1657 -10536 2057 -10530
rect 2293 -10536 2693 -10530
rect 3257 -10496 3660 -10490
rect 3257 -10530 3269 -10496
rect 3645 -10530 3660 -10496
rect 3890 -10490 4290 -10440
rect 4860 -10490 5260 -10440
rect 3890 -10496 4293 -10490
rect 3890 -10530 3905 -10496
rect 4281 -10530 4293 -10496
rect 3257 -10536 3657 -10530
rect 3893 -10536 4293 -10530
rect 4857 -10496 5260 -10490
rect 4857 -10530 4869 -10496
rect 5245 -10530 5260 -10496
rect 5490 -10490 5890 -10440
rect 6460 -10490 6860 -10440
rect 5490 -10496 5893 -10490
rect 5490 -10530 5505 -10496
rect 5881 -10530 5893 -10496
rect 4857 -10536 5257 -10530
rect 5493 -10536 5893 -10530
rect 6457 -10496 6860 -10490
rect 6457 -10530 6469 -10496
rect 6845 -10530 6860 -10496
rect 7090 -10490 7490 -10440
rect 8060 -10490 8460 -10440
rect 7090 -10496 7493 -10490
rect 7090 -10530 7105 -10496
rect 7481 -10530 7493 -10496
rect 6457 -10536 6857 -10530
rect 7093 -10536 7493 -10530
rect 8057 -10496 8460 -10490
rect 8057 -10530 8069 -10496
rect 8445 -10530 8460 -10496
rect 8690 -10490 9090 -10440
rect 9660 -10490 10060 -10440
rect 8690 -10496 9093 -10490
rect 8690 -10530 8705 -10496
rect 9081 -10530 9093 -10496
rect 8057 -10536 8457 -10530
rect 8693 -10536 9093 -10530
rect 9657 -10496 10060 -10490
rect 9657 -10530 9669 -10496
rect 10045 -10530 10060 -10496
rect 10290 -10490 10690 -10440
rect 11020 -10410 11160 -10400
rect 10290 -10496 10693 -10490
rect 10290 -10530 10305 -10496
rect 10681 -10530 10693 -10496
rect 9657 -10536 10057 -10530
rect 10293 -10536 10693 -10530
rect 11020 -10530 11030 -10410
rect 11150 -10490 13890 -10410
rect 15600 -10440 15610 -10320
rect 15730 -10330 15740 -10320
rect 16060 -10330 16450 -10268
rect 16700 -10330 17090 -10268
rect 15730 -10430 17090 -10330
rect 15730 -10440 15740 -10430
rect 15600 -10450 15740 -10440
rect 16060 -10490 16450 -10430
rect 16700 -10490 17090 -10430
rect 17200 -10320 17340 -10310
rect 17200 -10440 17210 -10320
rect 17330 -10330 17340 -10320
rect 17660 -10330 18050 -10268
rect 18300 -10330 18690 -10268
rect 17330 -10430 18690 -10330
rect 17330 -10440 17340 -10430
rect 17200 -10450 17340 -10440
rect 17660 -10490 18050 -10430
rect 18300 -10490 18690 -10430
rect 18800 -10320 18940 -10310
rect 18800 -10440 18810 -10320
rect 18930 -10330 18940 -10320
rect 19260 -10330 19650 -10268
rect 19900 -10330 20290 -10268
rect 18930 -10430 20290 -10330
rect 18930 -10440 18940 -10430
rect 18800 -10450 18940 -10440
rect 19260 -10490 19650 -10430
rect 19900 -10490 20290 -10430
rect 20400 -10320 20540 -10310
rect 20400 -10440 20410 -10320
rect 20530 -10330 20540 -10320
rect 20860 -10330 21250 -10268
rect 21500 -10330 21890 -10268
rect 20530 -10430 21890 -10330
rect 20530 -10440 20540 -10430
rect 20400 -10450 20540 -10440
rect 20860 -10490 21250 -10430
rect 21500 -10490 21890 -10430
rect 22000 -10320 22140 -10310
rect 22000 -10440 22010 -10320
rect 22130 -10330 22140 -10320
rect 22460 -10330 22850 -10268
rect 23100 -10330 23490 -10268
rect 22130 -10430 23490 -10330
rect 22130 -10440 22140 -10430
rect 22000 -10450 22140 -10440
rect 22460 -10490 22850 -10430
rect 23100 -10490 23490 -10430
rect 23600 -10320 23740 -10310
rect 23600 -10440 23610 -10320
rect 23730 -10330 23740 -10320
rect 24060 -10330 24450 -10268
rect 24700 -10330 25090 -10268
rect 23730 -10430 25090 -10330
rect 23730 -10440 23740 -10430
rect 23600 -10450 23740 -10440
rect 24060 -10490 24450 -10430
rect 24700 -10490 25090 -10430
rect 25200 -10320 25340 -10310
rect 25200 -10440 25210 -10320
rect 25330 -10330 25340 -10320
rect 25660 -10330 26050 -10268
rect 26300 -10330 26690 -10268
rect 25330 -10430 26690 -10330
rect 25330 -10440 25340 -10430
rect 25200 -10450 25340 -10440
rect 25660 -10490 26050 -10430
rect 26300 -10490 26690 -10430
rect 26800 -10320 26940 -10310
rect 26800 -10440 26810 -10320
rect 26930 -10330 26940 -10320
rect 27260 -10330 27650 -10268
rect 27900 -10330 28290 -10268
rect 26930 -10430 28290 -10330
rect 26930 -10440 26940 -10430
rect 26800 -10450 26940 -10440
rect 27260 -10490 27650 -10430
rect 27900 -10490 28290 -10430
rect 28400 -10320 28540 -10310
rect 28400 -10440 28410 -10320
rect 28530 -10330 28540 -10320
rect 28860 -10330 29250 -10268
rect 29500 -10330 29890 -10268
rect 28530 -10430 29890 -10330
rect 28530 -10440 28540 -10430
rect 28400 -10450 28540 -10440
rect 28860 -10490 29250 -10430
rect 29500 -10490 29890 -10430
rect 30000 -10320 30140 -10310
rect 30000 -10440 30010 -10320
rect 30130 -10330 30140 -10320
rect 30460 -10330 30850 -10268
rect 31100 -10330 31490 -10268
rect 30130 -10430 31490 -10330
rect 30130 -10440 30140 -10430
rect 30000 -10450 30140 -10440
rect 30460 -10490 30850 -10430
rect 31100 -10490 31490 -10430
rect 31600 -10320 31740 -10310
rect 31600 -10440 31610 -10320
rect 31730 -10330 31740 -10320
rect 32060 -10330 32450 -10268
rect 32700 -10330 33090 -10268
rect 33660 -10330 34050 -10268
rect 34300 -10330 34690 -10268
rect 35260 -10330 35650 -10268
rect 35900 -10330 36290 -10268
rect 31730 -10430 36290 -10330
rect 31730 -10440 31740 -10430
rect 31600 -10450 31740 -10440
rect 32060 -10490 32450 -10430
rect 32700 -10490 33090 -10430
rect 33660 -10490 34050 -10430
rect 34300 -10490 34690 -10430
rect 35260 -10490 35650 -10430
rect 35900 -10490 36290 -10430
rect 11150 -10496 13893 -10490
rect 11150 -10530 11269 -10496
rect 11645 -10530 11905 -10496
rect 12281 -10530 12869 -10496
rect 13245 -10530 13505 -10496
rect 13881 -10530 13893 -10496
rect 57 -11354 490 -11348
rect 57 -11360 69 -11354
rect 20 -11388 69 -11360
rect 445 -11388 490 -11354
rect 20 -11482 490 -11388
rect 1 -11488 490 -11482
rect 670 -11348 720 -10536
rect 11020 -10540 11160 -10530
rect 11257 -10536 11657 -10530
rect 11710 -10584 11840 -10530
rect 11893 -10536 12293 -10530
rect 12857 -10536 13257 -10530
rect 13310 -10584 13440 -10530
rect 13493 -10536 13893 -10530
rect 14457 -10496 14857 -10490
rect 14457 -10530 14469 -10496
rect 14845 -10530 14857 -10496
rect 14457 -10536 14857 -10530
rect 15093 -10496 15493 -10490
rect 15093 -10530 15105 -10496
rect 15481 -10530 15493 -10496
rect 15093 -10536 15493 -10530
rect 16057 -10496 16457 -10490
rect 16057 -10530 16069 -10496
rect 16445 -10530 16457 -10496
rect 16057 -10536 16457 -10530
rect 16693 -10496 17093 -10490
rect 16693 -10530 16705 -10496
rect 17081 -10530 17093 -10496
rect 16693 -10536 17093 -10530
rect 17657 -10496 18057 -10490
rect 17657 -10530 17669 -10496
rect 18045 -10530 18057 -10496
rect 17657 -10536 18057 -10530
rect 18293 -10496 18693 -10490
rect 18293 -10530 18305 -10496
rect 18681 -10530 18693 -10496
rect 18293 -10536 18693 -10530
rect 19257 -10496 19657 -10490
rect 19257 -10530 19269 -10496
rect 19645 -10530 19657 -10496
rect 19257 -10536 19657 -10530
rect 19893 -10496 20293 -10490
rect 19893 -10530 19905 -10496
rect 20281 -10530 20293 -10496
rect 19893 -10536 20293 -10530
rect 20857 -10496 21257 -10490
rect 20857 -10530 20869 -10496
rect 21245 -10530 21257 -10496
rect 20857 -10536 21257 -10530
rect 21493 -10496 21893 -10490
rect 21493 -10530 21505 -10496
rect 21881 -10530 21893 -10496
rect 21493 -10536 21893 -10530
rect 22457 -10496 22857 -10490
rect 22457 -10530 22469 -10496
rect 22845 -10530 22857 -10496
rect 22457 -10536 22857 -10530
rect 23093 -10496 23493 -10490
rect 23093 -10530 23105 -10496
rect 23481 -10530 23493 -10496
rect 23093 -10536 23493 -10530
rect 24057 -10496 24457 -10490
rect 24057 -10530 24069 -10496
rect 24445 -10530 24457 -10496
rect 24057 -10536 24457 -10530
rect 24693 -10496 25093 -10490
rect 24693 -10530 24705 -10496
rect 25081 -10530 25093 -10496
rect 24693 -10536 25093 -10530
rect 25657 -10496 26057 -10490
rect 25657 -10530 25669 -10496
rect 26045 -10530 26057 -10496
rect 25657 -10536 26057 -10530
rect 26293 -10496 26693 -10490
rect 26293 -10530 26305 -10496
rect 26681 -10530 26693 -10496
rect 26293 -10536 26693 -10530
rect 27257 -10496 27657 -10490
rect 27257 -10530 27269 -10496
rect 27645 -10530 27657 -10496
rect 27257 -10536 27657 -10530
rect 27893 -10496 28293 -10490
rect 27893 -10530 27905 -10496
rect 28281 -10530 28293 -10496
rect 27893 -10536 28293 -10530
rect 28857 -10496 29257 -10490
rect 28857 -10530 28869 -10496
rect 29245 -10530 29257 -10496
rect 28857 -10536 29257 -10530
rect 29493 -10496 29893 -10490
rect 29493 -10530 29505 -10496
rect 29881 -10530 29893 -10496
rect 29493 -10536 29893 -10530
rect 30457 -10496 30857 -10490
rect 30457 -10530 30469 -10496
rect 30845 -10530 30857 -10496
rect 30457 -10536 30857 -10530
rect 31093 -10496 31493 -10490
rect 31093 -10530 31105 -10496
rect 31481 -10530 31493 -10496
rect 31093 -10536 31493 -10530
rect 32057 -10496 32457 -10490
rect 32057 -10530 32069 -10496
rect 32445 -10530 32457 -10496
rect 32057 -10536 32457 -10530
rect 32693 -10496 33093 -10490
rect 32693 -10530 32705 -10496
rect 33081 -10530 33093 -10496
rect 32693 -10536 33093 -10530
rect 33657 -10496 34057 -10490
rect 33657 -10530 33669 -10496
rect 34045 -10530 34057 -10496
rect 33657 -10536 34057 -10530
rect 34293 -10496 34693 -10490
rect 34293 -10530 34305 -10496
rect 34681 -10530 34693 -10496
rect 34293 -10536 34693 -10530
rect 35257 -10496 35657 -10490
rect 35257 -10530 35269 -10496
rect 35645 -10530 35657 -10496
rect 35257 -10536 35657 -10530
rect 35893 -10496 36293 -10490
rect 35893 -10530 35905 -10496
rect 36281 -10530 36293 -10496
rect 35893 -10536 36293 -10530
rect 36857 -10496 37257 -10490
rect 36857 -10530 36869 -10496
rect 37245 -10530 37257 -10496
rect 36857 -10536 37257 -10530
rect 37493 -10496 37893 -10490
rect 37493 -10530 37505 -10496
rect 37881 -10530 37893 -10496
rect 37493 -10536 37893 -10530
rect 1134 -10596 1180 -10584
rect 1134 -11288 1140 -10596
rect 1174 -11288 1180 -10596
rect 1134 -11300 1180 -11288
rect 1570 -10596 1616 -10584
rect 1570 -11288 1576 -10596
rect 1610 -11288 1616 -10596
rect 1570 -11300 1616 -11288
rect 2098 -10596 2144 -10584
rect 2098 -11288 2104 -10596
rect 2138 -10600 2144 -10596
rect 2206 -10596 2252 -10584
rect 2206 -10600 2212 -10596
rect 2138 -10610 2212 -10600
rect 2138 -11280 2212 -11270
rect 2138 -11288 2144 -11280
rect 2098 -11300 2144 -11288
rect 2206 -11288 2212 -11280
rect 2246 -11288 2252 -10596
rect 2206 -11300 2252 -11288
rect 2734 -10596 2780 -10584
rect 2734 -11288 2740 -10596
rect 2774 -11288 2780 -10596
rect 2734 -11300 2780 -11288
rect 3170 -10596 3216 -10584
rect 3170 -11288 3176 -10596
rect 3210 -11288 3216 -10596
rect 3170 -11300 3216 -11288
rect 3698 -10596 3744 -10584
rect 3698 -11288 3704 -10596
rect 3738 -10600 3744 -10596
rect 3806 -10596 3852 -10584
rect 3806 -10600 3812 -10596
rect 3738 -10610 3812 -10600
rect 3738 -11280 3812 -11270
rect 3738 -11288 3744 -11280
rect 3698 -11300 3744 -11288
rect 3806 -11288 3812 -11280
rect 3846 -11288 3852 -10596
rect 3806 -11300 3852 -11288
rect 4334 -10596 4380 -10584
rect 4334 -11288 4340 -10596
rect 4374 -11288 4380 -10596
rect 4334 -11300 4380 -11288
rect 4770 -10596 4816 -10584
rect 4770 -11288 4776 -10596
rect 4810 -11288 4816 -10596
rect 4770 -11300 4816 -11288
rect 5298 -10596 5344 -10584
rect 5298 -11288 5304 -10596
rect 5338 -10600 5344 -10596
rect 5406 -10596 5452 -10584
rect 5406 -10600 5412 -10596
rect 5338 -10610 5412 -10600
rect 5338 -11280 5412 -11270
rect 5338 -11288 5344 -11280
rect 5298 -11300 5344 -11288
rect 5406 -11288 5412 -11280
rect 5446 -11288 5452 -10596
rect 5406 -11300 5452 -11288
rect 5934 -10596 5980 -10584
rect 5934 -11288 5940 -10596
rect 5974 -11288 5980 -10596
rect 5934 -11300 5980 -11288
rect 6370 -10596 6416 -10584
rect 6370 -11288 6376 -10596
rect 6410 -11288 6416 -10596
rect 6370 -11300 6416 -11288
rect 6898 -10596 6944 -10584
rect 6898 -11288 6904 -10596
rect 6938 -10600 6944 -10596
rect 7006 -10596 7052 -10584
rect 7006 -10600 7012 -10596
rect 6938 -10610 7012 -10600
rect 6938 -11280 7012 -11270
rect 6938 -11288 6944 -11280
rect 6898 -11300 6944 -11288
rect 7006 -11288 7012 -11280
rect 7046 -11288 7052 -10596
rect 7006 -11300 7052 -11288
rect 7534 -10596 7580 -10584
rect 7534 -11288 7540 -10596
rect 7574 -11288 7580 -10596
rect 7534 -11300 7580 -11288
rect 7970 -10596 8016 -10584
rect 7970 -11288 7976 -10596
rect 8010 -11288 8016 -10596
rect 7970 -11300 8016 -11288
rect 8498 -10596 8544 -10584
rect 8498 -11288 8504 -10596
rect 8538 -10600 8544 -10596
rect 8606 -10596 8652 -10584
rect 8606 -10600 8612 -10596
rect 8538 -10610 8612 -10600
rect 8538 -11280 8612 -11270
rect 8538 -11288 8544 -11280
rect 8498 -11300 8544 -11288
rect 8606 -11288 8612 -11280
rect 8646 -11288 8652 -10596
rect 8606 -11300 8652 -11288
rect 9134 -10596 9180 -10584
rect 9134 -11288 9140 -10596
rect 9174 -11288 9180 -10596
rect 9134 -11300 9180 -11288
rect 9570 -10596 9616 -10584
rect 9570 -11288 9576 -10596
rect 9610 -11288 9616 -10596
rect 9570 -11300 9616 -11288
rect 10098 -10596 10144 -10584
rect 10098 -11288 10104 -10596
rect 10138 -10600 10144 -10596
rect 10206 -10596 10252 -10584
rect 10206 -10600 10212 -10596
rect 10138 -10610 10212 -10600
rect 10138 -11280 10212 -11270
rect 10138 -11288 10144 -11280
rect 10098 -11300 10144 -11288
rect 10206 -11288 10212 -11280
rect 10246 -11288 10252 -10596
rect 10206 -11300 10252 -11288
rect 10734 -10596 10780 -10584
rect 10734 -11288 10740 -10596
rect 10774 -11288 10780 -10596
rect 10734 -11300 10780 -11288
rect 11170 -10596 11216 -10584
rect 11170 -11288 11176 -10596
rect 11210 -11288 11216 -10596
rect 11170 -11300 11216 -11288
rect 11698 -10596 11852 -10584
rect 11698 -11288 11704 -10596
rect 11738 -10610 11812 -10596
rect 11738 -11280 11812 -11270
rect 11738 -11288 11744 -11280
rect 11698 -11300 11744 -11288
rect 11806 -11288 11812 -11280
rect 11846 -11288 11852 -10596
rect 11806 -11300 11852 -11288
rect 12334 -10596 12380 -10584
rect 12334 -11288 12340 -10596
rect 12374 -11288 12380 -10596
rect 12334 -11300 12380 -11288
rect 12770 -10596 12816 -10584
rect 12770 -11288 12776 -10596
rect 12810 -11288 12816 -10596
rect 12770 -11300 12816 -11288
rect 13298 -10596 13452 -10584
rect 13298 -11288 13304 -10596
rect 13338 -10610 13412 -10596
rect 13338 -11280 13412 -11270
rect 13338 -11288 13344 -11280
rect 13298 -11300 13344 -11288
rect 13406 -11288 13412 -11280
rect 13446 -11288 13452 -10596
rect 13406 -11300 13452 -11288
rect 13934 -10596 13980 -10584
rect 13934 -11288 13940 -10596
rect 13974 -11288 13980 -10596
rect 13934 -11300 13980 -11288
rect 14370 -10596 14416 -10584
rect 14370 -11288 14376 -10596
rect 14410 -10880 14416 -10596
rect 14610 -10880 14740 -10536
rect 14898 -10596 14944 -10584
rect 14898 -10880 14904 -10596
rect 14410 -11030 14904 -10880
rect 14410 -11288 14416 -11030
rect 14370 -11300 14416 -11288
rect 14610 -11348 14740 -11030
rect 14898 -11288 14904 -11030
rect 14938 -10880 14944 -10596
rect 15006 -10596 15052 -10584
rect 15006 -10880 15012 -10596
rect 14938 -11030 15012 -10880
rect 14938 -11288 14944 -11030
rect 14898 -11300 14944 -11288
rect 15006 -11288 15012 -11030
rect 15046 -10880 15052 -10596
rect 15220 -10880 15350 -10536
rect 15534 -10596 15580 -10584
rect 15534 -10880 15540 -10596
rect 15046 -11030 15540 -10880
rect 15046 -11288 15052 -11030
rect 15006 -11300 15052 -11288
rect 15220 -11348 15350 -11030
rect 15534 -11288 15540 -11030
rect 15574 -11288 15580 -10596
rect 15534 -11300 15580 -11288
rect 15970 -10596 16016 -10584
rect 15970 -11288 15976 -10596
rect 16010 -11288 16016 -10596
rect 15970 -11300 16016 -11288
rect 16498 -10590 16544 -10584
rect 16606 -10590 16652 -10584
rect 16498 -10596 16652 -10590
rect 16498 -11288 16504 -10596
rect 16538 -10600 16612 -10596
rect 16538 -11288 16612 -11280
rect 16646 -11288 16652 -10596
rect 16498 -11290 16652 -11288
rect 16498 -11300 16544 -11290
rect 16606 -11300 16652 -11290
rect 17134 -10596 17180 -10584
rect 17134 -11288 17140 -10596
rect 17174 -11288 17180 -10596
rect 17134 -11300 17180 -11288
rect 17570 -10596 17616 -10584
rect 17570 -11288 17576 -10596
rect 17610 -11288 17616 -10596
rect 17570 -11300 17616 -11288
rect 18098 -10590 18144 -10584
rect 18206 -10590 18252 -10584
rect 18098 -10596 18252 -10590
rect 18098 -11288 18104 -10596
rect 18138 -10600 18212 -10596
rect 18138 -11288 18212 -11280
rect 18246 -11288 18252 -10596
rect 18098 -11290 18252 -11288
rect 18098 -11300 18144 -11290
rect 18206 -11300 18252 -11290
rect 18734 -10596 18780 -10584
rect 18734 -11288 18740 -10596
rect 18774 -11288 18780 -10596
rect 18734 -11300 18780 -11288
rect 19170 -10596 19216 -10584
rect 19170 -11288 19176 -10596
rect 19210 -11288 19216 -10596
rect 19170 -11300 19216 -11288
rect 19698 -10590 19744 -10584
rect 19806 -10590 19852 -10584
rect 19698 -10596 19852 -10590
rect 19698 -11288 19704 -10596
rect 19738 -10600 19812 -10596
rect 19738 -11288 19812 -11280
rect 19846 -11288 19852 -10596
rect 19698 -11290 19852 -11288
rect 19698 -11300 19744 -11290
rect 19806 -11300 19852 -11290
rect 20334 -10596 20380 -10584
rect 20334 -11288 20340 -10596
rect 20374 -11288 20380 -10596
rect 20334 -11300 20380 -11288
rect 20770 -10596 20816 -10584
rect 20770 -11288 20776 -10596
rect 20810 -11288 20816 -10596
rect 20770 -11300 20816 -11288
rect 21298 -10590 21344 -10584
rect 21406 -10590 21452 -10584
rect 21298 -10596 21452 -10590
rect 21298 -11288 21304 -10596
rect 21338 -10600 21412 -10596
rect 21338 -11288 21412 -11280
rect 21446 -11288 21452 -10596
rect 21298 -11290 21452 -11288
rect 21298 -11300 21344 -11290
rect 21406 -11300 21452 -11290
rect 21934 -10596 21980 -10584
rect 21934 -11288 21940 -10596
rect 21974 -11288 21980 -10596
rect 21934 -11300 21980 -11288
rect 22370 -10596 22416 -10584
rect 22370 -11288 22376 -10596
rect 22410 -11288 22416 -10596
rect 22370 -11300 22416 -11288
rect 22898 -10590 22944 -10584
rect 23006 -10590 23052 -10584
rect 22898 -10596 23052 -10590
rect 22898 -11288 22904 -10596
rect 22938 -10600 23012 -10596
rect 22938 -11288 23012 -11280
rect 23046 -11288 23052 -10596
rect 22898 -11290 23052 -11288
rect 22898 -11300 22944 -11290
rect 23006 -11300 23052 -11290
rect 23534 -10596 23580 -10584
rect 23534 -11288 23540 -10596
rect 23574 -11288 23580 -10596
rect 23534 -11300 23580 -11288
rect 23970 -10596 24016 -10584
rect 23970 -11288 23976 -10596
rect 24010 -11288 24016 -10596
rect 23970 -11300 24016 -11288
rect 24498 -10590 24544 -10584
rect 24606 -10590 24652 -10584
rect 24498 -10596 24652 -10590
rect 24498 -11288 24504 -10596
rect 24538 -10600 24612 -10596
rect 24538 -11288 24612 -11280
rect 24646 -11288 24652 -10596
rect 24498 -11290 24652 -11288
rect 24498 -11300 24544 -11290
rect 24606 -11300 24652 -11290
rect 25134 -10596 25180 -10584
rect 25134 -11288 25140 -10596
rect 25174 -11288 25180 -10596
rect 25134 -11300 25180 -11288
rect 25570 -10596 25616 -10584
rect 25570 -11288 25576 -10596
rect 25610 -11288 25616 -10596
rect 25570 -11300 25616 -11288
rect 26098 -10590 26144 -10584
rect 26206 -10590 26252 -10584
rect 26098 -10596 26252 -10590
rect 26098 -11288 26104 -10596
rect 26138 -10600 26212 -10596
rect 26138 -11288 26212 -11280
rect 26246 -11288 26252 -10596
rect 26098 -11290 26252 -11288
rect 26098 -11300 26144 -11290
rect 26206 -11300 26252 -11290
rect 26734 -10596 26780 -10584
rect 26734 -11288 26740 -10596
rect 26774 -11288 26780 -10596
rect 26734 -11300 26780 -11288
rect 27170 -10596 27216 -10584
rect 27170 -11288 27176 -10596
rect 27210 -11288 27216 -10596
rect 27170 -11300 27216 -11288
rect 27698 -10590 27744 -10584
rect 27806 -10590 27852 -10584
rect 27698 -10596 27852 -10590
rect 27698 -11288 27704 -10596
rect 27738 -10600 27812 -10596
rect 27738 -11288 27812 -11280
rect 27846 -11288 27852 -10596
rect 27698 -11290 27852 -11288
rect 27698 -11300 27744 -11290
rect 27806 -11300 27852 -11290
rect 28334 -10596 28380 -10584
rect 28334 -11288 28340 -10596
rect 28374 -11288 28380 -10596
rect 28334 -11300 28380 -11288
rect 28770 -10596 28816 -10584
rect 28770 -11288 28776 -10596
rect 28810 -11288 28816 -10596
rect 28770 -11300 28816 -11288
rect 29298 -10590 29344 -10584
rect 29406 -10590 29452 -10584
rect 29298 -10596 29452 -10590
rect 29298 -11288 29304 -10596
rect 29338 -10600 29412 -10596
rect 29338 -11288 29412 -11280
rect 29446 -11288 29452 -10596
rect 29298 -11290 29452 -11288
rect 29298 -11300 29344 -11290
rect 29406 -11300 29452 -11290
rect 29934 -10596 29980 -10584
rect 29934 -11288 29940 -10596
rect 29974 -11288 29980 -10596
rect 29934 -11300 29980 -11288
rect 30370 -10596 30416 -10584
rect 30370 -11288 30376 -10596
rect 30410 -11288 30416 -10596
rect 30370 -11300 30416 -11288
rect 30898 -10590 30944 -10584
rect 31006 -10590 31052 -10584
rect 30898 -10596 31052 -10590
rect 30898 -11288 30904 -10596
rect 30938 -10600 31012 -10596
rect 30938 -11288 31012 -11280
rect 31046 -11288 31052 -10596
rect 30898 -11290 31052 -11288
rect 30898 -11300 30944 -11290
rect 31006 -11300 31052 -11290
rect 31534 -10596 31580 -10584
rect 31534 -11288 31540 -10596
rect 31574 -11288 31580 -10596
rect 31534 -11300 31580 -11288
rect 31970 -10596 32016 -10584
rect 31970 -11288 31976 -10596
rect 32010 -11288 32016 -10596
rect 31970 -11300 32016 -11288
rect 32498 -10590 32544 -10584
rect 32606 -10590 32652 -10584
rect 32498 -10596 32652 -10590
rect 32498 -11288 32504 -10596
rect 32538 -10600 32612 -10596
rect 32538 -11288 32544 -11110
rect 32498 -11300 32544 -11288
rect 32606 -11288 32612 -11110
rect 32646 -11288 32652 -10596
rect 32606 -11300 32652 -11288
rect 33134 -10596 33180 -10584
rect 33134 -11288 33140 -10596
rect 33174 -11288 33180 -10596
rect 33134 -11300 33180 -11288
rect 33570 -10596 33616 -10584
rect 33570 -11288 33576 -10596
rect 33610 -11288 33616 -10596
rect 33570 -11300 33616 -11288
rect 34098 -10590 34144 -10584
rect 34206 -10590 34252 -10584
rect 34098 -10596 34252 -10590
rect 34098 -11288 34104 -10596
rect 34138 -10600 34212 -10596
rect 34138 -11288 34144 -11110
rect 34098 -11300 34144 -11288
rect 34206 -11288 34212 -11110
rect 34246 -11288 34252 -10596
rect 34206 -11300 34252 -11288
rect 34734 -10596 34780 -10584
rect 34734 -11288 34740 -10596
rect 34774 -11288 34780 -10596
rect 34734 -11300 34780 -11288
rect 35170 -10596 35216 -10584
rect 35170 -11288 35176 -10596
rect 35210 -11288 35216 -10596
rect 35170 -11300 35216 -11288
rect 35698 -10590 35744 -10584
rect 35806 -10590 35852 -10584
rect 35698 -10596 35852 -10590
rect 35698 -11288 35704 -10596
rect 35738 -10600 35812 -10596
rect 35738 -11288 35744 -11110
rect 35698 -11300 35744 -11288
rect 35806 -11288 35812 -11110
rect 35846 -11288 35852 -10596
rect 35806 -11300 35852 -11288
rect 36334 -10596 36380 -10584
rect 36334 -11288 36340 -10596
rect 36374 -11288 36380 -10596
rect 36334 -11300 36380 -11288
rect 36770 -10596 36816 -10584
rect 36770 -11288 36776 -10596
rect 36810 -11288 36816 -10596
rect 36770 -11300 36816 -11288
rect 37298 -10596 37344 -10584
rect 37298 -11288 37304 -10596
rect 37338 -11288 37344 -10596
rect 37298 -11300 37344 -11288
rect 37406 -10596 37452 -10584
rect 37406 -11288 37412 -10596
rect 37446 -11288 37452 -10596
rect 37406 -11300 37452 -11288
rect 37934 -10596 37980 -10584
rect 37934 -11288 37940 -10596
rect 37974 -11288 37980 -10596
rect 37934 -11300 37980 -11288
rect 35000 -11310 35140 -11300
rect 670 -11354 1093 -11348
rect 670 -11388 705 -11354
rect 1081 -11360 1093 -11354
rect 1657 -11354 2057 -11348
rect 1657 -11360 1669 -11354
rect 1081 -11388 1669 -11360
rect 2045 -11360 2057 -11354
rect 2293 -11354 2693 -11348
rect 2293 -11360 2305 -11354
rect 2045 -11388 2305 -11360
rect 2681 -11360 2693 -11354
rect 3257 -11354 3657 -11348
rect 3257 -11360 3269 -11354
rect 2681 -11388 3269 -11360
rect 3645 -11360 3657 -11354
rect 3893 -11354 4293 -11348
rect 3893 -11360 3905 -11354
rect 3645 -11388 3905 -11360
rect 4281 -11360 4293 -11354
rect 4857 -11354 5257 -11348
rect 4857 -11360 4869 -11354
rect 4281 -11388 4869 -11360
rect 5245 -11360 5257 -11354
rect 5493 -11354 5893 -11348
rect 5493 -11360 5505 -11354
rect 5245 -11388 5505 -11360
rect 5881 -11360 5893 -11354
rect 6457 -11354 6857 -11348
rect 6457 -11360 6469 -11354
rect 5881 -11388 6469 -11360
rect 6845 -11360 6857 -11354
rect 7093 -11354 7493 -11348
rect 7093 -11360 7105 -11354
rect 6845 -11388 7105 -11360
rect 7481 -11360 7493 -11354
rect 8057 -11354 8457 -11348
rect 8057 -11360 8069 -11354
rect 7481 -11388 8069 -11360
rect 8445 -11360 8457 -11354
rect 8693 -11354 9093 -11348
rect 8693 -11360 8705 -11354
rect 8445 -11388 8705 -11360
rect 9081 -11360 9093 -11354
rect 9657 -11354 10057 -11348
rect 9657 -11360 9669 -11354
rect 9081 -11388 9669 -11360
rect 10045 -11360 10057 -11354
rect 10293 -11354 10693 -11348
rect 10293 -11360 10305 -11354
rect 10045 -11388 10305 -11360
rect 10681 -11360 10693 -11354
rect 11257 -11354 11657 -11348
rect 11257 -11360 11269 -11354
rect 10681 -11388 11269 -11360
rect 11645 -11360 11657 -11354
rect 11893 -11354 12293 -11348
rect 11893 -11360 11905 -11354
rect 11645 -11388 11905 -11360
rect 12281 -11360 12293 -11354
rect 12857 -11354 13257 -11348
rect 12857 -11360 12869 -11354
rect 12281 -11388 12869 -11360
rect 13245 -11360 13257 -11354
rect 13493 -11354 13893 -11348
rect 13493 -11360 13505 -11354
rect 13245 -11388 13505 -11360
rect 13881 -11360 13893 -11354
rect 14457 -11354 14857 -11348
rect 14457 -11360 14469 -11354
rect 13881 -11388 14469 -11360
rect 14845 -11360 14857 -11354
rect 15093 -11354 15493 -11348
rect 15093 -11360 15105 -11354
rect 14845 -11388 15105 -11360
rect 15481 -11360 15493 -11354
rect 16057 -11354 16457 -11348
rect 16057 -11360 16069 -11354
rect 15481 -11388 16069 -11360
rect 16445 -11360 16457 -11354
rect 16693 -11354 17093 -11348
rect 16693 -11360 16705 -11354
rect 16445 -11388 16705 -11360
rect 17081 -11360 17093 -11354
rect 17657 -11354 18057 -11348
rect 17657 -11360 17669 -11354
rect 17081 -11388 17669 -11360
rect 18045 -11360 18057 -11354
rect 18293 -11354 18693 -11348
rect 18293 -11360 18305 -11354
rect 18045 -11388 18305 -11360
rect 18681 -11360 18693 -11354
rect 19257 -11354 19657 -11348
rect 19257 -11360 19269 -11354
rect 18681 -11388 19269 -11360
rect 19645 -11360 19657 -11354
rect 19893 -11354 20293 -11348
rect 19893 -11360 19905 -11354
rect 19645 -11388 19905 -11360
rect 20281 -11360 20293 -11354
rect 20857 -11354 21257 -11348
rect 20857 -11360 20869 -11354
rect 20281 -11388 20869 -11360
rect 21245 -11360 21257 -11354
rect 21493 -11354 21893 -11348
rect 21493 -11360 21505 -11354
rect 21245 -11388 21505 -11360
rect 21881 -11360 21893 -11354
rect 22457 -11354 22857 -11348
rect 22457 -11360 22469 -11354
rect 21881 -11388 22469 -11360
rect 22845 -11360 22857 -11354
rect 23093 -11354 23493 -11348
rect 23093 -11360 23105 -11354
rect 22845 -11388 23105 -11360
rect 23481 -11360 23493 -11354
rect 24057 -11354 24457 -11348
rect 24057 -11360 24069 -11354
rect 23481 -11388 24069 -11360
rect 24445 -11360 24457 -11354
rect 24693 -11354 25093 -11348
rect 24693 -11360 24705 -11354
rect 24445 -11388 24705 -11360
rect 25081 -11360 25093 -11354
rect 25657 -11354 26057 -11348
rect 25657 -11360 25669 -11354
rect 25081 -11388 25669 -11360
rect 26045 -11360 26057 -11354
rect 26293 -11354 26693 -11348
rect 26293 -11360 26305 -11354
rect 26045 -11388 26305 -11360
rect 26681 -11360 26693 -11354
rect 27257 -11354 27657 -11348
rect 27257 -11360 27269 -11354
rect 26681 -11388 27269 -11360
rect 27645 -11360 27657 -11354
rect 27893 -11354 28293 -11348
rect 27893 -11360 27905 -11354
rect 27645 -11388 27905 -11360
rect 28281 -11360 28293 -11354
rect 28857 -11354 29257 -11348
rect 28857 -11360 28869 -11354
rect 28281 -11388 28869 -11360
rect 29245 -11360 29257 -11354
rect 29493 -11354 29893 -11348
rect 29493 -11360 29505 -11354
rect 29245 -11388 29505 -11360
rect 29881 -11360 29893 -11354
rect 30457 -11354 30857 -11348
rect 30457 -11360 30469 -11354
rect 29881 -11388 30469 -11360
rect 30845 -11360 30857 -11354
rect 31093 -11354 31493 -11348
rect 31093 -11360 31105 -11354
rect 30845 -11388 31105 -11360
rect 31481 -11360 31493 -11354
rect 32057 -11350 32457 -11348
rect 32693 -11350 33093 -11348
rect 33657 -11350 34057 -11348
rect 34293 -11350 34693 -11348
rect 35000 -11350 35010 -11310
rect 32057 -11354 35010 -11350
rect 31481 -11388 31880 -11360
rect 670 -11488 31880 -11388
rect 32057 -11388 32069 -11354
rect 32445 -11388 32705 -11354
rect 33081 -11388 33669 -11354
rect 34045 -11388 34305 -11354
rect 34681 -11388 35010 -11354
rect 32057 -11394 35010 -11388
rect 32060 -11430 35010 -11394
rect 35130 -11350 35140 -11310
rect 35257 -11350 35657 -11348
rect 35893 -11350 36293 -11348
rect 35130 -11354 36293 -11350
rect 35130 -11388 35269 -11354
rect 35645 -11388 35905 -11354
rect 36281 -11388 36293 -11354
rect 35130 -11394 36293 -11388
rect 36857 -11354 37257 -11348
rect 36857 -11388 36869 -11354
rect 37245 -11388 37257 -11354
rect 36857 -11394 37257 -11388
rect 37493 -11354 37893 -11348
rect 37493 -11388 37505 -11354
rect 37881 -11388 37893 -11354
rect 37493 -11394 37893 -11388
rect 35130 -11430 36290 -11394
rect 32060 -11440 36290 -11430
rect 1 -11500 13 -11488
rect 0 -11522 13 -11500
rect 1137 -11522 1613 -11488
rect 2737 -11522 3213 -11488
rect 4337 -11522 4813 -11488
rect 5937 -11522 6413 -11488
rect 7537 -11522 8013 -11488
rect 9137 -11522 9613 -11488
rect 10737 -11522 11213 -11488
rect 12337 -11522 12813 -11488
rect 13937 -11522 14413 -11488
rect 15537 -11522 16013 -11488
rect 17137 -11522 17613 -11488
rect 18737 -11522 19213 -11488
rect 20337 -11522 20813 -11488
rect 21937 -11522 22413 -11488
rect 23537 -11522 24013 -11488
rect 25137 -11522 25613 -11488
rect 26737 -11522 27213 -11488
rect 28337 -11522 28813 -11488
rect 29937 -11522 30413 -11488
rect 31537 -11500 31880 -11488
rect 32001 -11488 33149 -11482
rect 32001 -11500 32013 -11488
rect 31537 -11522 32013 -11500
rect 33137 -11500 33149 -11488
rect 33601 -11488 34749 -11482
rect 33601 -11500 33613 -11488
rect 33137 -11522 33613 -11500
rect 34737 -11500 34749 -11488
rect 35201 -11488 36349 -11482
rect 35201 -11500 35213 -11488
rect 34737 -11522 35213 -11500
rect 36337 -11500 36349 -11488
rect 36801 -11488 37949 -11482
rect 36801 -11500 36813 -11488
rect 36337 -11522 36813 -11500
rect 37937 -11522 37949 -11488
rect 0 -11620 490 -11522
rect 440 -11764 490 -11620
rect 57 -11770 490 -11764
rect 57 -11804 69 -11770
rect 445 -11804 490 -11770
rect 57 -11810 490 -11804
rect -30 -11857 16 -11845
rect -30 -11975 -24 -11857
rect 10 -11975 16 -11857
rect -30 -11987 16 -11975
rect 440 -12022 490 -11810
rect 670 -11528 37949 -11522
rect 670 -11620 37940 -11528
rect 670 -11764 720 -11620
rect 1200 -11670 1340 -11660
rect 670 -11770 1093 -11764
rect 670 -11804 705 -11770
rect 1081 -11804 1093 -11770
rect 1200 -11790 1210 -11670
rect 1330 -11680 1340 -11670
rect 2800 -11670 2940 -11660
rect 2800 -11680 2810 -11670
rect 1330 -11770 2810 -11680
rect 1330 -11780 1669 -11770
rect 1330 -11790 1340 -11780
rect 1200 -11800 1340 -11790
rect 670 -11810 1093 -11804
rect 1657 -11804 1669 -11780
rect 2045 -11780 2305 -11770
rect 2045 -11804 2057 -11780
rect 1657 -11810 2057 -11804
rect 2293 -11804 2305 -11780
rect 2681 -11780 2810 -11770
rect 2681 -11804 2693 -11780
rect 2800 -11790 2810 -11780
rect 2930 -11680 2940 -11670
rect 4400 -11670 4540 -11660
rect 4400 -11680 4410 -11670
rect 2930 -11770 4410 -11680
rect 2930 -11780 3269 -11770
rect 2930 -11790 2940 -11780
rect 2800 -11800 2940 -11790
rect 2293 -11810 2693 -11804
rect 3257 -11804 3269 -11780
rect 3645 -11780 3905 -11770
rect 3645 -11804 3657 -11780
rect 3257 -11810 3657 -11804
rect 3893 -11804 3905 -11780
rect 4281 -11780 4410 -11770
rect 4281 -11804 4293 -11780
rect 4400 -11790 4410 -11780
rect 4530 -11680 4540 -11670
rect 6000 -11670 6140 -11660
rect 6000 -11680 6010 -11670
rect 4530 -11770 6010 -11680
rect 4530 -11780 4869 -11770
rect 4530 -11790 4540 -11780
rect 4400 -11800 4540 -11790
rect 3893 -11810 4293 -11804
rect 4857 -11804 4869 -11780
rect 5245 -11780 5505 -11770
rect 5245 -11804 5257 -11780
rect 4857 -11810 5257 -11804
rect 5493 -11804 5505 -11780
rect 5881 -11780 6010 -11770
rect 5881 -11804 5893 -11780
rect 6000 -11790 6010 -11780
rect 6130 -11680 6140 -11670
rect 7600 -11670 7740 -11660
rect 7600 -11680 7610 -11670
rect 6130 -11770 7610 -11680
rect 6130 -11780 6469 -11770
rect 6130 -11790 6140 -11780
rect 6000 -11800 6140 -11790
rect 5493 -11810 5893 -11804
rect 6457 -11804 6469 -11780
rect 6845 -11780 7105 -11770
rect 6845 -11804 6857 -11780
rect 6457 -11810 6857 -11804
rect 7093 -11804 7105 -11780
rect 7481 -11780 7610 -11770
rect 7481 -11804 7493 -11780
rect 7600 -11790 7610 -11780
rect 7730 -11680 7740 -11670
rect 9200 -11670 9340 -11660
rect 13300 -11670 13440 -11660
rect 14220 -11670 14360 -11660
rect 15820 -11670 15960 -11660
rect 9200 -11680 9210 -11670
rect 7730 -11770 9210 -11680
rect 7730 -11780 8069 -11770
rect 7730 -11790 7740 -11780
rect 7600 -11800 7740 -11790
rect 7093 -11810 7493 -11804
rect 8057 -11804 8069 -11780
rect 8445 -11780 8705 -11770
rect 8445 -11804 8457 -11780
rect 8057 -11810 8457 -11804
rect 8693 -11804 8705 -11780
rect 9081 -11780 9210 -11770
rect 9081 -11804 9093 -11780
rect 9200 -11790 9210 -11780
rect 9330 -11680 9340 -11670
rect 9330 -11770 10700 -11680
rect 12860 -11764 13310 -11670
rect 9330 -11780 9669 -11770
rect 9330 -11790 9340 -11780
rect 9200 -11800 9340 -11790
rect 8693 -11810 9093 -11804
rect 9657 -11804 9669 -11780
rect 10045 -11780 10305 -11770
rect 10045 -11804 10057 -11780
rect 9657 -11810 10057 -11804
rect 10293 -11804 10305 -11780
rect 10681 -11780 10700 -11770
rect 11257 -11770 11657 -11764
rect 10681 -11804 10693 -11780
rect 10293 -11810 10693 -11804
rect 11257 -11804 11269 -11770
rect 11645 -11804 11657 -11770
rect 11257 -11810 11657 -11804
rect 11893 -11770 12293 -11764
rect 11893 -11804 11905 -11770
rect 12281 -11804 12293 -11770
rect 11893 -11810 12293 -11804
rect 12857 -11770 13310 -11764
rect 12857 -11804 12869 -11770
rect 13245 -11790 13310 -11770
rect 13430 -11770 14230 -11670
rect 13430 -11790 13505 -11770
rect 13245 -11800 13505 -11790
rect 13245 -11804 13257 -11800
rect 12857 -11810 13257 -11804
rect 13493 -11804 13505 -11800
rect 13881 -11790 14230 -11770
rect 14350 -11764 15490 -11670
rect 14350 -11770 15493 -11764
rect 14350 -11790 14469 -11770
rect 13881 -11800 14469 -11790
rect 13881 -11804 13893 -11800
rect 13493 -11810 13893 -11804
rect 14457 -11804 14469 -11800
rect 14845 -11800 15105 -11770
rect 14845 -11804 14857 -11800
rect 14457 -11810 14857 -11804
rect 15093 -11804 15105 -11800
rect 15481 -11804 15493 -11770
rect 15820 -11790 15830 -11670
rect 15950 -11700 15960 -11670
rect 17420 -11670 17560 -11660
rect 15950 -11764 17090 -11700
rect 15950 -11770 17093 -11764
rect 15950 -11790 16069 -11770
rect 15820 -11800 16069 -11790
rect 15093 -11810 15493 -11804
rect 16057 -11804 16069 -11800
rect 16445 -11800 16705 -11770
rect 16445 -11804 16457 -11800
rect 16057 -11810 16457 -11804
rect 16693 -11804 16705 -11800
rect 17081 -11804 17093 -11770
rect 17420 -11790 17430 -11670
rect 17550 -11700 17560 -11670
rect 19020 -11670 19160 -11660
rect 17550 -11764 18690 -11700
rect 17550 -11770 18693 -11764
rect 17550 -11790 17669 -11770
rect 17420 -11800 17669 -11790
rect 16693 -11810 17093 -11804
rect 17657 -11804 17669 -11800
rect 18045 -11800 18305 -11770
rect 18045 -11804 18057 -11800
rect 17657 -11810 18057 -11804
rect 18293 -11804 18305 -11800
rect 18681 -11804 18693 -11770
rect 19020 -11790 19030 -11670
rect 19150 -11700 19160 -11670
rect 20620 -11670 20760 -11660
rect 19150 -11764 20290 -11700
rect 19150 -11770 20293 -11764
rect 19150 -11790 19269 -11770
rect 19020 -11800 19269 -11790
rect 18293 -11810 18693 -11804
rect 19257 -11804 19269 -11800
rect 19645 -11800 19905 -11770
rect 19645 -11804 19657 -11800
rect 19257 -11810 19657 -11804
rect 19893 -11804 19905 -11800
rect 20281 -11804 20293 -11770
rect 20620 -11790 20630 -11670
rect 20750 -11700 20760 -11670
rect 22220 -11670 22360 -11660
rect 20750 -11764 21890 -11700
rect 20750 -11770 21893 -11764
rect 20750 -11790 20869 -11770
rect 20620 -11800 20869 -11790
rect 19893 -11810 20293 -11804
rect 20857 -11804 20869 -11800
rect 21245 -11800 21505 -11770
rect 21245 -11804 21257 -11800
rect 20857 -11810 21257 -11804
rect 21493 -11804 21505 -11800
rect 21881 -11804 21893 -11770
rect 22220 -11790 22230 -11670
rect 22350 -11700 22360 -11670
rect 23820 -11670 23960 -11660
rect 22350 -11764 23490 -11700
rect 22350 -11770 23493 -11764
rect 22350 -11790 22469 -11770
rect 22220 -11800 22469 -11790
rect 21493 -11810 21893 -11804
rect 22457 -11804 22469 -11800
rect 22845 -11800 23105 -11770
rect 22845 -11804 22857 -11800
rect 22457 -11810 22857 -11804
rect 23093 -11804 23105 -11800
rect 23481 -11804 23493 -11770
rect 23820 -11790 23830 -11670
rect 23950 -11700 23960 -11670
rect 25420 -11670 25560 -11660
rect 23950 -11764 25090 -11700
rect 23950 -11770 25093 -11764
rect 23950 -11790 24069 -11770
rect 23820 -11800 24069 -11790
rect 23093 -11810 23493 -11804
rect 24057 -11804 24069 -11800
rect 24445 -11800 24705 -11770
rect 24445 -11804 24457 -11800
rect 24057 -11810 24457 -11804
rect 24693 -11804 24705 -11800
rect 25081 -11804 25093 -11770
rect 25420 -11790 25430 -11670
rect 25550 -11700 25560 -11670
rect 27020 -11670 27160 -11660
rect 25550 -11764 26680 -11700
rect 25550 -11770 26693 -11764
rect 25550 -11790 25669 -11770
rect 25420 -11800 25669 -11790
rect 24693 -11810 25093 -11804
rect 25657 -11804 25669 -11800
rect 26045 -11800 26305 -11770
rect 26045 -11804 26057 -11800
rect 25657 -11810 26057 -11804
rect 26293 -11804 26305 -11800
rect 26681 -11804 26693 -11770
rect 27020 -11790 27030 -11670
rect 27150 -11700 27160 -11670
rect 28620 -11670 28760 -11660
rect 27150 -11764 28290 -11700
rect 27150 -11770 28293 -11764
rect 27150 -11790 27269 -11770
rect 27020 -11800 27269 -11790
rect 26293 -11810 26693 -11804
rect 27257 -11804 27269 -11800
rect 27645 -11800 27905 -11770
rect 27645 -11804 27657 -11800
rect 27257 -11810 27657 -11804
rect 27893 -11804 27905 -11800
rect 28281 -11804 28293 -11770
rect 28620 -11790 28630 -11670
rect 28750 -11700 28760 -11670
rect 30220 -11670 30360 -11660
rect 28750 -11764 29890 -11700
rect 28750 -11770 29893 -11764
rect 28750 -11790 28869 -11770
rect 28620 -11800 28869 -11790
rect 27893 -11810 28293 -11804
rect 28857 -11804 28869 -11800
rect 29245 -11800 29505 -11770
rect 29245 -11804 29257 -11800
rect 28857 -11810 29257 -11804
rect 29493 -11804 29505 -11800
rect 29881 -11804 29893 -11770
rect 30220 -11790 30230 -11670
rect 30350 -11700 30360 -11670
rect 31820 -11670 31960 -11660
rect 30350 -11764 31490 -11700
rect 30350 -11770 31493 -11764
rect 30350 -11790 30469 -11770
rect 30220 -11800 30469 -11790
rect 29493 -11810 29893 -11804
rect 30457 -11804 30469 -11800
rect 30845 -11800 31105 -11770
rect 30845 -11804 30857 -11800
rect 30457 -11810 30857 -11804
rect 31093 -11804 31105 -11800
rect 31481 -11804 31493 -11770
rect 31820 -11790 31830 -11670
rect 31950 -11700 31960 -11670
rect 34800 -11670 34940 -11660
rect 34800 -11700 34810 -11670
rect 31950 -11770 34810 -11700
rect 31950 -11790 32069 -11770
rect 31820 -11800 32069 -11790
rect 31093 -11810 31493 -11804
rect 32057 -11804 32069 -11800
rect 32445 -11800 32705 -11770
rect 32445 -11804 32457 -11800
rect 32057 -11810 32457 -11804
rect 32693 -11804 32705 -11800
rect 33081 -11800 33669 -11770
rect 33081 -11804 33093 -11800
rect 32693 -11810 33093 -11804
rect 33657 -11804 33669 -11800
rect 34045 -11800 34305 -11770
rect 34045 -11804 34057 -11800
rect 33657 -11810 34057 -11804
rect 34293 -11804 34305 -11800
rect 34681 -11790 34810 -11770
rect 34930 -11700 34940 -11670
rect 34930 -11764 36280 -11700
rect 34930 -11770 36293 -11764
rect 34930 -11790 35269 -11770
rect 34681 -11800 35269 -11790
rect 34681 -11804 34693 -11800
rect 34293 -11810 34693 -11804
rect 35257 -11804 35269 -11800
rect 35645 -11800 35905 -11770
rect 35645 -11804 35657 -11800
rect 35257 -11810 35657 -11804
rect 35893 -11804 35905 -11800
rect 36281 -11804 36293 -11770
rect 35893 -11810 36293 -11804
rect 36857 -11770 37257 -11764
rect 36857 -11804 36869 -11770
rect 37245 -11804 37257 -11770
rect 36857 -11810 37257 -11804
rect 37493 -11770 37893 -11764
rect 37493 -11804 37505 -11770
rect 37881 -11804 37893 -11770
rect 37493 -11810 37893 -11804
rect 57 -12028 490 -12022
rect 57 -12062 69 -12028
rect 445 -12062 490 -12028
rect 57 -12068 490 -12062
rect 440 -12290 490 -12068
rect 57 -12296 490 -12290
rect 57 -12330 69 -12296
rect 445 -12330 490 -12296
rect 57 -12336 490 -12330
rect -30 -12396 16 -12384
rect -30 -13088 -24 -12396
rect 10 -13088 16 -12396
rect -30 -13100 16 -13088
rect 440 -13148 490 -12336
rect 670 -12022 720 -11810
rect 1134 -11857 1180 -11845
rect 1134 -11975 1140 -11857
rect 1174 -11975 1180 -11857
rect 1570 -11857 1616 -11845
rect 1570 -11860 1576 -11857
rect 1134 -11987 1180 -11975
rect 1560 -11975 1576 -11860
rect 1610 -11860 1616 -11857
rect 2098 -11857 2144 -11845
rect 2098 -11860 2104 -11857
rect 1610 -11975 2104 -11860
rect 2138 -11860 2144 -11857
rect 2206 -11857 2252 -11845
rect 2206 -11860 2212 -11857
rect 2138 -11975 2212 -11860
rect 2246 -11860 2252 -11857
rect 2734 -11857 2780 -11845
rect 2734 -11860 2740 -11857
rect 2246 -11975 2740 -11860
rect 2774 -11860 2780 -11857
rect 3170 -11857 3216 -11845
rect 3170 -11860 3176 -11857
rect 2774 -11975 3176 -11860
rect 3210 -11860 3216 -11857
rect 3698 -11857 3744 -11845
rect 3698 -11860 3704 -11857
rect 3210 -11975 3704 -11860
rect 3738 -11860 3744 -11857
rect 3806 -11857 3852 -11845
rect 3806 -11860 3812 -11857
rect 3738 -11975 3812 -11860
rect 3846 -11860 3852 -11857
rect 4334 -11857 4380 -11845
rect 4334 -11860 4340 -11857
rect 3846 -11975 4340 -11860
rect 4374 -11860 4380 -11857
rect 4770 -11857 4816 -11845
rect 4770 -11860 4776 -11857
rect 4374 -11975 4776 -11860
rect 4810 -11860 4816 -11857
rect 5298 -11857 5344 -11845
rect 5298 -11860 5304 -11857
rect 4810 -11975 5304 -11860
rect 5338 -11860 5344 -11857
rect 5406 -11857 5452 -11845
rect 5406 -11860 5412 -11857
rect 5338 -11975 5412 -11860
rect 5446 -11860 5452 -11857
rect 5934 -11857 5980 -11845
rect 5934 -11860 5940 -11857
rect 5446 -11975 5940 -11860
rect 5974 -11860 5980 -11857
rect 6370 -11857 6416 -11845
rect 6370 -11860 6376 -11857
rect 5974 -11975 6376 -11860
rect 6410 -11860 6416 -11857
rect 6898 -11857 6944 -11845
rect 6898 -11860 6904 -11857
rect 6410 -11975 6904 -11860
rect 6938 -11860 6944 -11857
rect 7006 -11857 7052 -11845
rect 7006 -11860 7012 -11857
rect 6938 -11975 7012 -11860
rect 7046 -11860 7052 -11857
rect 7534 -11857 7580 -11845
rect 7534 -11860 7540 -11857
rect 7046 -11975 7540 -11860
rect 7574 -11860 7580 -11857
rect 7970 -11857 8016 -11845
rect 7970 -11860 7976 -11857
rect 7574 -11975 7976 -11860
rect 8010 -11860 8016 -11857
rect 8498 -11857 8544 -11845
rect 8498 -11860 8504 -11857
rect 8010 -11975 8504 -11860
rect 8538 -11860 8544 -11857
rect 8606 -11857 8652 -11845
rect 8606 -11860 8612 -11857
rect 8538 -11975 8612 -11860
rect 8646 -11860 8652 -11857
rect 9134 -11857 9180 -11845
rect 9134 -11860 9140 -11857
rect 8646 -11975 9140 -11860
rect 9174 -11860 9180 -11857
rect 9570 -11857 9616 -11845
rect 9570 -11860 9576 -11857
rect 9174 -11975 9576 -11860
rect 9610 -11860 9616 -11857
rect 10098 -11857 10144 -11845
rect 10098 -11860 10104 -11857
rect 9610 -11975 10104 -11860
rect 10138 -11860 10144 -11857
rect 10206 -11857 10252 -11845
rect 10206 -11860 10212 -11857
rect 10138 -11975 10212 -11860
rect 10246 -11860 10252 -11857
rect 10734 -11850 10780 -11845
rect 10734 -11857 10940 -11850
rect 10734 -11860 10740 -11857
rect 10246 -11975 10740 -11860
rect 10774 -11860 10940 -11857
rect 11170 -11857 11216 -11845
rect 11170 -11860 11176 -11857
rect 10774 -11975 10810 -11860
rect 1560 -11980 10810 -11975
rect 10930 -11975 11176 -11860
rect 11210 -11860 11216 -11857
rect 11400 -11860 11520 -11810
rect 11698 -11857 11744 -11845
rect 11698 -11860 11704 -11857
rect 11210 -11975 11704 -11860
rect 11738 -11860 11744 -11857
rect 11806 -11857 11852 -11845
rect 11806 -11860 11812 -11857
rect 11738 -11975 11812 -11860
rect 11846 -11860 11852 -11857
rect 12040 -11860 12160 -11810
rect 12334 -11857 12380 -11845
rect 12334 -11860 12340 -11857
rect 11846 -11975 12340 -11860
rect 12374 -11860 12380 -11857
rect 12770 -11857 12816 -11845
rect 12770 -11860 12776 -11857
rect 12374 -11975 12776 -11860
rect 12810 -11860 12816 -11857
rect 13298 -11857 13344 -11845
rect 13298 -11860 13304 -11857
rect 12810 -11975 13304 -11860
rect 13338 -11860 13344 -11857
rect 13406 -11857 13452 -11845
rect 13406 -11860 13412 -11857
rect 13338 -11975 13412 -11860
rect 13446 -11860 13452 -11857
rect 13934 -11857 13980 -11845
rect 13934 -11860 13940 -11857
rect 13446 -11975 13940 -11860
rect 13974 -11860 13980 -11857
rect 14370 -11857 14416 -11845
rect 14370 -11860 14376 -11857
rect 13974 -11975 14376 -11860
rect 14410 -11860 14416 -11857
rect 14898 -11857 14944 -11845
rect 14898 -11860 14904 -11857
rect 14410 -11975 14904 -11860
rect 14938 -11860 14944 -11857
rect 15006 -11857 15052 -11845
rect 15006 -11860 15012 -11857
rect 14938 -11975 15012 -11860
rect 15046 -11860 15052 -11857
rect 15534 -11857 15580 -11845
rect 15534 -11860 15540 -11857
rect 15046 -11975 15540 -11860
rect 15574 -11860 15580 -11857
rect 15970 -11857 16016 -11845
rect 15970 -11860 15976 -11857
rect 15574 -11975 15976 -11860
rect 16010 -11860 16016 -11857
rect 16498 -11857 16544 -11845
rect 16498 -11860 16504 -11857
rect 16010 -11975 16504 -11860
rect 16538 -11860 16544 -11857
rect 16606 -11857 16652 -11845
rect 16606 -11860 16612 -11857
rect 16538 -11975 16612 -11860
rect 16646 -11860 16652 -11857
rect 17134 -11857 17180 -11845
rect 17134 -11860 17140 -11857
rect 16646 -11975 17140 -11860
rect 17174 -11860 17180 -11857
rect 17570 -11857 17616 -11845
rect 17570 -11860 17576 -11857
rect 17174 -11975 17576 -11860
rect 17610 -11860 17616 -11857
rect 18098 -11857 18144 -11845
rect 18098 -11860 18104 -11857
rect 17610 -11975 18104 -11860
rect 18138 -11860 18144 -11857
rect 18206 -11857 18252 -11845
rect 18206 -11860 18212 -11857
rect 18138 -11975 18212 -11860
rect 18246 -11860 18252 -11857
rect 18734 -11857 18780 -11845
rect 18734 -11860 18740 -11857
rect 18246 -11975 18740 -11860
rect 18774 -11860 18780 -11857
rect 19170 -11857 19216 -11845
rect 19170 -11860 19176 -11857
rect 18774 -11975 19176 -11860
rect 19210 -11860 19216 -11857
rect 19698 -11857 19744 -11845
rect 19698 -11860 19704 -11857
rect 19210 -11975 19704 -11860
rect 19738 -11860 19744 -11857
rect 19806 -11857 19852 -11845
rect 19806 -11860 19812 -11857
rect 19738 -11975 19812 -11860
rect 19846 -11860 19852 -11857
rect 20334 -11857 20380 -11845
rect 20334 -11860 20340 -11857
rect 19846 -11975 20340 -11860
rect 20374 -11860 20380 -11857
rect 20770 -11857 20816 -11845
rect 20770 -11860 20776 -11857
rect 20374 -11975 20776 -11860
rect 20810 -11860 20816 -11857
rect 21298 -11857 21344 -11845
rect 21298 -11860 21304 -11857
rect 20810 -11975 21304 -11860
rect 21338 -11860 21344 -11857
rect 21406 -11857 21452 -11845
rect 21406 -11860 21412 -11857
rect 21338 -11975 21412 -11860
rect 21446 -11860 21452 -11857
rect 21934 -11857 21980 -11845
rect 21934 -11860 21940 -11857
rect 21446 -11975 21940 -11860
rect 21974 -11860 21980 -11857
rect 22370 -11857 22416 -11845
rect 22370 -11860 22376 -11857
rect 21974 -11975 22376 -11860
rect 22410 -11860 22416 -11857
rect 22898 -11857 22944 -11845
rect 22898 -11860 22904 -11857
rect 22410 -11975 22904 -11860
rect 22938 -11860 22944 -11857
rect 23006 -11857 23052 -11845
rect 23006 -11860 23012 -11857
rect 22938 -11975 23012 -11860
rect 23046 -11860 23052 -11857
rect 23534 -11857 23580 -11845
rect 23534 -11860 23540 -11857
rect 23046 -11975 23540 -11860
rect 23574 -11860 23580 -11857
rect 23970 -11857 24016 -11845
rect 23970 -11860 23976 -11857
rect 23574 -11975 23976 -11860
rect 24010 -11860 24016 -11857
rect 24498 -11857 24544 -11845
rect 24498 -11860 24504 -11857
rect 24010 -11975 24504 -11860
rect 24538 -11860 24544 -11857
rect 24606 -11857 24652 -11845
rect 24606 -11860 24612 -11857
rect 24538 -11975 24612 -11860
rect 24646 -11860 24652 -11857
rect 25134 -11857 25180 -11845
rect 25134 -11860 25140 -11857
rect 24646 -11975 25140 -11860
rect 25174 -11860 25180 -11857
rect 25570 -11857 25616 -11845
rect 25570 -11860 25576 -11857
rect 25174 -11975 25576 -11860
rect 25610 -11860 25616 -11857
rect 26098 -11857 26144 -11845
rect 26098 -11860 26104 -11857
rect 25610 -11975 26104 -11860
rect 26138 -11860 26144 -11857
rect 26206 -11857 26252 -11845
rect 26206 -11860 26212 -11857
rect 26138 -11975 26212 -11860
rect 26246 -11860 26252 -11857
rect 26734 -11857 26780 -11845
rect 26734 -11860 26740 -11857
rect 26246 -11975 26740 -11860
rect 26774 -11860 26780 -11857
rect 27170 -11857 27216 -11845
rect 27170 -11860 27176 -11857
rect 26774 -11975 27176 -11860
rect 27210 -11860 27216 -11857
rect 27698 -11857 27744 -11845
rect 27698 -11860 27704 -11857
rect 27210 -11975 27704 -11860
rect 27738 -11860 27744 -11857
rect 27806 -11857 27852 -11845
rect 27806 -11860 27812 -11857
rect 27738 -11975 27812 -11860
rect 27846 -11860 27852 -11857
rect 28334 -11857 28380 -11845
rect 28334 -11860 28340 -11857
rect 27846 -11975 28340 -11860
rect 28374 -11860 28380 -11857
rect 28770 -11857 28816 -11845
rect 28770 -11860 28776 -11857
rect 28374 -11975 28776 -11860
rect 28810 -11860 28816 -11857
rect 29298 -11857 29344 -11845
rect 29298 -11860 29304 -11857
rect 28810 -11975 29304 -11860
rect 29338 -11860 29344 -11857
rect 29406 -11857 29452 -11845
rect 29406 -11860 29412 -11857
rect 29338 -11975 29412 -11860
rect 29446 -11860 29452 -11857
rect 29934 -11857 29980 -11845
rect 29934 -11860 29940 -11857
rect 29446 -11975 29940 -11860
rect 29974 -11860 29980 -11857
rect 30370 -11857 30416 -11837
rect 30370 -11860 30376 -11857
rect 29974 -11975 30376 -11860
rect 30410 -11860 30416 -11857
rect 30898 -11857 30944 -11837
rect 30898 -11860 30904 -11857
rect 30410 -11975 30904 -11860
rect 30938 -11860 30944 -11857
rect 31006 -11857 31052 -11837
rect 31006 -11860 31012 -11857
rect 30938 -11975 31012 -11860
rect 31046 -11860 31052 -11857
rect 31534 -11857 31580 -11845
rect 31534 -11860 31540 -11857
rect 31046 -11975 31540 -11860
rect 31574 -11860 31580 -11857
rect 31970 -11857 32016 -11845
rect 31970 -11860 31976 -11857
rect 31574 -11975 31976 -11860
rect 32010 -11860 32016 -11857
rect 32498 -11857 32544 -11845
rect 32498 -11860 32504 -11857
rect 32010 -11975 32504 -11860
rect 32538 -11860 32544 -11857
rect 32606 -11857 32652 -11845
rect 32606 -11860 32612 -11857
rect 32538 -11975 32612 -11860
rect 32646 -11860 32652 -11857
rect 33134 -11857 33180 -11845
rect 33134 -11860 33140 -11857
rect 32646 -11975 33140 -11860
rect 33174 -11860 33180 -11857
rect 33570 -11857 33616 -11845
rect 33570 -11860 33576 -11857
rect 33174 -11975 33576 -11860
rect 33610 -11860 33616 -11857
rect 34098 -11857 34144 -11845
rect 34098 -11860 34104 -11857
rect 33610 -11975 34104 -11860
rect 34138 -11860 34144 -11857
rect 34206 -11857 34252 -11845
rect 34206 -11860 34212 -11857
rect 34138 -11975 34212 -11860
rect 34246 -11860 34252 -11857
rect 34734 -11857 34780 -11845
rect 34734 -11860 34740 -11857
rect 34246 -11975 34740 -11860
rect 34774 -11860 34780 -11857
rect 35170 -11857 35216 -11845
rect 35170 -11860 35176 -11857
rect 34774 -11975 35176 -11860
rect 35210 -11860 35216 -11857
rect 35698 -11857 35744 -11845
rect 35698 -11860 35704 -11857
rect 35210 -11975 35704 -11860
rect 35738 -11860 35744 -11857
rect 35806 -11857 35852 -11845
rect 35806 -11860 35812 -11857
rect 35738 -11975 35812 -11860
rect 35846 -11860 35852 -11857
rect 36334 -11857 36380 -11845
rect 36334 -11860 36340 -11857
rect 35846 -11975 36340 -11860
rect 36374 -11975 36380 -11857
rect 10930 -11980 36380 -11975
rect 1570 -11987 1616 -11980
rect 2098 -11987 2144 -11980
rect 2206 -11987 2252 -11980
rect 2734 -11987 2780 -11980
rect 3170 -11987 3216 -11980
rect 3698 -11987 3744 -11980
rect 3806 -11987 3852 -11980
rect 4334 -11987 4380 -11980
rect 4770 -11987 4816 -11980
rect 5298 -11987 5344 -11980
rect 5406 -11987 5452 -11980
rect 5934 -11987 5980 -11980
rect 6370 -11987 6416 -11980
rect 6898 -11987 6944 -11980
rect 7006 -11987 7052 -11980
rect 7534 -11987 7580 -11980
rect 7970 -11987 8016 -11980
rect 8498 -11987 8544 -11980
rect 8606 -11987 8652 -11980
rect 9134 -11987 9180 -11980
rect 9570 -11987 9616 -11980
rect 10098 -11987 10144 -11980
rect 10206 -11987 10252 -11980
rect 10734 -11987 10940 -11980
rect 11170 -11987 11216 -11980
rect 10750 -11990 10940 -11987
rect 11400 -12022 11520 -11980
rect 11698 -11987 11744 -11980
rect 11806 -11987 11852 -11980
rect 12040 -12022 12160 -11980
rect 12334 -11987 12380 -11980
rect 12770 -11987 12816 -11980
rect 13298 -11987 13344 -11980
rect 13406 -11987 13452 -11980
rect 13934 -11987 13980 -11980
rect 14370 -11987 14416 -11980
rect 14898 -11987 14944 -11980
rect 15006 -11987 15052 -11980
rect 15534 -11987 15580 -11980
rect 15970 -11987 16016 -11980
rect 16498 -11987 16544 -11980
rect 16606 -11987 16652 -11980
rect 17134 -11987 17180 -11980
rect 17570 -11987 17616 -11980
rect 18098 -11987 18144 -11980
rect 18206 -11987 18252 -11980
rect 18734 -11987 18780 -11980
rect 19170 -11987 19216 -11980
rect 19698 -11987 19744 -11980
rect 19806 -11987 19852 -11980
rect 20334 -11987 20380 -11980
rect 20770 -11987 20816 -11980
rect 21298 -11987 21344 -11980
rect 21406 -11987 21452 -11980
rect 21934 -11987 21980 -11980
rect 22370 -11987 22416 -11980
rect 22898 -11987 22944 -11980
rect 23006 -11987 23052 -11980
rect 23534 -11987 23580 -11980
rect 23970 -11987 24016 -11980
rect 24498 -11987 24544 -11980
rect 24606 -11987 24652 -11980
rect 25134 -11987 25180 -11980
rect 25570 -11987 25616 -11980
rect 26098 -11987 26144 -11980
rect 26206 -11987 26252 -11980
rect 26734 -11987 26780 -11980
rect 27170 -11987 27216 -11980
rect 27698 -11987 27744 -11980
rect 27806 -11987 27852 -11980
rect 28334 -11987 28380 -11980
rect 28770 -11987 28816 -11980
rect 29298 -11987 29344 -11980
rect 29406 -11987 29452 -11980
rect 29934 -11987 29980 -11980
rect 30370 -11995 30416 -11980
rect 30898 -11995 30944 -11980
rect 31006 -11995 31052 -11980
rect 31534 -11987 31580 -11980
rect 31970 -11987 32016 -11980
rect 32498 -11987 32544 -11980
rect 32606 -11987 32652 -11980
rect 33134 -11987 33180 -11980
rect 33570 -11987 33616 -11980
rect 34098 -11987 34144 -11980
rect 34206 -11987 34252 -11980
rect 34734 -11987 34780 -11980
rect 35170 -11987 35216 -11980
rect 35698 -11987 35744 -11980
rect 35806 -11987 35852 -11980
rect 36334 -11987 36380 -11980
rect 36770 -11857 36816 -11845
rect 36770 -11975 36776 -11857
rect 36810 -11975 36816 -11857
rect 36770 -11987 36816 -11975
rect 37298 -11857 37344 -11845
rect 37298 -11975 37304 -11857
rect 37338 -11975 37344 -11857
rect 37298 -11987 37344 -11975
rect 37406 -11857 37452 -11845
rect 37406 -11975 37412 -11857
rect 37446 -11975 37452 -11857
rect 37406 -11987 37452 -11975
rect 37934 -11857 37980 -11845
rect 37934 -11975 37940 -11857
rect 37974 -11975 37980 -11857
rect 37934 -11987 37980 -11975
rect 670 -12028 1093 -12022
rect 670 -12062 705 -12028
rect 1081 -12062 1093 -12028
rect 670 -12068 1093 -12062
rect 1657 -12028 2057 -12022
rect 1657 -12062 1669 -12028
rect 2045 -12030 2057 -12028
rect 2293 -12028 2693 -12022
rect 2293 -12030 2305 -12028
rect 2045 -12062 2060 -12030
rect 1657 -12068 2060 -12062
rect 670 -12290 720 -12068
rect 1420 -12110 1560 -12100
rect 1420 -12230 1430 -12110
rect 1550 -12120 1560 -12110
rect 1660 -12120 2060 -12068
rect 2290 -12062 2305 -12030
rect 2681 -12062 2693 -12028
rect 2290 -12068 2693 -12062
rect 3257 -12028 3657 -12022
rect 3257 -12062 3269 -12028
rect 3645 -12030 3657 -12028
rect 3893 -12028 4293 -12022
rect 3893 -12030 3905 -12028
rect 3645 -12062 3660 -12030
rect 3257 -12068 3660 -12062
rect 2290 -12120 2690 -12068
rect 3020 -12110 3160 -12100
rect 3020 -12120 3030 -12110
rect 1550 -12220 3030 -12120
rect 1550 -12230 1560 -12220
rect 1420 -12240 1560 -12230
rect 1660 -12240 2690 -12220
rect 3020 -12230 3030 -12220
rect 3150 -12120 3160 -12110
rect 3260 -12120 3660 -12068
rect 3890 -12062 3905 -12030
rect 4281 -12062 4293 -12028
rect 3890 -12068 4293 -12062
rect 4857 -12028 5257 -12022
rect 4857 -12062 4869 -12028
rect 5245 -12030 5257 -12028
rect 5493 -12028 5893 -12022
rect 5493 -12030 5505 -12028
rect 5245 -12062 5260 -12030
rect 4857 -12068 5260 -12062
rect 3890 -12120 4290 -12068
rect 4620 -12110 4760 -12100
rect 4620 -12120 4630 -12110
rect 3150 -12220 4630 -12120
rect 3150 -12230 3160 -12220
rect 3020 -12240 3160 -12230
rect 3260 -12240 4290 -12220
rect 4620 -12230 4630 -12220
rect 4750 -12120 4760 -12110
rect 4860 -12120 5260 -12068
rect 5490 -12062 5505 -12030
rect 5881 -12062 5893 -12028
rect 5490 -12068 5893 -12062
rect 6457 -12028 6857 -12022
rect 6457 -12062 6469 -12028
rect 6845 -12030 6857 -12028
rect 7093 -12028 7493 -12022
rect 7093 -12030 7105 -12028
rect 6845 -12062 6860 -12030
rect 6457 -12068 6860 -12062
rect 5490 -12120 5890 -12068
rect 6220 -12110 6360 -12100
rect 6220 -12120 6230 -12110
rect 4750 -12220 6230 -12120
rect 4750 -12230 4760 -12220
rect 4620 -12240 4760 -12230
rect 4860 -12240 5890 -12220
rect 6220 -12230 6230 -12220
rect 6350 -12120 6360 -12110
rect 6460 -12120 6860 -12068
rect 7090 -12062 7105 -12030
rect 7481 -12062 7493 -12028
rect 7090 -12068 7493 -12062
rect 8057 -12028 8457 -12022
rect 8057 -12062 8069 -12028
rect 8445 -12030 8457 -12028
rect 8693 -12028 9093 -12022
rect 8693 -12030 8705 -12028
rect 8445 -12062 8460 -12030
rect 8057 -12068 8460 -12062
rect 7090 -12120 7490 -12068
rect 7820 -12110 7960 -12100
rect 7820 -12120 7830 -12110
rect 6350 -12220 7830 -12120
rect 6350 -12230 6360 -12220
rect 6220 -12240 6360 -12230
rect 6460 -12240 7490 -12220
rect 7820 -12230 7830 -12220
rect 7950 -12120 7960 -12110
rect 8060 -12120 8460 -12068
rect 8690 -12062 8705 -12030
rect 9081 -12062 9093 -12028
rect 8690 -12068 9093 -12062
rect 9657 -12028 10057 -12022
rect 9657 -12062 9669 -12028
rect 10045 -12030 10057 -12028
rect 10293 -12028 10693 -12022
rect 10293 -12030 10305 -12028
rect 10045 -12062 10060 -12030
rect 9657 -12068 10060 -12062
rect 8690 -12120 9090 -12068
rect 9420 -12110 9560 -12100
rect 9420 -12120 9430 -12110
rect 7950 -12220 9430 -12120
rect 7950 -12230 7960 -12220
rect 7820 -12240 7960 -12230
rect 8060 -12240 9090 -12220
rect 9420 -12230 9430 -12220
rect 9550 -12120 9560 -12110
rect 9660 -12120 10060 -12068
rect 10290 -12062 10305 -12030
rect 10681 -12062 10693 -12028
rect 10290 -12068 10693 -12062
rect 11257 -12028 11657 -12022
rect 11257 -12062 11269 -12028
rect 11645 -12062 11657 -12028
rect 11257 -12068 11657 -12062
rect 11893 -12028 12293 -12022
rect 11893 -12062 11905 -12028
rect 12281 -12062 12293 -12028
rect 11893 -12068 12293 -12062
rect 12857 -12028 13257 -12022
rect 12857 -12062 12869 -12028
rect 13245 -12030 13257 -12028
rect 13493 -12028 13893 -12022
rect 13493 -12030 13505 -12028
rect 13245 -12062 13260 -12030
rect 12857 -12068 13260 -12062
rect 10290 -12120 10690 -12068
rect 12860 -12120 13260 -12068
rect 13490 -12062 13505 -12030
rect 13881 -12062 13893 -12028
rect 13490 -12068 13893 -12062
rect 14457 -12028 14857 -12022
rect 14457 -12062 14469 -12028
rect 14845 -12030 14857 -12028
rect 15093 -12028 15493 -12022
rect 15093 -12030 15105 -12028
rect 14845 -12062 14860 -12030
rect 14457 -12068 14860 -12062
rect 13490 -12120 13890 -12068
rect 14460 -12120 14860 -12068
rect 15090 -12062 15105 -12030
rect 15481 -12062 15493 -12028
rect 15090 -12068 15493 -12062
rect 16057 -12028 16457 -12022
rect 16057 -12062 16069 -12028
rect 16445 -12062 16457 -12028
rect 16057 -12068 16457 -12062
rect 16693 -12028 17093 -12022
rect 16693 -12062 16705 -12028
rect 17081 -12062 17093 -12028
rect 16693 -12068 17093 -12062
rect 17657 -12028 18057 -12022
rect 17657 -12062 17669 -12028
rect 18045 -12062 18057 -12028
rect 17657 -12068 18057 -12062
rect 18293 -12028 18693 -12022
rect 18293 -12062 18305 -12028
rect 18681 -12062 18693 -12028
rect 18293 -12068 18693 -12062
rect 19257 -12028 19657 -12022
rect 19257 -12062 19269 -12028
rect 19645 -12062 19657 -12028
rect 19257 -12068 19657 -12062
rect 19893 -12028 20293 -12022
rect 19893 -12062 19905 -12028
rect 20281 -12062 20293 -12028
rect 19893 -12068 20293 -12062
rect 20857 -12028 21257 -12022
rect 20857 -12062 20869 -12028
rect 21245 -12062 21257 -12028
rect 20857 -12068 21257 -12062
rect 21493 -12028 21893 -12022
rect 21493 -12062 21505 -12028
rect 21881 -12062 21893 -12028
rect 21493 -12068 21893 -12062
rect 22457 -12028 22857 -12022
rect 22457 -12062 22469 -12028
rect 22845 -12062 22857 -12028
rect 22457 -12068 22857 -12062
rect 23093 -12028 23493 -12022
rect 23093 -12062 23105 -12028
rect 23481 -12062 23493 -12028
rect 23093 -12068 23493 -12062
rect 24057 -12028 24457 -12022
rect 24057 -12062 24069 -12028
rect 24445 -12062 24457 -12028
rect 24057 -12068 24457 -12062
rect 24693 -12028 25093 -12022
rect 24693 -12062 24705 -12028
rect 25081 -12062 25093 -12028
rect 24693 -12068 25093 -12062
rect 25657 -12028 26057 -12022
rect 25657 -12062 25669 -12028
rect 26045 -12062 26057 -12028
rect 25657 -12068 26057 -12062
rect 26293 -12028 26693 -12022
rect 26293 -12062 26305 -12028
rect 26681 -12062 26693 -12028
rect 26293 -12068 26693 -12062
rect 27257 -12028 27657 -12022
rect 27257 -12062 27269 -12028
rect 27645 -12062 27657 -12028
rect 27257 -12068 27657 -12062
rect 27893 -12028 28293 -12022
rect 27893 -12062 27905 -12028
rect 28281 -12062 28293 -12028
rect 27893 -12068 28293 -12062
rect 28857 -12028 29257 -12022
rect 28857 -12062 28869 -12028
rect 29245 -12062 29257 -12028
rect 28857 -12068 29257 -12062
rect 29493 -12028 29893 -12022
rect 29493 -12062 29505 -12028
rect 29881 -12062 29893 -12028
rect 29493 -12068 29893 -12062
rect 30457 -12028 30857 -12022
rect 30457 -12062 30469 -12028
rect 30845 -12062 30857 -12028
rect 30457 -12068 30857 -12062
rect 31093 -12028 31493 -12022
rect 31093 -12062 31105 -12028
rect 31481 -12062 31493 -12028
rect 31093 -12068 31493 -12062
rect 32057 -12028 32457 -12022
rect 32057 -12062 32069 -12028
rect 32445 -12062 32457 -12028
rect 32057 -12068 32457 -12062
rect 32693 -12028 33093 -12022
rect 32693 -12062 32705 -12028
rect 33081 -12062 33093 -12028
rect 32693 -12068 33093 -12062
rect 33657 -12028 34057 -12022
rect 33657 -12062 33669 -12028
rect 34045 -12062 34057 -12028
rect 33657 -12068 34057 -12062
rect 34293 -12028 34693 -12022
rect 34293 -12062 34305 -12028
rect 34681 -12062 34693 -12028
rect 34293 -12068 34693 -12062
rect 35257 -12028 35657 -12022
rect 35257 -12062 35269 -12028
rect 35645 -12062 35657 -12028
rect 35257 -12068 35657 -12062
rect 35893 -12028 36293 -12022
rect 35893 -12062 35905 -12028
rect 36281 -12062 36293 -12028
rect 35893 -12068 36293 -12062
rect 36857 -12028 37257 -12022
rect 36857 -12062 36869 -12028
rect 37245 -12062 37257 -12028
rect 36857 -12068 37257 -12062
rect 37493 -12028 37893 -12022
rect 37493 -12062 37505 -12028
rect 37881 -12062 37893 -12028
rect 37493 -12068 37893 -12062
rect 14900 -12100 15050 -12090
rect 14900 -12120 14910 -12100
rect 9550 -12220 10690 -12120
rect 9550 -12230 9560 -12220
rect 9420 -12240 9560 -12230
rect 9660 -12240 10690 -12220
rect 1660 -12290 2060 -12240
rect 670 -12296 1093 -12290
rect 670 -12330 705 -12296
rect 1081 -12330 1093 -12296
rect 670 -12336 1093 -12330
rect 1657 -12296 2060 -12290
rect 1657 -12330 1669 -12296
rect 2045 -12330 2060 -12296
rect 2290 -12290 2690 -12240
rect 3260 -12290 3660 -12240
rect 2290 -12296 2693 -12290
rect 2290 -12330 2305 -12296
rect 2681 -12330 2693 -12296
rect 1657 -12336 2057 -12330
rect 2293 -12336 2693 -12330
rect 3257 -12296 3660 -12290
rect 3257 -12330 3269 -12296
rect 3645 -12330 3660 -12296
rect 3890 -12290 4290 -12240
rect 4860 -12290 5260 -12240
rect 3890 -12296 4293 -12290
rect 3890 -12330 3905 -12296
rect 4281 -12330 4293 -12296
rect 3257 -12336 3657 -12330
rect 3893 -12336 4293 -12330
rect 4857 -12296 5260 -12290
rect 4857 -12330 4869 -12296
rect 5245 -12330 5260 -12296
rect 5490 -12290 5890 -12240
rect 6460 -12290 6860 -12240
rect 5490 -12296 5893 -12290
rect 5490 -12330 5505 -12296
rect 5881 -12330 5893 -12296
rect 4857 -12336 5257 -12330
rect 5493 -12336 5893 -12330
rect 6457 -12296 6860 -12290
rect 6457 -12330 6469 -12296
rect 6845 -12330 6860 -12296
rect 7090 -12290 7490 -12240
rect 8060 -12290 8460 -12240
rect 7090 -12296 7493 -12290
rect 7090 -12330 7105 -12296
rect 7481 -12330 7493 -12296
rect 6457 -12336 6857 -12330
rect 7093 -12336 7493 -12330
rect 8057 -12296 8460 -12290
rect 8057 -12330 8069 -12296
rect 8445 -12330 8460 -12296
rect 8690 -12290 9090 -12240
rect 9660 -12290 10060 -12240
rect 8690 -12296 9093 -12290
rect 8690 -12330 8705 -12296
rect 9081 -12330 9093 -12296
rect 8057 -12336 8457 -12330
rect 8693 -12336 9093 -12330
rect 9657 -12296 10060 -12290
rect 9657 -12330 9669 -12296
rect 10045 -12330 10060 -12296
rect 10290 -12290 10690 -12240
rect 11260 -12230 14910 -12120
rect 15040 -12120 15050 -12100
rect 15090 -12120 15490 -12068
rect 15040 -12230 15490 -12120
rect 11260 -12240 15490 -12230
rect 11260 -12290 12290 -12240
rect 12860 -12290 13260 -12240
rect 10290 -12296 10693 -12290
rect 10290 -12330 10305 -12296
rect 10681 -12330 10693 -12296
rect 9657 -12336 10057 -12330
rect 10293 -12336 10693 -12330
rect 11257 -12296 12293 -12290
rect 11257 -12330 11269 -12296
rect 11645 -12330 11905 -12296
rect 12281 -12330 12293 -12296
rect 11257 -12336 11657 -12330
rect 11893 -12336 12293 -12330
rect 12857 -12296 13260 -12290
rect 12857 -12330 12869 -12296
rect 13245 -12330 13260 -12296
rect 13490 -12290 13890 -12240
rect 14460 -12290 14860 -12240
rect 13490 -12296 13893 -12290
rect 13490 -12330 13505 -12296
rect 13881 -12330 13893 -12296
rect 12857 -12336 13257 -12330
rect 13493 -12336 13893 -12330
rect 14457 -12296 14860 -12290
rect 14457 -12330 14469 -12296
rect 14845 -12330 14860 -12296
rect 15090 -12290 15490 -12240
rect 15600 -12120 15740 -12110
rect 15600 -12240 15610 -12120
rect 15730 -12130 15740 -12120
rect 16060 -12130 16450 -12068
rect 16700 -12130 17090 -12068
rect 15730 -12230 17090 -12130
rect 15730 -12240 15740 -12230
rect 15600 -12250 15740 -12240
rect 16060 -12290 16450 -12230
rect 16700 -12290 17090 -12230
rect 17200 -12120 17340 -12110
rect 17200 -12240 17210 -12120
rect 17330 -12130 17340 -12120
rect 17660 -12130 18050 -12068
rect 18300 -12130 18690 -12068
rect 17330 -12230 18690 -12130
rect 17330 -12240 17340 -12230
rect 17200 -12250 17340 -12240
rect 17660 -12290 18050 -12230
rect 18300 -12290 18690 -12230
rect 18800 -12120 18940 -12110
rect 18800 -12240 18810 -12120
rect 18930 -12130 18940 -12120
rect 19260 -12130 19650 -12068
rect 19900 -12130 20290 -12068
rect 18930 -12230 20290 -12130
rect 18930 -12240 18940 -12230
rect 18800 -12250 18940 -12240
rect 19260 -12290 19650 -12230
rect 19900 -12290 20290 -12230
rect 20400 -12120 20540 -12110
rect 20400 -12240 20410 -12120
rect 20530 -12130 20540 -12120
rect 20860 -12130 21250 -12068
rect 21500 -12130 21890 -12068
rect 20530 -12230 21890 -12130
rect 20530 -12240 20540 -12230
rect 20400 -12250 20540 -12240
rect 20860 -12290 21250 -12230
rect 21500 -12290 21890 -12230
rect 22000 -12120 22140 -12110
rect 22000 -12240 22010 -12120
rect 22130 -12130 22140 -12120
rect 22460 -12130 22850 -12068
rect 23100 -12130 23490 -12068
rect 22130 -12230 23490 -12130
rect 22130 -12240 22140 -12230
rect 22000 -12250 22140 -12240
rect 22460 -12290 22850 -12230
rect 23100 -12290 23490 -12230
rect 23600 -12120 23740 -12110
rect 23600 -12240 23610 -12120
rect 23730 -12130 23740 -12120
rect 24060 -12130 24450 -12068
rect 24700 -12130 25090 -12068
rect 23730 -12230 25090 -12130
rect 23730 -12240 23740 -12230
rect 23600 -12250 23740 -12240
rect 24060 -12290 24450 -12230
rect 24700 -12290 25090 -12230
rect 25200 -12120 25340 -12110
rect 25200 -12240 25210 -12120
rect 25330 -12130 25340 -12120
rect 25660 -12130 26050 -12068
rect 26300 -12130 26690 -12068
rect 25330 -12230 26690 -12130
rect 25330 -12240 25340 -12230
rect 25200 -12250 25340 -12240
rect 25660 -12290 26050 -12230
rect 26300 -12290 26690 -12230
rect 26800 -12120 26940 -12110
rect 26800 -12240 26810 -12120
rect 26930 -12130 26940 -12120
rect 27260 -12130 27650 -12068
rect 27900 -12130 28290 -12068
rect 26930 -12230 28290 -12130
rect 26930 -12240 26940 -12230
rect 26800 -12250 26940 -12240
rect 27260 -12290 27650 -12230
rect 27900 -12290 28290 -12230
rect 28400 -12120 28540 -12110
rect 28400 -12240 28410 -12120
rect 28530 -12130 28540 -12120
rect 28860 -12130 29250 -12068
rect 29500 -12130 29890 -12068
rect 28530 -12230 29890 -12130
rect 28530 -12240 28540 -12230
rect 28400 -12250 28540 -12240
rect 28860 -12290 29250 -12230
rect 29500 -12290 29890 -12230
rect 30000 -12120 30140 -12110
rect 30000 -12240 30010 -12120
rect 30130 -12130 30140 -12120
rect 30460 -12130 30850 -12068
rect 31100 -12130 31490 -12068
rect 30130 -12230 31490 -12130
rect 30130 -12240 30140 -12230
rect 30000 -12250 30140 -12240
rect 30460 -12290 30850 -12230
rect 31100 -12290 31490 -12230
rect 31600 -12120 31740 -12110
rect 31600 -12240 31610 -12120
rect 31730 -12130 31740 -12120
rect 32060 -12130 32450 -12068
rect 32700 -12130 33090 -12068
rect 33660 -12130 34050 -12068
rect 34300 -12130 34690 -12068
rect 35260 -12130 35650 -12068
rect 35900 -12130 36290 -12068
rect 31730 -12230 36290 -12130
rect 31730 -12240 31740 -12230
rect 31600 -12250 31740 -12240
rect 32060 -12290 32450 -12230
rect 32700 -12290 33090 -12230
rect 33660 -12290 34050 -12230
rect 34300 -12290 34690 -12230
rect 35260 -12290 35650 -12230
rect 35900 -12290 36290 -12230
rect 15090 -12296 15493 -12290
rect 15090 -12330 15105 -12296
rect 15481 -12330 15493 -12296
rect 14457 -12336 14857 -12330
rect 15093 -12336 15493 -12330
rect 16057 -12296 16457 -12290
rect 16057 -12330 16069 -12296
rect 16445 -12330 16457 -12296
rect 16057 -12336 16457 -12330
rect 16693 -12296 17093 -12290
rect 16693 -12330 16705 -12296
rect 17081 -12330 17093 -12296
rect 16693 -12336 17093 -12330
rect 17657 -12296 18057 -12290
rect 17657 -12330 17669 -12296
rect 18045 -12330 18057 -12296
rect 17657 -12336 18057 -12330
rect 18293 -12296 18693 -12290
rect 18293 -12330 18305 -12296
rect 18681 -12330 18693 -12296
rect 18293 -12336 18693 -12330
rect 19257 -12296 19657 -12290
rect 19257 -12330 19269 -12296
rect 19645 -12330 19657 -12296
rect 19257 -12336 19657 -12330
rect 19893 -12296 20293 -12290
rect 19893 -12330 19905 -12296
rect 20281 -12330 20293 -12296
rect 19893 -12336 20293 -12330
rect 20857 -12296 21257 -12290
rect 20857 -12330 20869 -12296
rect 21245 -12330 21257 -12296
rect 20857 -12336 21257 -12330
rect 21493 -12296 21893 -12290
rect 21493 -12330 21505 -12296
rect 21881 -12330 21893 -12296
rect 21493 -12336 21893 -12330
rect 22457 -12296 22857 -12290
rect 22457 -12330 22469 -12296
rect 22845 -12330 22857 -12296
rect 22457 -12336 22857 -12330
rect 23093 -12296 23493 -12290
rect 23093 -12330 23105 -12296
rect 23481 -12330 23493 -12296
rect 23093 -12336 23493 -12330
rect 24057 -12296 24457 -12290
rect 24057 -12330 24069 -12296
rect 24445 -12330 24457 -12296
rect 24057 -12336 24457 -12330
rect 24693 -12296 25093 -12290
rect 24693 -12330 24705 -12296
rect 25081 -12330 25093 -12296
rect 24693 -12336 25093 -12330
rect 25657 -12296 26057 -12290
rect 25657 -12330 25669 -12296
rect 26045 -12330 26057 -12296
rect 25657 -12336 26057 -12330
rect 26293 -12296 26693 -12290
rect 26293 -12330 26305 -12296
rect 26681 -12330 26693 -12296
rect 26293 -12336 26693 -12330
rect 27257 -12296 27657 -12290
rect 27257 -12330 27269 -12296
rect 27645 -12330 27657 -12296
rect 27257 -12336 27657 -12330
rect 27893 -12296 28293 -12290
rect 27893 -12330 27905 -12296
rect 28281 -12330 28293 -12296
rect 27893 -12336 28293 -12330
rect 28857 -12296 29257 -12290
rect 28857 -12330 28869 -12296
rect 29245 -12330 29257 -12296
rect 28857 -12336 29257 -12330
rect 29493 -12296 29893 -12290
rect 29493 -12330 29505 -12296
rect 29881 -12330 29893 -12296
rect 29493 -12336 29893 -12330
rect 30457 -12296 30857 -12290
rect 30457 -12330 30469 -12296
rect 30845 -12330 30857 -12296
rect 30457 -12336 30857 -12330
rect 31093 -12296 31493 -12290
rect 31093 -12330 31105 -12296
rect 31481 -12330 31493 -12296
rect 31093 -12336 31493 -12330
rect 32057 -12296 32457 -12290
rect 32057 -12330 32069 -12296
rect 32445 -12330 32457 -12296
rect 32057 -12336 32457 -12330
rect 32693 -12296 33093 -12290
rect 32693 -12330 32705 -12296
rect 33081 -12330 33093 -12296
rect 32693 -12336 33093 -12330
rect 33657 -12296 34057 -12290
rect 33657 -12330 33669 -12296
rect 34045 -12330 34057 -12296
rect 33657 -12336 34057 -12330
rect 34293 -12296 34693 -12290
rect 34293 -12330 34305 -12296
rect 34681 -12330 34693 -12296
rect 34293 -12336 34693 -12330
rect 35257 -12296 35657 -12290
rect 35257 -12330 35269 -12296
rect 35645 -12330 35657 -12296
rect 35257 -12336 35657 -12330
rect 35893 -12296 36293 -12290
rect 35893 -12330 35905 -12296
rect 36281 -12330 36293 -12296
rect 35893 -12336 36293 -12330
rect 36857 -12296 37257 -12290
rect 36857 -12330 36869 -12296
rect 37245 -12330 37257 -12296
rect 36857 -12336 37257 -12330
rect 37493 -12296 37893 -12290
rect 37493 -12330 37505 -12296
rect 37881 -12330 37893 -12296
rect 37493 -12336 37893 -12330
rect 57 -13154 490 -13148
rect 57 -13180 69 -13154
rect 0 -13188 69 -13180
rect 445 -13188 490 -13154
rect 0 -13288 490 -13188
rect 670 -13148 720 -12336
rect 1134 -12396 1180 -12384
rect 1134 -13088 1140 -12396
rect 1174 -13088 1180 -12396
rect 1134 -13100 1180 -13088
rect 1570 -12396 1616 -12384
rect 1570 -13088 1576 -12396
rect 1610 -13088 1616 -12396
rect 1570 -13100 1616 -13088
rect 2098 -12396 2144 -12384
rect 2098 -13088 2104 -12396
rect 2138 -12400 2144 -12396
rect 2206 -12396 2252 -12384
rect 2206 -12400 2212 -12396
rect 2138 -12410 2212 -12400
rect 2138 -13080 2212 -13070
rect 2138 -13088 2144 -13080
rect 2098 -13100 2144 -13088
rect 2206 -13088 2212 -13080
rect 2246 -13088 2252 -12396
rect 2206 -13100 2252 -13088
rect 2734 -12396 2780 -12384
rect 2734 -13088 2740 -12396
rect 2774 -13088 2780 -12396
rect 2734 -13100 2780 -13088
rect 3170 -12396 3216 -12384
rect 3170 -13088 3176 -12396
rect 3210 -13088 3216 -12396
rect 3170 -13100 3216 -13088
rect 3698 -12396 3744 -12384
rect 3698 -13088 3704 -12396
rect 3738 -12400 3744 -12396
rect 3806 -12396 3852 -12384
rect 3806 -12400 3812 -12396
rect 3738 -12410 3812 -12400
rect 3738 -13080 3812 -13070
rect 3738 -13088 3744 -13080
rect 3698 -13100 3744 -13088
rect 3806 -13088 3812 -13080
rect 3846 -13088 3852 -12396
rect 3806 -13100 3852 -13088
rect 4334 -12396 4380 -12384
rect 4334 -13088 4340 -12396
rect 4374 -13088 4380 -12396
rect 4334 -13100 4380 -13088
rect 4770 -12396 4816 -12384
rect 4770 -13088 4776 -12396
rect 4810 -13088 4816 -12396
rect 4770 -13100 4816 -13088
rect 5298 -12396 5344 -12384
rect 5298 -13088 5304 -12396
rect 5338 -12400 5344 -12396
rect 5406 -12396 5452 -12384
rect 5406 -12400 5412 -12396
rect 5338 -12410 5412 -12400
rect 5338 -13080 5412 -13070
rect 5338 -13088 5344 -13080
rect 5298 -13100 5344 -13088
rect 5406 -13088 5412 -13080
rect 5446 -13088 5452 -12396
rect 5406 -13100 5452 -13088
rect 5934 -12396 5980 -12384
rect 5934 -13088 5940 -12396
rect 5974 -13088 5980 -12396
rect 5934 -13100 5980 -13088
rect 6370 -12396 6416 -12384
rect 6370 -13088 6376 -12396
rect 6410 -13088 6416 -12396
rect 6370 -13100 6416 -13088
rect 6898 -12396 6944 -12384
rect 6898 -13088 6904 -12396
rect 6938 -12400 6944 -12396
rect 7006 -12396 7052 -12384
rect 7006 -12400 7012 -12396
rect 6938 -12410 7012 -12400
rect 6938 -13080 7012 -13070
rect 6938 -13088 6944 -13080
rect 6898 -13100 6944 -13088
rect 7006 -13088 7012 -13080
rect 7046 -13088 7052 -12396
rect 7006 -13100 7052 -13088
rect 7534 -12396 7580 -12384
rect 7534 -13088 7540 -12396
rect 7574 -13088 7580 -12396
rect 7534 -13100 7580 -13088
rect 7970 -12396 8016 -12384
rect 7970 -13088 7976 -12396
rect 8010 -13088 8016 -12396
rect 7970 -13100 8016 -13088
rect 8498 -12396 8544 -12384
rect 8498 -13088 8504 -12396
rect 8538 -12400 8544 -12396
rect 8606 -12396 8652 -12384
rect 8606 -12400 8612 -12396
rect 8538 -12410 8612 -12400
rect 8538 -13080 8612 -13070
rect 8538 -13088 8544 -13080
rect 8498 -13100 8544 -13088
rect 8606 -13088 8612 -13080
rect 8646 -13088 8652 -12396
rect 8606 -13100 8652 -13088
rect 9134 -12396 9180 -12384
rect 9134 -13088 9140 -12396
rect 9174 -13088 9180 -12396
rect 9134 -13100 9180 -13088
rect 9570 -12396 9616 -12384
rect 9570 -13088 9576 -12396
rect 9610 -13088 9616 -12396
rect 9570 -13100 9616 -13088
rect 10098 -12396 10144 -12384
rect 10098 -13088 10104 -12396
rect 10138 -12400 10144 -12396
rect 10206 -12396 10252 -12384
rect 10206 -12400 10212 -12396
rect 10138 -12410 10212 -12400
rect 10138 -13080 10212 -13070
rect 10138 -13088 10144 -13080
rect 10098 -13100 10144 -13088
rect 10206 -13088 10212 -13080
rect 10246 -13088 10252 -12396
rect 10206 -13100 10252 -13088
rect 10734 -12396 10780 -12384
rect 10734 -13088 10740 -12396
rect 10774 -13088 10780 -12396
rect 10734 -13100 10780 -13088
rect 11170 -12396 11216 -12384
rect 11170 -13088 11176 -12396
rect 11210 -13088 11216 -12396
rect 11170 -13100 11216 -13088
rect 11698 -12396 11744 -12384
rect 11698 -13088 11704 -12396
rect 11738 -12400 11744 -12396
rect 11806 -12396 11852 -12384
rect 11806 -12400 11812 -12396
rect 11738 -12410 11812 -12400
rect 11738 -13080 11812 -13070
rect 11738 -13088 11744 -13080
rect 11698 -13100 11744 -13088
rect 11806 -13088 11812 -13080
rect 11846 -13088 11852 -12396
rect 11806 -13100 11852 -13088
rect 12334 -12396 12380 -12384
rect 12334 -13088 12340 -12396
rect 12374 -13088 12380 -12396
rect 12334 -13100 12380 -13088
rect 12770 -12396 12816 -12384
rect 12770 -13088 12776 -12396
rect 12810 -13088 12816 -12396
rect 12770 -13100 12816 -13088
rect 13298 -12396 13344 -12384
rect 13298 -13088 13304 -12396
rect 13338 -12400 13344 -12396
rect 13406 -12396 13452 -12384
rect 13406 -12400 13412 -12396
rect 13338 -12410 13412 -12400
rect 13338 -13080 13412 -13070
rect 13338 -13088 13344 -13080
rect 13298 -13100 13344 -13088
rect 13406 -13088 13412 -13080
rect 13446 -13088 13452 -12396
rect 13406 -13100 13452 -13088
rect 13934 -12396 13980 -12384
rect 13934 -13088 13940 -12396
rect 13974 -13088 13980 -12396
rect 13934 -13100 13980 -13088
rect 14370 -12396 14416 -12384
rect 14370 -13088 14376 -12396
rect 14410 -13088 14416 -12396
rect 14370 -13100 14416 -13088
rect 14898 -12396 14944 -12384
rect 14898 -13088 14904 -12396
rect 14938 -12400 14944 -12396
rect 15006 -12396 15052 -12384
rect 15006 -12400 15012 -12396
rect 14938 -12410 15012 -12400
rect 14938 -13080 15012 -13070
rect 14938 -13088 14944 -13080
rect 14898 -13100 14944 -13088
rect 15006 -13088 15012 -13080
rect 15046 -13088 15052 -12396
rect 15006 -13100 15052 -13088
rect 15534 -12396 15580 -12384
rect 15534 -13088 15540 -12396
rect 15574 -13088 15580 -12396
rect 15534 -13100 15580 -13088
rect 15970 -12396 16016 -12384
rect 15970 -13088 15976 -12396
rect 16010 -13088 16016 -12396
rect 15970 -13100 16016 -13088
rect 16498 -12390 16544 -12384
rect 16606 -12390 16652 -12384
rect 16498 -12396 16652 -12390
rect 16498 -13088 16504 -12396
rect 16538 -12400 16612 -12396
rect 16538 -13088 16612 -13080
rect 16646 -13088 16652 -12396
rect 16498 -13090 16652 -13088
rect 16498 -13100 16544 -13090
rect 16606 -13100 16652 -13090
rect 17134 -12396 17180 -12384
rect 17134 -13088 17140 -12396
rect 17174 -13088 17180 -12396
rect 17134 -13100 17180 -13088
rect 17570 -12396 17616 -12384
rect 17570 -13088 17576 -12396
rect 17610 -13088 17616 -12396
rect 17570 -13100 17616 -13088
rect 18098 -12390 18144 -12384
rect 18206 -12390 18252 -12384
rect 18098 -12396 18252 -12390
rect 18098 -13088 18104 -12396
rect 18138 -12400 18212 -12396
rect 18138 -13088 18212 -13080
rect 18246 -13088 18252 -12396
rect 18098 -13090 18252 -13088
rect 18098 -13100 18144 -13090
rect 18206 -13100 18252 -13090
rect 18734 -12396 18780 -12384
rect 18734 -13088 18740 -12396
rect 18774 -13088 18780 -12396
rect 18734 -13100 18780 -13088
rect 19170 -12396 19216 -12384
rect 19170 -13088 19176 -12396
rect 19210 -13088 19216 -12396
rect 19170 -13100 19216 -13088
rect 19698 -12390 19744 -12384
rect 19806 -12390 19852 -12384
rect 19698 -12396 19852 -12390
rect 19698 -13088 19704 -12396
rect 19738 -12400 19812 -12396
rect 19738 -13088 19812 -13080
rect 19846 -13088 19852 -12396
rect 19698 -13090 19852 -13088
rect 19698 -13100 19744 -13090
rect 19806 -13100 19852 -13090
rect 20334 -12396 20380 -12384
rect 20334 -13088 20340 -12396
rect 20374 -13088 20380 -12396
rect 20334 -13100 20380 -13088
rect 20770 -12396 20816 -12384
rect 20770 -13088 20776 -12396
rect 20810 -13088 20816 -12396
rect 20770 -13100 20816 -13088
rect 21298 -12390 21344 -12384
rect 21406 -12390 21452 -12384
rect 21298 -12396 21452 -12390
rect 21298 -13088 21304 -12396
rect 21338 -12400 21412 -12396
rect 21338 -13088 21412 -13080
rect 21446 -13088 21452 -12396
rect 21298 -13090 21452 -13088
rect 21298 -13100 21344 -13090
rect 21406 -13100 21452 -13090
rect 21934 -12396 21980 -12384
rect 21934 -13088 21940 -12396
rect 21974 -13088 21980 -12396
rect 21934 -13100 21980 -13088
rect 22370 -12396 22416 -12384
rect 22370 -13088 22376 -12396
rect 22410 -13088 22416 -12396
rect 22370 -13100 22416 -13088
rect 22898 -12390 22944 -12384
rect 23006 -12390 23052 -12384
rect 22898 -12396 23052 -12390
rect 22898 -13088 22904 -12396
rect 22938 -12400 23012 -12396
rect 22938 -13088 23012 -13080
rect 23046 -13088 23052 -12396
rect 22898 -13090 23052 -13088
rect 22898 -13100 22944 -13090
rect 23006 -13100 23052 -13090
rect 23534 -12396 23580 -12384
rect 23534 -13088 23540 -12396
rect 23574 -13088 23580 -12396
rect 23534 -13100 23580 -13088
rect 23970 -12396 24016 -12384
rect 23970 -13088 23976 -12396
rect 24010 -13088 24016 -12396
rect 23970 -13100 24016 -13088
rect 24498 -12390 24544 -12384
rect 24606 -12390 24652 -12384
rect 24498 -12396 24652 -12390
rect 24498 -13088 24504 -12396
rect 24538 -12400 24612 -12396
rect 24538 -13088 24612 -13080
rect 24646 -13088 24652 -12396
rect 24498 -13090 24652 -13088
rect 24498 -13100 24544 -13090
rect 24606 -13100 24652 -13090
rect 25134 -12396 25180 -12384
rect 25134 -13088 25140 -12396
rect 25174 -13088 25180 -12396
rect 25134 -13100 25180 -13088
rect 25570 -12396 25616 -12384
rect 25570 -13088 25576 -12396
rect 25610 -13088 25616 -12396
rect 25570 -13100 25616 -13088
rect 26098 -12390 26144 -12384
rect 26206 -12390 26252 -12384
rect 26098 -12396 26252 -12390
rect 26098 -13088 26104 -12396
rect 26138 -12400 26212 -12396
rect 26138 -13088 26212 -13080
rect 26246 -13088 26252 -12396
rect 26098 -13090 26252 -13088
rect 26098 -13100 26144 -13090
rect 26206 -13100 26252 -13090
rect 26734 -12396 26780 -12384
rect 26734 -13088 26740 -12396
rect 26774 -13088 26780 -12396
rect 26734 -13100 26780 -13088
rect 27170 -12396 27216 -12384
rect 27170 -13088 27176 -12396
rect 27210 -13088 27216 -12396
rect 27170 -13100 27216 -13088
rect 27698 -12390 27744 -12384
rect 27806 -12390 27852 -12384
rect 27698 -12396 27852 -12390
rect 27698 -13088 27704 -12396
rect 27738 -12400 27812 -12396
rect 27738 -13088 27812 -13080
rect 27846 -13088 27852 -12396
rect 27698 -13090 27852 -13088
rect 27698 -13100 27744 -13090
rect 27806 -13100 27852 -13090
rect 28334 -12396 28380 -12384
rect 28334 -13088 28340 -12396
rect 28374 -13088 28380 -12396
rect 28334 -13100 28380 -13088
rect 28770 -12396 28816 -12384
rect 28770 -13088 28776 -12396
rect 28810 -13088 28816 -12396
rect 28770 -13100 28816 -13088
rect 29298 -12390 29344 -12384
rect 29406 -12390 29452 -12384
rect 29298 -12396 29452 -12390
rect 29298 -13088 29304 -12396
rect 29338 -12400 29412 -12396
rect 29338 -13088 29412 -13080
rect 29446 -13088 29452 -12396
rect 29298 -13090 29452 -13088
rect 29298 -13100 29344 -13090
rect 29406 -13100 29452 -13090
rect 29934 -12396 29980 -12384
rect 29934 -13088 29940 -12396
rect 29974 -13088 29980 -12396
rect 29934 -13100 29980 -13088
rect 30370 -12396 30416 -12384
rect 30370 -13088 30376 -12396
rect 30410 -13088 30416 -12396
rect 30370 -13100 30416 -13088
rect 30898 -12390 30944 -12384
rect 31006 -12390 31052 -12384
rect 30898 -12396 31052 -12390
rect 30898 -13088 30904 -12396
rect 30938 -12400 31012 -12396
rect 30938 -13088 31012 -13080
rect 31046 -13088 31052 -12396
rect 30898 -13090 31052 -13088
rect 30898 -13100 30944 -13090
rect 31006 -13100 31052 -13090
rect 31534 -12396 31580 -12384
rect 31534 -13088 31540 -12396
rect 31574 -13088 31580 -12396
rect 31534 -13100 31580 -13088
rect 31970 -12396 32016 -12384
rect 31970 -13088 31976 -12396
rect 32010 -13088 32016 -12396
rect 31970 -13100 32016 -13088
rect 32498 -12390 32544 -12384
rect 32606 -12390 32652 -12384
rect 32498 -12396 32652 -12390
rect 32498 -13088 32504 -12396
rect 32538 -12400 32612 -12396
rect 32538 -13088 32544 -12910
rect 32498 -13100 32544 -13088
rect 32606 -13088 32612 -12910
rect 32646 -13088 32652 -12396
rect 32606 -13100 32652 -13088
rect 33134 -12396 33180 -12384
rect 33134 -13088 33140 -12396
rect 33174 -13088 33180 -12396
rect 33134 -13100 33180 -13088
rect 33570 -12396 33616 -12384
rect 33570 -13088 33576 -12396
rect 33610 -13088 33616 -12396
rect 33570 -13100 33616 -13088
rect 34098 -12390 34144 -12384
rect 34206 -12390 34252 -12384
rect 34098 -12396 34252 -12390
rect 34098 -13088 34104 -12396
rect 34138 -12400 34212 -12396
rect 34138 -13088 34144 -12910
rect 34098 -13100 34144 -13088
rect 34206 -13088 34212 -12910
rect 34246 -13088 34252 -12396
rect 34206 -13100 34252 -13088
rect 34734 -12396 34780 -12384
rect 34734 -13088 34740 -12396
rect 34774 -13088 34780 -12396
rect 34734 -13100 34780 -13088
rect 35170 -12396 35216 -12384
rect 35170 -13088 35176 -12396
rect 35210 -13088 35216 -12396
rect 35170 -13100 35216 -13088
rect 35698 -12390 35744 -12384
rect 35806 -12390 35852 -12384
rect 35698 -12396 35852 -12390
rect 35698 -13088 35704 -12396
rect 35738 -12400 35812 -12396
rect 35738 -13088 35744 -12910
rect 35698 -13100 35744 -13088
rect 35806 -13088 35812 -12910
rect 35846 -13088 35852 -12396
rect 35806 -13100 35852 -13088
rect 36334 -12396 36380 -12384
rect 36334 -13088 36340 -12396
rect 36374 -13088 36380 -12396
rect 36334 -13100 36380 -13088
rect 36770 -12396 36816 -12384
rect 36770 -13088 36776 -12396
rect 36810 -13088 36816 -12396
rect 36770 -13100 36816 -13088
rect 37298 -12396 37344 -12384
rect 37298 -13088 37304 -12396
rect 37338 -13088 37344 -12396
rect 37298 -13100 37344 -13088
rect 37406 -12396 37452 -12384
rect 37406 -13088 37412 -12396
rect 37446 -13088 37452 -12396
rect 37406 -13100 37452 -13088
rect 37934 -12396 37980 -12384
rect 37934 -13088 37940 -12396
rect 37974 -13088 37980 -12396
rect 37934 -13100 37980 -13088
rect 35000 -13110 35140 -13100
rect 670 -13154 1093 -13148
rect 670 -13188 705 -13154
rect 1081 -13180 1093 -13154
rect 1657 -13154 2057 -13148
rect 1657 -13180 1669 -13154
rect 1081 -13188 1669 -13180
rect 2045 -13180 2057 -13154
rect 2293 -13154 2693 -13148
rect 2293 -13180 2305 -13154
rect 2045 -13188 2305 -13180
rect 2681 -13180 2693 -13154
rect 3257 -13154 3657 -13148
rect 3257 -13180 3269 -13154
rect 2681 -13188 3269 -13180
rect 3645 -13180 3657 -13154
rect 3893 -13154 4293 -13148
rect 3893 -13180 3905 -13154
rect 3645 -13188 3905 -13180
rect 4281 -13180 4293 -13154
rect 4857 -13154 5257 -13148
rect 4857 -13180 4869 -13154
rect 4281 -13188 4869 -13180
rect 5245 -13180 5257 -13154
rect 5493 -13154 5893 -13148
rect 5493 -13180 5505 -13154
rect 5245 -13188 5505 -13180
rect 5881 -13180 5893 -13154
rect 6457 -13154 6857 -13148
rect 6457 -13180 6469 -13154
rect 5881 -13188 6469 -13180
rect 6845 -13180 6857 -13154
rect 7093 -13154 7493 -13148
rect 7093 -13180 7105 -13154
rect 6845 -13188 7105 -13180
rect 7481 -13180 7493 -13154
rect 8057 -13154 8457 -13148
rect 8057 -13180 8069 -13154
rect 7481 -13188 8069 -13180
rect 8445 -13180 8457 -13154
rect 8693 -13154 9093 -13148
rect 8693 -13180 8705 -13154
rect 8445 -13188 8705 -13180
rect 9081 -13180 9093 -13154
rect 9657 -13154 10057 -13148
rect 9657 -13180 9669 -13154
rect 9081 -13188 9669 -13180
rect 10045 -13180 10057 -13154
rect 10293 -13154 10693 -13148
rect 10293 -13180 10305 -13154
rect 10045 -13188 10305 -13180
rect 10681 -13180 10693 -13154
rect 11257 -13150 11657 -13148
rect 11893 -13150 12293 -13148
rect 11257 -13154 11270 -13150
rect 11650 -13154 12300 -13150
rect 10681 -13188 11080 -13180
rect 670 -13288 11080 -13188
rect 11257 -13188 11269 -13154
rect 11650 -13188 11905 -13154
rect 12281 -13188 12300 -13154
rect 12857 -13154 13257 -13148
rect 12857 -13180 12869 -13154
rect 11257 -13194 11270 -13188
rect 11260 -13210 11270 -13194
rect 11650 -13210 12300 -13188
rect 12720 -13188 12869 -13180
rect 13245 -13180 13257 -13154
rect 13493 -13154 13893 -13148
rect 13493 -13180 13505 -13154
rect 13245 -13188 13505 -13180
rect 13881 -13180 13893 -13154
rect 14457 -13154 14857 -13148
rect 14457 -13180 14469 -13154
rect 13881 -13188 14469 -13180
rect 14845 -13180 14857 -13154
rect 15093 -13154 15493 -13148
rect 15093 -13180 15105 -13154
rect 14845 -13188 15105 -13180
rect 15481 -13180 15493 -13154
rect 16057 -13154 16457 -13148
rect 16057 -13180 16069 -13154
rect 15481 -13188 16069 -13180
rect 16445 -13180 16457 -13154
rect 16693 -13154 17093 -13148
rect 16693 -13180 16705 -13154
rect 16445 -13188 16705 -13180
rect 17081 -13180 17093 -13154
rect 17657 -13154 18057 -13148
rect 17657 -13180 17669 -13154
rect 17081 -13188 17669 -13180
rect 18045 -13180 18057 -13154
rect 18293 -13154 18693 -13148
rect 18293 -13180 18305 -13154
rect 18045 -13188 18305 -13180
rect 18681 -13180 18693 -13154
rect 19257 -13154 19657 -13148
rect 19257 -13180 19269 -13154
rect 18681 -13188 19269 -13180
rect 19645 -13180 19657 -13154
rect 19893 -13154 20293 -13148
rect 19893 -13180 19905 -13154
rect 19645 -13188 19905 -13180
rect 20281 -13180 20293 -13154
rect 20857 -13154 21257 -13148
rect 20857 -13180 20869 -13154
rect 20281 -13188 20869 -13180
rect 21245 -13180 21257 -13154
rect 21493 -13154 21893 -13148
rect 21493 -13180 21505 -13154
rect 21245 -13188 21505 -13180
rect 21881 -13180 21893 -13154
rect 22457 -13154 22857 -13148
rect 22457 -13180 22469 -13154
rect 21881 -13188 22469 -13180
rect 22845 -13180 22857 -13154
rect 23093 -13154 23493 -13148
rect 23093 -13180 23105 -13154
rect 22845 -13188 23105 -13180
rect 23481 -13180 23493 -13154
rect 24057 -13154 24457 -13148
rect 24057 -13180 24069 -13154
rect 23481 -13188 24069 -13180
rect 24445 -13180 24457 -13154
rect 24693 -13154 25093 -13148
rect 24693 -13180 24705 -13154
rect 24445 -13188 24705 -13180
rect 25081 -13180 25093 -13154
rect 25657 -13154 26057 -13148
rect 25657 -13180 25669 -13154
rect 25081 -13188 25669 -13180
rect 26045 -13180 26057 -13154
rect 26293 -13154 26693 -13148
rect 26293 -13180 26305 -13154
rect 26045 -13188 26305 -13180
rect 26681 -13180 26693 -13154
rect 27257 -13154 27657 -13148
rect 27257 -13180 27269 -13154
rect 26681 -13188 27269 -13180
rect 27645 -13180 27657 -13154
rect 27893 -13154 28293 -13148
rect 27893 -13180 27905 -13154
rect 27645 -13188 27905 -13180
rect 28281 -13180 28293 -13154
rect 28857 -13154 29257 -13148
rect 28857 -13180 28869 -13154
rect 28281 -13188 28869 -13180
rect 29245 -13180 29257 -13154
rect 29493 -13154 29893 -13148
rect 29493 -13180 29505 -13154
rect 29245 -13188 29505 -13180
rect 29881 -13180 29893 -13154
rect 30457 -13154 30857 -13148
rect 30457 -13180 30469 -13154
rect 29881 -13188 30469 -13180
rect 30845 -13180 30857 -13154
rect 31093 -13154 31493 -13148
rect 31093 -13180 31105 -13154
rect 30845 -13188 31105 -13180
rect 31481 -13180 31493 -13154
rect 32057 -13150 32457 -13148
rect 32693 -13150 33093 -13148
rect 33657 -13150 34057 -13148
rect 34293 -13150 34693 -13148
rect 35000 -13150 35010 -13110
rect 32057 -13154 35010 -13150
rect 31481 -13188 31860 -13180
rect 0 -13322 13 -13288
rect 1137 -13322 1613 -13288
rect 2737 -13322 3213 -13288
rect 4337 -13322 4813 -13288
rect 5937 -13322 6413 -13288
rect 7537 -13322 8013 -13288
rect 9137 -13322 9613 -13288
rect 10737 -13300 11080 -13288
rect 11201 -13288 12349 -13282
rect 11201 -13300 11213 -13288
rect 10737 -13322 11213 -13300
rect 12337 -13300 12349 -13288
rect 12720 -13288 31860 -13188
rect 32057 -13188 32069 -13154
rect 32445 -13188 32705 -13154
rect 33081 -13188 33669 -13154
rect 34045 -13188 34305 -13154
rect 34681 -13188 35010 -13154
rect 32057 -13194 35010 -13188
rect 32060 -13230 35010 -13194
rect 35130 -13150 35140 -13110
rect 35257 -13150 35657 -13148
rect 35893 -13150 36293 -13148
rect 35130 -13154 36293 -13150
rect 35130 -13188 35269 -13154
rect 35645 -13188 35905 -13154
rect 36281 -13188 36293 -13154
rect 35130 -13194 36293 -13188
rect 36857 -13154 37257 -13148
rect 36857 -13188 36869 -13154
rect 37245 -13188 37257 -13154
rect 36857 -13194 37257 -13188
rect 37493 -13154 37893 -13148
rect 37493 -13188 37505 -13154
rect 37881 -13188 37893 -13154
rect 37493 -13194 37893 -13188
rect 35130 -13230 36290 -13194
rect 32060 -13240 36290 -13230
rect 12720 -13300 12813 -13288
rect 12337 -13322 12813 -13300
rect 13937 -13322 14413 -13288
rect 15537 -13322 16013 -13288
rect 17137 -13322 17613 -13288
rect 18737 -13322 19213 -13288
rect 20337 -13322 20813 -13288
rect 21937 -13322 22413 -13288
rect 23537 -13322 24013 -13288
rect 25137 -13322 25613 -13288
rect 26737 -13322 27213 -13288
rect 28337 -13322 28813 -13288
rect 29937 -13322 30413 -13288
rect 31537 -13300 31860 -13288
rect 32001 -13288 33149 -13282
rect 32001 -13300 32013 -13288
rect 31537 -13322 32013 -13300
rect 33137 -13300 33149 -13288
rect 33601 -13288 34749 -13282
rect 33601 -13300 33613 -13288
rect 33137 -13322 33613 -13300
rect 34737 -13300 34749 -13288
rect 35201 -13288 36349 -13282
rect 35201 -13300 35213 -13288
rect 34737 -13322 35213 -13300
rect 36337 -13300 36349 -13288
rect 36801 -13288 37949 -13282
rect 36801 -13300 36813 -13288
rect 36337 -13322 36813 -13300
rect 37937 -13322 37949 -13288
rect 0 -13420 490 -13322
rect 440 -13564 490 -13420
rect 57 -13570 490 -13564
rect 57 -13604 69 -13570
rect 445 -13604 490 -13570
rect 57 -13610 490 -13604
rect -30 -13657 16 -13645
rect -30 -13775 -24 -13657
rect 10 -13775 16 -13657
rect -30 -13787 16 -13775
rect 440 -13822 490 -13610
rect 670 -13328 37949 -13322
rect 670 -13420 37940 -13328
rect 670 -13564 720 -13420
rect 1200 -13470 1340 -13460
rect 670 -13570 1093 -13564
rect 670 -13604 705 -13570
rect 1081 -13604 1093 -13570
rect 1200 -13590 1210 -13470
rect 1330 -13480 1340 -13470
rect 2800 -13470 2940 -13460
rect 2800 -13480 2810 -13470
rect 1330 -13570 2810 -13480
rect 1330 -13580 1669 -13570
rect 1330 -13590 1340 -13580
rect 1200 -13600 1340 -13590
rect 670 -13610 1093 -13604
rect 1657 -13604 1669 -13580
rect 2045 -13580 2305 -13570
rect 2045 -13604 2057 -13580
rect 1657 -13610 2057 -13604
rect 2293 -13604 2305 -13580
rect 2681 -13580 2810 -13570
rect 2681 -13604 2693 -13580
rect 2800 -13590 2810 -13580
rect 2930 -13480 2940 -13470
rect 4400 -13470 4540 -13460
rect 4400 -13480 4410 -13470
rect 2930 -13570 4410 -13480
rect 2930 -13580 3269 -13570
rect 2930 -13590 2940 -13580
rect 2800 -13600 2940 -13590
rect 2293 -13610 2693 -13604
rect 3257 -13604 3269 -13580
rect 3645 -13580 3905 -13570
rect 3645 -13604 3657 -13580
rect 3257 -13610 3657 -13604
rect 3893 -13604 3905 -13580
rect 4281 -13580 4410 -13570
rect 4281 -13604 4293 -13580
rect 4400 -13590 4410 -13580
rect 4530 -13480 4540 -13470
rect 6000 -13470 6140 -13460
rect 6000 -13480 6010 -13470
rect 4530 -13570 6010 -13480
rect 4530 -13580 4869 -13570
rect 4530 -13590 4540 -13580
rect 4400 -13600 4540 -13590
rect 3893 -13610 4293 -13604
rect 4857 -13604 4869 -13580
rect 5245 -13580 5505 -13570
rect 5245 -13604 5257 -13580
rect 4857 -13610 5257 -13604
rect 5493 -13604 5505 -13580
rect 5881 -13580 6010 -13570
rect 5881 -13604 5893 -13580
rect 6000 -13590 6010 -13580
rect 6130 -13480 6140 -13470
rect 7600 -13470 7740 -13460
rect 7600 -13480 7610 -13470
rect 6130 -13570 7610 -13480
rect 6130 -13580 6469 -13570
rect 6130 -13590 6140 -13580
rect 6000 -13600 6140 -13590
rect 5493 -13610 5893 -13604
rect 6457 -13604 6469 -13580
rect 6845 -13580 7105 -13570
rect 6845 -13604 6857 -13580
rect 6457 -13610 6857 -13604
rect 7093 -13604 7105 -13580
rect 7481 -13580 7610 -13570
rect 7481 -13604 7493 -13580
rect 7600 -13590 7610 -13580
rect 7730 -13480 7740 -13470
rect 9200 -13470 9340 -13460
rect 15820 -13470 15960 -13460
rect 9200 -13480 9210 -13470
rect 7730 -13570 9210 -13480
rect 7730 -13580 8069 -13570
rect 7730 -13590 7740 -13580
rect 7600 -13600 7740 -13590
rect 7093 -13610 7493 -13604
rect 8057 -13604 8069 -13580
rect 8445 -13580 8705 -13570
rect 8445 -13604 8457 -13580
rect 8057 -13610 8457 -13604
rect 8693 -13604 8705 -13580
rect 9081 -13580 9210 -13570
rect 9081 -13604 9093 -13580
rect 9200 -13590 9210 -13580
rect 9330 -13480 9340 -13470
rect 14000 -13480 14140 -13470
rect 9330 -13570 10700 -13480
rect 14000 -13520 14010 -13480
rect 12860 -13564 14010 -13520
rect 9330 -13580 9669 -13570
rect 9330 -13590 9340 -13580
rect 9200 -13600 9340 -13590
rect 8693 -13610 9093 -13604
rect 9657 -13604 9669 -13580
rect 10045 -13580 10305 -13570
rect 10045 -13604 10057 -13580
rect 9657 -13610 10057 -13604
rect 10293 -13604 10305 -13580
rect 10681 -13580 10700 -13570
rect 11257 -13570 11657 -13564
rect 10681 -13604 10693 -13580
rect 10293 -13610 10693 -13604
rect 11257 -13604 11269 -13570
rect 11645 -13604 11657 -13570
rect 11257 -13610 11657 -13604
rect 11893 -13570 12293 -13564
rect 11893 -13604 11905 -13570
rect 12281 -13604 12293 -13570
rect 11893 -13610 12293 -13604
rect 12857 -13570 14010 -13564
rect 12857 -13604 12869 -13570
rect 13245 -13600 13505 -13570
rect 13245 -13604 13257 -13600
rect 12857 -13610 13257 -13604
rect 13493 -13604 13505 -13600
rect 13881 -13600 14010 -13570
rect 14130 -13520 14140 -13480
rect 14130 -13564 15490 -13520
rect 14130 -13570 15493 -13564
rect 14130 -13600 14469 -13570
rect 13881 -13604 13893 -13600
rect 13493 -13610 13893 -13604
rect 14000 -13610 14140 -13600
rect 14457 -13604 14469 -13600
rect 14845 -13600 15105 -13570
rect 14845 -13604 14857 -13600
rect 14457 -13610 14857 -13604
rect 15093 -13604 15105 -13600
rect 15481 -13604 15493 -13570
rect 15820 -13590 15830 -13470
rect 15950 -13500 15960 -13470
rect 17420 -13470 17560 -13460
rect 15950 -13564 17090 -13500
rect 15950 -13570 17093 -13564
rect 15950 -13590 16069 -13570
rect 15820 -13600 16069 -13590
rect 15093 -13610 15493 -13604
rect 16057 -13604 16069 -13600
rect 16445 -13600 16705 -13570
rect 16445 -13604 16457 -13600
rect 16057 -13610 16457 -13604
rect 16693 -13604 16705 -13600
rect 17081 -13604 17093 -13570
rect 17420 -13590 17430 -13470
rect 17550 -13500 17560 -13470
rect 19020 -13470 19160 -13460
rect 17550 -13564 18690 -13500
rect 17550 -13570 18693 -13564
rect 17550 -13590 17669 -13570
rect 17420 -13600 17669 -13590
rect 16693 -13610 17093 -13604
rect 17657 -13604 17669 -13600
rect 18045 -13600 18305 -13570
rect 18045 -13604 18057 -13600
rect 17657 -13610 18057 -13604
rect 18293 -13604 18305 -13600
rect 18681 -13604 18693 -13570
rect 19020 -13590 19030 -13470
rect 19150 -13500 19160 -13470
rect 20620 -13470 20760 -13460
rect 19150 -13564 20290 -13500
rect 19150 -13570 20293 -13564
rect 19150 -13590 19269 -13570
rect 19020 -13600 19269 -13590
rect 18293 -13610 18693 -13604
rect 19257 -13604 19269 -13600
rect 19645 -13600 19905 -13570
rect 19645 -13604 19657 -13600
rect 19257 -13610 19657 -13604
rect 19893 -13604 19905 -13600
rect 20281 -13604 20293 -13570
rect 20620 -13590 20630 -13470
rect 20750 -13500 20760 -13470
rect 22220 -13470 22360 -13460
rect 20750 -13564 21890 -13500
rect 20750 -13570 21893 -13564
rect 20750 -13590 20869 -13570
rect 20620 -13600 20869 -13590
rect 19893 -13610 20293 -13604
rect 20857 -13604 20869 -13600
rect 21245 -13600 21505 -13570
rect 21245 -13604 21257 -13600
rect 20857 -13610 21257 -13604
rect 21493 -13604 21505 -13600
rect 21881 -13604 21893 -13570
rect 22220 -13590 22230 -13470
rect 22350 -13500 22360 -13470
rect 23820 -13470 23960 -13460
rect 22350 -13564 23490 -13500
rect 22350 -13570 23493 -13564
rect 22350 -13590 22469 -13570
rect 22220 -13600 22469 -13590
rect 21493 -13610 21893 -13604
rect 22457 -13604 22469 -13600
rect 22845 -13600 23105 -13570
rect 22845 -13604 22857 -13600
rect 22457 -13610 22857 -13604
rect 23093 -13604 23105 -13600
rect 23481 -13604 23493 -13570
rect 23820 -13590 23830 -13470
rect 23950 -13500 23960 -13470
rect 25420 -13470 25560 -13460
rect 23950 -13564 25090 -13500
rect 23950 -13570 25093 -13564
rect 23950 -13590 24069 -13570
rect 23820 -13600 24069 -13590
rect 23093 -13610 23493 -13604
rect 24057 -13604 24069 -13600
rect 24445 -13600 24705 -13570
rect 24445 -13604 24457 -13600
rect 24057 -13610 24457 -13604
rect 24693 -13604 24705 -13600
rect 25081 -13604 25093 -13570
rect 25420 -13590 25430 -13470
rect 25550 -13500 25560 -13470
rect 27020 -13470 27160 -13460
rect 25550 -13564 26680 -13500
rect 25550 -13570 26693 -13564
rect 25550 -13590 25669 -13570
rect 25420 -13600 25669 -13590
rect 24693 -13610 25093 -13604
rect 25657 -13604 25669 -13600
rect 26045 -13600 26305 -13570
rect 26045 -13604 26057 -13600
rect 25657 -13610 26057 -13604
rect 26293 -13604 26305 -13600
rect 26681 -13604 26693 -13570
rect 27020 -13590 27030 -13470
rect 27150 -13500 27160 -13470
rect 28620 -13470 28760 -13460
rect 27150 -13564 28290 -13500
rect 27150 -13570 28293 -13564
rect 27150 -13590 27269 -13570
rect 27020 -13600 27269 -13590
rect 26293 -13610 26693 -13604
rect 27257 -13604 27269 -13600
rect 27645 -13600 27905 -13570
rect 27645 -13604 27657 -13600
rect 27257 -13610 27657 -13604
rect 27893 -13604 27905 -13600
rect 28281 -13604 28293 -13570
rect 28620 -13590 28630 -13470
rect 28750 -13500 28760 -13470
rect 30220 -13470 30360 -13460
rect 28750 -13564 29890 -13500
rect 28750 -13570 29893 -13564
rect 28750 -13590 28869 -13570
rect 28620 -13600 28869 -13590
rect 27893 -13610 28293 -13604
rect 28857 -13604 28869 -13600
rect 29245 -13600 29505 -13570
rect 29245 -13604 29257 -13600
rect 28857 -13610 29257 -13604
rect 29493 -13604 29505 -13600
rect 29881 -13604 29893 -13570
rect 30220 -13590 30230 -13470
rect 30350 -13500 30360 -13470
rect 31820 -13470 31960 -13460
rect 30350 -13564 31490 -13500
rect 30350 -13570 31493 -13564
rect 30350 -13590 30469 -13570
rect 30220 -13600 30469 -13590
rect 29493 -13610 29893 -13604
rect 30457 -13604 30469 -13600
rect 30845 -13600 31105 -13570
rect 30845 -13604 30857 -13600
rect 30457 -13610 30857 -13604
rect 31093 -13604 31105 -13600
rect 31481 -13604 31493 -13570
rect 31820 -13590 31830 -13470
rect 31950 -13500 31960 -13470
rect 34800 -13470 34940 -13460
rect 34800 -13500 34810 -13470
rect 31950 -13570 34810 -13500
rect 31950 -13590 32069 -13570
rect 31820 -13600 32069 -13590
rect 31093 -13610 31493 -13604
rect 32057 -13604 32069 -13600
rect 32445 -13600 32705 -13570
rect 32445 -13604 32457 -13600
rect 32057 -13610 32457 -13604
rect 32693 -13604 32705 -13600
rect 33081 -13600 33669 -13570
rect 33081 -13604 33093 -13600
rect 32693 -13610 33093 -13604
rect 33657 -13604 33669 -13600
rect 34045 -13600 34305 -13570
rect 34045 -13604 34057 -13600
rect 33657 -13610 34057 -13604
rect 34293 -13604 34305 -13600
rect 34681 -13590 34810 -13570
rect 34930 -13500 34940 -13470
rect 34930 -13564 36280 -13500
rect 34930 -13570 36293 -13564
rect 34930 -13590 35269 -13570
rect 34681 -13600 35269 -13590
rect 34681 -13604 34693 -13600
rect 34293 -13610 34693 -13604
rect 35257 -13604 35269 -13600
rect 35645 -13600 35905 -13570
rect 35645 -13604 35657 -13600
rect 35257 -13610 35657 -13604
rect 35893 -13604 35905 -13600
rect 36281 -13604 36293 -13570
rect 35893 -13610 36293 -13604
rect 36857 -13570 37257 -13564
rect 36857 -13604 36869 -13570
rect 37245 -13604 37257 -13570
rect 36857 -13610 37257 -13604
rect 37493 -13570 37893 -13564
rect 37493 -13604 37505 -13570
rect 37881 -13604 37893 -13570
rect 37493 -13610 37893 -13604
rect 57 -13828 490 -13822
rect 57 -13862 69 -13828
rect 445 -13862 490 -13828
rect 57 -13868 490 -13862
rect 440 -14090 490 -13868
rect 57 -14096 490 -14090
rect 57 -14130 69 -14096
rect 445 -14130 490 -14096
rect 57 -14136 490 -14130
rect -30 -14196 16 -14184
rect -30 -14888 -24 -14196
rect 10 -14888 16 -14196
rect -30 -14900 16 -14888
rect 440 -14948 490 -14136
rect 670 -13822 720 -13610
rect 1134 -13657 1180 -13645
rect 1134 -13775 1140 -13657
rect 1174 -13775 1180 -13657
rect 1570 -13657 1616 -13645
rect 1570 -13660 1576 -13657
rect 1134 -13787 1180 -13775
rect 1560 -13775 1576 -13660
rect 1610 -13660 1616 -13657
rect 2098 -13657 2144 -13645
rect 2098 -13660 2104 -13657
rect 1610 -13775 2104 -13660
rect 2138 -13660 2144 -13657
rect 2206 -13657 2252 -13645
rect 2206 -13660 2212 -13657
rect 2138 -13775 2212 -13660
rect 2246 -13660 2252 -13657
rect 2734 -13657 2780 -13645
rect 2734 -13660 2740 -13657
rect 2246 -13775 2740 -13660
rect 2774 -13660 2780 -13657
rect 3170 -13657 3216 -13645
rect 3170 -13660 3176 -13657
rect 2774 -13775 3176 -13660
rect 3210 -13660 3216 -13657
rect 3698 -13657 3744 -13645
rect 3698 -13660 3704 -13657
rect 3210 -13775 3704 -13660
rect 3738 -13660 3744 -13657
rect 3806 -13657 3852 -13645
rect 3806 -13660 3812 -13657
rect 3738 -13775 3812 -13660
rect 3846 -13660 3852 -13657
rect 4334 -13657 4380 -13645
rect 4334 -13660 4340 -13657
rect 3846 -13775 4340 -13660
rect 4374 -13660 4380 -13657
rect 4770 -13657 4816 -13645
rect 4770 -13660 4776 -13657
rect 4374 -13775 4776 -13660
rect 4810 -13660 4816 -13657
rect 5298 -13657 5344 -13645
rect 5298 -13660 5304 -13657
rect 4810 -13775 5304 -13660
rect 5338 -13660 5344 -13657
rect 5406 -13657 5452 -13645
rect 5406 -13660 5412 -13657
rect 5338 -13775 5412 -13660
rect 5446 -13660 5452 -13657
rect 5934 -13657 5980 -13645
rect 5934 -13660 5940 -13657
rect 5446 -13775 5940 -13660
rect 5974 -13660 5980 -13657
rect 6370 -13657 6416 -13645
rect 6370 -13660 6376 -13657
rect 5974 -13775 6376 -13660
rect 6410 -13660 6416 -13657
rect 6898 -13657 6944 -13645
rect 6898 -13660 6904 -13657
rect 6410 -13775 6904 -13660
rect 6938 -13660 6944 -13657
rect 7006 -13657 7052 -13645
rect 7006 -13660 7012 -13657
rect 6938 -13775 7012 -13660
rect 7046 -13660 7052 -13657
rect 7534 -13657 7580 -13645
rect 7534 -13660 7540 -13657
rect 7046 -13775 7540 -13660
rect 7574 -13660 7580 -13657
rect 7970 -13657 8016 -13645
rect 7970 -13660 7976 -13657
rect 7574 -13775 7976 -13660
rect 8010 -13660 8016 -13657
rect 8498 -13657 8544 -13645
rect 8498 -13660 8504 -13657
rect 8010 -13775 8504 -13660
rect 8538 -13660 8544 -13657
rect 8606 -13657 8652 -13645
rect 8606 -13660 8612 -13657
rect 8538 -13775 8612 -13660
rect 8646 -13660 8652 -13657
rect 9134 -13657 9180 -13645
rect 9134 -13660 9140 -13657
rect 8646 -13775 9140 -13660
rect 9174 -13660 9180 -13657
rect 9570 -13657 9616 -13645
rect 9570 -13660 9576 -13657
rect 9174 -13775 9576 -13660
rect 9610 -13660 9616 -13657
rect 10098 -13657 10144 -13645
rect 10098 -13660 10104 -13657
rect 9610 -13775 10104 -13660
rect 10138 -13660 10144 -13657
rect 10206 -13657 10252 -13645
rect 10206 -13660 10212 -13657
rect 10138 -13775 10212 -13660
rect 10246 -13660 10252 -13657
rect 10734 -13650 10780 -13645
rect 10734 -13657 10940 -13650
rect 10734 -13660 10740 -13657
rect 10246 -13775 10740 -13660
rect 10774 -13660 10940 -13657
rect 11170 -13657 11216 -13645
rect 11170 -13660 11176 -13657
rect 10774 -13775 10810 -13660
rect 1560 -13780 10810 -13775
rect 10930 -13775 11176 -13660
rect 11210 -13660 11216 -13657
rect 11400 -13660 11520 -13610
rect 11698 -13657 11744 -13645
rect 11698 -13660 11704 -13657
rect 11210 -13775 11704 -13660
rect 11738 -13660 11744 -13657
rect 11806 -13657 11852 -13645
rect 11806 -13660 11812 -13657
rect 11738 -13775 11812 -13660
rect 11846 -13660 11852 -13657
rect 12040 -13660 12160 -13610
rect 12334 -13657 12380 -13645
rect 12334 -13660 12340 -13657
rect 11846 -13775 12340 -13660
rect 12374 -13660 12380 -13657
rect 12770 -13657 12816 -13645
rect 12770 -13660 12776 -13657
rect 12374 -13775 12776 -13660
rect 12810 -13660 12816 -13657
rect 13298 -13657 13344 -13645
rect 13298 -13660 13304 -13657
rect 12810 -13775 13304 -13660
rect 13338 -13660 13344 -13657
rect 13406 -13657 13452 -13645
rect 13406 -13660 13412 -13657
rect 13338 -13775 13412 -13660
rect 13446 -13660 13452 -13657
rect 13934 -13657 13980 -13645
rect 13934 -13660 13940 -13657
rect 13446 -13775 13940 -13660
rect 13974 -13660 13980 -13657
rect 14370 -13657 14416 -13645
rect 14370 -13660 14376 -13657
rect 13974 -13775 14376 -13660
rect 14410 -13660 14416 -13657
rect 14898 -13657 14944 -13645
rect 14898 -13660 14904 -13657
rect 14410 -13775 14904 -13660
rect 14938 -13660 14944 -13657
rect 15006 -13657 15052 -13645
rect 15006 -13660 15012 -13657
rect 14938 -13775 15012 -13660
rect 15046 -13660 15052 -13657
rect 15534 -13657 15580 -13645
rect 15534 -13660 15540 -13657
rect 15046 -13775 15540 -13660
rect 15574 -13660 15580 -13657
rect 15970 -13657 16016 -13645
rect 15970 -13660 15976 -13657
rect 15574 -13775 15976 -13660
rect 16010 -13660 16016 -13657
rect 16498 -13657 16544 -13645
rect 16498 -13660 16504 -13657
rect 16010 -13775 16504 -13660
rect 16538 -13660 16544 -13657
rect 16606 -13657 16652 -13645
rect 16606 -13660 16612 -13657
rect 16538 -13775 16612 -13660
rect 16646 -13660 16652 -13657
rect 17134 -13657 17180 -13645
rect 17134 -13660 17140 -13657
rect 16646 -13775 17140 -13660
rect 17174 -13660 17180 -13657
rect 17570 -13657 17616 -13645
rect 17570 -13660 17576 -13657
rect 17174 -13775 17576 -13660
rect 17610 -13660 17616 -13657
rect 18098 -13657 18144 -13645
rect 18098 -13660 18104 -13657
rect 17610 -13775 18104 -13660
rect 18138 -13660 18144 -13657
rect 18206 -13657 18252 -13645
rect 18206 -13660 18212 -13657
rect 18138 -13775 18212 -13660
rect 18246 -13660 18252 -13657
rect 18734 -13657 18780 -13645
rect 18734 -13660 18740 -13657
rect 18246 -13775 18740 -13660
rect 18774 -13660 18780 -13657
rect 19170 -13657 19216 -13645
rect 19170 -13660 19176 -13657
rect 18774 -13775 19176 -13660
rect 19210 -13660 19216 -13657
rect 19698 -13657 19744 -13645
rect 19698 -13660 19704 -13657
rect 19210 -13775 19704 -13660
rect 19738 -13660 19744 -13657
rect 19806 -13657 19852 -13645
rect 19806 -13660 19812 -13657
rect 19738 -13775 19812 -13660
rect 19846 -13660 19852 -13657
rect 20334 -13657 20380 -13645
rect 20334 -13660 20340 -13657
rect 19846 -13775 20340 -13660
rect 20374 -13660 20380 -13657
rect 20770 -13657 20816 -13645
rect 20770 -13660 20776 -13657
rect 20374 -13775 20776 -13660
rect 20810 -13660 20816 -13657
rect 21298 -13657 21344 -13645
rect 21298 -13660 21304 -13657
rect 20810 -13775 21304 -13660
rect 21338 -13660 21344 -13657
rect 21406 -13657 21452 -13645
rect 21406 -13660 21412 -13657
rect 21338 -13775 21412 -13660
rect 21446 -13660 21452 -13657
rect 21934 -13657 21980 -13645
rect 21934 -13660 21940 -13657
rect 21446 -13775 21940 -13660
rect 21974 -13660 21980 -13657
rect 22370 -13657 22416 -13645
rect 22370 -13660 22376 -13657
rect 21974 -13775 22376 -13660
rect 22410 -13660 22416 -13657
rect 22898 -13657 22944 -13645
rect 22898 -13660 22904 -13657
rect 22410 -13775 22904 -13660
rect 22938 -13660 22944 -13657
rect 23006 -13657 23052 -13645
rect 23006 -13660 23012 -13657
rect 22938 -13775 23012 -13660
rect 23046 -13660 23052 -13657
rect 23534 -13657 23580 -13645
rect 23534 -13660 23540 -13657
rect 23046 -13775 23540 -13660
rect 23574 -13660 23580 -13657
rect 23970 -13657 24016 -13645
rect 23970 -13660 23976 -13657
rect 23574 -13775 23976 -13660
rect 24010 -13660 24016 -13657
rect 24498 -13657 24544 -13645
rect 24498 -13660 24504 -13657
rect 24010 -13775 24504 -13660
rect 24538 -13660 24544 -13657
rect 24606 -13657 24652 -13645
rect 24606 -13660 24612 -13657
rect 24538 -13775 24612 -13660
rect 24646 -13660 24652 -13657
rect 25134 -13657 25180 -13645
rect 25134 -13660 25140 -13657
rect 24646 -13775 25140 -13660
rect 25174 -13660 25180 -13657
rect 25570 -13657 25616 -13645
rect 25570 -13660 25576 -13657
rect 25174 -13775 25576 -13660
rect 25610 -13660 25616 -13657
rect 26098 -13657 26144 -13645
rect 26098 -13660 26104 -13657
rect 25610 -13775 26104 -13660
rect 26138 -13660 26144 -13657
rect 26206 -13657 26252 -13645
rect 26206 -13660 26212 -13657
rect 26138 -13775 26212 -13660
rect 26246 -13660 26252 -13657
rect 26734 -13657 26780 -13645
rect 26734 -13660 26740 -13657
rect 26246 -13775 26740 -13660
rect 26774 -13660 26780 -13657
rect 27170 -13657 27216 -13645
rect 27170 -13660 27176 -13657
rect 26774 -13775 27176 -13660
rect 27210 -13660 27216 -13657
rect 27698 -13657 27744 -13645
rect 27698 -13660 27704 -13657
rect 27210 -13775 27704 -13660
rect 27738 -13660 27744 -13657
rect 27806 -13657 27852 -13645
rect 27806 -13660 27812 -13657
rect 27738 -13775 27812 -13660
rect 27846 -13660 27852 -13657
rect 28334 -13657 28380 -13645
rect 28334 -13660 28340 -13657
rect 27846 -13775 28340 -13660
rect 28374 -13660 28380 -13657
rect 28770 -13657 28816 -13645
rect 28770 -13660 28776 -13657
rect 28374 -13775 28776 -13660
rect 28810 -13660 28816 -13657
rect 29298 -13657 29344 -13645
rect 29298 -13660 29304 -13657
rect 28810 -13775 29304 -13660
rect 29338 -13660 29344 -13657
rect 29406 -13657 29452 -13645
rect 29406 -13660 29412 -13657
rect 29338 -13775 29412 -13660
rect 29446 -13660 29452 -13657
rect 29934 -13657 29980 -13645
rect 29934 -13660 29940 -13657
rect 29446 -13775 29940 -13660
rect 29974 -13660 29980 -13657
rect 30370 -13657 30416 -13637
rect 30370 -13660 30376 -13657
rect 29974 -13775 30376 -13660
rect 30410 -13660 30416 -13657
rect 30898 -13657 30944 -13637
rect 30898 -13660 30904 -13657
rect 30410 -13775 30904 -13660
rect 30938 -13660 30944 -13657
rect 31006 -13657 31052 -13637
rect 31006 -13660 31012 -13657
rect 30938 -13775 31012 -13660
rect 31046 -13660 31052 -13657
rect 31534 -13657 31580 -13645
rect 31534 -13660 31540 -13657
rect 31046 -13775 31540 -13660
rect 31574 -13660 31580 -13657
rect 31970 -13657 32016 -13645
rect 31970 -13660 31976 -13657
rect 31574 -13775 31976 -13660
rect 32010 -13660 32016 -13657
rect 32498 -13657 32544 -13645
rect 32498 -13660 32504 -13657
rect 32010 -13775 32504 -13660
rect 32538 -13660 32544 -13657
rect 32606 -13657 32652 -13645
rect 32606 -13660 32612 -13657
rect 32538 -13775 32612 -13660
rect 32646 -13660 32652 -13657
rect 33134 -13657 33180 -13645
rect 33134 -13660 33140 -13657
rect 32646 -13775 33140 -13660
rect 33174 -13660 33180 -13657
rect 33570 -13657 33616 -13645
rect 33570 -13660 33576 -13657
rect 33174 -13775 33576 -13660
rect 33610 -13660 33616 -13657
rect 34098 -13657 34144 -13645
rect 34098 -13660 34104 -13657
rect 33610 -13775 34104 -13660
rect 34138 -13660 34144 -13657
rect 34206 -13657 34252 -13645
rect 34206 -13660 34212 -13657
rect 34138 -13775 34212 -13660
rect 34246 -13660 34252 -13657
rect 34734 -13657 34780 -13645
rect 34734 -13660 34740 -13657
rect 34246 -13775 34740 -13660
rect 34774 -13660 34780 -13657
rect 35170 -13657 35216 -13645
rect 35170 -13660 35176 -13657
rect 34774 -13775 35176 -13660
rect 35210 -13660 35216 -13657
rect 35698 -13657 35744 -13645
rect 35698 -13660 35704 -13657
rect 35210 -13775 35704 -13660
rect 35738 -13660 35744 -13657
rect 35806 -13657 35852 -13645
rect 35806 -13660 35812 -13657
rect 35738 -13775 35812 -13660
rect 35846 -13660 35852 -13657
rect 36334 -13657 36380 -13645
rect 36334 -13660 36340 -13657
rect 35846 -13775 36340 -13660
rect 36374 -13775 36380 -13657
rect 10930 -13780 36380 -13775
rect 1570 -13787 1616 -13780
rect 2098 -13787 2144 -13780
rect 2206 -13787 2252 -13780
rect 2734 -13787 2780 -13780
rect 3170 -13787 3216 -13780
rect 3698 -13787 3744 -13780
rect 3806 -13787 3852 -13780
rect 4334 -13787 4380 -13780
rect 4770 -13787 4816 -13780
rect 5298 -13787 5344 -13780
rect 5406 -13787 5452 -13780
rect 5934 -13787 5980 -13780
rect 6370 -13787 6416 -13780
rect 6898 -13787 6944 -13780
rect 7006 -13787 7052 -13780
rect 7534 -13787 7580 -13780
rect 7970 -13787 8016 -13780
rect 8498 -13787 8544 -13780
rect 8606 -13787 8652 -13780
rect 9134 -13787 9180 -13780
rect 9570 -13787 9616 -13780
rect 10098 -13787 10144 -13780
rect 10206 -13787 10252 -13780
rect 10734 -13787 10940 -13780
rect 11170 -13787 11216 -13780
rect 10750 -13790 10940 -13787
rect 11400 -13822 11520 -13780
rect 11698 -13787 11744 -13780
rect 11806 -13787 11852 -13780
rect 12040 -13822 12160 -13780
rect 12334 -13787 12380 -13780
rect 12770 -13787 12816 -13780
rect 13298 -13787 13344 -13780
rect 13406 -13787 13452 -13780
rect 13934 -13787 13980 -13780
rect 14370 -13787 14416 -13780
rect 14898 -13787 14944 -13780
rect 15006 -13787 15052 -13780
rect 15534 -13787 15580 -13780
rect 15970 -13787 16016 -13780
rect 16498 -13787 16544 -13780
rect 16606 -13787 16652 -13780
rect 17134 -13787 17180 -13780
rect 17570 -13787 17616 -13780
rect 18098 -13787 18144 -13780
rect 18206 -13787 18252 -13780
rect 18734 -13787 18780 -13780
rect 19170 -13787 19216 -13780
rect 19698 -13787 19744 -13780
rect 19806 -13787 19852 -13780
rect 20334 -13787 20380 -13780
rect 20770 -13787 20816 -13780
rect 21298 -13787 21344 -13780
rect 21406 -13787 21452 -13780
rect 21934 -13787 21980 -13780
rect 22370 -13787 22416 -13780
rect 22898 -13787 22944 -13780
rect 23006 -13787 23052 -13780
rect 23534 -13787 23580 -13780
rect 23970 -13787 24016 -13780
rect 24498 -13787 24544 -13780
rect 24606 -13787 24652 -13780
rect 25134 -13787 25180 -13780
rect 25570 -13787 25616 -13780
rect 26098 -13787 26144 -13780
rect 26206 -13787 26252 -13780
rect 26734 -13787 26780 -13780
rect 27170 -13787 27216 -13780
rect 27698 -13787 27744 -13780
rect 27806 -13787 27852 -13780
rect 28334 -13787 28380 -13780
rect 28770 -13787 28816 -13780
rect 29298 -13787 29344 -13780
rect 29406 -13787 29452 -13780
rect 29934 -13787 29980 -13780
rect 30370 -13795 30416 -13780
rect 30898 -13795 30944 -13780
rect 31006 -13795 31052 -13780
rect 31534 -13787 31580 -13780
rect 31970 -13787 32016 -13780
rect 32498 -13787 32544 -13780
rect 32606 -13787 32652 -13780
rect 33134 -13787 33180 -13780
rect 33570 -13787 33616 -13780
rect 34098 -13787 34144 -13780
rect 34206 -13787 34252 -13780
rect 34734 -13787 34780 -13780
rect 35170 -13787 35216 -13780
rect 35698 -13787 35744 -13780
rect 35806 -13787 35852 -13780
rect 36334 -13787 36380 -13780
rect 36770 -13657 36816 -13645
rect 36770 -13775 36776 -13657
rect 36810 -13775 36816 -13657
rect 36770 -13787 36816 -13775
rect 37298 -13657 37344 -13645
rect 37298 -13775 37304 -13657
rect 37338 -13775 37344 -13657
rect 37298 -13787 37344 -13775
rect 37406 -13657 37452 -13645
rect 37406 -13775 37412 -13657
rect 37446 -13775 37452 -13657
rect 37406 -13787 37452 -13775
rect 37934 -13657 37980 -13645
rect 37934 -13775 37940 -13657
rect 37974 -13775 37980 -13657
rect 37934 -13787 37980 -13775
rect 670 -13828 1093 -13822
rect 670 -13862 705 -13828
rect 1081 -13862 1093 -13828
rect 670 -13868 1093 -13862
rect 1657 -13828 2057 -13822
rect 1657 -13862 1669 -13828
rect 2045 -13830 2057 -13828
rect 2293 -13828 2693 -13822
rect 2293 -13830 2305 -13828
rect 2045 -13862 2060 -13830
rect 1657 -13868 2060 -13862
rect 670 -14090 720 -13868
rect 1420 -13910 1560 -13900
rect 1420 -14030 1430 -13910
rect 1550 -13920 1560 -13910
rect 1660 -13920 2060 -13868
rect 2290 -13862 2305 -13830
rect 2681 -13862 2693 -13828
rect 2290 -13868 2693 -13862
rect 3257 -13828 3657 -13822
rect 3257 -13862 3269 -13828
rect 3645 -13830 3657 -13828
rect 3893 -13828 4293 -13822
rect 3893 -13830 3905 -13828
rect 3645 -13862 3660 -13830
rect 3257 -13868 3660 -13862
rect 2290 -13920 2690 -13868
rect 3020 -13910 3160 -13900
rect 3020 -13920 3030 -13910
rect 1550 -14020 3030 -13920
rect 1550 -14030 1560 -14020
rect 1420 -14040 1560 -14030
rect 1660 -14040 2690 -14020
rect 3020 -14030 3030 -14020
rect 3150 -13920 3160 -13910
rect 3260 -13920 3660 -13868
rect 3890 -13862 3905 -13830
rect 4281 -13862 4293 -13828
rect 3890 -13868 4293 -13862
rect 4857 -13828 5257 -13822
rect 4857 -13862 4869 -13828
rect 5245 -13830 5257 -13828
rect 5493 -13828 5893 -13822
rect 5493 -13830 5505 -13828
rect 5245 -13862 5260 -13830
rect 4857 -13868 5260 -13862
rect 3890 -13920 4290 -13868
rect 4620 -13910 4760 -13900
rect 4620 -13920 4630 -13910
rect 3150 -14020 4630 -13920
rect 3150 -14030 3160 -14020
rect 3020 -14040 3160 -14030
rect 3260 -14040 4290 -14020
rect 4620 -14030 4630 -14020
rect 4750 -13920 4760 -13910
rect 4860 -13920 5260 -13868
rect 5490 -13862 5505 -13830
rect 5881 -13862 5893 -13828
rect 5490 -13868 5893 -13862
rect 6457 -13828 6857 -13822
rect 6457 -13862 6469 -13828
rect 6845 -13830 6857 -13828
rect 7093 -13828 7493 -13822
rect 7093 -13830 7105 -13828
rect 6845 -13862 6860 -13830
rect 6457 -13868 6860 -13862
rect 5490 -13920 5890 -13868
rect 6220 -13910 6360 -13900
rect 6220 -13920 6230 -13910
rect 4750 -14020 6230 -13920
rect 4750 -14030 4760 -14020
rect 4620 -14040 4760 -14030
rect 4860 -14040 5890 -14020
rect 6220 -14030 6230 -14020
rect 6350 -13920 6360 -13910
rect 6460 -13920 6860 -13868
rect 7090 -13862 7105 -13830
rect 7481 -13862 7493 -13828
rect 7090 -13868 7493 -13862
rect 8057 -13828 8457 -13822
rect 8057 -13862 8069 -13828
rect 8445 -13830 8457 -13828
rect 8693 -13828 9093 -13822
rect 8693 -13830 8705 -13828
rect 8445 -13862 8460 -13830
rect 8057 -13868 8460 -13862
rect 7090 -13920 7490 -13868
rect 7820 -13910 7960 -13900
rect 7820 -13920 7830 -13910
rect 6350 -14020 7830 -13920
rect 6350 -14030 6360 -14020
rect 6220 -14040 6360 -14030
rect 6460 -14040 7490 -14020
rect 7820 -14030 7830 -14020
rect 7950 -13920 7960 -13910
rect 8060 -13920 8460 -13868
rect 8690 -13862 8705 -13830
rect 9081 -13862 9093 -13828
rect 8690 -13868 9093 -13862
rect 9657 -13828 10057 -13822
rect 9657 -13862 9669 -13828
rect 10045 -13830 10057 -13828
rect 10293 -13828 10693 -13822
rect 10293 -13830 10305 -13828
rect 10045 -13862 10060 -13830
rect 9657 -13868 10060 -13862
rect 8690 -13920 9090 -13868
rect 9420 -13910 9560 -13900
rect 9420 -13920 9430 -13910
rect 7950 -14020 9430 -13920
rect 7950 -14030 7960 -14020
rect 7820 -14040 7960 -14030
rect 8060 -14040 9090 -14020
rect 9420 -14030 9430 -14020
rect 9550 -13920 9560 -13910
rect 9660 -13920 10060 -13868
rect 10290 -13862 10305 -13830
rect 10681 -13862 10693 -13828
rect 10290 -13868 10693 -13862
rect 11257 -13828 11657 -13822
rect 11257 -13862 11269 -13828
rect 11645 -13862 11657 -13828
rect 11257 -13868 11657 -13862
rect 11893 -13828 12293 -13822
rect 11893 -13862 11905 -13828
rect 12281 -13862 12293 -13828
rect 11893 -13868 12293 -13862
rect 12857 -13828 13257 -13822
rect 12857 -13862 12869 -13828
rect 13245 -13830 13257 -13828
rect 13493 -13828 13893 -13822
rect 13493 -13830 13505 -13828
rect 13245 -13862 13260 -13830
rect 12857 -13868 13260 -13862
rect 10290 -13920 10690 -13868
rect 9550 -14020 10690 -13920
rect 9550 -14030 9560 -14020
rect 9420 -14040 9560 -14030
rect 9660 -14040 10690 -14020
rect 1660 -14090 2060 -14040
rect 670 -14096 1093 -14090
rect 670 -14130 705 -14096
rect 1081 -14130 1093 -14096
rect 670 -14136 1093 -14130
rect 1657 -14096 2060 -14090
rect 1657 -14130 1669 -14096
rect 2045 -14130 2060 -14096
rect 2290 -14090 2690 -14040
rect 3260 -14090 3660 -14040
rect 2290 -14096 2693 -14090
rect 2290 -14130 2305 -14096
rect 2681 -14130 2693 -14096
rect 1657 -14136 2057 -14130
rect 2293 -14136 2693 -14130
rect 3257 -14096 3660 -14090
rect 3257 -14130 3269 -14096
rect 3645 -14130 3660 -14096
rect 3890 -14090 4290 -14040
rect 4860 -14090 5260 -14040
rect 3890 -14096 4293 -14090
rect 3890 -14130 3905 -14096
rect 4281 -14130 4293 -14096
rect 3257 -14136 3657 -14130
rect 3893 -14136 4293 -14130
rect 4857 -14096 5260 -14090
rect 4857 -14130 4869 -14096
rect 5245 -14130 5260 -14096
rect 5490 -14090 5890 -14040
rect 6460 -14090 6860 -14040
rect 5490 -14096 5893 -14090
rect 5490 -14130 5505 -14096
rect 5881 -14130 5893 -14096
rect 4857 -14136 5257 -14130
rect 5493 -14136 5893 -14130
rect 6457 -14096 6860 -14090
rect 6457 -14130 6469 -14096
rect 6845 -14130 6860 -14096
rect 7090 -14090 7490 -14040
rect 8060 -14090 8460 -14040
rect 7090 -14096 7493 -14090
rect 7090 -14130 7105 -14096
rect 7481 -14130 7493 -14096
rect 6457 -14136 6857 -14130
rect 7093 -14136 7493 -14130
rect 8057 -14096 8460 -14090
rect 8057 -14130 8069 -14096
rect 8445 -14130 8460 -14096
rect 8690 -14090 9090 -14040
rect 9660 -14090 10060 -14040
rect 8690 -14096 9093 -14090
rect 8690 -14130 8705 -14096
rect 9081 -14130 9093 -14096
rect 8057 -14136 8457 -14130
rect 8693 -14136 9093 -14130
rect 9657 -14096 10060 -14090
rect 9657 -14130 9669 -14096
rect 10045 -14130 10060 -14096
rect 10290 -14090 10690 -14040
rect 12860 -13920 13260 -13868
rect 13490 -13862 13505 -13830
rect 13881 -13862 13893 -13828
rect 13490 -13868 13893 -13862
rect 14457 -13828 14857 -13822
rect 14457 -13862 14469 -13828
rect 14845 -13830 14857 -13828
rect 15093 -13828 15493 -13822
rect 15093 -13830 15105 -13828
rect 14845 -13862 14860 -13830
rect 14457 -13868 14860 -13862
rect 13490 -13920 13890 -13868
rect 14460 -13920 14860 -13868
rect 15090 -13862 15105 -13830
rect 15481 -13862 15493 -13828
rect 15090 -13868 15493 -13862
rect 16057 -13828 16457 -13822
rect 16057 -13862 16069 -13828
rect 16445 -13862 16457 -13828
rect 16057 -13868 16457 -13862
rect 16693 -13828 17093 -13822
rect 16693 -13862 16705 -13828
rect 17081 -13862 17093 -13828
rect 16693 -13868 17093 -13862
rect 17657 -13828 18057 -13822
rect 17657 -13862 17669 -13828
rect 18045 -13862 18057 -13828
rect 17657 -13868 18057 -13862
rect 18293 -13828 18693 -13822
rect 18293 -13862 18305 -13828
rect 18681 -13862 18693 -13828
rect 18293 -13868 18693 -13862
rect 19257 -13828 19657 -13822
rect 19257 -13862 19269 -13828
rect 19645 -13862 19657 -13828
rect 19257 -13868 19657 -13862
rect 19893 -13828 20293 -13822
rect 19893 -13862 19905 -13828
rect 20281 -13862 20293 -13828
rect 19893 -13868 20293 -13862
rect 20857 -13828 21257 -13822
rect 20857 -13862 20869 -13828
rect 21245 -13862 21257 -13828
rect 20857 -13868 21257 -13862
rect 21493 -13828 21893 -13822
rect 21493 -13862 21505 -13828
rect 21881 -13862 21893 -13828
rect 21493 -13868 21893 -13862
rect 22457 -13828 22857 -13822
rect 22457 -13862 22469 -13828
rect 22845 -13862 22857 -13828
rect 22457 -13868 22857 -13862
rect 23093 -13828 23493 -13822
rect 23093 -13862 23105 -13828
rect 23481 -13862 23493 -13828
rect 23093 -13868 23493 -13862
rect 24057 -13828 24457 -13822
rect 24057 -13862 24069 -13828
rect 24445 -13862 24457 -13828
rect 24057 -13868 24457 -13862
rect 24693 -13828 25093 -13822
rect 24693 -13862 24705 -13828
rect 25081 -13862 25093 -13828
rect 24693 -13868 25093 -13862
rect 25657 -13828 26057 -13822
rect 25657 -13862 25669 -13828
rect 26045 -13862 26057 -13828
rect 25657 -13868 26057 -13862
rect 26293 -13828 26693 -13822
rect 26293 -13862 26305 -13828
rect 26681 -13862 26693 -13828
rect 26293 -13868 26693 -13862
rect 27257 -13828 27657 -13822
rect 27257 -13862 27269 -13828
rect 27645 -13862 27657 -13828
rect 27257 -13868 27657 -13862
rect 27893 -13828 28293 -13822
rect 27893 -13862 27905 -13828
rect 28281 -13862 28293 -13828
rect 27893 -13868 28293 -13862
rect 28857 -13828 29257 -13822
rect 28857 -13862 28869 -13828
rect 29245 -13862 29257 -13828
rect 28857 -13868 29257 -13862
rect 29493 -13828 29893 -13822
rect 29493 -13862 29505 -13828
rect 29881 -13862 29893 -13828
rect 29493 -13868 29893 -13862
rect 30457 -13828 30857 -13822
rect 30457 -13862 30469 -13828
rect 30845 -13862 30857 -13828
rect 30457 -13868 30857 -13862
rect 31093 -13828 31493 -13822
rect 31093 -13862 31105 -13828
rect 31481 -13862 31493 -13828
rect 31093 -13868 31493 -13862
rect 32057 -13828 32457 -13822
rect 32057 -13862 32069 -13828
rect 32445 -13862 32457 -13828
rect 32057 -13868 32457 -13862
rect 32693 -13828 33093 -13822
rect 32693 -13862 32705 -13828
rect 33081 -13862 33093 -13828
rect 32693 -13868 33093 -13862
rect 33657 -13828 34057 -13822
rect 33657 -13862 33669 -13828
rect 34045 -13862 34057 -13828
rect 33657 -13868 34057 -13862
rect 34293 -13828 34693 -13822
rect 34293 -13862 34305 -13828
rect 34681 -13862 34693 -13828
rect 34293 -13868 34693 -13862
rect 35257 -13828 35657 -13822
rect 35257 -13862 35269 -13828
rect 35645 -13862 35657 -13828
rect 35257 -13868 35657 -13862
rect 35893 -13828 36293 -13822
rect 35893 -13862 35905 -13828
rect 36281 -13862 36293 -13828
rect 35893 -13868 36293 -13862
rect 36857 -13828 37257 -13822
rect 36857 -13862 36869 -13828
rect 37245 -13862 37257 -13828
rect 36857 -13868 37257 -13862
rect 37493 -13828 37893 -13822
rect 37493 -13862 37505 -13828
rect 37881 -13862 37893 -13828
rect 37493 -13868 37893 -13862
rect 15090 -13920 15490 -13868
rect 12860 -14040 15490 -13920
rect 11260 -14060 12290 -14050
rect 11260 -14090 11270 -14060
rect 10290 -14096 10693 -14090
rect 10290 -14130 10305 -14096
rect 10681 -14130 10693 -14096
rect 9657 -14136 10057 -14130
rect 10293 -14136 10693 -14130
rect 11257 -14096 11270 -14090
rect 11650 -14090 12290 -14060
rect 12860 -14090 13260 -14040
rect 11650 -14096 12293 -14090
rect 11257 -14130 11269 -14096
rect 11650 -14120 11905 -14096
rect 11645 -14130 11660 -14120
rect 11893 -14130 11905 -14120
rect 12281 -14130 12293 -14096
rect 11257 -14136 11657 -14130
rect 11893 -14136 12293 -14130
rect 12857 -14096 13260 -14090
rect 12857 -14130 12869 -14096
rect 13245 -14130 13260 -14096
rect 13490 -14090 13890 -14040
rect 14460 -14090 14860 -14040
rect 13490 -14096 13893 -14090
rect 13490 -14130 13505 -14096
rect 13881 -14130 13893 -14096
rect 12857 -14136 13257 -14130
rect 13493 -14136 13893 -14130
rect 14457 -14096 14860 -14090
rect 14457 -14130 14469 -14096
rect 14845 -14130 14860 -14096
rect 15090 -14090 15490 -14040
rect 15600 -13920 15740 -13910
rect 15600 -14040 15610 -13920
rect 15730 -13930 15740 -13920
rect 16060 -13930 16450 -13868
rect 16700 -13930 17090 -13868
rect 15730 -14030 17090 -13930
rect 15730 -14040 15740 -14030
rect 15600 -14050 15740 -14040
rect 16060 -14090 16450 -14030
rect 16700 -14090 17090 -14030
rect 17200 -13920 17340 -13910
rect 17200 -14040 17210 -13920
rect 17330 -13930 17340 -13920
rect 17660 -13930 18050 -13868
rect 18300 -13930 18690 -13868
rect 17330 -14030 18690 -13930
rect 17330 -14040 17340 -14030
rect 17200 -14050 17340 -14040
rect 17660 -14090 18050 -14030
rect 18300 -14090 18690 -14030
rect 18800 -13920 18940 -13910
rect 18800 -14040 18810 -13920
rect 18930 -13930 18940 -13920
rect 19260 -13930 19650 -13868
rect 19900 -13930 20290 -13868
rect 18930 -14030 20290 -13930
rect 18930 -14040 18940 -14030
rect 18800 -14050 18940 -14040
rect 19260 -14090 19650 -14030
rect 19900 -14090 20290 -14030
rect 20400 -13920 20540 -13910
rect 20400 -14040 20410 -13920
rect 20530 -13930 20540 -13920
rect 20860 -13930 21250 -13868
rect 21500 -13930 21890 -13868
rect 20530 -14030 21890 -13930
rect 20530 -14040 20540 -14030
rect 20400 -14050 20540 -14040
rect 20860 -14090 21250 -14030
rect 21500 -14090 21890 -14030
rect 22000 -13920 22140 -13910
rect 22000 -14040 22010 -13920
rect 22130 -13930 22140 -13920
rect 22460 -13930 22850 -13868
rect 23100 -13930 23490 -13868
rect 22130 -14030 23490 -13930
rect 22130 -14040 22140 -14030
rect 22000 -14050 22140 -14040
rect 22460 -14090 22850 -14030
rect 23100 -14090 23490 -14030
rect 23600 -13920 23740 -13910
rect 23600 -14040 23610 -13920
rect 23730 -13930 23740 -13920
rect 24060 -13930 24450 -13868
rect 24700 -13930 25090 -13868
rect 23730 -14030 25090 -13930
rect 23730 -14040 23740 -14030
rect 23600 -14050 23740 -14040
rect 24060 -14090 24450 -14030
rect 24700 -14090 25090 -14030
rect 25200 -13920 25340 -13910
rect 25200 -14040 25210 -13920
rect 25330 -13930 25340 -13920
rect 25660 -13930 26050 -13868
rect 26300 -13930 26690 -13868
rect 25330 -14030 26690 -13930
rect 25330 -14040 25340 -14030
rect 25200 -14050 25340 -14040
rect 25660 -14090 26050 -14030
rect 26300 -14090 26690 -14030
rect 26800 -13920 26940 -13910
rect 26800 -14040 26810 -13920
rect 26930 -13930 26940 -13920
rect 27260 -13930 27650 -13868
rect 27900 -13930 28290 -13868
rect 26930 -14030 28290 -13930
rect 26930 -14040 26940 -14030
rect 26800 -14050 26940 -14040
rect 27260 -14090 27650 -14030
rect 27900 -14090 28290 -14030
rect 28400 -13920 28540 -13910
rect 28400 -14040 28410 -13920
rect 28530 -13930 28540 -13920
rect 28860 -13930 29250 -13868
rect 29500 -13930 29890 -13868
rect 28530 -14030 29890 -13930
rect 28530 -14040 28540 -14030
rect 28400 -14050 28540 -14040
rect 28860 -14090 29250 -14030
rect 29500 -14090 29890 -14030
rect 30000 -13920 30140 -13910
rect 30000 -14040 30010 -13920
rect 30130 -13930 30140 -13920
rect 30460 -13930 30850 -13868
rect 31100 -13930 31490 -13868
rect 30130 -14030 31490 -13930
rect 30130 -14040 30140 -14030
rect 30000 -14050 30140 -14040
rect 30460 -14090 30850 -14030
rect 31100 -14090 31490 -14030
rect 31600 -13920 31740 -13910
rect 31600 -14040 31610 -13920
rect 31730 -13930 31740 -13920
rect 32060 -13930 32450 -13868
rect 32700 -13930 33090 -13868
rect 33660 -13930 34050 -13868
rect 34300 -13930 34690 -13868
rect 35260 -13930 35650 -13868
rect 35900 -13930 36290 -13868
rect 31730 -14030 36290 -13930
rect 31730 -14040 31740 -14030
rect 31600 -14050 31740 -14040
rect 32060 -14090 32450 -14030
rect 32700 -14090 33090 -14030
rect 33660 -14090 34050 -14030
rect 34300 -14090 34690 -14030
rect 35260 -14090 35650 -14030
rect 35900 -14090 36290 -14030
rect 15090 -14096 15493 -14090
rect 15090 -14130 15105 -14096
rect 15481 -14130 15493 -14096
rect 14457 -14136 14857 -14130
rect 15093 -14136 15493 -14130
rect 16057 -14096 16457 -14090
rect 16057 -14130 16069 -14096
rect 16445 -14130 16457 -14096
rect 16057 -14136 16457 -14130
rect 16693 -14096 17093 -14090
rect 16693 -14130 16705 -14096
rect 17081 -14130 17093 -14096
rect 16693 -14136 17093 -14130
rect 17657 -14096 18057 -14090
rect 17657 -14130 17669 -14096
rect 18045 -14130 18057 -14096
rect 17657 -14136 18057 -14130
rect 18293 -14096 18693 -14090
rect 18293 -14130 18305 -14096
rect 18681 -14130 18693 -14096
rect 18293 -14136 18693 -14130
rect 19257 -14096 19657 -14090
rect 19257 -14130 19269 -14096
rect 19645 -14130 19657 -14096
rect 19257 -14136 19657 -14130
rect 19893 -14096 20293 -14090
rect 19893 -14130 19905 -14096
rect 20281 -14130 20293 -14096
rect 19893 -14136 20293 -14130
rect 20857 -14096 21257 -14090
rect 20857 -14130 20869 -14096
rect 21245 -14130 21257 -14096
rect 20857 -14136 21257 -14130
rect 21493 -14096 21893 -14090
rect 21493 -14130 21505 -14096
rect 21881 -14130 21893 -14096
rect 21493 -14136 21893 -14130
rect 22457 -14096 22857 -14090
rect 22457 -14130 22469 -14096
rect 22845 -14130 22857 -14096
rect 22457 -14136 22857 -14130
rect 23093 -14096 23493 -14090
rect 23093 -14130 23105 -14096
rect 23481 -14130 23493 -14096
rect 23093 -14136 23493 -14130
rect 24057 -14096 24457 -14090
rect 24057 -14130 24069 -14096
rect 24445 -14130 24457 -14096
rect 24057 -14136 24457 -14130
rect 24693 -14096 25093 -14090
rect 24693 -14130 24705 -14096
rect 25081 -14130 25093 -14096
rect 24693 -14136 25093 -14130
rect 25657 -14096 26057 -14090
rect 25657 -14130 25669 -14096
rect 26045 -14130 26057 -14096
rect 25657 -14136 26057 -14130
rect 26293 -14096 26693 -14090
rect 26293 -14130 26305 -14096
rect 26681 -14130 26693 -14096
rect 26293 -14136 26693 -14130
rect 27257 -14096 27657 -14090
rect 27257 -14130 27269 -14096
rect 27645 -14130 27657 -14096
rect 27257 -14136 27657 -14130
rect 27893 -14096 28293 -14090
rect 27893 -14130 27905 -14096
rect 28281 -14130 28293 -14096
rect 27893 -14136 28293 -14130
rect 28857 -14096 29257 -14090
rect 28857 -14130 28869 -14096
rect 29245 -14130 29257 -14096
rect 28857 -14136 29257 -14130
rect 29493 -14096 29893 -14090
rect 29493 -14130 29505 -14096
rect 29881 -14130 29893 -14096
rect 29493 -14136 29893 -14130
rect 30457 -14096 30857 -14090
rect 30457 -14130 30469 -14096
rect 30845 -14130 30857 -14096
rect 30457 -14136 30857 -14130
rect 31093 -14096 31493 -14090
rect 31093 -14130 31105 -14096
rect 31481 -14130 31493 -14096
rect 31093 -14136 31493 -14130
rect 32057 -14096 32457 -14090
rect 32057 -14130 32069 -14096
rect 32445 -14130 32457 -14096
rect 32057 -14136 32457 -14130
rect 32693 -14096 33093 -14090
rect 32693 -14130 32705 -14096
rect 33081 -14130 33093 -14096
rect 32693 -14136 33093 -14130
rect 33657 -14096 34057 -14090
rect 33657 -14130 33669 -14096
rect 34045 -14130 34057 -14096
rect 33657 -14136 34057 -14130
rect 34293 -14096 34693 -14090
rect 34293 -14130 34305 -14096
rect 34681 -14130 34693 -14096
rect 34293 -14136 34693 -14130
rect 35257 -14096 35657 -14090
rect 35257 -14130 35269 -14096
rect 35645 -14130 35657 -14096
rect 35257 -14136 35657 -14130
rect 35893 -14096 36293 -14090
rect 35893 -14130 35905 -14096
rect 36281 -14130 36293 -14096
rect 35893 -14136 36293 -14130
rect 36857 -14096 37257 -14090
rect 36857 -14130 36869 -14096
rect 37245 -14130 37257 -14096
rect 36857 -14136 37257 -14130
rect 37493 -14096 37893 -14090
rect 37493 -14130 37505 -14096
rect 37881 -14130 37893 -14096
rect 37493 -14136 37893 -14130
rect 57 -14954 490 -14948
rect 57 -14980 69 -14954
rect 0 -14988 69 -14980
rect 445 -14988 490 -14954
rect 0 -15088 490 -14988
rect 670 -14948 720 -14136
rect 1134 -14196 1180 -14184
rect 1134 -14888 1140 -14196
rect 1174 -14888 1180 -14196
rect 1134 -14900 1180 -14888
rect 1570 -14196 1616 -14184
rect 1570 -14888 1576 -14196
rect 1610 -14888 1616 -14196
rect 1570 -14900 1616 -14888
rect 2098 -14196 2144 -14184
rect 2098 -14888 2104 -14196
rect 2138 -14200 2144 -14196
rect 2206 -14196 2252 -14184
rect 2206 -14200 2212 -14196
rect 2138 -14210 2212 -14200
rect 2138 -14880 2212 -14870
rect 2138 -14888 2144 -14880
rect 2098 -14900 2144 -14888
rect 2206 -14888 2212 -14880
rect 2246 -14888 2252 -14196
rect 2206 -14900 2252 -14888
rect 2734 -14196 2780 -14184
rect 2734 -14888 2740 -14196
rect 2774 -14888 2780 -14196
rect 2734 -14900 2780 -14888
rect 3170 -14196 3216 -14184
rect 3170 -14888 3176 -14196
rect 3210 -14888 3216 -14196
rect 3170 -14900 3216 -14888
rect 3698 -14196 3744 -14184
rect 3698 -14888 3704 -14196
rect 3738 -14200 3744 -14196
rect 3806 -14196 3852 -14184
rect 3806 -14200 3812 -14196
rect 3738 -14210 3812 -14200
rect 3738 -14880 3812 -14870
rect 3738 -14888 3744 -14880
rect 3698 -14900 3744 -14888
rect 3806 -14888 3812 -14880
rect 3846 -14888 3852 -14196
rect 3806 -14900 3852 -14888
rect 4334 -14196 4380 -14184
rect 4334 -14888 4340 -14196
rect 4374 -14888 4380 -14196
rect 4334 -14900 4380 -14888
rect 4770 -14196 4816 -14184
rect 4770 -14888 4776 -14196
rect 4810 -14888 4816 -14196
rect 4770 -14900 4816 -14888
rect 5298 -14196 5344 -14184
rect 5298 -14888 5304 -14196
rect 5338 -14200 5344 -14196
rect 5406 -14196 5452 -14184
rect 5406 -14200 5412 -14196
rect 5338 -14210 5412 -14200
rect 5338 -14880 5412 -14870
rect 5338 -14888 5344 -14880
rect 5298 -14900 5344 -14888
rect 5406 -14888 5412 -14880
rect 5446 -14888 5452 -14196
rect 5406 -14900 5452 -14888
rect 5934 -14196 5980 -14184
rect 5934 -14888 5940 -14196
rect 5974 -14888 5980 -14196
rect 5934 -14900 5980 -14888
rect 6370 -14196 6416 -14184
rect 6370 -14888 6376 -14196
rect 6410 -14888 6416 -14196
rect 6370 -14900 6416 -14888
rect 6898 -14196 6944 -14184
rect 6898 -14888 6904 -14196
rect 6938 -14200 6944 -14196
rect 7006 -14196 7052 -14184
rect 7006 -14200 7012 -14196
rect 6938 -14210 7012 -14200
rect 6938 -14880 7012 -14870
rect 6938 -14888 6944 -14880
rect 6898 -14900 6944 -14888
rect 7006 -14888 7012 -14880
rect 7046 -14888 7052 -14196
rect 7006 -14900 7052 -14888
rect 7534 -14196 7580 -14184
rect 7534 -14888 7540 -14196
rect 7574 -14888 7580 -14196
rect 7534 -14900 7580 -14888
rect 7970 -14196 8016 -14184
rect 7970 -14888 7976 -14196
rect 8010 -14888 8016 -14196
rect 7970 -14900 8016 -14888
rect 8498 -14196 8544 -14184
rect 8498 -14888 8504 -14196
rect 8538 -14200 8544 -14196
rect 8606 -14196 8652 -14184
rect 8606 -14200 8612 -14196
rect 8538 -14210 8612 -14200
rect 8538 -14880 8612 -14870
rect 8538 -14888 8544 -14880
rect 8498 -14900 8544 -14888
rect 8606 -14888 8612 -14880
rect 8646 -14888 8652 -14196
rect 8606 -14900 8652 -14888
rect 9134 -14196 9180 -14184
rect 9134 -14888 9140 -14196
rect 9174 -14888 9180 -14196
rect 9134 -14900 9180 -14888
rect 9570 -14196 9616 -14184
rect 9570 -14888 9576 -14196
rect 9610 -14888 9616 -14196
rect 9570 -14900 9616 -14888
rect 10098 -14196 10144 -14184
rect 10098 -14888 10104 -14196
rect 10138 -14200 10144 -14196
rect 10206 -14196 10252 -14184
rect 10206 -14200 10212 -14196
rect 10138 -14210 10212 -14200
rect 10138 -14880 10212 -14870
rect 10138 -14888 10144 -14880
rect 10098 -14900 10144 -14888
rect 10206 -14888 10212 -14880
rect 10246 -14888 10252 -14196
rect 10206 -14900 10252 -14888
rect 10734 -14196 10780 -14184
rect 10734 -14888 10740 -14196
rect 10774 -14888 10780 -14196
rect 10734 -14900 10780 -14888
rect 11170 -14196 11216 -14184
rect 11170 -14888 11176 -14196
rect 11210 -14888 11216 -14196
rect 11170 -14900 11216 -14888
rect 11698 -14196 11744 -14184
rect 11698 -14888 11704 -14196
rect 11738 -14200 11744 -14196
rect 11806 -14196 11852 -14184
rect 11806 -14200 11812 -14196
rect 11738 -14210 11812 -14200
rect 11738 -14880 11812 -14870
rect 11738 -14888 11744 -14880
rect 11698 -14900 11744 -14888
rect 11806 -14888 11812 -14880
rect 11846 -14888 11852 -14196
rect 11806 -14900 11852 -14888
rect 12334 -14196 12380 -14184
rect 12334 -14888 12340 -14196
rect 12374 -14888 12380 -14196
rect 12334 -14900 12380 -14888
rect 12770 -14196 12816 -14184
rect 12770 -14888 12776 -14196
rect 12810 -14888 12816 -14196
rect 12770 -14900 12816 -14888
rect 13298 -14196 13344 -14184
rect 13298 -14888 13304 -14196
rect 13338 -14200 13344 -14196
rect 13406 -14196 13452 -14184
rect 13406 -14200 13412 -14196
rect 13338 -14210 13412 -14200
rect 13338 -14880 13412 -14870
rect 13338 -14888 13344 -14880
rect 13298 -14900 13344 -14888
rect 13406 -14888 13412 -14880
rect 13446 -14888 13452 -14196
rect 13406 -14900 13452 -14888
rect 13934 -14196 13980 -14184
rect 13934 -14888 13940 -14196
rect 13974 -14888 13980 -14196
rect 13934 -14900 13980 -14888
rect 14370 -14196 14416 -14184
rect 14370 -14888 14376 -14196
rect 14410 -14888 14416 -14196
rect 14370 -14900 14416 -14888
rect 14898 -14196 14944 -14184
rect 14898 -14888 14904 -14196
rect 14938 -14200 14944 -14196
rect 15006 -14196 15052 -14184
rect 15006 -14200 15012 -14196
rect 14938 -14210 15012 -14200
rect 14938 -14880 15012 -14870
rect 14938 -14888 14944 -14880
rect 14898 -14900 14944 -14888
rect 15006 -14888 15012 -14880
rect 15046 -14888 15052 -14196
rect 15006 -14900 15052 -14888
rect 15534 -14196 15580 -14184
rect 15534 -14888 15540 -14196
rect 15574 -14888 15580 -14196
rect 15534 -14900 15580 -14888
rect 15970 -14196 16016 -14184
rect 15970 -14888 15976 -14196
rect 16010 -14888 16016 -14196
rect 15970 -14900 16016 -14888
rect 16498 -14190 16544 -14184
rect 16606 -14190 16652 -14184
rect 16498 -14196 16652 -14190
rect 16498 -14888 16504 -14196
rect 16538 -14200 16612 -14196
rect 16538 -14888 16612 -14880
rect 16646 -14888 16652 -14196
rect 16498 -14890 16652 -14888
rect 16498 -14900 16544 -14890
rect 16606 -14900 16652 -14890
rect 17134 -14196 17180 -14184
rect 17134 -14888 17140 -14196
rect 17174 -14888 17180 -14196
rect 17134 -14900 17180 -14888
rect 17570 -14196 17616 -14184
rect 17570 -14888 17576 -14196
rect 17610 -14888 17616 -14196
rect 17570 -14900 17616 -14888
rect 18098 -14190 18144 -14184
rect 18206 -14190 18252 -14184
rect 18098 -14196 18252 -14190
rect 18098 -14888 18104 -14196
rect 18138 -14200 18212 -14196
rect 18138 -14888 18212 -14880
rect 18246 -14888 18252 -14196
rect 18098 -14890 18252 -14888
rect 18098 -14900 18144 -14890
rect 18206 -14900 18252 -14890
rect 18734 -14196 18780 -14184
rect 18734 -14888 18740 -14196
rect 18774 -14888 18780 -14196
rect 18734 -14900 18780 -14888
rect 19170 -14196 19216 -14184
rect 19170 -14888 19176 -14196
rect 19210 -14888 19216 -14196
rect 19170 -14900 19216 -14888
rect 19698 -14190 19744 -14184
rect 19806 -14190 19852 -14184
rect 19698 -14196 19852 -14190
rect 19698 -14888 19704 -14196
rect 19738 -14200 19812 -14196
rect 19738 -14888 19812 -14880
rect 19846 -14888 19852 -14196
rect 19698 -14890 19852 -14888
rect 19698 -14900 19744 -14890
rect 19806 -14900 19852 -14890
rect 20334 -14196 20380 -14184
rect 20334 -14888 20340 -14196
rect 20374 -14888 20380 -14196
rect 20334 -14900 20380 -14888
rect 20770 -14196 20816 -14184
rect 20770 -14888 20776 -14196
rect 20810 -14888 20816 -14196
rect 20770 -14900 20816 -14888
rect 21298 -14190 21344 -14184
rect 21406 -14190 21452 -14184
rect 21298 -14196 21452 -14190
rect 21298 -14888 21304 -14196
rect 21338 -14200 21412 -14196
rect 21338 -14888 21412 -14880
rect 21446 -14888 21452 -14196
rect 21298 -14890 21452 -14888
rect 21298 -14900 21344 -14890
rect 21406 -14900 21452 -14890
rect 21934 -14196 21980 -14184
rect 21934 -14888 21940 -14196
rect 21974 -14888 21980 -14196
rect 21934 -14900 21980 -14888
rect 22370 -14196 22416 -14184
rect 22370 -14888 22376 -14196
rect 22410 -14888 22416 -14196
rect 22370 -14900 22416 -14888
rect 22898 -14190 22944 -14184
rect 23006 -14190 23052 -14184
rect 22898 -14196 23052 -14190
rect 22898 -14888 22904 -14196
rect 22938 -14200 23012 -14196
rect 22938 -14888 23012 -14880
rect 23046 -14888 23052 -14196
rect 22898 -14890 23052 -14888
rect 22898 -14900 22944 -14890
rect 23006 -14900 23052 -14890
rect 23534 -14196 23580 -14184
rect 23534 -14888 23540 -14196
rect 23574 -14888 23580 -14196
rect 23534 -14900 23580 -14888
rect 23970 -14196 24016 -14184
rect 23970 -14888 23976 -14196
rect 24010 -14888 24016 -14196
rect 23970 -14900 24016 -14888
rect 24498 -14190 24544 -14184
rect 24606 -14190 24652 -14184
rect 24498 -14196 24652 -14190
rect 24498 -14888 24504 -14196
rect 24538 -14200 24612 -14196
rect 24538 -14888 24612 -14880
rect 24646 -14888 24652 -14196
rect 24498 -14890 24652 -14888
rect 24498 -14900 24544 -14890
rect 24606 -14900 24652 -14890
rect 25134 -14196 25180 -14184
rect 25134 -14888 25140 -14196
rect 25174 -14888 25180 -14196
rect 25134 -14900 25180 -14888
rect 25570 -14196 25616 -14184
rect 25570 -14888 25576 -14196
rect 25610 -14888 25616 -14196
rect 25570 -14900 25616 -14888
rect 26098 -14190 26144 -14184
rect 26206 -14190 26252 -14184
rect 26098 -14196 26252 -14190
rect 26098 -14888 26104 -14196
rect 26138 -14200 26212 -14196
rect 26138 -14888 26212 -14880
rect 26246 -14888 26252 -14196
rect 26098 -14890 26252 -14888
rect 26098 -14900 26144 -14890
rect 26206 -14900 26252 -14890
rect 26734 -14196 26780 -14184
rect 26734 -14888 26740 -14196
rect 26774 -14888 26780 -14196
rect 26734 -14900 26780 -14888
rect 27170 -14196 27216 -14184
rect 27170 -14888 27176 -14196
rect 27210 -14888 27216 -14196
rect 27170 -14900 27216 -14888
rect 27698 -14190 27744 -14184
rect 27806 -14190 27852 -14184
rect 27698 -14196 27852 -14190
rect 27698 -14888 27704 -14196
rect 27738 -14200 27812 -14196
rect 27738 -14888 27812 -14880
rect 27846 -14888 27852 -14196
rect 27698 -14890 27852 -14888
rect 27698 -14900 27744 -14890
rect 27806 -14900 27852 -14890
rect 28334 -14196 28380 -14184
rect 28334 -14888 28340 -14196
rect 28374 -14888 28380 -14196
rect 28334 -14900 28380 -14888
rect 28770 -14196 28816 -14184
rect 28770 -14888 28776 -14196
rect 28810 -14888 28816 -14196
rect 28770 -14900 28816 -14888
rect 29298 -14190 29344 -14184
rect 29406 -14190 29452 -14184
rect 29298 -14196 29452 -14190
rect 29298 -14888 29304 -14196
rect 29338 -14200 29412 -14196
rect 29338 -14888 29412 -14880
rect 29446 -14888 29452 -14196
rect 29298 -14890 29452 -14888
rect 29298 -14900 29344 -14890
rect 29406 -14900 29452 -14890
rect 29934 -14196 29980 -14184
rect 29934 -14888 29940 -14196
rect 29974 -14888 29980 -14196
rect 29934 -14900 29980 -14888
rect 30370 -14196 30416 -14184
rect 30370 -14888 30376 -14196
rect 30410 -14888 30416 -14196
rect 30370 -14900 30416 -14888
rect 30898 -14190 30944 -14184
rect 31006 -14190 31052 -14184
rect 30898 -14196 31052 -14190
rect 30898 -14888 30904 -14196
rect 30938 -14200 31012 -14196
rect 30938 -14888 31012 -14880
rect 31046 -14888 31052 -14196
rect 30898 -14890 31052 -14888
rect 30898 -14900 30944 -14890
rect 31006 -14900 31052 -14890
rect 31534 -14196 31580 -14184
rect 31534 -14888 31540 -14196
rect 31574 -14888 31580 -14196
rect 31534 -14900 31580 -14888
rect 31970 -14196 32016 -14184
rect 31970 -14888 31976 -14196
rect 32010 -14888 32016 -14196
rect 31970 -14900 32016 -14888
rect 32498 -14190 32544 -14184
rect 32606 -14190 32652 -14184
rect 32498 -14196 32652 -14190
rect 32498 -14888 32504 -14196
rect 32538 -14200 32612 -14196
rect 32538 -14888 32544 -14710
rect 32498 -14900 32544 -14888
rect 32606 -14888 32612 -14710
rect 32646 -14888 32652 -14196
rect 32606 -14900 32652 -14888
rect 33134 -14196 33180 -14184
rect 33134 -14888 33140 -14196
rect 33174 -14888 33180 -14196
rect 33134 -14900 33180 -14888
rect 33570 -14196 33616 -14184
rect 33570 -14888 33576 -14196
rect 33610 -14888 33616 -14196
rect 33570 -14900 33616 -14888
rect 34098 -14190 34144 -14184
rect 34206 -14190 34252 -14184
rect 34098 -14196 34252 -14190
rect 34098 -14888 34104 -14196
rect 34138 -14200 34212 -14196
rect 34138 -14888 34144 -14710
rect 34098 -14900 34144 -14888
rect 34206 -14888 34212 -14710
rect 34246 -14888 34252 -14196
rect 34206 -14900 34252 -14888
rect 34734 -14196 34780 -14184
rect 34734 -14888 34740 -14196
rect 34774 -14888 34780 -14196
rect 34734 -14900 34780 -14888
rect 35170 -14196 35216 -14184
rect 35170 -14888 35176 -14196
rect 35210 -14888 35216 -14196
rect 35170 -14900 35216 -14888
rect 35698 -14190 35744 -14184
rect 35806 -14190 35852 -14184
rect 35698 -14196 35852 -14190
rect 35698 -14888 35704 -14196
rect 35738 -14200 35812 -14196
rect 35738 -14888 35744 -14710
rect 35698 -14900 35744 -14888
rect 35806 -14888 35812 -14710
rect 35846 -14888 35852 -14196
rect 35806 -14900 35852 -14888
rect 36334 -14196 36380 -14184
rect 36334 -14888 36340 -14196
rect 36374 -14888 36380 -14196
rect 36334 -14900 36380 -14888
rect 36770 -14196 36816 -14184
rect 36770 -14888 36776 -14196
rect 36810 -14888 36816 -14196
rect 36770 -14900 36816 -14888
rect 37298 -14196 37344 -14184
rect 37298 -14888 37304 -14196
rect 37338 -14888 37344 -14196
rect 37298 -14900 37344 -14888
rect 37406 -14196 37452 -14184
rect 37406 -14888 37412 -14196
rect 37446 -14888 37452 -14196
rect 37406 -14900 37452 -14888
rect 37934 -14196 37980 -14184
rect 37934 -14888 37940 -14196
rect 37974 -14888 37980 -14196
rect 37934 -14900 37980 -14888
rect 35000 -14910 35140 -14900
rect 670 -14954 1093 -14948
rect 670 -14988 705 -14954
rect 1081 -14980 1093 -14954
rect 1657 -14954 2057 -14948
rect 1657 -14980 1669 -14954
rect 1081 -14988 1669 -14980
rect 2045 -14980 2057 -14954
rect 2293 -14954 2693 -14948
rect 2293 -14980 2305 -14954
rect 2045 -14988 2305 -14980
rect 2681 -14980 2693 -14954
rect 3257 -14954 3657 -14948
rect 3257 -14980 3269 -14954
rect 2681 -14988 3269 -14980
rect 3645 -14980 3657 -14954
rect 3893 -14954 4293 -14948
rect 3893 -14980 3905 -14954
rect 3645 -14988 3905 -14980
rect 4281 -14980 4293 -14954
rect 4857 -14954 5257 -14948
rect 4857 -14980 4869 -14954
rect 4281 -14988 4869 -14980
rect 5245 -14980 5257 -14954
rect 5493 -14954 5893 -14948
rect 5493 -14980 5505 -14954
rect 5245 -14988 5505 -14980
rect 5881 -14980 5893 -14954
rect 6457 -14954 6857 -14948
rect 6457 -14980 6469 -14954
rect 5881 -14988 6469 -14980
rect 6845 -14980 6857 -14954
rect 7093 -14954 7493 -14948
rect 7093 -14980 7105 -14954
rect 6845 -14988 7105 -14980
rect 7481 -14980 7493 -14954
rect 8057 -14954 8457 -14948
rect 8057 -14980 8069 -14954
rect 7481 -14988 8069 -14980
rect 8445 -14980 8457 -14954
rect 8693 -14954 9093 -14948
rect 8693 -14980 8705 -14954
rect 8445 -14988 8705 -14980
rect 9081 -14980 9093 -14954
rect 9657 -14954 10057 -14948
rect 9657 -14980 9669 -14954
rect 9081 -14988 9669 -14980
rect 10045 -14980 10057 -14954
rect 10293 -14954 10693 -14948
rect 10293 -14980 10305 -14954
rect 10045 -14988 10305 -14980
rect 10681 -14980 10693 -14954
rect 11257 -14954 11657 -14948
rect 11257 -14980 11269 -14954
rect 10681 -14988 11269 -14980
rect 11645 -14980 11657 -14954
rect 11893 -14954 12293 -14948
rect 11893 -14980 11905 -14954
rect 11645 -14988 11905 -14980
rect 12281 -14980 12293 -14954
rect 12857 -14954 13257 -14948
rect 12857 -14980 12869 -14954
rect 12281 -14988 12869 -14980
rect 13245 -14980 13257 -14954
rect 13493 -14954 13893 -14948
rect 13493 -14980 13505 -14954
rect 13245 -14988 13505 -14980
rect 13881 -14980 13893 -14954
rect 14457 -14954 14857 -14948
rect 14457 -14980 14469 -14954
rect 13881 -14988 14469 -14980
rect 14845 -14980 14857 -14954
rect 15093 -14954 15493 -14948
rect 15093 -14980 15105 -14954
rect 14845 -14988 15105 -14980
rect 15481 -14980 15493 -14954
rect 16057 -14954 16457 -14948
rect 16057 -14980 16069 -14954
rect 15481 -14988 16069 -14980
rect 16445 -14980 16457 -14954
rect 16693 -14954 17093 -14948
rect 16693 -14980 16705 -14954
rect 16445 -14988 16705 -14980
rect 17081 -14980 17093 -14954
rect 17657 -14954 18057 -14948
rect 17657 -14980 17669 -14954
rect 17081 -14988 17669 -14980
rect 18045 -14980 18057 -14954
rect 18293 -14954 18693 -14948
rect 18293 -14980 18305 -14954
rect 18045 -14988 18305 -14980
rect 18681 -14980 18693 -14954
rect 19257 -14954 19657 -14948
rect 19257 -14980 19269 -14954
rect 18681 -14988 19269 -14980
rect 19645 -14980 19657 -14954
rect 19893 -14954 20293 -14948
rect 19893 -14980 19905 -14954
rect 19645 -14988 19905 -14980
rect 20281 -14980 20293 -14954
rect 20857 -14954 21257 -14948
rect 20857 -14980 20869 -14954
rect 20281 -14988 20869 -14980
rect 21245 -14980 21257 -14954
rect 21493 -14954 21893 -14948
rect 21493 -14980 21505 -14954
rect 21245 -14988 21505 -14980
rect 21881 -14980 21893 -14954
rect 22457 -14954 22857 -14948
rect 22457 -14980 22469 -14954
rect 21881 -14988 22469 -14980
rect 22845 -14980 22857 -14954
rect 23093 -14954 23493 -14948
rect 23093 -14980 23105 -14954
rect 22845 -14988 23105 -14980
rect 23481 -14980 23493 -14954
rect 24057 -14954 24457 -14948
rect 24057 -14980 24069 -14954
rect 23481 -14988 24069 -14980
rect 24445 -14980 24457 -14954
rect 24693 -14954 25093 -14948
rect 24693 -14980 24705 -14954
rect 24445 -14988 24705 -14980
rect 25081 -14980 25093 -14954
rect 25657 -14954 26057 -14948
rect 25657 -14980 25669 -14954
rect 25081 -14988 25669 -14980
rect 26045 -14980 26057 -14954
rect 26293 -14954 26693 -14948
rect 26293 -14980 26305 -14954
rect 26045 -14988 26305 -14980
rect 26681 -14980 26693 -14954
rect 27257 -14954 27657 -14948
rect 27257 -14980 27269 -14954
rect 26681 -14988 27269 -14980
rect 27645 -14980 27657 -14954
rect 27893 -14954 28293 -14948
rect 27893 -14980 27905 -14954
rect 27645 -14988 27905 -14980
rect 28281 -14980 28293 -14954
rect 28857 -14954 29257 -14948
rect 28857 -14980 28869 -14954
rect 28281 -14988 28869 -14980
rect 29245 -14980 29257 -14954
rect 29493 -14954 29893 -14948
rect 29493 -14980 29505 -14954
rect 29245 -14988 29505 -14980
rect 29881 -14980 29893 -14954
rect 30457 -14954 30857 -14948
rect 30457 -14980 30469 -14954
rect 29881 -14988 30469 -14980
rect 30845 -14980 30857 -14954
rect 31093 -14954 31493 -14948
rect 31093 -14980 31105 -14954
rect 30845 -14988 31105 -14980
rect 31481 -14980 31493 -14954
rect 32057 -14950 32457 -14948
rect 32693 -14950 33093 -14948
rect 33657 -14950 34057 -14948
rect 34293 -14950 34693 -14948
rect 35000 -14950 35010 -14910
rect 32057 -14954 35010 -14950
rect 31481 -14988 31800 -14980
rect 670 -15088 31800 -14988
rect 32057 -14988 32069 -14954
rect 32445 -14988 32705 -14954
rect 33081 -14988 33669 -14954
rect 34045 -14988 34305 -14954
rect 34681 -14988 35010 -14954
rect 32057 -14994 35010 -14988
rect 32060 -15030 35010 -14994
rect 35130 -14950 35140 -14910
rect 35257 -14950 35657 -14948
rect 35893 -14950 36293 -14948
rect 35130 -14954 36293 -14950
rect 35130 -14988 35269 -14954
rect 35645 -14988 35905 -14954
rect 36281 -14988 36293 -14954
rect 35130 -14994 36293 -14988
rect 36857 -14954 37257 -14948
rect 36857 -14988 36869 -14954
rect 37245 -14988 37257 -14954
rect 36857 -14994 37257 -14988
rect 37493 -14954 37893 -14948
rect 37493 -14988 37505 -14954
rect 37881 -14988 37893 -14954
rect 37493 -14994 37893 -14988
rect 35130 -15030 36290 -14994
rect 32060 -15040 36290 -15030
rect 0 -15122 13 -15088
rect 1137 -15122 1613 -15088
rect 2737 -15122 3213 -15088
rect 4337 -15122 4813 -15088
rect 5937 -15122 6413 -15088
rect 7537 -15122 8013 -15088
rect 9137 -15122 9613 -15088
rect 10737 -15122 11213 -15088
rect 12337 -15122 12813 -15088
rect 13937 -15122 14413 -15088
rect 15537 -15122 16013 -15088
rect 17137 -15122 17613 -15088
rect 18737 -15122 19213 -15088
rect 20337 -15122 20813 -15088
rect 21937 -15122 22413 -15088
rect 23537 -15122 24013 -15088
rect 25137 -15122 25613 -15088
rect 26737 -15122 27213 -15088
rect 28337 -15122 28813 -15088
rect 29937 -15122 30413 -15088
rect 31537 -15100 31800 -15088
rect 32001 -15088 33149 -15082
rect 32001 -15100 32013 -15088
rect 31537 -15122 32013 -15100
rect 33137 -15100 33149 -15088
rect 33601 -15088 34749 -15082
rect 33601 -15100 33613 -15088
rect 33137 -15122 33613 -15100
rect 34737 -15100 34749 -15088
rect 35201 -15088 36349 -15082
rect 35201 -15100 35213 -15088
rect 34737 -15122 35213 -15100
rect 36337 -15100 36349 -15088
rect 36801 -15088 37949 -15082
rect 36801 -15100 36813 -15088
rect 36337 -15122 36813 -15100
rect 37937 -15122 37949 -15088
rect 0 -15220 490 -15122
rect 440 -15364 490 -15220
rect 57 -15370 490 -15364
rect 57 -15404 69 -15370
rect 445 -15404 490 -15370
rect 57 -15410 490 -15404
rect -30 -15457 16 -15445
rect -30 -15575 -24 -15457
rect 10 -15575 16 -15457
rect -30 -15587 16 -15575
rect 440 -15622 490 -15410
rect 670 -15128 37949 -15122
rect 670 -15220 37940 -15128
rect 670 -15364 720 -15220
rect 1200 -15270 1340 -15260
rect 670 -15370 1093 -15364
rect 670 -15404 705 -15370
rect 1081 -15404 1093 -15370
rect 1200 -15390 1210 -15270
rect 1330 -15280 1340 -15270
rect 2800 -15270 2940 -15260
rect 2800 -15280 2810 -15270
rect 1330 -15370 2810 -15280
rect 1330 -15380 1669 -15370
rect 1330 -15390 1340 -15380
rect 1200 -15400 1340 -15390
rect 670 -15410 1093 -15404
rect 1657 -15404 1669 -15380
rect 2045 -15380 2305 -15370
rect 2045 -15404 2057 -15380
rect 1657 -15410 2057 -15404
rect 2293 -15404 2305 -15380
rect 2681 -15380 2810 -15370
rect 2681 -15404 2693 -15380
rect 2800 -15390 2810 -15380
rect 2930 -15280 2940 -15270
rect 4400 -15270 4540 -15260
rect 4400 -15280 4410 -15270
rect 2930 -15370 4410 -15280
rect 2930 -15380 3269 -15370
rect 2930 -15390 2940 -15380
rect 2800 -15400 2940 -15390
rect 2293 -15410 2693 -15404
rect 3257 -15404 3269 -15380
rect 3645 -15380 3905 -15370
rect 3645 -15404 3657 -15380
rect 3257 -15410 3657 -15404
rect 3893 -15404 3905 -15380
rect 4281 -15380 4410 -15370
rect 4281 -15404 4293 -15380
rect 4400 -15390 4410 -15380
rect 4530 -15280 4540 -15270
rect 6000 -15270 6140 -15260
rect 6000 -15280 6010 -15270
rect 4530 -15370 6010 -15280
rect 4530 -15380 4869 -15370
rect 4530 -15390 4540 -15380
rect 4400 -15400 4540 -15390
rect 3893 -15410 4293 -15404
rect 4857 -15404 4869 -15380
rect 5245 -15380 5505 -15370
rect 5245 -15404 5257 -15380
rect 4857 -15410 5257 -15404
rect 5493 -15404 5505 -15380
rect 5881 -15380 6010 -15370
rect 5881 -15404 5893 -15380
rect 6000 -15390 6010 -15380
rect 6130 -15280 6140 -15270
rect 7600 -15270 7740 -15260
rect 7600 -15280 7610 -15270
rect 6130 -15370 7610 -15280
rect 6130 -15380 6469 -15370
rect 6130 -15390 6140 -15380
rect 6000 -15400 6140 -15390
rect 5493 -15410 5893 -15404
rect 6457 -15404 6469 -15380
rect 6845 -15380 7105 -15370
rect 6845 -15404 6857 -15380
rect 6457 -15410 6857 -15404
rect 7093 -15404 7105 -15380
rect 7481 -15380 7610 -15370
rect 7481 -15404 7493 -15380
rect 7600 -15390 7610 -15380
rect 7730 -15280 7740 -15270
rect 9200 -15270 9340 -15260
rect 9200 -15280 9210 -15270
rect 7730 -15370 9210 -15280
rect 7730 -15380 8069 -15370
rect 7730 -15390 7740 -15380
rect 7600 -15400 7740 -15390
rect 7093 -15410 7493 -15404
rect 8057 -15404 8069 -15380
rect 8445 -15380 8705 -15370
rect 8445 -15404 8457 -15380
rect 8057 -15410 8457 -15404
rect 8693 -15404 8705 -15380
rect 9081 -15380 9210 -15370
rect 9081 -15404 9093 -15380
rect 9200 -15390 9210 -15380
rect 9330 -15280 9340 -15270
rect 15820 -15270 15960 -15260
rect 9330 -15370 10700 -15280
rect 13320 -15290 13440 -15280
rect 13320 -15320 13330 -15290
rect 12860 -15364 13330 -15320
rect 9330 -15380 9669 -15370
rect 9330 -15390 9340 -15380
rect 9200 -15400 9340 -15390
rect 8693 -15410 9093 -15404
rect 9657 -15404 9669 -15380
rect 10045 -15380 10305 -15370
rect 10045 -15404 10057 -15380
rect 9657 -15410 10057 -15404
rect 10293 -15404 10305 -15380
rect 10681 -15380 10700 -15370
rect 11257 -15370 11657 -15364
rect 10681 -15404 10693 -15380
rect 10293 -15410 10693 -15404
rect 11257 -15404 11269 -15370
rect 11645 -15404 11657 -15370
rect 11257 -15410 11657 -15404
rect 11893 -15370 12293 -15364
rect 11893 -15404 11905 -15370
rect 12281 -15404 12293 -15370
rect 11893 -15410 12293 -15404
rect 12857 -15370 13330 -15364
rect 12857 -15404 12869 -15370
rect 13245 -15390 13330 -15370
rect 13430 -15320 13440 -15290
rect 14920 -15290 15040 -15280
rect 14010 -15310 14130 -15300
rect 14010 -15320 14020 -15310
rect 13430 -15370 14020 -15320
rect 13430 -15390 13505 -15370
rect 13245 -15400 13505 -15390
rect 13245 -15404 13257 -15400
rect 12857 -15410 13257 -15404
rect 13493 -15404 13505 -15400
rect 13881 -15400 14020 -15370
rect 13881 -15404 13893 -15400
rect 13493 -15410 13893 -15404
rect 14010 -15410 14020 -15400
rect 14120 -15320 14130 -15310
rect 14920 -15320 14930 -15290
rect 14120 -15370 14930 -15320
rect 14120 -15400 14469 -15370
rect 14120 -15410 14130 -15400
rect 14457 -15404 14469 -15400
rect 14845 -15390 14930 -15370
rect 15030 -15320 15040 -15290
rect 15030 -15364 15490 -15320
rect 15030 -15370 15493 -15364
rect 15030 -15390 15105 -15370
rect 14845 -15400 15105 -15390
rect 14845 -15404 14857 -15400
rect 14457 -15410 14857 -15404
rect 15093 -15404 15105 -15400
rect 15481 -15404 15493 -15370
rect 15820 -15390 15830 -15270
rect 15950 -15300 15960 -15270
rect 17420 -15270 17560 -15260
rect 15950 -15364 17090 -15300
rect 15950 -15370 17093 -15364
rect 15950 -15390 16069 -15370
rect 15820 -15400 16069 -15390
rect 15093 -15410 15493 -15404
rect 16057 -15404 16069 -15400
rect 16445 -15400 16705 -15370
rect 16445 -15404 16457 -15400
rect 16057 -15410 16457 -15404
rect 16693 -15404 16705 -15400
rect 17081 -15404 17093 -15370
rect 17420 -15390 17430 -15270
rect 17550 -15300 17560 -15270
rect 19020 -15270 19160 -15260
rect 17550 -15364 18690 -15300
rect 17550 -15370 18693 -15364
rect 17550 -15390 17669 -15370
rect 17420 -15400 17669 -15390
rect 16693 -15410 17093 -15404
rect 17657 -15404 17669 -15400
rect 18045 -15400 18305 -15370
rect 18045 -15404 18057 -15400
rect 17657 -15410 18057 -15404
rect 18293 -15404 18305 -15400
rect 18681 -15404 18693 -15370
rect 19020 -15390 19030 -15270
rect 19150 -15300 19160 -15270
rect 20620 -15270 20760 -15260
rect 19150 -15364 20290 -15300
rect 19150 -15370 20293 -15364
rect 19150 -15390 19269 -15370
rect 19020 -15400 19269 -15390
rect 18293 -15410 18693 -15404
rect 19257 -15404 19269 -15400
rect 19645 -15400 19905 -15370
rect 19645 -15404 19657 -15400
rect 19257 -15410 19657 -15404
rect 19893 -15404 19905 -15400
rect 20281 -15404 20293 -15370
rect 20620 -15390 20630 -15270
rect 20750 -15300 20760 -15270
rect 22220 -15270 22360 -15260
rect 20750 -15364 21890 -15300
rect 20750 -15370 21893 -15364
rect 20750 -15390 20869 -15370
rect 20620 -15400 20869 -15390
rect 19893 -15410 20293 -15404
rect 20857 -15404 20869 -15400
rect 21245 -15400 21505 -15370
rect 21245 -15404 21257 -15400
rect 20857 -15410 21257 -15404
rect 21493 -15404 21505 -15400
rect 21881 -15404 21893 -15370
rect 22220 -15390 22230 -15270
rect 22350 -15300 22360 -15270
rect 23820 -15270 23960 -15260
rect 22350 -15364 23490 -15300
rect 22350 -15370 23493 -15364
rect 22350 -15390 22469 -15370
rect 22220 -15400 22469 -15390
rect 21493 -15410 21893 -15404
rect 22457 -15404 22469 -15400
rect 22845 -15400 23105 -15370
rect 22845 -15404 22857 -15400
rect 22457 -15410 22857 -15404
rect 23093 -15404 23105 -15400
rect 23481 -15404 23493 -15370
rect 23820 -15390 23830 -15270
rect 23950 -15300 23960 -15270
rect 27020 -15270 27160 -15260
rect 27020 -15300 27030 -15270
rect 23950 -15364 25090 -15300
rect 25660 -15364 27030 -15300
rect 23950 -15370 25093 -15364
rect 23950 -15390 24069 -15370
rect 23820 -15400 24069 -15390
rect 23093 -15410 23493 -15404
rect 24057 -15404 24069 -15400
rect 24445 -15400 24705 -15370
rect 24445 -15404 24457 -15400
rect 24057 -15410 24457 -15404
rect 24693 -15404 24705 -15400
rect 25081 -15404 25093 -15370
rect 24693 -15410 25093 -15404
rect 25657 -15370 27030 -15364
rect 25657 -15404 25669 -15370
rect 26045 -15400 26305 -15370
rect 26045 -15404 26057 -15400
rect 25657 -15410 26057 -15404
rect 26293 -15404 26305 -15400
rect 26681 -15390 27030 -15370
rect 27150 -15300 27160 -15270
rect 28620 -15270 28760 -15260
rect 27150 -15364 28290 -15300
rect 27150 -15370 28293 -15364
rect 27150 -15390 27269 -15370
rect 26681 -15400 27269 -15390
rect 26681 -15404 26693 -15400
rect 26293 -15410 26693 -15404
rect 27257 -15404 27269 -15400
rect 27645 -15400 27905 -15370
rect 27645 -15404 27657 -15400
rect 27257 -15410 27657 -15404
rect 27893 -15404 27905 -15400
rect 28281 -15404 28293 -15370
rect 28620 -15390 28630 -15270
rect 28750 -15300 28760 -15270
rect 31840 -15280 31980 -15270
rect 28750 -15364 31490 -15300
rect 28750 -15370 31493 -15364
rect 28750 -15390 28869 -15370
rect 28620 -15400 28869 -15390
rect 27893 -15410 28293 -15404
rect 28857 -15404 28869 -15400
rect 29245 -15400 29505 -15370
rect 29245 -15404 29257 -15400
rect 28857 -15410 29257 -15404
rect 29493 -15404 29505 -15400
rect 29881 -15400 30469 -15370
rect 29881 -15404 29893 -15400
rect 29493 -15410 29893 -15404
rect 30457 -15404 30469 -15400
rect 30845 -15400 31105 -15370
rect 30845 -15404 30857 -15400
rect 30457 -15410 30857 -15404
rect 31093 -15404 31105 -15400
rect 31481 -15404 31493 -15370
rect 31093 -15410 31493 -15404
rect 31840 -15400 31850 -15280
rect 31970 -15300 31980 -15280
rect 31970 -15364 36290 -15300
rect 31970 -15370 36293 -15364
rect 31970 -15400 32069 -15370
rect 31840 -15410 31980 -15400
rect 32057 -15404 32069 -15400
rect 32445 -15400 32705 -15370
rect 32445 -15404 32457 -15400
rect 32057 -15410 32457 -15404
rect 32693 -15404 32705 -15400
rect 33081 -15400 33669 -15370
rect 33081 -15404 33093 -15400
rect 32693 -15410 33093 -15404
rect 33657 -15404 33669 -15400
rect 34045 -15400 34305 -15370
rect 34045 -15404 34057 -15400
rect 33657 -15410 34057 -15404
rect 34293 -15404 34305 -15400
rect 34681 -15400 35269 -15370
rect 34681 -15404 34693 -15400
rect 34293 -15410 34693 -15404
rect 35257 -15404 35269 -15400
rect 35645 -15400 35905 -15370
rect 35645 -15404 35657 -15400
rect 35257 -15410 35657 -15404
rect 35893 -15404 35905 -15400
rect 36281 -15404 36293 -15370
rect 35893 -15410 36293 -15404
rect 36857 -15370 37257 -15364
rect 36857 -15404 36869 -15370
rect 37245 -15404 37257 -15370
rect 36857 -15410 37257 -15404
rect 37493 -15370 37893 -15364
rect 37493 -15404 37505 -15370
rect 37881 -15404 37893 -15370
rect 37493 -15410 37893 -15404
rect 57 -15628 490 -15622
rect 57 -15662 69 -15628
rect 445 -15662 490 -15628
rect 57 -15668 490 -15662
rect 440 -15890 490 -15668
rect 57 -15896 490 -15890
rect 57 -15930 69 -15896
rect 445 -15930 490 -15896
rect 57 -15936 490 -15930
rect -30 -15996 16 -15984
rect -30 -16688 -24 -15996
rect 10 -16688 16 -15996
rect -30 -16700 16 -16688
rect 440 -16748 490 -15936
rect 670 -15622 720 -15410
rect 1134 -15457 1180 -15445
rect 1134 -15575 1140 -15457
rect 1174 -15575 1180 -15457
rect 1570 -15457 1616 -15445
rect 1570 -15460 1576 -15457
rect 1134 -15587 1180 -15575
rect 1560 -15575 1576 -15460
rect 1610 -15460 1616 -15457
rect 2098 -15457 2144 -15445
rect 2098 -15460 2104 -15457
rect 1610 -15575 2104 -15460
rect 2138 -15460 2144 -15457
rect 2206 -15457 2252 -15445
rect 2206 -15460 2212 -15457
rect 2138 -15575 2212 -15460
rect 2246 -15460 2252 -15457
rect 2734 -15457 2780 -15445
rect 2734 -15460 2740 -15457
rect 2246 -15575 2740 -15460
rect 2774 -15460 2780 -15457
rect 3170 -15457 3216 -15445
rect 3170 -15460 3176 -15457
rect 2774 -15575 3176 -15460
rect 3210 -15460 3216 -15457
rect 3698 -15457 3744 -15445
rect 3698 -15460 3704 -15457
rect 3210 -15575 3704 -15460
rect 3738 -15460 3744 -15457
rect 3806 -15457 3852 -15445
rect 3806 -15460 3812 -15457
rect 3738 -15575 3812 -15460
rect 3846 -15460 3852 -15457
rect 4334 -15457 4380 -15445
rect 4334 -15460 4340 -15457
rect 3846 -15575 4340 -15460
rect 4374 -15460 4380 -15457
rect 4770 -15457 4816 -15445
rect 4770 -15460 4776 -15457
rect 4374 -15575 4776 -15460
rect 4810 -15460 4816 -15457
rect 5298 -15457 5344 -15445
rect 5298 -15460 5304 -15457
rect 4810 -15575 5304 -15460
rect 5338 -15460 5344 -15457
rect 5406 -15457 5452 -15445
rect 5406 -15460 5412 -15457
rect 5338 -15575 5412 -15460
rect 5446 -15460 5452 -15457
rect 5934 -15457 5980 -15445
rect 5934 -15460 5940 -15457
rect 5446 -15575 5940 -15460
rect 5974 -15460 5980 -15457
rect 6370 -15457 6416 -15445
rect 6370 -15460 6376 -15457
rect 5974 -15575 6376 -15460
rect 6410 -15460 6416 -15457
rect 6898 -15457 6944 -15445
rect 6898 -15460 6904 -15457
rect 6410 -15575 6904 -15460
rect 6938 -15460 6944 -15457
rect 7006 -15457 7052 -15445
rect 7006 -15460 7012 -15457
rect 6938 -15575 7012 -15460
rect 7046 -15460 7052 -15457
rect 7534 -15457 7580 -15445
rect 7534 -15460 7540 -15457
rect 7046 -15575 7540 -15460
rect 7574 -15460 7580 -15457
rect 7970 -15457 8016 -15445
rect 7970 -15460 7976 -15457
rect 7574 -15575 7976 -15460
rect 8010 -15460 8016 -15457
rect 8498 -15457 8544 -15445
rect 8498 -15460 8504 -15457
rect 8010 -15575 8504 -15460
rect 8538 -15460 8544 -15457
rect 8606 -15457 8652 -15445
rect 8606 -15460 8612 -15457
rect 8538 -15575 8612 -15460
rect 8646 -15460 8652 -15457
rect 9134 -15457 9180 -15445
rect 9134 -15460 9140 -15457
rect 8646 -15575 9140 -15460
rect 9174 -15460 9180 -15457
rect 9570 -15457 9616 -15445
rect 9570 -15460 9576 -15457
rect 9174 -15575 9576 -15460
rect 9610 -15460 9616 -15457
rect 10098 -15457 10144 -15445
rect 10098 -15460 10104 -15457
rect 9610 -15575 10104 -15460
rect 10138 -15460 10144 -15457
rect 10206 -15457 10252 -15445
rect 10206 -15460 10212 -15457
rect 10138 -15575 10212 -15460
rect 10246 -15460 10252 -15457
rect 10734 -15450 10780 -15445
rect 10734 -15457 10940 -15450
rect 10734 -15460 10740 -15457
rect 10246 -15575 10740 -15460
rect 10774 -15460 10940 -15457
rect 11170 -15457 11216 -15445
rect 11170 -15460 11176 -15457
rect 10774 -15575 10810 -15460
rect 1560 -15580 10810 -15575
rect 10930 -15575 11176 -15460
rect 11210 -15460 11216 -15457
rect 11400 -15460 11520 -15410
rect 11698 -15457 11744 -15445
rect 11698 -15460 11704 -15457
rect 11210 -15575 11704 -15460
rect 11738 -15460 11744 -15457
rect 11806 -15457 11852 -15445
rect 11806 -15460 11812 -15457
rect 11738 -15575 11812 -15460
rect 11846 -15460 11852 -15457
rect 12040 -15460 12160 -15410
rect 14010 -15420 14130 -15410
rect 12334 -15457 12380 -15445
rect 12334 -15460 12340 -15457
rect 11846 -15575 12340 -15460
rect 12374 -15460 12380 -15457
rect 12770 -15457 12816 -15445
rect 12770 -15460 12776 -15457
rect 12374 -15575 12776 -15460
rect 12810 -15460 12816 -15457
rect 13298 -15457 13344 -15445
rect 13298 -15460 13304 -15457
rect 12810 -15575 13304 -15460
rect 13338 -15460 13344 -15457
rect 13406 -15457 13452 -15445
rect 13406 -15460 13412 -15457
rect 13338 -15575 13412 -15460
rect 13446 -15460 13452 -15457
rect 13934 -15457 13980 -15445
rect 13934 -15460 13940 -15457
rect 13446 -15575 13940 -15460
rect 13974 -15460 13980 -15457
rect 14370 -15457 14416 -15445
rect 14370 -15460 14376 -15457
rect 13974 -15575 14376 -15460
rect 14410 -15460 14416 -15457
rect 14898 -15457 14944 -15445
rect 14898 -15460 14904 -15457
rect 14410 -15575 14904 -15460
rect 14938 -15460 14944 -15457
rect 15006 -15457 15052 -15445
rect 15006 -15460 15012 -15457
rect 14938 -15575 15012 -15460
rect 15046 -15460 15052 -15457
rect 15534 -15457 15580 -15445
rect 15534 -15460 15540 -15457
rect 15046 -15575 15540 -15460
rect 15574 -15460 15580 -15457
rect 15970 -15457 16016 -15445
rect 15970 -15460 15976 -15457
rect 15574 -15575 15976 -15460
rect 16010 -15460 16016 -15457
rect 16498 -15457 16544 -15445
rect 16498 -15460 16504 -15457
rect 16010 -15575 16504 -15460
rect 16538 -15460 16544 -15457
rect 16606 -15457 16652 -15445
rect 16606 -15460 16612 -15457
rect 16538 -15575 16612 -15460
rect 16646 -15460 16652 -15457
rect 17134 -15457 17180 -15445
rect 17134 -15460 17140 -15457
rect 16646 -15575 17140 -15460
rect 17174 -15460 17180 -15457
rect 17570 -15457 17616 -15445
rect 17570 -15460 17576 -15457
rect 17174 -15575 17576 -15460
rect 17610 -15460 17616 -15457
rect 18098 -15457 18144 -15445
rect 18098 -15460 18104 -15457
rect 17610 -15575 18104 -15460
rect 18138 -15460 18144 -15457
rect 18206 -15457 18252 -15445
rect 18206 -15460 18212 -15457
rect 18138 -15575 18212 -15460
rect 18246 -15460 18252 -15457
rect 18734 -15457 18780 -15445
rect 18734 -15460 18740 -15457
rect 18246 -15575 18740 -15460
rect 18774 -15460 18780 -15457
rect 19170 -15457 19216 -15445
rect 19170 -15460 19176 -15457
rect 18774 -15575 19176 -15460
rect 19210 -15460 19216 -15457
rect 19698 -15457 19744 -15445
rect 19698 -15460 19704 -15457
rect 19210 -15575 19704 -15460
rect 19738 -15460 19744 -15457
rect 19806 -15457 19852 -15445
rect 19806 -15460 19812 -15457
rect 19738 -15575 19812 -15460
rect 19846 -15460 19852 -15457
rect 20334 -15457 20380 -15445
rect 20334 -15460 20340 -15457
rect 19846 -15575 20340 -15460
rect 20374 -15460 20380 -15457
rect 20770 -15457 20816 -15445
rect 20770 -15460 20776 -15457
rect 20374 -15575 20776 -15460
rect 20810 -15460 20816 -15457
rect 21298 -15457 21344 -15445
rect 21298 -15460 21304 -15457
rect 20810 -15575 21304 -15460
rect 21338 -15460 21344 -15457
rect 21406 -15457 21452 -15445
rect 21406 -15460 21412 -15457
rect 21338 -15575 21412 -15460
rect 21446 -15460 21452 -15457
rect 21934 -15457 21980 -15445
rect 21934 -15460 21940 -15457
rect 21446 -15575 21940 -15460
rect 21974 -15460 21980 -15457
rect 22370 -15457 22416 -15445
rect 22370 -15460 22376 -15457
rect 21974 -15575 22376 -15460
rect 22410 -15460 22416 -15457
rect 22898 -15457 22944 -15445
rect 22898 -15460 22904 -15457
rect 22410 -15575 22904 -15460
rect 22938 -15460 22944 -15457
rect 23006 -15457 23052 -15445
rect 23006 -15460 23012 -15457
rect 22938 -15575 23012 -15460
rect 23046 -15460 23052 -15457
rect 23534 -15457 23580 -15445
rect 23534 -15460 23540 -15457
rect 23046 -15575 23540 -15460
rect 23574 -15460 23580 -15457
rect 23970 -15457 24016 -15445
rect 23970 -15460 23976 -15457
rect 23574 -15575 23976 -15460
rect 24010 -15460 24016 -15457
rect 24498 -15457 24544 -15445
rect 24498 -15460 24504 -15457
rect 24010 -15575 24504 -15460
rect 24538 -15460 24544 -15457
rect 24606 -15457 24652 -15445
rect 24606 -15460 24612 -15457
rect 24538 -15575 24612 -15460
rect 24646 -15460 24652 -15457
rect 25134 -15457 25180 -15445
rect 25134 -15460 25140 -15457
rect 24646 -15575 25140 -15460
rect 25174 -15460 25180 -15457
rect 25570 -15457 25616 -15445
rect 25570 -15460 25576 -15457
rect 25174 -15575 25576 -15460
rect 25610 -15460 25616 -15457
rect 26098 -15457 26144 -15445
rect 26098 -15460 26104 -15457
rect 25610 -15575 26104 -15460
rect 26138 -15460 26144 -15457
rect 26206 -15457 26252 -15445
rect 26206 -15460 26212 -15457
rect 26138 -15575 26212 -15460
rect 26246 -15460 26252 -15457
rect 26734 -15457 26780 -15445
rect 26734 -15460 26740 -15457
rect 26246 -15575 26740 -15460
rect 26774 -15460 26780 -15457
rect 27170 -15457 27216 -15445
rect 27170 -15460 27176 -15457
rect 26774 -15575 27176 -15460
rect 27210 -15460 27216 -15457
rect 27698 -15457 27744 -15445
rect 27698 -15460 27704 -15457
rect 27210 -15575 27704 -15460
rect 27738 -15460 27744 -15457
rect 27806 -15457 27852 -15445
rect 27806 -15460 27812 -15457
rect 27738 -15575 27812 -15460
rect 27846 -15460 27852 -15457
rect 28334 -15457 28380 -15445
rect 28334 -15460 28340 -15457
rect 27846 -15575 28340 -15460
rect 28374 -15460 28380 -15457
rect 28770 -15457 28816 -15445
rect 28770 -15460 28776 -15457
rect 28374 -15575 28776 -15460
rect 28810 -15460 28816 -15457
rect 29298 -15457 29344 -15445
rect 29298 -15460 29304 -15457
rect 28810 -15575 29304 -15460
rect 29338 -15460 29344 -15457
rect 29406 -15457 29452 -15445
rect 29406 -15460 29412 -15457
rect 29338 -15575 29412 -15460
rect 29446 -15460 29452 -15457
rect 29934 -15457 29980 -15445
rect 29934 -15460 29940 -15457
rect 29446 -15575 29940 -15460
rect 29974 -15460 29980 -15457
rect 30370 -15457 30416 -15445
rect 30370 -15460 30376 -15457
rect 29974 -15575 30376 -15460
rect 30410 -15460 30416 -15457
rect 30898 -15457 30944 -15445
rect 30898 -15460 30904 -15457
rect 30410 -15575 30904 -15460
rect 30938 -15460 30944 -15457
rect 31006 -15457 31052 -15445
rect 31006 -15460 31012 -15457
rect 30938 -15575 31012 -15460
rect 31046 -15460 31052 -15457
rect 31534 -15457 31580 -15445
rect 31534 -15460 31540 -15457
rect 31046 -15575 31540 -15460
rect 31574 -15460 31580 -15457
rect 31970 -15457 32016 -15445
rect 31970 -15460 31976 -15457
rect 31574 -15575 31976 -15460
rect 32010 -15460 32016 -15457
rect 32498 -15457 32544 -15445
rect 32498 -15460 32504 -15457
rect 32010 -15575 32504 -15460
rect 32538 -15460 32544 -15457
rect 32606 -15457 32652 -15445
rect 32606 -15460 32612 -15457
rect 32538 -15575 32612 -15460
rect 32646 -15460 32652 -15457
rect 33134 -15457 33180 -15445
rect 33134 -15460 33140 -15457
rect 32646 -15575 33140 -15460
rect 33174 -15460 33180 -15457
rect 33570 -15457 33616 -15445
rect 33570 -15460 33576 -15457
rect 33174 -15575 33576 -15460
rect 33610 -15460 33616 -15457
rect 34098 -15457 34144 -15445
rect 34098 -15460 34104 -15457
rect 33610 -15575 34104 -15460
rect 34138 -15460 34144 -15457
rect 34206 -15457 34252 -15445
rect 34206 -15460 34212 -15457
rect 34138 -15575 34212 -15460
rect 34246 -15460 34252 -15457
rect 34734 -15457 34780 -15445
rect 34734 -15460 34740 -15457
rect 34246 -15575 34740 -15460
rect 34774 -15460 34780 -15457
rect 35170 -15457 35216 -15445
rect 35170 -15460 35176 -15457
rect 34774 -15575 35176 -15460
rect 35210 -15460 35216 -15457
rect 35698 -15457 35744 -15445
rect 35698 -15460 35704 -15457
rect 35210 -15575 35704 -15460
rect 35738 -15460 35744 -15457
rect 35806 -15457 35852 -15445
rect 35806 -15460 35812 -15457
rect 35738 -15575 35812 -15460
rect 35846 -15460 35852 -15457
rect 36334 -15457 36380 -15445
rect 36334 -15460 36340 -15457
rect 35846 -15575 36340 -15460
rect 36374 -15575 36380 -15457
rect 10930 -15580 36380 -15575
rect 1570 -15587 1616 -15580
rect 2098 -15587 2144 -15580
rect 2206 -15587 2252 -15580
rect 2734 -15587 2780 -15580
rect 3170 -15587 3216 -15580
rect 3698 -15587 3744 -15580
rect 3806 -15587 3852 -15580
rect 4334 -15587 4380 -15580
rect 4770 -15587 4816 -15580
rect 5298 -15587 5344 -15580
rect 5406 -15587 5452 -15580
rect 5934 -15587 5980 -15580
rect 6370 -15587 6416 -15580
rect 6898 -15587 6944 -15580
rect 7006 -15587 7052 -15580
rect 7534 -15587 7580 -15580
rect 7970 -15587 8016 -15580
rect 8498 -15587 8544 -15580
rect 8606 -15587 8652 -15580
rect 9134 -15587 9180 -15580
rect 9570 -15587 9616 -15580
rect 10098 -15587 10144 -15580
rect 10206 -15587 10252 -15580
rect 10734 -15587 10940 -15580
rect 11170 -15587 11216 -15580
rect 10750 -15590 10940 -15587
rect 11400 -15622 11520 -15580
rect 11698 -15587 11744 -15580
rect 11806 -15587 11852 -15580
rect 12040 -15622 12160 -15580
rect 12334 -15587 12380 -15580
rect 12770 -15587 12816 -15580
rect 13298 -15587 13344 -15580
rect 13406 -15587 13452 -15580
rect 13934 -15587 13980 -15580
rect 14370 -15587 14416 -15580
rect 14898 -15587 14944 -15580
rect 15006 -15587 15052 -15580
rect 15534 -15587 15580 -15580
rect 15970 -15587 16016 -15580
rect 16498 -15587 16544 -15580
rect 16606 -15587 16652 -15580
rect 17134 -15587 17180 -15580
rect 17570 -15587 17616 -15580
rect 18098 -15587 18144 -15580
rect 18206 -15587 18252 -15580
rect 18734 -15587 18780 -15580
rect 19170 -15587 19216 -15580
rect 19698 -15587 19744 -15580
rect 19806 -15587 19852 -15580
rect 20334 -15587 20380 -15580
rect 20770 -15587 20816 -15580
rect 21298 -15587 21344 -15580
rect 21406 -15587 21452 -15580
rect 21934 -15587 21980 -15580
rect 22370 -15587 22416 -15580
rect 22898 -15587 22944 -15580
rect 23006 -15587 23052 -15580
rect 23534 -15587 23580 -15580
rect 23970 -15587 24016 -15580
rect 24498 -15587 24544 -15580
rect 24606 -15587 24652 -15580
rect 25134 -15587 25180 -15580
rect 25570 -15587 25616 -15580
rect 26098 -15587 26144 -15580
rect 26206 -15587 26252 -15580
rect 26734 -15587 26780 -15580
rect 27170 -15587 27216 -15580
rect 27698 -15587 27744 -15580
rect 27806 -15587 27852 -15580
rect 28334 -15587 28380 -15580
rect 28770 -15587 28816 -15580
rect 29298 -15587 29344 -15580
rect 29406 -15587 29452 -15580
rect 29934 -15587 29980 -15580
rect 30370 -15587 30416 -15580
rect 30898 -15587 30944 -15580
rect 31006 -15587 31052 -15580
rect 31534 -15587 31580 -15580
rect 31970 -15587 32016 -15580
rect 32498 -15587 32544 -15580
rect 32606 -15587 32652 -15580
rect 33134 -15587 33180 -15580
rect 33570 -15587 33616 -15580
rect 34098 -15587 34144 -15580
rect 34206 -15587 34252 -15580
rect 34734 -15587 34780 -15580
rect 35170 -15587 35216 -15580
rect 35698 -15587 35744 -15580
rect 35806 -15587 35852 -15580
rect 36334 -15587 36380 -15580
rect 36770 -15457 36816 -15445
rect 36770 -15575 36776 -15457
rect 36810 -15575 36816 -15457
rect 36770 -15587 36816 -15575
rect 37298 -15457 37344 -15445
rect 37298 -15575 37304 -15457
rect 37338 -15575 37344 -15457
rect 37298 -15587 37344 -15575
rect 37406 -15457 37452 -15445
rect 37406 -15575 37412 -15457
rect 37446 -15575 37452 -15457
rect 37406 -15587 37452 -15575
rect 37934 -15457 37980 -15445
rect 37934 -15575 37940 -15457
rect 37974 -15575 37980 -15457
rect 37934 -15587 37980 -15575
rect 670 -15628 1093 -15622
rect 670 -15662 705 -15628
rect 1081 -15662 1093 -15628
rect 670 -15668 1093 -15662
rect 1657 -15628 2057 -15622
rect 1657 -15662 1669 -15628
rect 2045 -15630 2057 -15628
rect 2293 -15628 2693 -15622
rect 2293 -15630 2305 -15628
rect 2045 -15662 2060 -15630
rect 1657 -15668 2060 -15662
rect 670 -15890 720 -15668
rect 1420 -15710 1560 -15700
rect 1420 -15830 1430 -15710
rect 1550 -15720 1560 -15710
rect 1660 -15720 2060 -15668
rect 2290 -15662 2305 -15630
rect 2681 -15662 2693 -15628
rect 2290 -15668 2693 -15662
rect 3257 -15628 3657 -15622
rect 3257 -15662 3269 -15628
rect 3645 -15630 3657 -15628
rect 3893 -15628 4293 -15622
rect 3893 -15630 3905 -15628
rect 3645 -15662 3660 -15630
rect 3257 -15668 3660 -15662
rect 2290 -15720 2690 -15668
rect 3020 -15710 3160 -15700
rect 3020 -15720 3030 -15710
rect 1550 -15820 3030 -15720
rect 1550 -15830 1560 -15820
rect 1420 -15840 1560 -15830
rect 1660 -15840 2690 -15820
rect 3020 -15830 3030 -15820
rect 3150 -15720 3160 -15710
rect 3260 -15720 3660 -15668
rect 3890 -15662 3905 -15630
rect 4281 -15662 4293 -15628
rect 3890 -15668 4293 -15662
rect 4857 -15628 5257 -15622
rect 4857 -15662 4869 -15628
rect 5245 -15630 5257 -15628
rect 5493 -15628 5893 -15622
rect 5493 -15630 5505 -15628
rect 5245 -15662 5260 -15630
rect 4857 -15668 5260 -15662
rect 3890 -15720 4290 -15668
rect 4620 -15710 4760 -15700
rect 4620 -15720 4630 -15710
rect 3150 -15820 4630 -15720
rect 3150 -15830 3160 -15820
rect 3020 -15840 3160 -15830
rect 3260 -15840 4290 -15820
rect 4620 -15830 4630 -15820
rect 4750 -15720 4760 -15710
rect 4860 -15720 5260 -15668
rect 5490 -15662 5505 -15630
rect 5881 -15662 5893 -15628
rect 5490 -15668 5893 -15662
rect 6457 -15628 6857 -15622
rect 6457 -15662 6469 -15628
rect 6845 -15630 6857 -15628
rect 7093 -15628 7493 -15622
rect 7093 -15630 7105 -15628
rect 6845 -15662 6860 -15630
rect 6457 -15668 6860 -15662
rect 5490 -15720 5890 -15668
rect 6220 -15710 6360 -15700
rect 6220 -15720 6230 -15710
rect 4750 -15820 6230 -15720
rect 4750 -15830 4760 -15820
rect 4620 -15840 4760 -15830
rect 4860 -15840 5890 -15820
rect 6220 -15830 6230 -15820
rect 6350 -15720 6360 -15710
rect 6460 -15720 6860 -15668
rect 7090 -15662 7105 -15630
rect 7481 -15662 7493 -15628
rect 7090 -15668 7493 -15662
rect 8057 -15628 8457 -15622
rect 8057 -15662 8069 -15628
rect 8445 -15630 8457 -15628
rect 8693 -15628 9093 -15622
rect 8693 -15630 8705 -15628
rect 8445 -15662 8460 -15630
rect 8057 -15668 8460 -15662
rect 7090 -15720 7490 -15668
rect 7820 -15710 7960 -15700
rect 7820 -15720 7830 -15710
rect 6350 -15820 7830 -15720
rect 6350 -15830 6360 -15820
rect 6220 -15840 6360 -15830
rect 6460 -15840 7490 -15820
rect 7820 -15830 7830 -15820
rect 7950 -15720 7960 -15710
rect 8060 -15720 8460 -15668
rect 8690 -15662 8705 -15630
rect 9081 -15662 9093 -15628
rect 8690 -15668 9093 -15662
rect 9657 -15628 10057 -15622
rect 9657 -15662 9669 -15628
rect 10045 -15630 10057 -15628
rect 10293 -15628 10693 -15622
rect 10293 -15630 10305 -15628
rect 10045 -15662 10060 -15630
rect 9657 -15668 10060 -15662
rect 8690 -15720 9090 -15668
rect 9420 -15710 9560 -15700
rect 9420 -15720 9430 -15710
rect 7950 -15820 9430 -15720
rect 7950 -15830 7960 -15820
rect 7820 -15840 7960 -15830
rect 8060 -15840 9090 -15820
rect 9420 -15830 9430 -15820
rect 9550 -15720 9560 -15710
rect 9660 -15720 10060 -15668
rect 10290 -15662 10305 -15630
rect 10681 -15662 10693 -15628
rect 10290 -15668 10693 -15662
rect 11257 -15628 11657 -15622
rect 11257 -15662 11269 -15628
rect 11645 -15662 11657 -15628
rect 11257 -15668 11657 -15662
rect 11893 -15628 12293 -15622
rect 11893 -15662 11905 -15628
rect 12281 -15662 12293 -15628
rect 11893 -15668 12293 -15662
rect 12857 -15628 13257 -15622
rect 12857 -15662 12869 -15628
rect 13245 -15630 13257 -15628
rect 13493 -15628 13893 -15622
rect 13493 -15630 13505 -15628
rect 13245 -15662 13260 -15630
rect 12857 -15668 13260 -15662
rect 10290 -15720 10690 -15668
rect 9550 -15820 10690 -15720
rect 9550 -15830 9560 -15820
rect 9420 -15840 9560 -15830
rect 9660 -15840 10690 -15820
rect 1660 -15890 2060 -15840
rect 670 -15896 1093 -15890
rect 670 -15930 705 -15896
rect 1081 -15930 1093 -15896
rect 670 -15936 1093 -15930
rect 1657 -15896 2060 -15890
rect 1657 -15930 1669 -15896
rect 2045 -15930 2060 -15896
rect 2290 -15890 2690 -15840
rect 3260 -15890 3660 -15840
rect 2290 -15896 2693 -15890
rect 2290 -15930 2305 -15896
rect 2681 -15930 2693 -15896
rect 1657 -15936 2057 -15930
rect 2293 -15936 2693 -15930
rect 3257 -15896 3660 -15890
rect 3257 -15930 3269 -15896
rect 3645 -15930 3660 -15896
rect 3890 -15890 4290 -15840
rect 4860 -15890 5260 -15840
rect 3890 -15896 4293 -15890
rect 3890 -15930 3905 -15896
rect 4281 -15930 4293 -15896
rect 3257 -15936 3657 -15930
rect 3893 -15936 4293 -15930
rect 4857 -15896 5260 -15890
rect 4857 -15930 4869 -15896
rect 5245 -15930 5260 -15896
rect 5490 -15890 5890 -15840
rect 6460 -15890 6860 -15840
rect 5490 -15896 5893 -15890
rect 5490 -15930 5505 -15896
rect 5881 -15930 5893 -15896
rect 4857 -15936 5257 -15930
rect 5493 -15936 5893 -15930
rect 6457 -15896 6860 -15890
rect 6457 -15930 6469 -15896
rect 6845 -15930 6860 -15896
rect 7090 -15890 7490 -15840
rect 8060 -15890 8460 -15840
rect 7090 -15896 7493 -15890
rect 7090 -15930 7105 -15896
rect 7481 -15930 7493 -15896
rect 6457 -15936 6857 -15930
rect 7093 -15936 7493 -15930
rect 8057 -15896 8460 -15890
rect 8057 -15930 8069 -15896
rect 8445 -15930 8460 -15896
rect 8690 -15890 9090 -15840
rect 9660 -15890 10060 -15840
rect 8690 -15896 9093 -15890
rect 8690 -15930 8705 -15896
rect 9081 -15930 9093 -15896
rect 8057 -15936 8457 -15930
rect 8693 -15936 9093 -15930
rect 9657 -15896 10060 -15890
rect 9657 -15930 9669 -15896
rect 10045 -15930 10060 -15896
rect 10290 -15890 10690 -15840
rect 12860 -15710 13260 -15668
rect 13490 -15662 13505 -15630
rect 13881 -15662 13893 -15628
rect 13490 -15668 13893 -15662
rect 14457 -15628 14857 -15622
rect 14457 -15662 14469 -15628
rect 14845 -15630 14857 -15628
rect 15093 -15628 15493 -15622
rect 15093 -15630 15105 -15628
rect 14845 -15662 14860 -15630
rect 14457 -15668 14860 -15662
rect 13490 -15710 13890 -15668
rect 14460 -15710 14860 -15668
rect 15090 -15662 15105 -15630
rect 15481 -15662 15493 -15628
rect 15090 -15668 15493 -15662
rect 16057 -15628 16457 -15622
rect 16057 -15662 16069 -15628
rect 16445 -15662 16457 -15628
rect 16057 -15668 16457 -15662
rect 16693 -15628 17093 -15622
rect 16693 -15662 16705 -15628
rect 17081 -15662 17093 -15628
rect 16693 -15668 17093 -15662
rect 17657 -15628 18057 -15622
rect 17657 -15662 17669 -15628
rect 18045 -15662 18057 -15628
rect 17657 -15668 18057 -15662
rect 18293 -15628 18693 -15622
rect 18293 -15662 18305 -15628
rect 18681 -15662 18693 -15628
rect 18293 -15668 18693 -15662
rect 19257 -15628 19657 -15622
rect 19257 -15662 19269 -15628
rect 19645 -15662 19657 -15628
rect 19257 -15668 19657 -15662
rect 19893 -15628 20293 -15622
rect 19893 -15662 19905 -15628
rect 20281 -15662 20293 -15628
rect 19893 -15668 20293 -15662
rect 20857 -15628 21257 -15622
rect 20857 -15662 20869 -15628
rect 21245 -15662 21257 -15628
rect 20857 -15668 21257 -15662
rect 21493 -15628 21893 -15622
rect 21493 -15662 21505 -15628
rect 21881 -15662 21893 -15628
rect 21493 -15668 21893 -15662
rect 22457 -15628 22857 -15622
rect 22457 -15662 22469 -15628
rect 22845 -15662 22857 -15628
rect 22457 -15668 22857 -15662
rect 23093 -15628 23493 -15622
rect 23093 -15662 23105 -15628
rect 23481 -15662 23493 -15628
rect 23093 -15668 23493 -15662
rect 24057 -15628 24457 -15622
rect 24057 -15662 24069 -15628
rect 24445 -15662 24457 -15628
rect 24057 -15668 24457 -15662
rect 24693 -15628 25093 -15622
rect 24693 -15662 24705 -15628
rect 25081 -15662 25093 -15628
rect 24693 -15668 25093 -15662
rect 25657 -15628 26057 -15622
rect 25657 -15662 25669 -15628
rect 26045 -15662 26057 -15628
rect 25657 -15668 26057 -15662
rect 26293 -15628 26693 -15622
rect 26293 -15662 26305 -15628
rect 26681 -15662 26693 -15628
rect 26293 -15668 26693 -15662
rect 27257 -15628 27657 -15622
rect 27257 -15662 27269 -15628
rect 27645 -15662 27657 -15628
rect 27257 -15668 27657 -15662
rect 27893 -15628 28293 -15622
rect 27893 -15662 27905 -15628
rect 28281 -15662 28293 -15628
rect 27893 -15668 28293 -15662
rect 28857 -15628 29257 -15622
rect 28857 -15662 28869 -15628
rect 29245 -15662 29257 -15628
rect 28857 -15668 29257 -15662
rect 29493 -15628 29893 -15622
rect 29493 -15662 29505 -15628
rect 29881 -15662 29893 -15628
rect 29493 -15668 29893 -15662
rect 30457 -15628 30857 -15622
rect 30457 -15662 30469 -15628
rect 30845 -15662 30857 -15628
rect 30457 -15668 30857 -15662
rect 31093 -15628 31493 -15622
rect 31093 -15662 31105 -15628
rect 31481 -15662 31493 -15628
rect 31093 -15668 31493 -15662
rect 32057 -15628 32457 -15622
rect 32057 -15662 32069 -15628
rect 32445 -15662 32457 -15628
rect 32057 -15668 32457 -15662
rect 32693 -15628 33093 -15622
rect 32693 -15662 32705 -15628
rect 33081 -15662 33093 -15628
rect 32693 -15668 33093 -15662
rect 33657 -15628 34057 -15622
rect 33657 -15662 33669 -15628
rect 34045 -15662 34057 -15628
rect 33657 -15668 34057 -15662
rect 34293 -15628 34693 -15622
rect 34293 -15662 34305 -15628
rect 34681 -15662 34693 -15628
rect 34293 -15668 34693 -15662
rect 35257 -15628 35657 -15622
rect 35257 -15662 35269 -15628
rect 35645 -15662 35657 -15628
rect 35257 -15668 35657 -15662
rect 35893 -15628 36293 -15622
rect 35893 -15662 35905 -15628
rect 36281 -15662 36293 -15628
rect 35893 -15668 36293 -15662
rect 36857 -15628 37257 -15622
rect 36857 -15662 36869 -15628
rect 37245 -15662 37257 -15628
rect 36857 -15668 37257 -15662
rect 37493 -15628 37893 -15622
rect 37493 -15662 37505 -15628
rect 37881 -15662 37893 -15628
rect 37493 -15668 37893 -15662
rect 12860 -15720 15050 -15710
rect 15090 -15720 15490 -15668
rect 12860 -15830 15490 -15720
rect 12860 -15840 13890 -15830
rect 12860 -15890 13260 -15840
rect 10290 -15896 10693 -15890
rect 10290 -15930 10305 -15896
rect 10681 -15930 10693 -15896
rect 9657 -15936 10057 -15930
rect 10293 -15936 10693 -15930
rect 11257 -15896 11657 -15890
rect 11257 -15930 11269 -15896
rect 11645 -15930 11657 -15896
rect 11257 -15936 11657 -15930
rect 11893 -15896 12293 -15890
rect 11893 -15930 11905 -15896
rect 12281 -15930 12293 -15896
rect 11893 -15936 12293 -15930
rect 12857 -15896 13260 -15890
rect 12857 -15930 12869 -15896
rect 13245 -15930 13260 -15896
rect 13490 -15890 13890 -15840
rect 14460 -15840 15490 -15830
rect 14460 -15890 14860 -15840
rect 13490 -15896 13893 -15890
rect 13490 -15930 13505 -15896
rect 13881 -15930 13893 -15896
rect 12857 -15936 13257 -15930
rect 13493 -15936 13893 -15930
rect 14457 -15896 14860 -15890
rect 14457 -15930 14469 -15896
rect 14845 -15930 14860 -15896
rect 15090 -15890 15490 -15840
rect 15600 -15720 15740 -15710
rect 15600 -15840 15610 -15720
rect 15730 -15730 15740 -15720
rect 16060 -15730 16450 -15668
rect 16700 -15730 17090 -15668
rect 15730 -15830 17090 -15730
rect 15730 -15840 15740 -15830
rect 15600 -15850 15740 -15840
rect 16060 -15890 16450 -15830
rect 16700 -15890 17090 -15830
rect 17200 -15720 17340 -15710
rect 17200 -15840 17210 -15720
rect 17330 -15730 17340 -15720
rect 17660 -15730 18050 -15668
rect 18300 -15730 18690 -15668
rect 17330 -15830 18690 -15730
rect 17330 -15840 17340 -15830
rect 17200 -15850 17340 -15840
rect 17660 -15890 18050 -15830
rect 18300 -15890 18690 -15830
rect 18800 -15720 18940 -15710
rect 18800 -15840 18810 -15720
rect 18930 -15730 18940 -15720
rect 19260 -15730 19650 -15668
rect 19900 -15730 20290 -15668
rect 18930 -15830 20290 -15730
rect 18930 -15840 18940 -15830
rect 18800 -15850 18940 -15840
rect 19260 -15890 19650 -15830
rect 19900 -15890 20290 -15830
rect 20400 -15720 20540 -15710
rect 20400 -15840 20410 -15720
rect 20530 -15730 20540 -15720
rect 20860 -15730 21250 -15668
rect 21500 -15730 21890 -15668
rect 20530 -15830 21890 -15730
rect 20530 -15840 20540 -15830
rect 20400 -15850 20540 -15840
rect 20860 -15890 21250 -15830
rect 21500 -15890 21890 -15830
rect 22000 -15720 22140 -15710
rect 22000 -15840 22010 -15720
rect 22130 -15730 22140 -15720
rect 22460 -15730 22850 -15668
rect 23100 -15730 23490 -15668
rect 22130 -15830 23490 -15730
rect 22130 -15840 22140 -15830
rect 22000 -15850 22140 -15840
rect 22460 -15890 22850 -15830
rect 23100 -15890 23490 -15830
rect 23600 -15720 23740 -15710
rect 23600 -15840 23610 -15720
rect 23730 -15730 23740 -15720
rect 24060 -15730 24450 -15668
rect 24700 -15730 25090 -15668
rect 23730 -15830 25090 -15730
rect 23730 -15840 23740 -15830
rect 23600 -15850 23740 -15840
rect 24060 -15890 24450 -15830
rect 24700 -15890 25090 -15830
rect 25660 -15730 26050 -15668
rect 26300 -15730 26690 -15668
rect 26800 -15720 26940 -15710
rect 26800 -15730 26810 -15720
rect 25660 -15830 26810 -15730
rect 25660 -15890 26050 -15830
rect 26300 -15890 26690 -15830
rect 26800 -15840 26810 -15830
rect 26930 -15730 26940 -15720
rect 27260 -15730 27650 -15668
rect 27900 -15730 28290 -15668
rect 26930 -15830 28290 -15730
rect 26930 -15840 26940 -15830
rect 26800 -15850 26940 -15840
rect 27260 -15890 27650 -15830
rect 27900 -15890 28290 -15830
rect 28400 -15720 28540 -15710
rect 28400 -15840 28410 -15720
rect 28530 -15730 28540 -15720
rect 28860 -15730 29250 -15668
rect 29500 -15730 29890 -15668
rect 30460 -15730 30850 -15668
rect 31100 -15730 31490 -15668
rect 28530 -15830 31490 -15730
rect 28530 -15840 28540 -15830
rect 28400 -15850 28540 -15840
rect 28860 -15890 29250 -15830
rect 29500 -15890 29890 -15830
rect 30460 -15890 30850 -15830
rect 31100 -15890 31490 -15830
rect 31580 -15720 31720 -15710
rect 31580 -15840 31590 -15720
rect 31710 -15730 31720 -15720
rect 32060 -15730 32450 -15668
rect 32700 -15730 33090 -15668
rect 33660 -15730 34050 -15668
rect 34300 -15730 34690 -15668
rect 35260 -15730 35650 -15668
rect 35900 -15730 36290 -15668
rect 31710 -15830 36290 -15730
rect 31710 -15840 31720 -15830
rect 31580 -15850 31720 -15840
rect 32060 -15890 32450 -15830
rect 32700 -15890 33090 -15830
rect 33660 -15890 34050 -15830
rect 34300 -15890 34690 -15830
rect 35260 -15890 35650 -15830
rect 35900 -15890 36290 -15830
rect 15090 -15896 15493 -15890
rect 15090 -15930 15105 -15896
rect 15481 -15930 15493 -15896
rect 14457 -15936 14857 -15930
rect 15093 -15936 15493 -15930
rect 16057 -15896 16457 -15890
rect 16057 -15930 16069 -15896
rect 16445 -15930 16457 -15896
rect 16057 -15936 16457 -15930
rect 16693 -15896 17093 -15890
rect 16693 -15930 16705 -15896
rect 17081 -15930 17093 -15896
rect 16693 -15936 17093 -15930
rect 17657 -15896 18057 -15890
rect 17657 -15930 17669 -15896
rect 18045 -15930 18057 -15896
rect 17657 -15936 18057 -15930
rect 18293 -15896 18693 -15890
rect 18293 -15930 18305 -15896
rect 18681 -15930 18693 -15896
rect 18293 -15936 18693 -15930
rect 19257 -15896 19657 -15890
rect 19257 -15930 19269 -15896
rect 19645 -15930 19657 -15896
rect 19257 -15936 19657 -15930
rect 19893 -15896 20293 -15890
rect 19893 -15930 19905 -15896
rect 20281 -15930 20293 -15896
rect 19893 -15936 20293 -15930
rect 20857 -15896 21257 -15890
rect 20857 -15930 20869 -15896
rect 21245 -15930 21257 -15896
rect 20857 -15936 21257 -15930
rect 21493 -15896 21893 -15890
rect 21493 -15930 21505 -15896
rect 21881 -15930 21893 -15896
rect 21493 -15936 21893 -15930
rect 22457 -15896 22857 -15890
rect 22457 -15930 22469 -15896
rect 22845 -15930 22857 -15896
rect 22457 -15936 22857 -15930
rect 23093 -15896 23493 -15890
rect 23093 -15930 23105 -15896
rect 23481 -15930 23493 -15896
rect 23093 -15936 23493 -15930
rect 24057 -15896 24457 -15890
rect 24057 -15930 24069 -15896
rect 24445 -15930 24457 -15896
rect 24057 -15936 24457 -15930
rect 24693 -15896 25093 -15890
rect 24693 -15930 24705 -15896
rect 25081 -15930 25093 -15896
rect 24693 -15936 25093 -15930
rect 25657 -15896 26057 -15890
rect 25657 -15930 25669 -15896
rect 26045 -15930 26057 -15896
rect 25657 -15936 26057 -15930
rect 26293 -15896 26693 -15890
rect 26293 -15930 26305 -15896
rect 26681 -15930 26693 -15896
rect 26293 -15936 26693 -15930
rect 27257 -15896 27657 -15890
rect 27257 -15930 27269 -15896
rect 27645 -15930 27657 -15896
rect 27257 -15936 27657 -15930
rect 27893 -15896 28293 -15890
rect 27893 -15930 27905 -15896
rect 28281 -15930 28293 -15896
rect 27893 -15936 28293 -15930
rect 28857 -15896 29257 -15890
rect 28857 -15930 28869 -15896
rect 29245 -15930 29257 -15896
rect 28857 -15936 29257 -15930
rect 29493 -15896 29893 -15890
rect 29493 -15930 29505 -15896
rect 29881 -15930 29893 -15896
rect 29493 -15936 29893 -15930
rect 30457 -15896 30857 -15890
rect 30457 -15930 30469 -15896
rect 30845 -15930 30857 -15896
rect 30457 -15936 30857 -15930
rect 31093 -15896 31493 -15890
rect 31093 -15930 31105 -15896
rect 31481 -15930 31493 -15896
rect 31093 -15936 31493 -15930
rect 32057 -15896 32457 -15890
rect 32057 -15930 32069 -15896
rect 32445 -15930 32457 -15896
rect 32057 -15936 32457 -15930
rect 32693 -15896 33093 -15890
rect 32693 -15930 32705 -15896
rect 33081 -15930 33093 -15896
rect 32693 -15936 33093 -15930
rect 33657 -15896 34057 -15890
rect 33657 -15930 33669 -15896
rect 34045 -15930 34057 -15896
rect 33657 -15936 34057 -15930
rect 34293 -15896 34693 -15890
rect 34293 -15930 34305 -15896
rect 34681 -15930 34693 -15896
rect 34293 -15936 34693 -15930
rect 35257 -15896 35657 -15890
rect 35257 -15930 35269 -15896
rect 35645 -15930 35657 -15896
rect 35257 -15936 35657 -15930
rect 35893 -15896 36293 -15890
rect 35893 -15930 35905 -15896
rect 36281 -15930 36293 -15896
rect 35893 -15936 36293 -15930
rect 36857 -15896 37257 -15890
rect 36857 -15930 36869 -15896
rect 37245 -15930 37257 -15896
rect 36857 -15936 37257 -15930
rect 37493 -15896 37893 -15890
rect 37493 -15930 37505 -15896
rect 37881 -15930 37893 -15896
rect 37493 -15936 37893 -15930
rect 57 -16754 490 -16748
rect 57 -16760 69 -16754
rect 0 -16788 69 -16760
rect 445 -16788 490 -16754
rect 0 -16888 490 -16788
rect 670 -16748 720 -15936
rect 1134 -15996 1180 -15984
rect 1134 -16688 1140 -15996
rect 1174 -16688 1180 -15996
rect 1134 -16700 1180 -16688
rect 1570 -15996 1616 -15984
rect 1570 -16688 1576 -15996
rect 1610 -16688 1616 -15996
rect 1570 -16700 1616 -16688
rect 2098 -15996 2144 -15984
rect 2098 -16688 2104 -15996
rect 2138 -16000 2144 -15996
rect 2206 -15996 2252 -15984
rect 2206 -16000 2212 -15996
rect 2138 -16010 2212 -16000
rect 2138 -16680 2212 -16670
rect 2138 -16688 2144 -16680
rect 2098 -16700 2144 -16688
rect 2206 -16688 2212 -16680
rect 2246 -16688 2252 -15996
rect 2206 -16700 2252 -16688
rect 2734 -15996 2780 -15984
rect 2734 -16688 2740 -15996
rect 2774 -16688 2780 -15996
rect 2734 -16700 2780 -16688
rect 3170 -15996 3216 -15984
rect 3170 -16688 3176 -15996
rect 3210 -16688 3216 -15996
rect 3170 -16700 3216 -16688
rect 3698 -15996 3744 -15984
rect 3698 -16688 3704 -15996
rect 3738 -16000 3744 -15996
rect 3806 -15996 3852 -15984
rect 3806 -16000 3812 -15996
rect 3738 -16010 3812 -16000
rect 3738 -16680 3812 -16670
rect 3738 -16688 3744 -16680
rect 3698 -16700 3744 -16688
rect 3806 -16688 3812 -16680
rect 3846 -16688 3852 -15996
rect 3806 -16700 3852 -16688
rect 4334 -15996 4380 -15984
rect 4334 -16688 4340 -15996
rect 4374 -16688 4380 -15996
rect 4334 -16700 4380 -16688
rect 4770 -15996 4816 -15984
rect 4770 -16688 4776 -15996
rect 4810 -16688 4816 -15996
rect 4770 -16700 4816 -16688
rect 5298 -15996 5344 -15984
rect 5298 -16688 5304 -15996
rect 5338 -16000 5344 -15996
rect 5406 -15996 5452 -15984
rect 5406 -16000 5412 -15996
rect 5338 -16010 5412 -16000
rect 5338 -16680 5412 -16670
rect 5338 -16688 5344 -16680
rect 5298 -16700 5344 -16688
rect 5406 -16688 5412 -16680
rect 5446 -16688 5452 -15996
rect 5406 -16700 5452 -16688
rect 5934 -15996 5980 -15984
rect 5934 -16688 5940 -15996
rect 5974 -16688 5980 -15996
rect 5934 -16700 5980 -16688
rect 6370 -15996 6416 -15984
rect 6370 -16688 6376 -15996
rect 6410 -16688 6416 -15996
rect 6370 -16700 6416 -16688
rect 6898 -15996 6944 -15984
rect 6898 -16688 6904 -15996
rect 6938 -16000 6944 -15996
rect 7006 -15996 7052 -15984
rect 7006 -16000 7012 -15996
rect 6938 -16010 7012 -16000
rect 6938 -16680 7012 -16670
rect 6938 -16688 6944 -16680
rect 6898 -16700 6944 -16688
rect 7006 -16688 7012 -16680
rect 7046 -16688 7052 -15996
rect 7006 -16700 7052 -16688
rect 7534 -15996 7580 -15984
rect 7534 -16688 7540 -15996
rect 7574 -16688 7580 -15996
rect 7534 -16700 7580 -16688
rect 7970 -15996 8016 -15984
rect 7970 -16688 7976 -15996
rect 8010 -16688 8016 -15996
rect 7970 -16700 8016 -16688
rect 8498 -15996 8544 -15984
rect 8498 -16688 8504 -15996
rect 8538 -16000 8544 -15996
rect 8606 -15996 8652 -15984
rect 8606 -16000 8612 -15996
rect 8538 -16010 8612 -16000
rect 8538 -16680 8612 -16670
rect 8538 -16688 8544 -16680
rect 8498 -16700 8544 -16688
rect 8606 -16688 8612 -16680
rect 8646 -16688 8652 -15996
rect 8606 -16700 8652 -16688
rect 9134 -15996 9180 -15984
rect 9134 -16688 9140 -15996
rect 9174 -16688 9180 -15996
rect 9134 -16700 9180 -16688
rect 9570 -15996 9616 -15984
rect 9570 -16688 9576 -15996
rect 9610 -16688 9616 -15996
rect 9570 -16700 9616 -16688
rect 10098 -15996 10144 -15984
rect 10098 -16688 10104 -15996
rect 10138 -16000 10144 -15996
rect 10206 -15996 10252 -15984
rect 10206 -16000 10212 -15996
rect 10138 -16010 10212 -16000
rect 10138 -16680 10212 -16670
rect 10138 -16688 10144 -16680
rect 10098 -16700 10144 -16688
rect 10206 -16688 10212 -16680
rect 10246 -16688 10252 -15996
rect 10206 -16700 10252 -16688
rect 10734 -15996 10780 -15984
rect 10734 -16688 10740 -15996
rect 10774 -16688 10780 -15996
rect 10734 -16700 10780 -16688
rect 11170 -15996 11216 -15984
rect 11170 -16688 11176 -15996
rect 11210 -16290 11216 -15996
rect 11420 -16290 11500 -15936
rect 11698 -15996 11744 -15984
rect 11698 -16290 11704 -15996
rect 11210 -16410 11704 -16290
rect 11210 -16688 11216 -16410
rect 11170 -16700 11216 -16688
rect 11420 -16748 11500 -16410
rect 11698 -16688 11704 -16410
rect 11738 -16290 11744 -15996
rect 11806 -15996 11852 -15984
rect 11806 -16290 11812 -15996
rect 11738 -16410 11812 -16290
rect 11738 -16688 11744 -16410
rect 11698 -16700 11744 -16688
rect 11806 -16688 11812 -16410
rect 11846 -16290 11852 -15996
rect 12040 -16290 12120 -15936
rect 12334 -15996 12380 -15984
rect 12334 -16290 12340 -15996
rect 11846 -16410 12340 -16290
rect 11846 -16688 11852 -16410
rect 11806 -16700 11852 -16688
rect 12040 -16748 12120 -16410
rect 12334 -16688 12340 -16410
rect 12374 -16688 12380 -15996
rect 12334 -16700 12380 -16688
rect 12770 -15996 12816 -15984
rect 12770 -16688 12776 -15996
rect 12810 -16688 12816 -15996
rect 12770 -16700 12816 -16688
rect 13298 -15996 13344 -15984
rect 13298 -16688 13304 -15996
rect 13338 -16000 13344 -15996
rect 13406 -15996 13452 -15984
rect 13406 -16000 13412 -15996
rect 13338 -16010 13412 -16000
rect 13338 -16680 13412 -16670
rect 13338 -16688 13344 -16680
rect 13298 -16700 13344 -16688
rect 13406 -16688 13412 -16680
rect 13446 -16688 13452 -15996
rect 13406 -16700 13452 -16688
rect 13934 -15996 13980 -15984
rect 13934 -16688 13940 -15996
rect 13974 -16688 13980 -15996
rect 13934 -16700 13980 -16688
rect 14370 -15996 14416 -15984
rect 14370 -16688 14376 -15996
rect 14410 -16688 14416 -15996
rect 14370 -16700 14416 -16688
rect 14898 -15996 14944 -15984
rect 14898 -16688 14904 -15996
rect 14938 -16000 14944 -15996
rect 15006 -15996 15052 -15984
rect 15006 -16000 15012 -15996
rect 14938 -16010 15012 -16000
rect 14938 -16680 15012 -16670
rect 14938 -16688 14944 -16680
rect 14898 -16700 14944 -16688
rect 15006 -16688 15012 -16680
rect 15046 -16688 15052 -15996
rect 15006 -16700 15052 -16688
rect 15534 -15996 15580 -15984
rect 15534 -16688 15540 -15996
rect 15574 -16688 15580 -15996
rect 15534 -16700 15580 -16688
rect 15970 -15996 16016 -15984
rect 15970 -16688 15976 -15996
rect 16010 -16688 16016 -15996
rect 15970 -16700 16016 -16688
rect 16498 -15990 16544 -15984
rect 16606 -15990 16652 -15984
rect 16498 -15996 16652 -15990
rect 16498 -16688 16504 -15996
rect 16538 -16000 16612 -15996
rect 16538 -16688 16612 -16680
rect 16646 -16688 16652 -15996
rect 16498 -16690 16652 -16688
rect 16498 -16700 16544 -16690
rect 16606 -16700 16652 -16690
rect 17134 -15996 17180 -15984
rect 17134 -16688 17140 -15996
rect 17174 -16688 17180 -15996
rect 17134 -16700 17180 -16688
rect 17570 -15996 17616 -15984
rect 17570 -16688 17576 -15996
rect 17610 -16688 17616 -15996
rect 17570 -16700 17616 -16688
rect 18098 -15990 18144 -15984
rect 18206 -15990 18252 -15984
rect 18098 -15996 18252 -15990
rect 18098 -16688 18104 -15996
rect 18138 -16000 18212 -15996
rect 18138 -16688 18212 -16680
rect 18246 -16688 18252 -15996
rect 18098 -16690 18252 -16688
rect 18098 -16700 18144 -16690
rect 18206 -16700 18252 -16690
rect 18734 -15996 18780 -15984
rect 18734 -16688 18740 -15996
rect 18774 -16688 18780 -15996
rect 18734 -16700 18780 -16688
rect 19170 -15996 19216 -15984
rect 19170 -16688 19176 -15996
rect 19210 -16688 19216 -15996
rect 19170 -16700 19216 -16688
rect 19698 -15990 19744 -15984
rect 19806 -15990 19852 -15984
rect 19698 -15996 19852 -15990
rect 19698 -16688 19704 -15996
rect 19738 -16000 19812 -15996
rect 19738 -16688 19812 -16680
rect 19846 -16688 19852 -15996
rect 19698 -16690 19852 -16688
rect 19698 -16700 19744 -16690
rect 19806 -16700 19852 -16690
rect 20334 -15996 20380 -15984
rect 20334 -16688 20340 -15996
rect 20374 -16688 20380 -15996
rect 20334 -16700 20380 -16688
rect 20770 -15996 20816 -15984
rect 20770 -16688 20776 -15996
rect 20810 -16688 20816 -15996
rect 20770 -16700 20816 -16688
rect 21298 -15990 21344 -15984
rect 21406 -15990 21452 -15984
rect 21298 -15996 21452 -15990
rect 21298 -16688 21304 -15996
rect 21338 -16000 21412 -15996
rect 21338 -16688 21412 -16680
rect 21446 -16688 21452 -15996
rect 21298 -16690 21452 -16688
rect 21298 -16700 21344 -16690
rect 21406 -16700 21452 -16690
rect 21934 -15996 21980 -15984
rect 21934 -16688 21940 -15996
rect 21974 -16688 21980 -15996
rect 21934 -16700 21980 -16688
rect 22370 -15996 22416 -15984
rect 22370 -16688 22376 -15996
rect 22410 -16688 22416 -15996
rect 22370 -16700 22416 -16688
rect 22898 -15990 22944 -15984
rect 23006 -15990 23052 -15984
rect 22898 -15996 23052 -15990
rect 22898 -16688 22904 -15996
rect 22938 -16000 23012 -15996
rect 22938 -16688 23012 -16680
rect 23046 -16688 23052 -15996
rect 22898 -16690 23052 -16688
rect 22898 -16700 22944 -16690
rect 23006 -16700 23052 -16690
rect 23534 -15996 23580 -15984
rect 23534 -16688 23540 -15996
rect 23574 -16688 23580 -15996
rect 23534 -16700 23580 -16688
rect 23970 -15996 24016 -15984
rect 23970 -16688 23976 -15996
rect 24010 -16688 24016 -15996
rect 23970 -16700 24016 -16688
rect 24498 -15990 24544 -15984
rect 24606 -15990 24652 -15984
rect 24498 -15996 24652 -15990
rect 24498 -16688 24504 -15996
rect 24538 -16000 24612 -15996
rect 24538 -16688 24612 -16680
rect 24646 -16688 24652 -15996
rect 24498 -16690 24652 -16688
rect 24498 -16700 24544 -16690
rect 24606 -16700 24652 -16690
rect 25134 -15996 25180 -15984
rect 25134 -16688 25140 -15996
rect 25174 -16688 25180 -15996
rect 25134 -16700 25180 -16688
rect 25570 -15996 25616 -15984
rect 25570 -16688 25576 -15996
rect 25610 -16688 25616 -15996
rect 25570 -16700 25616 -16688
rect 26098 -15990 26144 -15984
rect 26206 -15990 26252 -15984
rect 26098 -15996 26252 -15990
rect 26098 -16688 26104 -15996
rect 26138 -16000 26212 -15996
rect 26138 -16688 26212 -16680
rect 26246 -16688 26252 -15996
rect 26098 -16690 26252 -16688
rect 26098 -16700 26144 -16690
rect 26206 -16700 26252 -16690
rect 26734 -15996 26780 -15984
rect 26734 -16688 26740 -15996
rect 26774 -16688 26780 -15996
rect 26734 -16700 26780 -16688
rect 27170 -15996 27216 -15984
rect 27170 -16688 27176 -15996
rect 27210 -16688 27216 -15996
rect 27170 -16700 27216 -16688
rect 27698 -15990 27744 -15984
rect 27806 -15990 27852 -15984
rect 27698 -15996 27852 -15990
rect 27698 -16688 27704 -15996
rect 27738 -16000 27812 -15996
rect 27738 -16688 27812 -16680
rect 27846 -16688 27852 -15996
rect 27698 -16690 27852 -16688
rect 27698 -16700 27744 -16690
rect 27806 -16700 27852 -16690
rect 28334 -15996 28380 -15984
rect 28334 -16688 28340 -15996
rect 28374 -16688 28380 -15996
rect 28334 -16700 28380 -16688
rect 28770 -15996 28816 -15984
rect 28770 -16688 28776 -15996
rect 28810 -16688 28816 -15996
rect 28770 -16700 28816 -16688
rect 29298 -15990 29344 -15984
rect 29406 -15990 29452 -15984
rect 29298 -15996 29452 -15990
rect 29298 -16688 29304 -15996
rect 29338 -16000 29412 -15996
rect 29338 -16688 29412 -16680
rect 29446 -16688 29452 -15996
rect 29298 -16690 29452 -16688
rect 29298 -16700 29344 -16690
rect 29406 -16700 29452 -16690
rect 29934 -15996 29980 -15984
rect 29934 -16688 29940 -15996
rect 29974 -16688 29980 -15996
rect 29934 -16700 29980 -16688
rect 30370 -15996 30416 -15984
rect 30370 -16688 30376 -15996
rect 30410 -16688 30416 -15996
rect 30370 -16700 30416 -16688
rect 30898 -15990 30944 -15984
rect 31006 -15990 31052 -15984
rect 30898 -15996 31052 -15990
rect 30898 -16688 30904 -15996
rect 30938 -16000 31012 -15996
rect 30938 -16688 31012 -16680
rect 31046 -16688 31052 -15996
rect 30898 -16690 31052 -16688
rect 30898 -16700 30944 -16690
rect 31006 -16700 31052 -16690
rect 31534 -15996 31580 -15984
rect 31534 -16688 31540 -15996
rect 31574 -16688 31580 -15996
rect 31534 -16700 31580 -16688
rect 31970 -15996 32016 -15984
rect 31970 -16688 31976 -15996
rect 32010 -16688 32016 -15996
rect 31970 -16700 32016 -16688
rect 32498 -15990 32544 -15984
rect 32606 -15990 32652 -15984
rect 32498 -15996 32652 -15990
rect 32498 -16688 32504 -15996
rect 32538 -16000 32612 -15996
rect 32538 -16688 32612 -16680
rect 32646 -16688 32652 -15996
rect 32498 -16690 32652 -16688
rect 32498 -16700 32544 -16690
rect 32606 -16700 32652 -16690
rect 33134 -15996 33180 -15984
rect 33134 -16688 33140 -15996
rect 33174 -16688 33180 -15996
rect 33134 -16700 33180 -16688
rect 33570 -15996 33616 -15984
rect 33570 -16688 33576 -15996
rect 33610 -16688 33616 -15996
rect 33570 -16700 33616 -16688
rect 34098 -15990 34144 -15984
rect 34206 -15990 34252 -15984
rect 34098 -15996 34252 -15990
rect 34098 -16688 34104 -15996
rect 34138 -16000 34212 -15996
rect 34138 -16688 34212 -16680
rect 34246 -16688 34252 -15996
rect 34098 -16690 34252 -16688
rect 34098 -16700 34144 -16690
rect 34206 -16700 34252 -16690
rect 34734 -15996 34780 -15984
rect 34734 -16688 34740 -15996
rect 34774 -16688 34780 -15996
rect 34734 -16700 34780 -16688
rect 35170 -15996 35216 -15984
rect 35170 -16688 35176 -15996
rect 35210 -16688 35216 -15996
rect 35170 -16700 35216 -16688
rect 35698 -15990 35744 -15984
rect 35806 -15990 35852 -15984
rect 35698 -15996 35852 -15990
rect 35698 -16688 35704 -15996
rect 35738 -16000 35812 -15996
rect 35738 -16688 35812 -16680
rect 35846 -16688 35852 -15996
rect 35698 -16690 35852 -16688
rect 35698 -16700 35744 -16690
rect 35806 -16700 35852 -16690
rect 36334 -15996 36380 -15984
rect 36334 -16688 36340 -15996
rect 36374 -16688 36380 -15996
rect 36334 -16700 36380 -16688
rect 36770 -15996 36816 -15984
rect 36770 -16688 36776 -15996
rect 36810 -16688 36816 -15996
rect 36770 -16700 36816 -16688
rect 37298 -15996 37344 -15984
rect 37298 -16688 37304 -15996
rect 37338 -16688 37344 -15996
rect 37298 -16700 37344 -16688
rect 37406 -15996 37452 -15984
rect 37406 -16688 37412 -15996
rect 37446 -16688 37452 -15996
rect 37406 -16700 37452 -16688
rect 37934 -15996 37980 -15984
rect 37934 -16688 37940 -15996
rect 37974 -16688 37980 -15996
rect 37934 -16700 37980 -16688
rect 670 -16754 1093 -16748
rect 670 -16788 705 -16754
rect 1081 -16760 1093 -16754
rect 1657 -16754 2057 -16748
rect 1657 -16760 1669 -16754
rect 1081 -16788 1669 -16760
rect 2045 -16760 2057 -16754
rect 2293 -16754 2693 -16748
rect 2293 -16760 2305 -16754
rect 2045 -16788 2305 -16760
rect 2681 -16760 2693 -16754
rect 3257 -16754 3657 -16748
rect 3257 -16760 3269 -16754
rect 2681 -16788 3269 -16760
rect 3645 -16760 3657 -16754
rect 3893 -16754 4293 -16748
rect 3893 -16760 3905 -16754
rect 3645 -16788 3905 -16760
rect 4281 -16760 4293 -16754
rect 4857 -16754 5257 -16748
rect 4857 -16760 4869 -16754
rect 4281 -16788 4869 -16760
rect 5245 -16760 5257 -16754
rect 5493 -16754 5893 -16748
rect 5493 -16760 5505 -16754
rect 5245 -16788 5505 -16760
rect 5881 -16760 5893 -16754
rect 6457 -16754 6857 -16748
rect 6457 -16760 6469 -16754
rect 5881 -16788 6469 -16760
rect 6845 -16760 6857 -16754
rect 7093 -16754 7493 -16748
rect 7093 -16760 7105 -16754
rect 6845 -16788 7105 -16760
rect 7481 -16760 7493 -16754
rect 8057 -16754 8457 -16748
rect 8057 -16760 8069 -16754
rect 7481 -16788 8069 -16760
rect 8445 -16760 8457 -16754
rect 8693 -16754 9093 -16748
rect 8693 -16760 8705 -16754
rect 8445 -16788 8705 -16760
rect 9081 -16760 9093 -16754
rect 9657 -16754 10057 -16748
rect 9657 -16760 9669 -16754
rect 9081 -16788 9669 -16760
rect 10045 -16760 10057 -16754
rect 10293 -16754 10693 -16748
rect 10293 -16760 10305 -16754
rect 10045 -16788 10305 -16760
rect 10681 -16760 10693 -16754
rect 11257 -16754 11657 -16748
rect 11257 -16760 11269 -16754
rect 10681 -16788 11269 -16760
rect 11645 -16760 11657 -16754
rect 11893 -16754 12293 -16748
rect 11893 -16760 11905 -16754
rect 11645 -16788 11905 -16760
rect 12281 -16760 12293 -16754
rect 12857 -16754 13257 -16748
rect 12857 -16760 12869 -16754
rect 12281 -16788 12869 -16760
rect 13245 -16760 13257 -16754
rect 13493 -16754 13893 -16748
rect 13493 -16760 13505 -16754
rect 13245 -16788 13505 -16760
rect 13881 -16760 13893 -16754
rect 14457 -16754 14857 -16748
rect 14457 -16760 14469 -16754
rect 13881 -16788 14469 -16760
rect 14845 -16760 14857 -16754
rect 15093 -16754 15493 -16748
rect 15093 -16760 15105 -16754
rect 14845 -16788 15105 -16760
rect 15481 -16760 15493 -16754
rect 16057 -16754 16457 -16748
rect 16057 -16760 16069 -16754
rect 15481 -16788 16069 -16760
rect 16445 -16760 16457 -16754
rect 16693 -16754 17093 -16748
rect 16693 -16760 16705 -16754
rect 16445 -16788 16705 -16760
rect 17081 -16760 17093 -16754
rect 17657 -16754 18057 -16748
rect 17657 -16760 17669 -16754
rect 17081 -16788 17669 -16760
rect 18045 -16760 18057 -16754
rect 18293 -16754 18693 -16748
rect 18293 -16760 18305 -16754
rect 18045 -16788 18305 -16760
rect 18681 -16760 18693 -16754
rect 19257 -16754 19657 -16748
rect 19257 -16760 19269 -16754
rect 18681 -16788 19269 -16760
rect 19645 -16760 19657 -16754
rect 19893 -16754 20293 -16748
rect 19893 -16760 19905 -16754
rect 19645 -16788 19905 -16760
rect 20281 -16760 20293 -16754
rect 20857 -16754 21257 -16748
rect 20857 -16760 20869 -16754
rect 20281 -16788 20869 -16760
rect 21245 -16760 21257 -16754
rect 21493 -16754 21893 -16748
rect 21493 -16760 21505 -16754
rect 21245 -16788 21505 -16760
rect 21881 -16760 21893 -16754
rect 22457 -16754 22857 -16748
rect 22457 -16760 22469 -16754
rect 21881 -16788 22469 -16760
rect 22845 -16760 22857 -16754
rect 23093 -16754 23493 -16748
rect 23093 -16760 23105 -16754
rect 22845 -16788 23105 -16760
rect 23481 -16760 23493 -16754
rect 24057 -16754 24457 -16748
rect 24057 -16760 24069 -16754
rect 23481 -16788 24069 -16760
rect 24445 -16760 24457 -16754
rect 24693 -16754 25093 -16748
rect 24693 -16760 24705 -16754
rect 24445 -16788 24705 -16760
rect 25081 -16760 25093 -16754
rect 25657 -16754 26057 -16748
rect 25657 -16760 25669 -16754
rect 25081 -16788 25669 -16760
rect 26045 -16760 26057 -16754
rect 26293 -16754 26693 -16748
rect 26293 -16760 26305 -16754
rect 26045 -16788 26305 -16760
rect 26681 -16760 26693 -16754
rect 27257 -16754 27657 -16748
rect 27257 -16760 27269 -16754
rect 26681 -16788 27269 -16760
rect 27645 -16760 27657 -16754
rect 27893 -16754 28293 -16748
rect 27893 -16760 27905 -16754
rect 27645 -16788 27905 -16760
rect 28281 -16760 28293 -16754
rect 28857 -16754 29257 -16748
rect 28857 -16760 28869 -16754
rect 28281 -16788 28869 -16760
rect 29245 -16760 29257 -16754
rect 29493 -16754 29893 -16748
rect 29493 -16760 29505 -16754
rect 29245 -16788 29505 -16760
rect 29881 -16760 29893 -16754
rect 30457 -16754 30857 -16748
rect 30457 -16760 30469 -16754
rect 29881 -16788 30469 -16760
rect 30845 -16760 30857 -16754
rect 31093 -16754 31493 -16748
rect 31093 -16760 31105 -16754
rect 30845 -16788 31105 -16760
rect 31481 -16760 31493 -16754
rect 32057 -16754 32457 -16748
rect 32057 -16760 32069 -16754
rect 31481 -16788 32069 -16760
rect 32445 -16760 32457 -16754
rect 32693 -16754 33093 -16748
rect 32693 -16760 32705 -16754
rect 32445 -16788 32705 -16760
rect 33081 -16760 33093 -16754
rect 33657 -16754 34057 -16748
rect 33657 -16760 33669 -16754
rect 33081 -16788 33669 -16760
rect 34045 -16760 34057 -16754
rect 34293 -16754 34693 -16748
rect 34293 -16760 34305 -16754
rect 34045 -16788 34305 -16760
rect 34681 -16760 34693 -16754
rect 35257 -16754 35657 -16748
rect 35257 -16760 35269 -16754
rect 34681 -16788 35269 -16760
rect 35645 -16760 35657 -16754
rect 35893 -16754 36293 -16748
rect 35893 -16760 35905 -16754
rect 35645 -16788 35905 -16760
rect 36281 -16760 36293 -16754
rect 36857 -16754 37257 -16748
rect 36857 -16760 36869 -16754
rect 36281 -16788 36869 -16760
rect 37245 -16760 37257 -16754
rect 37493 -16754 37893 -16748
rect 37493 -16760 37505 -16754
rect 37245 -16788 37505 -16760
rect 37881 -16788 37893 -16754
rect 670 -16794 37893 -16788
rect 670 -16882 37880 -16794
rect 670 -16888 37949 -16882
rect 0 -16922 13 -16888
rect 1137 -16922 1613 -16888
rect 2737 -16922 3213 -16888
rect 4337 -16922 4813 -16888
rect 5937 -16922 6413 -16888
rect 7537 -16922 8013 -16888
rect 9137 -16922 9613 -16888
rect 10737 -16922 11213 -16888
rect 12337 -16922 12813 -16888
rect 13937 -16922 14413 -16888
rect 15537 -16922 16013 -16888
rect 17137 -16922 17613 -16888
rect 18737 -16922 19213 -16888
rect 20337 -16922 20813 -16888
rect 21937 -16922 22413 -16888
rect 23537 -16922 24013 -16888
rect 25137 -16922 25613 -16888
rect 26737 -16922 27213 -16888
rect 28337 -16922 28813 -16888
rect 29937 -16922 30413 -16888
rect 31537 -16922 32013 -16888
rect 33137 -16922 33613 -16888
rect 34737 -16922 35213 -16888
rect 36337 -16922 36813 -16888
rect 37937 -16922 37949 -16888
rect 0 -17020 490 -16922
rect 440 -17164 490 -17020
rect 57 -17170 490 -17164
rect 57 -17204 69 -17170
rect 445 -17204 490 -17170
rect 57 -17210 490 -17204
rect -30 -17257 16 -17245
rect -30 -17375 -24 -17257
rect 10 -17375 16 -17257
rect -30 -17387 16 -17375
rect 440 -17422 490 -17210
rect 670 -16928 37949 -16922
rect 670 -17020 37940 -16928
rect 670 -17164 720 -17020
rect 1200 -17070 1340 -17060
rect 670 -17170 1093 -17164
rect 670 -17204 705 -17170
rect 1081 -17204 1093 -17170
rect 1200 -17190 1210 -17070
rect 1330 -17080 1340 -17070
rect 2800 -17070 2940 -17060
rect 2800 -17080 2810 -17070
rect 1330 -17170 2810 -17080
rect 1330 -17180 1669 -17170
rect 1330 -17190 1340 -17180
rect 1200 -17200 1340 -17190
rect 670 -17210 1093 -17204
rect 1657 -17204 1669 -17180
rect 2045 -17180 2305 -17170
rect 2045 -17204 2057 -17180
rect 1657 -17210 2057 -17204
rect 2293 -17204 2305 -17180
rect 2681 -17180 2810 -17170
rect 2681 -17204 2693 -17180
rect 2800 -17190 2810 -17180
rect 2930 -17080 2940 -17070
rect 4400 -17070 4540 -17060
rect 4400 -17080 4410 -17070
rect 2930 -17170 4410 -17080
rect 2930 -17180 3269 -17170
rect 2930 -17190 2940 -17180
rect 2800 -17200 2940 -17190
rect 2293 -17210 2693 -17204
rect 3257 -17204 3269 -17180
rect 3645 -17180 3905 -17170
rect 3645 -17204 3657 -17180
rect 3257 -17210 3657 -17204
rect 3893 -17204 3905 -17180
rect 4281 -17180 4410 -17170
rect 4281 -17204 4293 -17180
rect 4400 -17190 4410 -17180
rect 4530 -17080 4540 -17070
rect 6000 -17070 6140 -17060
rect 6000 -17080 6010 -17070
rect 4530 -17170 6010 -17080
rect 4530 -17180 4869 -17170
rect 4530 -17190 4540 -17180
rect 4400 -17200 4540 -17190
rect 3893 -17210 4293 -17204
rect 4857 -17204 4869 -17180
rect 5245 -17180 5505 -17170
rect 5245 -17204 5257 -17180
rect 4857 -17210 5257 -17204
rect 5493 -17204 5505 -17180
rect 5881 -17180 6010 -17170
rect 5881 -17204 5893 -17180
rect 6000 -17190 6010 -17180
rect 6130 -17080 6140 -17070
rect 7600 -17070 7740 -17060
rect 7600 -17080 7610 -17070
rect 6130 -17170 7610 -17080
rect 6130 -17180 6469 -17170
rect 6130 -17190 6140 -17180
rect 6000 -17200 6140 -17190
rect 5493 -17210 5893 -17204
rect 6457 -17204 6469 -17180
rect 6845 -17180 7105 -17170
rect 6845 -17204 6857 -17180
rect 6457 -17210 6857 -17204
rect 7093 -17204 7105 -17180
rect 7481 -17180 7610 -17170
rect 7481 -17204 7493 -17180
rect 7600 -17190 7610 -17180
rect 7730 -17080 7740 -17070
rect 9200 -17070 9340 -17060
rect 15820 -17070 15960 -17060
rect 9200 -17080 9210 -17070
rect 7730 -17170 9210 -17080
rect 7730 -17180 8069 -17170
rect 7730 -17190 7740 -17180
rect 7600 -17200 7740 -17190
rect 7093 -17210 7493 -17204
rect 8057 -17204 8069 -17180
rect 8445 -17180 8705 -17170
rect 8445 -17204 8457 -17180
rect 8057 -17210 8457 -17204
rect 8693 -17204 8705 -17180
rect 9081 -17180 9210 -17170
rect 9081 -17204 9093 -17180
rect 9200 -17190 9210 -17180
rect 9330 -17080 9340 -17070
rect 12620 -17080 12760 -17070
rect 9330 -17170 10700 -17080
rect 9330 -17180 9669 -17170
rect 9330 -17190 9340 -17180
rect 9200 -17200 9340 -17190
rect 8693 -17210 9093 -17204
rect 9657 -17204 9669 -17180
rect 10045 -17180 10305 -17170
rect 10045 -17204 10057 -17180
rect 9657 -17210 10057 -17204
rect 10293 -17204 10305 -17180
rect 10681 -17180 10700 -17170
rect 11257 -17170 11657 -17164
rect 10681 -17204 10693 -17180
rect 10293 -17210 10693 -17204
rect 11257 -17204 11269 -17170
rect 11645 -17204 11657 -17170
rect 11257 -17210 11657 -17204
rect 11893 -17170 12293 -17164
rect 11893 -17204 11905 -17170
rect 12281 -17204 12293 -17170
rect 11893 -17210 12293 -17204
rect 12620 -17200 12630 -17080
rect 12750 -17110 12760 -17080
rect 12750 -17164 15490 -17110
rect 12750 -17170 15493 -17164
rect 12750 -17200 12869 -17170
rect 12620 -17210 12760 -17200
rect 12857 -17204 12869 -17200
rect 13245 -17200 13505 -17170
rect 13245 -17204 13257 -17200
rect 12857 -17210 13257 -17204
rect 13493 -17204 13505 -17200
rect 13881 -17200 14469 -17170
rect 13881 -17204 13893 -17200
rect 13493 -17210 13893 -17204
rect 14457 -17204 14469 -17200
rect 14845 -17200 15105 -17170
rect 14845 -17204 14857 -17200
rect 14457 -17210 14857 -17204
rect 15093 -17204 15105 -17200
rect 15481 -17204 15493 -17170
rect 15820 -17190 15830 -17070
rect 15950 -17100 15960 -17070
rect 17420 -17070 17560 -17060
rect 15950 -17164 17090 -17100
rect 15950 -17170 17093 -17164
rect 15950 -17190 16069 -17170
rect 15820 -17200 16069 -17190
rect 15093 -17210 15493 -17204
rect 16057 -17204 16069 -17200
rect 16445 -17200 16705 -17170
rect 16445 -17204 16457 -17200
rect 16057 -17210 16457 -17204
rect 16693 -17204 16705 -17200
rect 17081 -17204 17093 -17170
rect 17420 -17190 17430 -17070
rect 17550 -17100 17560 -17070
rect 19020 -17070 19160 -17060
rect 17550 -17164 18690 -17100
rect 17550 -17170 18693 -17164
rect 17550 -17190 17669 -17170
rect 17420 -17200 17669 -17190
rect 16693 -17210 17093 -17204
rect 17657 -17204 17669 -17200
rect 18045 -17200 18305 -17170
rect 18045 -17204 18057 -17200
rect 17657 -17210 18057 -17204
rect 18293 -17204 18305 -17200
rect 18681 -17204 18693 -17170
rect 19020 -17190 19030 -17070
rect 19150 -17100 19160 -17070
rect 20620 -17070 20760 -17060
rect 19150 -17164 20290 -17100
rect 19150 -17170 20293 -17164
rect 19150 -17190 19269 -17170
rect 19020 -17200 19269 -17190
rect 18293 -17210 18693 -17204
rect 19257 -17204 19269 -17200
rect 19645 -17200 19905 -17170
rect 19645 -17204 19657 -17200
rect 19257 -17210 19657 -17204
rect 19893 -17204 19905 -17200
rect 20281 -17204 20293 -17170
rect 20620 -17190 20630 -17070
rect 20750 -17100 20760 -17070
rect 22220 -17070 22360 -17060
rect 20750 -17164 21890 -17100
rect 20750 -17170 21893 -17164
rect 20750 -17190 20869 -17170
rect 20620 -17200 20869 -17190
rect 19893 -17210 20293 -17204
rect 20857 -17204 20869 -17200
rect 21245 -17200 21505 -17170
rect 21245 -17204 21257 -17200
rect 20857 -17210 21257 -17204
rect 21493 -17204 21505 -17200
rect 21881 -17204 21893 -17170
rect 22220 -17190 22230 -17070
rect 22350 -17100 22360 -17070
rect 23820 -17070 23960 -17060
rect 22350 -17164 23490 -17100
rect 22350 -17170 23493 -17164
rect 22350 -17190 22469 -17170
rect 22220 -17200 22469 -17190
rect 21493 -17210 21893 -17204
rect 22457 -17204 22469 -17200
rect 22845 -17200 23105 -17170
rect 22845 -17204 22857 -17200
rect 22457 -17210 22857 -17204
rect 23093 -17204 23105 -17200
rect 23481 -17204 23493 -17170
rect 23820 -17190 23830 -17070
rect 23950 -17100 23960 -17070
rect 27020 -17070 27160 -17060
rect 27020 -17100 27030 -17070
rect 23950 -17164 25090 -17100
rect 25660 -17164 27030 -17100
rect 23950 -17170 25093 -17164
rect 23950 -17190 24069 -17170
rect 23820 -17200 24069 -17190
rect 23093 -17210 23493 -17204
rect 24057 -17204 24069 -17200
rect 24445 -17200 24705 -17170
rect 24445 -17204 24457 -17200
rect 24057 -17210 24457 -17204
rect 24693 -17204 24705 -17200
rect 25081 -17204 25093 -17170
rect 24693 -17210 25093 -17204
rect 25657 -17170 27030 -17164
rect 25657 -17204 25669 -17170
rect 26045 -17200 26305 -17170
rect 26045 -17204 26057 -17200
rect 25657 -17210 26057 -17204
rect 26293 -17204 26305 -17200
rect 26681 -17190 27030 -17170
rect 27150 -17100 27160 -17070
rect 28620 -17070 28760 -17060
rect 27150 -17164 28290 -17100
rect 27150 -17170 28293 -17164
rect 27150 -17190 27269 -17170
rect 26681 -17200 27269 -17190
rect 26681 -17204 26693 -17200
rect 26293 -17210 26693 -17204
rect 27257 -17204 27269 -17200
rect 27645 -17200 27905 -17170
rect 27645 -17204 27657 -17200
rect 27257 -17210 27657 -17204
rect 27893 -17204 27905 -17200
rect 28281 -17204 28293 -17170
rect 28620 -17190 28630 -17070
rect 28750 -17100 28760 -17070
rect 31840 -17080 31980 -17070
rect 28750 -17164 31490 -17100
rect 28750 -17170 31493 -17164
rect 28750 -17190 28869 -17170
rect 28620 -17200 28869 -17190
rect 27893 -17210 28293 -17204
rect 28857 -17204 28869 -17200
rect 29245 -17200 29505 -17170
rect 29245 -17204 29257 -17200
rect 28857 -17210 29257 -17204
rect 29493 -17204 29505 -17200
rect 29881 -17200 30469 -17170
rect 29881 -17204 29893 -17200
rect 29493 -17210 29893 -17204
rect 30457 -17204 30469 -17200
rect 30845 -17200 31105 -17170
rect 30845 -17204 30857 -17200
rect 30457 -17210 30857 -17204
rect 31093 -17204 31105 -17200
rect 31481 -17204 31493 -17170
rect 31093 -17210 31493 -17204
rect 31840 -17200 31850 -17080
rect 31970 -17100 31980 -17080
rect 31970 -17164 36290 -17100
rect 31970 -17170 36293 -17164
rect 31970 -17200 32069 -17170
rect 31840 -17210 31980 -17200
rect 32057 -17204 32069 -17200
rect 32445 -17200 32705 -17170
rect 32445 -17204 32457 -17200
rect 32057 -17210 32457 -17204
rect 32693 -17204 32705 -17200
rect 33081 -17200 33669 -17170
rect 33081 -17204 33093 -17200
rect 32693 -17210 33093 -17204
rect 33657 -17204 33669 -17200
rect 34045 -17200 34305 -17170
rect 34045 -17204 34057 -17200
rect 33657 -17210 34057 -17204
rect 34293 -17204 34305 -17200
rect 34681 -17200 35269 -17170
rect 34681 -17204 34693 -17200
rect 34293 -17210 34693 -17204
rect 35257 -17204 35269 -17200
rect 35645 -17200 35905 -17170
rect 35645 -17204 35657 -17200
rect 35257 -17210 35657 -17204
rect 35893 -17204 35905 -17200
rect 36281 -17204 36293 -17170
rect 35893 -17210 36293 -17204
rect 36857 -17170 37257 -17164
rect 36857 -17204 36869 -17170
rect 37245 -17204 37257 -17170
rect 36857 -17210 37257 -17204
rect 37493 -17170 37893 -17164
rect 37493 -17204 37505 -17170
rect 37881 -17204 37893 -17170
rect 37493 -17210 37893 -17204
rect 57 -17428 490 -17422
rect 57 -17462 69 -17428
rect 445 -17462 490 -17428
rect 57 -17468 490 -17462
rect 440 -17690 490 -17468
rect 57 -17696 490 -17690
rect 57 -17730 69 -17696
rect 445 -17730 490 -17696
rect 57 -17736 490 -17730
rect -30 -17796 16 -17784
rect -30 -18488 -24 -17796
rect 10 -18488 16 -17796
rect -30 -18500 16 -18488
rect 440 -18548 490 -17736
rect 670 -17422 720 -17210
rect 1134 -17257 1180 -17245
rect 1134 -17375 1140 -17257
rect 1174 -17375 1180 -17257
rect 1570 -17257 1616 -17245
rect 1570 -17260 1576 -17257
rect 1134 -17387 1180 -17375
rect 1560 -17375 1576 -17260
rect 1610 -17260 1616 -17257
rect 2098 -17257 2144 -17245
rect 2098 -17260 2104 -17257
rect 1610 -17375 2104 -17260
rect 2138 -17260 2144 -17257
rect 2206 -17257 2252 -17245
rect 2206 -17260 2212 -17257
rect 2138 -17375 2212 -17260
rect 2246 -17260 2252 -17257
rect 2734 -17257 2780 -17245
rect 2734 -17260 2740 -17257
rect 2246 -17375 2740 -17260
rect 2774 -17260 2780 -17257
rect 3170 -17257 3216 -17245
rect 3170 -17260 3176 -17257
rect 2774 -17375 3176 -17260
rect 3210 -17260 3216 -17257
rect 3698 -17257 3744 -17245
rect 3698 -17260 3704 -17257
rect 3210 -17375 3704 -17260
rect 3738 -17260 3744 -17257
rect 3806 -17257 3852 -17245
rect 3806 -17260 3812 -17257
rect 3738 -17375 3812 -17260
rect 3846 -17260 3852 -17257
rect 4334 -17257 4380 -17245
rect 4334 -17260 4340 -17257
rect 3846 -17375 4340 -17260
rect 4374 -17260 4380 -17257
rect 4770 -17257 4816 -17245
rect 4770 -17260 4776 -17257
rect 4374 -17375 4776 -17260
rect 4810 -17260 4816 -17257
rect 5298 -17257 5344 -17245
rect 5298 -17260 5304 -17257
rect 4810 -17375 5304 -17260
rect 5338 -17260 5344 -17257
rect 5406 -17257 5452 -17245
rect 5406 -17260 5412 -17257
rect 5338 -17375 5412 -17260
rect 5446 -17260 5452 -17257
rect 5934 -17257 5980 -17245
rect 5934 -17260 5940 -17257
rect 5446 -17375 5940 -17260
rect 5974 -17260 5980 -17257
rect 6370 -17257 6416 -17245
rect 6370 -17260 6376 -17257
rect 5974 -17375 6376 -17260
rect 6410 -17260 6416 -17257
rect 6898 -17257 6944 -17245
rect 6898 -17260 6904 -17257
rect 6410 -17375 6904 -17260
rect 6938 -17260 6944 -17257
rect 7006 -17257 7052 -17245
rect 7006 -17260 7012 -17257
rect 6938 -17375 7012 -17260
rect 7046 -17260 7052 -17257
rect 7534 -17257 7580 -17245
rect 7534 -17260 7540 -17257
rect 7046 -17375 7540 -17260
rect 7574 -17260 7580 -17257
rect 7970 -17257 8016 -17245
rect 7970 -17260 7976 -17257
rect 7574 -17375 7976 -17260
rect 8010 -17260 8016 -17257
rect 8498 -17257 8544 -17245
rect 8498 -17260 8504 -17257
rect 8010 -17375 8504 -17260
rect 8538 -17260 8544 -17257
rect 8606 -17257 8652 -17245
rect 8606 -17260 8612 -17257
rect 8538 -17375 8612 -17260
rect 8646 -17260 8652 -17257
rect 9134 -17257 9180 -17245
rect 9134 -17260 9140 -17257
rect 8646 -17375 9140 -17260
rect 9174 -17260 9180 -17257
rect 9570 -17257 9616 -17245
rect 9570 -17260 9576 -17257
rect 9174 -17375 9576 -17260
rect 9610 -17260 9616 -17257
rect 10098 -17257 10144 -17245
rect 10098 -17260 10104 -17257
rect 9610 -17375 10104 -17260
rect 10138 -17260 10144 -17257
rect 10206 -17257 10252 -17245
rect 10206 -17260 10212 -17257
rect 10138 -17375 10212 -17260
rect 10246 -17260 10252 -17257
rect 10734 -17250 10780 -17245
rect 10734 -17257 10940 -17250
rect 10734 -17260 10740 -17257
rect 10246 -17375 10740 -17260
rect 10774 -17260 10940 -17257
rect 11170 -17257 11216 -17245
rect 11170 -17260 11176 -17257
rect 10774 -17375 10810 -17260
rect 1560 -17380 10810 -17375
rect 10930 -17375 11176 -17260
rect 11210 -17260 11216 -17257
rect 11380 -17260 11500 -17210
rect 11698 -17257 11744 -17245
rect 11698 -17260 11704 -17257
rect 11210 -17375 11704 -17260
rect 11738 -17260 11744 -17257
rect 11806 -17257 11852 -17245
rect 11806 -17260 11812 -17257
rect 11738 -17375 11812 -17260
rect 11846 -17260 11852 -17257
rect 12040 -17260 12160 -17210
rect 12334 -17257 12380 -17245
rect 12334 -17260 12340 -17257
rect 11846 -17375 12340 -17260
rect 12374 -17260 12380 -17257
rect 12770 -17257 12816 -17245
rect 12770 -17260 12776 -17257
rect 12374 -17375 12776 -17260
rect 12810 -17260 12816 -17257
rect 13298 -17257 13344 -17245
rect 13298 -17260 13304 -17257
rect 12810 -17375 13304 -17260
rect 13338 -17260 13344 -17257
rect 13406 -17257 13452 -17245
rect 13406 -17260 13412 -17257
rect 13338 -17375 13412 -17260
rect 13446 -17260 13452 -17257
rect 13934 -17257 13980 -17245
rect 13934 -17260 13940 -17257
rect 13446 -17375 13940 -17260
rect 13974 -17260 13980 -17257
rect 14370 -17257 14416 -17245
rect 14370 -17260 14376 -17257
rect 13974 -17375 14376 -17260
rect 14410 -17260 14416 -17257
rect 14898 -17257 14944 -17245
rect 14898 -17260 14904 -17257
rect 14410 -17375 14904 -17260
rect 14938 -17260 14944 -17257
rect 15006 -17257 15052 -17245
rect 15006 -17260 15012 -17257
rect 14938 -17375 15012 -17260
rect 15046 -17260 15052 -17257
rect 15534 -17257 15580 -17245
rect 15534 -17260 15540 -17257
rect 15046 -17375 15540 -17260
rect 15574 -17260 15580 -17257
rect 15970 -17257 16016 -17245
rect 15970 -17260 15976 -17257
rect 15574 -17375 15976 -17260
rect 16010 -17260 16016 -17257
rect 16498 -17257 16544 -17245
rect 16498 -17260 16504 -17257
rect 16010 -17375 16504 -17260
rect 16538 -17260 16544 -17257
rect 16606 -17257 16652 -17245
rect 16606 -17260 16612 -17257
rect 16538 -17375 16612 -17260
rect 16646 -17260 16652 -17257
rect 17134 -17257 17180 -17245
rect 17134 -17260 17140 -17257
rect 16646 -17375 17140 -17260
rect 17174 -17260 17180 -17257
rect 17570 -17257 17616 -17245
rect 17570 -17260 17576 -17257
rect 17174 -17375 17576 -17260
rect 17610 -17260 17616 -17257
rect 18098 -17257 18144 -17245
rect 18098 -17260 18104 -17257
rect 17610 -17375 18104 -17260
rect 18138 -17260 18144 -17257
rect 18206 -17257 18252 -17245
rect 18206 -17260 18212 -17257
rect 18138 -17375 18212 -17260
rect 18246 -17260 18252 -17257
rect 18734 -17257 18780 -17245
rect 18734 -17260 18740 -17257
rect 18246 -17375 18740 -17260
rect 18774 -17260 18780 -17257
rect 19170 -17257 19216 -17245
rect 19170 -17260 19176 -17257
rect 18774 -17375 19176 -17260
rect 19210 -17260 19216 -17257
rect 19698 -17257 19744 -17245
rect 19698 -17260 19704 -17257
rect 19210 -17375 19704 -17260
rect 19738 -17260 19744 -17257
rect 19806 -17257 19852 -17245
rect 19806 -17260 19812 -17257
rect 19738 -17375 19812 -17260
rect 19846 -17260 19852 -17257
rect 20334 -17257 20380 -17245
rect 20334 -17260 20340 -17257
rect 19846 -17375 20340 -17260
rect 20374 -17260 20380 -17257
rect 20770 -17257 20816 -17245
rect 20770 -17260 20776 -17257
rect 20374 -17375 20776 -17260
rect 20810 -17260 20816 -17257
rect 21298 -17257 21344 -17245
rect 21298 -17260 21304 -17257
rect 20810 -17375 21304 -17260
rect 21338 -17260 21344 -17257
rect 21406 -17257 21452 -17245
rect 21406 -17260 21412 -17257
rect 21338 -17375 21412 -17260
rect 21446 -17260 21452 -17257
rect 21934 -17257 21980 -17245
rect 21934 -17260 21940 -17257
rect 21446 -17375 21940 -17260
rect 21974 -17260 21980 -17257
rect 22370 -17257 22416 -17245
rect 22370 -17260 22376 -17257
rect 21974 -17375 22376 -17260
rect 22410 -17260 22416 -17257
rect 22898 -17257 22944 -17245
rect 22898 -17260 22904 -17257
rect 22410 -17375 22904 -17260
rect 22938 -17260 22944 -17257
rect 23006 -17257 23052 -17245
rect 23006 -17260 23012 -17257
rect 22938 -17375 23012 -17260
rect 23046 -17260 23052 -17257
rect 23534 -17257 23580 -17245
rect 23534 -17260 23540 -17257
rect 23046 -17375 23540 -17260
rect 23574 -17260 23580 -17257
rect 23970 -17257 24016 -17245
rect 23970 -17260 23976 -17257
rect 23574 -17375 23976 -17260
rect 24010 -17260 24016 -17257
rect 24498 -17257 24544 -17245
rect 24498 -17260 24504 -17257
rect 24010 -17375 24504 -17260
rect 24538 -17260 24544 -17257
rect 24606 -17257 24652 -17245
rect 24606 -17260 24612 -17257
rect 24538 -17375 24612 -17260
rect 24646 -17260 24652 -17257
rect 25134 -17257 25180 -17245
rect 25134 -17260 25140 -17257
rect 24646 -17375 25140 -17260
rect 25174 -17260 25180 -17257
rect 25570 -17257 25616 -17245
rect 25570 -17260 25576 -17257
rect 25174 -17375 25576 -17260
rect 25610 -17260 25616 -17257
rect 26098 -17257 26144 -17245
rect 26098 -17260 26104 -17257
rect 25610 -17375 26104 -17260
rect 26138 -17260 26144 -17257
rect 26206 -17257 26252 -17245
rect 26206 -17260 26212 -17257
rect 26138 -17375 26212 -17260
rect 26246 -17260 26252 -17257
rect 26734 -17257 26780 -17245
rect 26734 -17260 26740 -17257
rect 26246 -17375 26740 -17260
rect 26774 -17260 26780 -17257
rect 27170 -17257 27216 -17245
rect 27170 -17260 27176 -17257
rect 26774 -17375 27176 -17260
rect 27210 -17260 27216 -17257
rect 27698 -17257 27744 -17245
rect 27698 -17260 27704 -17257
rect 27210 -17375 27704 -17260
rect 27738 -17260 27744 -17257
rect 27806 -17257 27852 -17245
rect 27806 -17260 27812 -17257
rect 27738 -17375 27812 -17260
rect 27846 -17260 27852 -17257
rect 28334 -17257 28380 -17245
rect 28334 -17260 28340 -17257
rect 27846 -17375 28340 -17260
rect 28374 -17260 28380 -17257
rect 28770 -17257 28816 -17245
rect 28770 -17260 28776 -17257
rect 28374 -17375 28776 -17260
rect 28810 -17260 28816 -17257
rect 29298 -17257 29344 -17245
rect 29298 -17260 29304 -17257
rect 28810 -17375 29304 -17260
rect 29338 -17260 29344 -17257
rect 29406 -17257 29452 -17245
rect 29406 -17260 29412 -17257
rect 29338 -17375 29412 -17260
rect 29446 -17260 29452 -17257
rect 29934 -17257 29980 -17245
rect 29934 -17260 29940 -17257
rect 29446 -17375 29940 -17260
rect 29974 -17260 29980 -17257
rect 30370 -17257 30416 -17245
rect 30370 -17260 30376 -17257
rect 29974 -17375 30376 -17260
rect 30410 -17260 30416 -17257
rect 30898 -17257 30944 -17245
rect 30898 -17260 30904 -17257
rect 30410 -17375 30904 -17260
rect 30938 -17260 30944 -17257
rect 31006 -17257 31052 -17245
rect 31006 -17260 31012 -17257
rect 30938 -17375 31012 -17260
rect 31046 -17260 31052 -17257
rect 31534 -17257 31580 -17245
rect 31534 -17260 31540 -17257
rect 31046 -17375 31540 -17260
rect 31574 -17260 31580 -17257
rect 31970 -17257 32016 -17245
rect 31970 -17260 31976 -17257
rect 31574 -17375 31976 -17260
rect 32010 -17260 32016 -17257
rect 32498 -17257 32544 -17245
rect 32498 -17260 32504 -17257
rect 32010 -17375 32504 -17260
rect 32538 -17260 32544 -17257
rect 32606 -17257 32652 -17245
rect 32606 -17260 32612 -17257
rect 32538 -17375 32612 -17260
rect 32646 -17260 32652 -17257
rect 33134 -17257 33180 -17245
rect 33134 -17260 33140 -17257
rect 32646 -17375 33140 -17260
rect 33174 -17260 33180 -17257
rect 33570 -17257 33616 -17245
rect 33570 -17260 33576 -17257
rect 33174 -17375 33576 -17260
rect 33610 -17260 33616 -17257
rect 34098 -17257 34144 -17245
rect 34098 -17260 34104 -17257
rect 33610 -17375 34104 -17260
rect 34138 -17260 34144 -17257
rect 34206 -17257 34252 -17245
rect 34206 -17260 34212 -17257
rect 34138 -17375 34212 -17260
rect 34246 -17260 34252 -17257
rect 34734 -17257 34780 -17245
rect 34734 -17260 34740 -17257
rect 34246 -17375 34740 -17260
rect 34774 -17260 34780 -17257
rect 35170 -17257 35216 -17245
rect 35170 -17260 35176 -17257
rect 34774 -17375 35176 -17260
rect 35210 -17260 35216 -17257
rect 35698 -17257 35744 -17245
rect 35698 -17260 35704 -17257
rect 35210 -17375 35704 -17260
rect 35738 -17260 35744 -17257
rect 35806 -17257 35852 -17245
rect 35806 -17260 35812 -17257
rect 35738 -17375 35812 -17260
rect 35846 -17260 35852 -17257
rect 36334 -17257 36380 -17245
rect 36334 -17260 36340 -17257
rect 35846 -17375 36340 -17260
rect 36374 -17375 36380 -17257
rect 10930 -17380 36380 -17375
rect 1570 -17387 1616 -17380
rect 2098 -17387 2144 -17380
rect 2206 -17387 2252 -17380
rect 2734 -17387 2780 -17380
rect 3170 -17387 3216 -17380
rect 3698 -17387 3744 -17380
rect 3806 -17387 3852 -17380
rect 4334 -17387 4380 -17380
rect 4770 -17387 4816 -17380
rect 5298 -17387 5344 -17380
rect 5406 -17387 5452 -17380
rect 5934 -17387 5980 -17380
rect 6370 -17387 6416 -17380
rect 6898 -17387 6944 -17380
rect 7006 -17387 7052 -17380
rect 7534 -17387 7580 -17380
rect 7970 -17387 8016 -17380
rect 8498 -17387 8544 -17380
rect 8606 -17387 8652 -17380
rect 9134 -17387 9180 -17380
rect 9570 -17387 9616 -17380
rect 10098 -17387 10144 -17380
rect 10206 -17387 10252 -17380
rect 10734 -17387 10940 -17380
rect 11170 -17387 11216 -17380
rect 10750 -17390 10940 -17387
rect 11380 -17422 11500 -17380
rect 11698 -17387 11744 -17380
rect 11806 -17387 11852 -17380
rect 12040 -17422 12160 -17380
rect 12334 -17387 12380 -17380
rect 12770 -17387 12816 -17380
rect 13298 -17387 13344 -17380
rect 13406 -17387 13452 -17380
rect 13934 -17387 13980 -17380
rect 14370 -17387 14416 -17380
rect 14898 -17387 14944 -17380
rect 15006 -17387 15052 -17380
rect 15534 -17387 15580 -17380
rect 15970 -17387 16016 -17380
rect 16498 -17387 16544 -17380
rect 16606 -17387 16652 -17380
rect 17134 -17387 17180 -17380
rect 17570 -17387 17616 -17380
rect 18098 -17387 18144 -17380
rect 18206 -17387 18252 -17380
rect 18734 -17387 18780 -17380
rect 19170 -17387 19216 -17380
rect 19698 -17387 19744 -17380
rect 19806 -17387 19852 -17380
rect 20334 -17387 20380 -17380
rect 20770 -17387 20816 -17380
rect 21298 -17387 21344 -17380
rect 21406 -17387 21452 -17380
rect 21934 -17387 21980 -17380
rect 22370 -17387 22416 -17380
rect 22898 -17387 22944 -17380
rect 23006 -17387 23052 -17380
rect 23534 -17387 23580 -17380
rect 23970 -17387 24016 -17380
rect 24498 -17387 24544 -17380
rect 24606 -17387 24652 -17380
rect 25134 -17387 25180 -17380
rect 25570 -17387 25616 -17380
rect 26098 -17387 26144 -17380
rect 26206 -17387 26252 -17380
rect 26734 -17387 26780 -17380
rect 27170 -17387 27216 -17380
rect 27698 -17387 27744 -17380
rect 27806 -17387 27852 -17380
rect 28334 -17387 28380 -17380
rect 28770 -17387 28816 -17380
rect 29298 -17387 29344 -17380
rect 29406 -17387 29452 -17380
rect 29934 -17387 29980 -17380
rect 30370 -17387 30416 -17380
rect 30898 -17387 30944 -17380
rect 31006 -17387 31052 -17380
rect 31534 -17387 31580 -17380
rect 31970 -17387 32016 -17380
rect 32498 -17387 32544 -17380
rect 32606 -17387 32652 -17380
rect 33134 -17387 33180 -17380
rect 33570 -17387 33616 -17380
rect 34098 -17387 34144 -17380
rect 34206 -17387 34252 -17380
rect 34734 -17387 34780 -17380
rect 35170 -17387 35216 -17380
rect 35698 -17387 35744 -17380
rect 35806 -17387 35852 -17380
rect 36334 -17387 36380 -17380
rect 36770 -17257 36816 -17245
rect 36770 -17375 36776 -17257
rect 36810 -17375 36816 -17257
rect 36770 -17387 36816 -17375
rect 37298 -17257 37344 -17245
rect 37298 -17375 37304 -17257
rect 37338 -17375 37344 -17257
rect 37298 -17387 37344 -17375
rect 37406 -17257 37452 -17245
rect 37406 -17375 37412 -17257
rect 37446 -17375 37452 -17257
rect 37406 -17387 37452 -17375
rect 37934 -17257 37980 -17245
rect 37934 -17375 37940 -17257
rect 37974 -17375 37980 -17257
rect 37934 -17387 37980 -17375
rect 670 -17428 1093 -17422
rect 670 -17462 705 -17428
rect 1081 -17462 1093 -17428
rect 670 -17468 1093 -17462
rect 1657 -17428 2057 -17422
rect 1657 -17462 1669 -17428
rect 2045 -17430 2057 -17428
rect 2293 -17428 2693 -17422
rect 2293 -17430 2305 -17428
rect 2045 -17462 2060 -17430
rect 1657 -17468 2060 -17462
rect 670 -17690 720 -17468
rect 1420 -17510 1560 -17500
rect 1420 -17630 1430 -17510
rect 1550 -17520 1560 -17510
rect 1660 -17520 2060 -17468
rect 2290 -17462 2305 -17430
rect 2681 -17462 2693 -17428
rect 2290 -17468 2693 -17462
rect 3257 -17428 3657 -17422
rect 3257 -17462 3269 -17428
rect 3645 -17430 3657 -17428
rect 3893 -17428 4293 -17422
rect 3893 -17430 3905 -17428
rect 3645 -17462 3660 -17430
rect 3257 -17468 3660 -17462
rect 2290 -17520 2690 -17468
rect 3020 -17510 3160 -17500
rect 3020 -17520 3030 -17510
rect 1550 -17620 3030 -17520
rect 1550 -17630 1560 -17620
rect 1420 -17640 1560 -17630
rect 1660 -17640 2690 -17620
rect 3020 -17630 3030 -17620
rect 3150 -17520 3160 -17510
rect 3260 -17520 3660 -17468
rect 3890 -17462 3905 -17430
rect 4281 -17462 4293 -17428
rect 3890 -17468 4293 -17462
rect 4857 -17428 5257 -17422
rect 4857 -17462 4869 -17428
rect 5245 -17430 5257 -17428
rect 5493 -17428 5893 -17422
rect 5493 -17430 5505 -17428
rect 5245 -17462 5260 -17430
rect 4857 -17468 5260 -17462
rect 3890 -17520 4290 -17468
rect 4620 -17510 4760 -17500
rect 4620 -17520 4630 -17510
rect 3150 -17620 4630 -17520
rect 3150 -17630 3160 -17620
rect 3020 -17640 3160 -17630
rect 3260 -17640 4290 -17620
rect 4620 -17630 4630 -17620
rect 4750 -17520 4760 -17510
rect 4860 -17520 5260 -17468
rect 5490 -17462 5505 -17430
rect 5881 -17462 5893 -17428
rect 5490 -17468 5893 -17462
rect 6457 -17428 6857 -17422
rect 6457 -17462 6469 -17428
rect 6845 -17430 6857 -17428
rect 7093 -17428 7493 -17422
rect 7093 -17430 7105 -17428
rect 6845 -17462 6860 -17430
rect 6457 -17468 6860 -17462
rect 5490 -17520 5890 -17468
rect 6220 -17510 6360 -17500
rect 6220 -17520 6230 -17510
rect 4750 -17620 6230 -17520
rect 4750 -17630 4760 -17620
rect 4620 -17640 4760 -17630
rect 4860 -17640 5890 -17620
rect 6220 -17630 6230 -17620
rect 6350 -17520 6360 -17510
rect 6460 -17520 6860 -17468
rect 7090 -17462 7105 -17430
rect 7481 -17462 7493 -17428
rect 7090 -17468 7493 -17462
rect 8057 -17428 8457 -17422
rect 8057 -17462 8069 -17428
rect 8445 -17430 8457 -17428
rect 8693 -17428 9093 -17422
rect 8693 -17430 8705 -17428
rect 8445 -17462 8460 -17430
rect 8057 -17468 8460 -17462
rect 7090 -17520 7490 -17468
rect 7820 -17510 7960 -17500
rect 7820 -17520 7830 -17510
rect 6350 -17620 7830 -17520
rect 6350 -17630 6360 -17620
rect 6220 -17640 6360 -17630
rect 6460 -17640 7490 -17620
rect 7820 -17630 7830 -17620
rect 7950 -17520 7960 -17510
rect 8060 -17520 8460 -17468
rect 8690 -17462 8705 -17430
rect 9081 -17462 9093 -17428
rect 8690 -17468 9093 -17462
rect 9657 -17428 10057 -17422
rect 9657 -17462 9669 -17428
rect 10045 -17430 10057 -17428
rect 10293 -17428 10693 -17422
rect 10293 -17430 10305 -17428
rect 10045 -17462 10060 -17430
rect 9657 -17468 10060 -17462
rect 8690 -17520 9090 -17468
rect 9420 -17510 9560 -17500
rect 9420 -17520 9430 -17510
rect 7950 -17620 9430 -17520
rect 7950 -17630 7960 -17620
rect 7820 -17640 7960 -17630
rect 8060 -17640 9090 -17620
rect 9420 -17630 9430 -17620
rect 9550 -17520 9560 -17510
rect 9660 -17520 10060 -17468
rect 10290 -17462 10305 -17430
rect 10681 -17462 10693 -17428
rect 10290 -17468 10693 -17462
rect 11257 -17428 11657 -17422
rect 11257 -17462 11269 -17428
rect 11645 -17462 11657 -17428
rect 11257 -17468 11657 -17462
rect 11893 -17428 12293 -17422
rect 11893 -17462 11905 -17428
rect 12281 -17462 12293 -17428
rect 11893 -17468 12293 -17462
rect 12857 -17428 13257 -17422
rect 12857 -17462 12869 -17428
rect 13245 -17430 13257 -17428
rect 13493 -17428 13893 -17422
rect 13493 -17430 13505 -17428
rect 13245 -17462 13260 -17430
rect 12857 -17468 13260 -17462
rect 10290 -17520 10690 -17468
rect 9550 -17620 10690 -17520
rect 9550 -17630 9560 -17620
rect 9420 -17640 9560 -17630
rect 9660 -17640 10690 -17620
rect 1660 -17690 2060 -17640
rect 670 -17696 1093 -17690
rect 670 -17730 705 -17696
rect 1081 -17730 1093 -17696
rect 670 -17736 1093 -17730
rect 1657 -17696 2060 -17690
rect 1657 -17730 1669 -17696
rect 2045 -17730 2060 -17696
rect 2290 -17690 2690 -17640
rect 3260 -17690 3660 -17640
rect 2290 -17696 2693 -17690
rect 2290 -17730 2305 -17696
rect 2681 -17730 2693 -17696
rect 1657 -17736 2057 -17730
rect 2293 -17736 2693 -17730
rect 3257 -17696 3660 -17690
rect 3257 -17730 3269 -17696
rect 3645 -17730 3660 -17696
rect 3890 -17690 4290 -17640
rect 4860 -17690 5260 -17640
rect 3890 -17696 4293 -17690
rect 3890 -17730 3905 -17696
rect 4281 -17730 4293 -17696
rect 3257 -17736 3657 -17730
rect 3893 -17736 4293 -17730
rect 4857 -17696 5260 -17690
rect 4857 -17730 4869 -17696
rect 5245 -17730 5260 -17696
rect 5490 -17690 5890 -17640
rect 6460 -17690 6860 -17640
rect 5490 -17696 5893 -17690
rect 5490 -17730 5505 -17696
rect 5881 -17730 5893 -17696
rect 4857 -17736 5257 -17730
rect 5493 -17736 5893 -17730
rect 6457 -17696 6860 -17690
rect 6457 -17730 6469 -17696
rect 6845 -17730 6860 -17696
rect 7090 -17690 7490 -17640
rect 8060 -17690 8460 -17640
rect 7090 -17696 7493 -17690
rect 7090 -17730 7105 -17696
rect 7481 -17730 7493 -17696
rect 6457 -17736 6857 -17730
rect 7093 -17736 7493 -17730
rect 8057 -17696 8460 -17690
rect 8057 -17730 8069 -17696
rect 8445 -17730 8460 -17696
rect 8690 -17690 9090 -17640
rect 9660 -17690 10060 -17640
rect 8690 -17696 9093 -17690
rect 8690 -17730 8705 -17696
rect 9081 -17730 9093 -17696
rect 8057 -17736 8457 -17730
rect 8693 -17736 9093 -17730
rect 9657 -17696 10060 -17690
rect 9657 -17730 9669 -17696
rect 10045 -17730 10060 -17696
rect 10290 -17690 10690 -17640
rect 12860 -17520 13260 -17468
rect 13490 -17462 13505 -17430
rect 13881 -17462 13893 -17428
rect 13490 -17468 13893 -17462
rect 14457 -17428 14857 -17422
rect 14457 -17462 14469 -17428
rect 14845 -17430 14857 -17428
rect 15093 -17428 15493 -17422
rect 15093 -17430 15105 -17428
rect 14845 -17462 14860 -17430
rect 14457 -17468 14860 -17462
rect 13490 -17520 13890 -17468
rect 14460 -17520 14860 -17468
rect 15090 -17462 15105 -17430
rect 15481 -17462 15493 -17428
rect 15090 -17468 15493 -17462
rect 16057 -17428 16457 -17422
rect 16057 -17462 16069 -17428
rect 16445 -17462 16457 -17428
rect 16057 -17468 16457 -17462
rect 16693 -17428 17093 -17422
rect 16693 -17462 16705 -17428
rect 17081 -17462 17093 -17428
rect 16693 -17468 17093 -17462
rect 17657 -17428 18057 -17422
rect 17657 -17462 17669 -17428
rect 18045 -17462 18057 -17428
rect 17657 -17468 18057 -17462
rect 18293 -17428 18693 -17422
rect 18293 -17462 18305 -17428
rect 18681 -17462 18693 -17428
rect 18293 -17468 18693 -17462
rect 19257 -17428 19657 -17422
rect 19257 -17462 19269 -17428
rect 19645 -17462 19657 -17428
rect 19257 -17468 19657 -17462
rect 19893 -17428 20293 -17422
rect 19893 -17462 19905 -17428
rect 20281 -17462 20293 -17428
rect 19893 -17468 20293 -17462
rect 20857 -17428 21257 -17422
rect 20857 -17462 20869 -17428
rect 21245 -17462 21257 -17428
rect 20857 -17468 21257 -17462
rect 21493 -17428 21893 -17422
rect 21493 -17462 21505 -17428
rect 21881 -17462 21893 -17428
rect 21493 -17468 21893 -17462
rect 22457 -17428 22857 -17422
rect 22457 -17462 22469 -17428
rect 22845 -17462 22857 -17428
rect 22457 -17468 22857 -17462
rect 23093 -17428 23493 -17422
rect 23093 -17462 23105 -17428
rect 23481 -17462 23493 -17428
rect 23093 -17468 23493 -17462
rect 24057 -17428 24457 -17422
rect 24057 -17462 24069 -17428
rect 24445 -17462 24457 -17428
rect 24057 -17468 24457 -17462
rect 24693 -17428 25093 -17422
rect 24693 -17462 24705 -17428
rect 25081 -17462 25093 -17428
rect 24693 -17468 25093 -17462
rect 25657 -17428 26057 -17422
rect 25657 -17462 25669 -17428
rect 26045 -17462 26057 -17428
rect 25657 -17468 26057 -17462
rect 26293 -17428 26693 -17422
rect 26293 -17462 26305 -17428
rect 26681 -17462 26693 -17428
rect 26293 -17468 26693 -17462
rect 27257 -17428 27657 -17422
rect 27257 -17462 27269 -17428
rect 27645 -17462 27657 -17428
rect 27257 -17468 27657 -17462
rect 27893 -17428 28293 -17422
rect 27893 -17462 27905 -17428
rect 28281 -17462 28293 -17428
rect 27893 -17468 28293 -17462
rect 28857 -17428 29257 -17422
rect 28857 -17462 28869 -17428
rect 29245 -17462 29257 -17428
rect 28857 -17468 29257 -17462
rect 29493 -17428 29893 -17422
rect 29493 -17462 29505 -17428
rect 29881 -17462 29893 -17428
rect 29493 -17468 29893 -17462
rect 30457 -17428 30857 -17422
rect 30457 -17462 30469 -17428
rect 30845 -17462 30857 -17428
rect 30457 -17468 30857 -17462
rect 31093 -17428 31493 -17422
rect 31093 -17462 31105 -17428
rect 31481 -17462 31493 -17428
rect 31093 -17468 31493 -17462
rect 32057 -17428 32457 -17422
rect 32057 -17462 32069 -17428
rect 32445 -17462 32457 -17428
rect 32057 -17468 32457 -17462
rect 32693 -17428 33093 -17422
rect 32693 -17462 32705 -17428
rect 33081 -17462 33093 -17428
rect 32693 -17468 33093 -17462
rect 33657 -17428 34057 -17422
rect 33657 -17462 33669 -17428
rect 34045 -17462 34057 -17428
rect 33657 -17468 34057 -17462
rect 34293 -17428 34693 -17422
rect 34293 -17462 34305 -17428
rect 34681 -17462 34693 -17428
rect 34293 -17468 34693 -17462
rect 35257 -17428 35657 -17422
rect 35257 -17462 35269 -17428
rect 35645 -17462 35657 -17428
rect 35257 -17468 35657 -17462
rect 35893 -17428 36293 -17422
rect 35893 -17462 35905 -17428
rect 36281 -17462 36293 -17428
rect 35893 -17468 36293 -17462
rect 36857 -17428 37257 -17422
rect 36857 -17462 36869 -17428
rect 37245 -17462 37257 -17428
rect 36857 -17468 37257 -17462
rect 37493 -17428 37893 -17422
rect 37493 -17462 37505 -17428
rect 37881 -17462 37893 -17428
rect 37493 -17468 37893 -17462
rect 15090 -17520 15490 -17468
rect 12860 -17640 15490 -17520
rect 12860 -17690 13260 -17640
rect 10290 -17696 10693 -17690
rect 10290 -17730 10305 -17696
rect 10681 -17730 10693 -17696
rect 9657 -17736 10057 -17730
rect 10293 -17736 10693 -17730
rect 11257 -17696 11657 -17690
rect 11257 -17730 11269 -17696
rect 11645 -17730 11657 -17696
rect 11257 -17736 11657 -17730
rect 11893 -17696 12293 -17690
rect 11893 -17730 11905 -17696
rect 12281 -17730 12293 -17696
rect 11893 -17736 12293 -17730
rect 12857 -17696 13260 -17690
rect 12857 -17730 12869 -17696
rect 13245 -17730 13260 -17696
rect 13490 -17690 13890 -17640
rect 14460 -17690 14860 -17640
rect 13490 -17696 13893 -17690
rect 13490 -17730 13505 -17696
rect 13881 -17730 13893 -17696
rect 12857 -17736 13257 -17730
rect 13493 -17736 13893 -17730
rect 14457 -17696 14860 -17690
rect 14457 -17730 14469 -17696
rect 14845 -17730 14860 -17696
rect 15090 -17690 15490 -17640
rect 15600 -17520 15740 -17510
rect 15600 -17640 15610 -17520
rect 15730 -17530 15740 -17520
rect 16060 -17530 16450 -17468
rect 16700 -17530 17090 -17468
rect 15730 -17630 17090 -17530
rect 15730 -17640 15740 -17630
rect 15600 -17650 15740 -17640
rect 16060 -17690 16450 -17630
rect 16700 -17690 17090 -17630
rect 17200 -17520 17340 -17510
rect 17200 -17640 17210 -17520
rect 17330 -17530 17340 -17520
rect 17660 -17530 18050 -17468
rect 18300 -17530 18690 -17468
rect 17330 -17630 18690 -17530
rect 17330 -17640 17340 -17630
rect 17200 -17650 17340 -17640
rect 17660 -17690 18050 -17630
rect 18300 -17690 18690 -17630
rect 18800 -17520 18940 -17510
rect 18800 -17640 18810 -17520
rect 18930 -17530 18940 -17520
rect 19260 -17530 19650 -17468
rect 19900 -17530 20290 -17468
rect 18930 -17630 20290 -17530
rect 18930 -17640 18940 -17630
rect 18800 -17650 18940 -17640
rect 19260 -17690 19650 -17630
rect 19900 -17690 20290 -17630
rect 20400 -17520 20540 -17510
rect 20400 -17640 20410 -17520
rect 20530 -17530 20540 -17520
rect 20860 -17530 21250 -17468
rect 21500 -17530 21890 -17468
rect 20530 -17630 21890 -17530
rect 20530 -17640 20540 -17630
rect 20400 -17650 20540 -17640
rect 20860 -17690 21250 -17630
rect 21500 -17690 21890 -17630
rect 22000 -17520 22140 -17510
rect 22000 -17640 22010 -17520
rect 22130 -17530 22140 -17520
rect 22460 -17530 22850 -17468
rect 23100 -17530 23490 -17468
rect 22130 -17630 23490 -17530
rect 22130 -17640 22140 -17630
rect 22000 -17650 22140 -17640
rect 22460 -17690 22850 -17630
rect 23100 -17690 23490 -17630
rect 23600 -17520 23740 -17510
rect 23600 -17640 23610 -17520
rect 23730 -17530 23740 -17520
rect 24060 -17530 24450 -17468
rect 24700 -17530 25090 -17468
rect 23730 -17630 25090 -17530
rect 23730 -17640 23740 -17630
rect 23600 -17650 23740 -17640
rect 24060 -17690 24450 -17630
rect 24700 -17690 25090 -17630
rect 25660 -17530 26050 -17468
rect 26300 -17530 26690 -17468
rect 26800 -17520 26940 -17510
rect 26800 -17530 26810 -17520
rect 25660 -17630 26810 -17530
rect 25660 -17690 26050 -17630
rect 26300 -17690 26690 -17630
rect 26800 -17640 26810 -17630
rect 26930 -17530 26940 -17520
rect 27260 -17530 27650 -17468
rect 27900 -17530 28290 -17468
rect 26930 -17630 28290 -17530
rect 26930 -17640 26940 -17630
rect 26800 -17650 26940 -17640
rect 27260 -17690 27650 -17630
rect 27900 -17690 28290 -17630
rect 28400 -17520 28540 -17510
rect 28400 -17640 28410 -17520
rect 28530 -17530 28540 -17520
rect 28860 -17530 29250 -17468
rect 29500 -17530 29890 -17468
rect 30460 -17530 30850 -17468
rect 31100 -17530 31490 -17468
rect 28530 -17630 31490 -17530
rect 28530 -17640 28540 -17630
rect 28400 -17650 28540 -17640
rect 28860 -17690 29250 -17630
rect 29500 -17690 29890 -17630
rect 30460 -17690 30850 -17630
rect 31100 -17690 31490 -17630
rect 31580 -17520 31720 -17510
rect 31580 -17640 31590 -17520
rect 31710 -17540 31720 -17520
rect 32060 -17530 32450 -17468
rect 32700 -17530 33090 -17468
rect 33660 -17530 34050 -17468
rect 34300 -17530 34690 -17468
rect 35260 -17530 35650 -17468
rect 35900 -17530 36290 -17468
rect 32060 -17540 36290 -17530
rect 31710 -17630 36290 -17540
rect 31710 -17640 31720 -17630
rect 31580 -17650 31720 -17640
rect 32060 -17690 32450 -17630
rect 32700 -17690 33090 -17630
rect 33660 -17690 34050 -17630
rect 34300 -17690 34690 -17630
rect 35260 -17690 35650 -17630
rect 35900 -17690 36290 -17630
rect 15090 -17696 15493 -17690
rect 15090 -17730 15105 -17696
rect 15481 -17730 15493 -17696
rect 14457 -17736 14857 -17730
rect 15093 -17736 15493 -17730
rect 16057 -17696 16457 -17690
rect 16057 -17730 16069 -17696
rect 16445 -17730 16457 -17696
rect 16057 -17736 16457 -17730
rect 16693 -17696 17093 -17690
rect 16693 -17730 16705 -17696
rect 17081 -17730 17093 -17696
rect 16693 -17736 17093 -17730
rect 17657 -17696 18057 -17690
rect 17657 -17730 17669 -17696
rect 18045 -17730 18057 -17696
rect 17657 -17736 18057 -17730
rect 18293 -17696 18693 -17690
rect 18293 -17730 18305 -17696
rect 18681 -17730 18693 -17696
rect 18293 -17736 18693 -17730
rect 19257 -17696 19657 -17690
rect 19257 -17730 19269 -17696
rect 19645 -17730 19657 -17696
rect 19257 -17736 19657 -17730
rect 19893 -17696 20293 -17690
rect 19893 -17730 19905 -17696
rect 20281 -17730 20293 -17696
rect 19893 -17736 20293 -17730
rect 20857 -17696 21257 -17690
rect 20857 -17730 20869 -17696
rect 21245 -17730 21257 -17696
rect 20857 -17736 21257 -17730
rect 21493 -17696 21893 -17690
rect 21493 -17730 21505 -17696
rect 21881 -17730 21893 -17696
rect 21493 -17736 21893 -17730
rect 22457 -17696 22857 -17690
rect 22457 -17730 22469 -17696
rect 22845 -17730 22857 -17696
rect 22457 -17736 22857 -17730
rect 23093 -17696 23493 -17690
rect 23093 -17730 23105 -17696
rect 23481 -17730 23493 -17696
rect 23093 -17736 23493 -17730
rect 24057 -17696 24457 -17690
rect 24057 -17730 24069 -17696
rect 24445 -17730 24457 -17696
rect 24057 -17736 24457 -17730
rect 24693 -17696 25093 -17690
rect 24693 -17730 24705 -17696
rect 25081 -17730 25093 -17696
rect 24693 -17736 25093 -17730
rect 25657 -17696 26057 -17690
rect 25657 -17730 25669 -17696
rect 26045 -17730 26057 -17696
rect 25657 -17736 26057 -17730
rect 26293 -17696 26693 -17690
rect 26293 -17730 26305 -17696
rect 26681 -17730 26693 -17696
rect 26293 -17736 26693 -17730
rect 27257 -17696 27657 -17690
rect 27257 -17730 27269 -17696
rect 27645 -17730 27657 -17696
rect 27257 -17736 27657 -17730
rect 27893 -17696 28293 -17690
rect 27893 -17730 27905 -17696
rect 28281 -17730 28293 -17696
rect 27893 -17736 28293 -17730
rect 28857 -17696 29257 -17690
rect 28857 -17730 28869 -17696
rect 29245 -17730 29257 -17696
rect 28857 -17736 29257 -17730
rect 29493 -17696 29893 -17690
rect 29493 -17730 29505 -17696
rect 29881 -17730 29893 -17696
rect 29493 -17736 29893 -17730
rect 30457 -17696 30857 -17690
rect 30457 -17730 30469 -17696
rect 30845 -17730 30857 -17696
rect 30457 -17736 30857 -17730
rect 31093 -17696 31493 -17690
rect 31093 -17730 31105 -17696
rect 31481 -17730 31493 -17696
rect 31093 -17736 31493 -17730
rect 32057 -17696 32457 -17690
rect 32057 -17730 32069 -17696
rect 32445 -17730 32457 -17696
rect 32057 -17736 32457 -17730
rect 32693 -17696 33093 -17690
rect 32693 -17730 32705 -17696
rect 33081 -17730 33093 -17696
rect 32693 -17736 33093 -17730
rect 33657 -17696 34057 -17690
rect 33657 -17730 33669 -17696
rect 34045 -17730 34057 -17696
rect 33657 -17736 34057 -17730
rect 34293 -17696 34693 -17690
rect 34293 -17730 34305 -17696
rect 34681 -17730 34693 -17696
rect 34293 -17736 34693 -17730
rect 35257 -17696 35657 -17690
rect 35257 -17730 35269 -17696
rect 35645 -17730 35657 -17696
rect 35257 -17736 35657 -17730
rect 35893 -17696 36293 -17690
rect 35893 -17730 35905 -17696
rect 36281 -17730 36293 -17696
rect 35893 -17736 36293 -17730
rect 36857 -17696 37257 -17690
rect 36857 -17730 36869 -17696
rect 37245 -17730 37257 -17696
rect 36857 -17736 37257 -17730
rect 37493 -17696 37893 -17690
rect 37493 -17730 37505 -17696
rect 37881 -17730 37893 -17696
rect 37493 -17736 37893 -17730
rect 57 -18554 490 -18548
rect 57 -18560 69 -18554
rect 0 -18588 69 -18560
rect 445 -18588 490 -18554
rect 0 -18688 490 -18588
rect 670 -18548 720 -17736
rect 1134 -17796 1180 -17784
rect 1134 -18488 1140 -17796
rect 1174 -18488 1180 -17796
rect 1134 -18500 1180 -18488
rect 1570 -17796 1616 -17784
rect 1570 -18488 1576 -17796
rect 1610 -18488 1616 -17796
rect 1570 -18500 1616 -18488
rect 2098 -17796 2144 -17784
rect 2098 -18488 2104 -17796
rect 2138 -17800 2144 -17796
rect 2206 -17796 2252 -17784
rect 2206 -17800 2212 -17796
rect 2138 -17810 2212 -17800
rect 2138 -18480 2212 -18470
rect 2138 -18488 2144 -18480
rect 2098 -18500 2144 -18488
rect 2206 -18488 2212 -18480
rect 2246 -18488 2252 -17796
rect 2206 -18500 2252 -18488
rect 2734 -17796 2780 -17784
rect 2734 -18488 2740 -17796
rect 2774 -18488 2780 -17796
rect 2734 -18500 2780 -18488
rect 3170 -17796 3216 -17784
rect 3170 -18488 3176 -17796
rect 3210 -18488 3216 -17796
rect 3170 -18500 3216 -18488
rect 3698 -17796 3744 -17784
rect 3698 -18488 3704 -17796
rect 3738 -17800 3744 -17796
rect 3806 -17796 3852 -17784
rect 3806 -17800 3812 -17796
rect 3738 -17810 3812 -17800
rect 3738 -18480 3812 -18470
rect 3738 -18488 3744 -18480
rect 3698 -18500 3744 -18488
rect 3806 -18488 3812 -18480
rect 3846 -18488 3852 -17796
rect 3806 -18500 3852 -18488
rect 4334 -17796 4380 -17784
rect 4334 -18488 4340 -17796
rect 4374 -18488 4380 -17796
rect 4334 -18500 4380 -18488
rect 4770 -17796 4816 -17784
rect 4770 -18488 4776 -17796
rect 4810 -18488 4816 -17796
rect 4770 -18500 4816 -18488
rect 5298 -17796 5344 -17784
rect 5298 -18488 5304 -17796
rect 5338 -17800 5344 -17796
rect 5406 -17796 5452 -17784
rect 5406 -17800 5412 -17796
rect 5338 -17810 5412 -17800
rect 5338 -18480 5412 -18470
rect 5338 -18488 5344 -18480
rect 5298 -18500 5344 -18488
rect 5406 -18488 5412 -18480
rect 5446 -18488 5452 -17796
rect 5406 -18500 5452 -18488
rect 5934 -17796 5980 -17784
rect 5934 -18488 5940 -17796
rect 5974 -18488 5980 -17796
rect 5934 -18500 5980 -18488
rect 6370 -17796 6416 -17784
rect 6370 -18488 6376 -17796
rect 6410 -18488 6416 -17796
rect 6370 -18500 6416 -18488
rect 6898 -17796 6944 -17784
rect 6898 -18488 6904 -17796
rect 6938 -17800 6944 -17796
rect 7006 -17796 7052 -17784
rect 7006 -17800 7012 -17796
rect 6938 -17810 7012 -17800
rect 6938 -18480 7012 -18470
rect 6938 -18488 6944 -18480
rect 6898 -18500 6944 -18488
rect 7006 -18488 7012 -18480
rect 7046 -18488 7052 -17796
rect 7006 -18500 7052 -18488
rect 7534 -17796 7580 -17784
rect 7534 -18488 7540 -17796
rect 7574 -18488 7580 -17796
rect 7534 -18500 7580 -18488
rect 7970 -17796 8016 -17784
rect 7970 -18488 7976 -17796
rect 8010 -18488 8016 -17796
rect 7970 -18500 8016 -18488
rect 8498 -17796 8544 -17784
rect 8498 -18488 8504 -17796
rect 8538 -17800 8544 -17796
rect 8606 -17796 8652 -17784
rect 8606 -17800 8612 -17796
rect 8538 -17810 8612 -17800
rect 8538 -18480 8612 -18470
rect 8538 -18488 8544 -18480
rect 8498 -18500 8544 -18488
rect 8606 -18488 8612 -18480
rect 8646 -18488 8652 -17796
rect 8606 -18500 8652 -18488
rect 9134 -17796 9180 -17784
rect 9134 -18488 9140 -17796
rect 9174 -18488 9180 -17796
rect 9134 -18500 9180 -18488
rect 9570 -17796 9616 -17784
rect 9570 -18488 9576 -17796
rect 9610 -18488 9616 -17796
rect 9570 -18500 9616 -18488
rect 10098 -17796 10144 -17784
rect 10098 -18488 10104 -17796
rect 10138 -17800 10144 -17796
rect 10206 -17796 10252 -17784
rect 10206 -17800 10212 -17796
rect 10138 -17810 10212 -17800
rect 10138 -18480 10212 -18470
rect 10138 -18488 10144 -18480
rect 10098 -18500 10144 -18488
rect 10206 -18488 10212 -18480
rect 10246 -18488 10252 -17796
rect 10206 -18500 10252 -18488
rect 10734 -17796 10780 -17784
rect 10734 -18488 10740 -17796
rect 10774 -18488 10780 -17796
rect 10734 -18500 10780 -18488
rect 11170 -17796 11216 -17784
rect 11170 -18488 11176 -17796
rect 11210 -18070 11216 -17796
rect 11400 -18070 11510 -17736
rect 11698 -17796 11744 -17784
rect 11698 -18070 11704 -17796
rect 11210 -18220 11704 -18070
rect 11210 -18488 11216 -18220
rect 11170 -18500 11216 -18488
rect 11400 -18548 11510 -18220
rect 11698 -18488 11704 -18220
rect 11738 -18070 11744 -17796
rect 11806 -17796 11852 -17784
rect 11806 -18070 11812 -17796
rect 11738 -18220 11812 -18070
rect 11738 -18488 11744 -18220
rect 11698 -18500 11744 -18488
rect 11806 -18488 11812 -18220
rect 11846 -18070 11852 -17796
rect 12040 -18070 12150 -17736
rect 12334 -17796 12380 -17784
rect 12334 -18070 12340 -17796
rect 11846 -18220 12340 -18070
rect 11846 -18488 11852 -18220
rect 11806 -18500 11852 -18488
rect 12040 -18548 12150 -18220
rect 12334 -18488 12340 -18220
rect 12374 -18488 12380 -17796
rect 12334 -18500 12380 -18488
rect 12770 -17796 12816 -17784
rect 12770 -18488 12776 -17796
rect 12810 -18488 12816 -17796
rect 12770 -18500 12816 -18488
rect 13298 -17796 13344 -17784
rect 13298 -18488 13304 -17796
rect 13338 -17800 13344 -17796
rect 13406 -17796 13452 -17784
rect 13406 -17800 13412 -17796
rect 13338 -17810 13412 -17800
rect 13338 -18480 13412 -18470
rect 13338 -18488 13344 -18480
rect 13298 -18500 13344 -18488
rect 13406 -18488 13412 -18480
rect 13446 -18488 13452 -17796
rect 13406 -18500 13452 -18488
rect 13934 -17796 13980 -17784
rect 13934 -18488 13940 -17796
rect 13974 -18488 13980 -17796
rect 13934 -18500 13980 -18488
rect 14370 -17796 14416 -17784
rect 14370 -18488 14376 -17796
rect 14410 -18488 14416 -17796
rect 14370 -18500 14416 -18488
rect 14898 -17796 14944 -17784
rect 14898 -18488 14904 -17796
rect 14938 -17800 14944 -17796
rect 15006 -17796 15052 -17784
rect 15006 -17800 15012 -17796
rect 14938 -17810 15012 -17800
rect 14938 -18480 15012 -18470
rect 14938 -18488 14944 -18480
rect 14898 -18500 14944 -18488
rect 15006 -18488 15012 -18480
rect 15046 -18488 15052 -17796
rect 15006 -18500 15052 -18488
rect 15534 -17796 15580 -17784
rect 15534 -18488 15540 -17796
rect 15574 -18488 15580 -17796
rect 15534 -18500 15580 -18488
rect 15970 -17796 16016 -17784
rect 15970 -18488 15976 -17796
rect 16010 -18488 16016 -17796
rect 15970 -18500 16016 -18488
rect 16498 -17790 16544 -17784
rect 16606 -17790 16652 -17784
rect 16498 -17796 16652 -17790
rect 16498 -18488 16504 -17796
rect 16538 -17800 16612 -17796
rect 16538 -18488 16612 -18480
rect 16646 -18488 16652 -17796
rect 16498 -18490 16652 -18488
rect 16498 -18500 16544 -18490
rect 16606 -18500 16652 -18490
rect 17134 -17796 17180 -17784
rect 17134 -18488 17140 -17796
rect 17174 -18488 17180 -17796
rect 17134 -18500 17180 -18488
rect 17570 -17796 17616 -17784
rect 17570 -18488 17576 -17796
rect 17610 -18488 17616 -17796
rect 17570 -18500 17616 -18488
rect 18098 -17790 18144 -17784
rect 18206 -17790 18252 -17784
rect 18098 -17796 18252 -17790
rect 18098 -18488 18104 -17796
rect 18138 -17800 18212 -17796
rect 18138 -18488 18212 -18480
rect 18246 -18488 18252 -17796
rect 18098 -18490 18252 -18488
rect 18098 -18500 18144 -18490
rect 18206 -18500 18252 -18490
rect 18734 -17796 18780 -17784
rect 18734 -18488 18740 -17796
rect 18774 -18488 18780 -17796
rect 18734 -18500 18780 -18488
rect 19170 -17796 19216 -17784
rect 19170 -18488 19176 -17796
rect 19210 -18488 19216 -17796
rect 19170 -18500 19216 -18488
rect 19698 -17790 19744 -17784
rect 19806 -17790 19852 -17784
rect 19698 -17796 19852 -17790
rect 19698 -18488 19704 -17796
rect 19738 -17800 19812 -17796
rect 19738 -18488 19812 -18480
rect 19846 -18488 19852 -17796
rect 19698 -18490 19852 -18488
rect 19698 -18500 19744 -18490
rect 19806 -18500 19852 -18490
rect 20334 -17796 20380 -17784
rect 20334 -18488 20340 -17796
rect 20374 -18488 20380 -17796
rect 20334 -18500 20380 -18488
rect 20770 -17796 20816 -17784
rect 20770 -18488 20776 -17796
rect 20810 -18488 20816 -17796
rect 20770 -18500 20816 -18488
rect 21298 -17790 21344 -17784
rect 21406 -17790 21452 -17784
rect 21298 -17796 21452 -17790
rect 21298 -18488 21304 -17796
rect 21338 -17800 21412 -17796
rect 21338 -18488 21412 -18480
rect 21446 -18488 21452 -17796
rect 21298 -18490 21452 -18488
rect 21298 -18500 21344 -18490
rect 21406 -18500 21452 -18490
rect 21934 -17796 21980 -17784
rect 21934 -18488 21940 -17796
rect 21974 -18488 21980 -17796
rect 21934 -18500 21980 -18488
rect 22370 -17796 22416 -17784
rect 22370 -18488 22376 -17796
rect 22410 -18488 22416 -17796
rect 22370 -18500 22416 -18488
rect 22898 -17790 22944 -17784
rect 23006 -17790 23052 -17784
rect 22898 -17796 23052 -17790
rect 22898 -18488 22904 -17796
rect 22938 -17800 23012 -17796
rect 22938 -18488 23012 -18480
rect 23046 -18488 23052 -17796
rect 22898 -18490 23052 -18488
rect 22898 -18500 22944 -18490
rect 23006 -18500 23052 -18490
rect 23534 -17796 23580 -17784
rect 23534 -18488 23540 -17796
rect 23574 -18488 23580 -17796
rect 23534 -18500 23580 -18488
rect 23970 -17796 24016 -17784
rect 23970 -18488 23976 -17796
rect 24010 -18488 24016 -17796
rect 23970 -18500 24016 -18488
rect 24498 -17790 24544 -17784
rect 24606 -17790 24652 -17784
rect 24498 -17796 24652 -17790
rect 24498 -18488 24504 -17796
rect 24538 -17800 24612 -17796
rect 24538 -18488 24612 -18480
rect 24646 -18488 24652 -17796
rect 24498 -18490 24652 -18488
rect 24498 -18500 24544 -18490
rect 24606 -18500 24652 -18490
rect 25134 -17796 25180 -17784
rect 25134 -18488 25140 -17796
rect 25174 -18488 25180 -17796
rect 25134 -18500 25180 -18488
rect 25570 -17796 25616 -17784
rect 25570 -18488 25576 -17796
rect 25610 -18488 25616 -17796
rect 25570 -18500 25616 -18488
rect 26098 -17790 26144 -17784
rect 26206 -17790 26252 -17784
rect 26098 -17796 26252 -17790
rect 26098 -18488 26104 -17796
rect 26138 -17800 26212 -17796
rect 26138 -18488 26212 -18480
rect 26246 -18488 26252 -17796
rect 26098 -18490 26252 -18488
rect 26098 -18500 26144 -18490
rect 26206 -18500 26252 -18490
rect 26734 -17796 26780 -17784
rect 26734 -18488 26740 -17796
rect 26774 -18488 26780 -17796
rect 26734 -18500 26780 -18488
rect 27170 -17796 27216 -17784
rect 27170 -18488 27176 -17796
rect 27210 -18488 27216 -17796
rect 27170 -18500 27216 -18488
rect 27698 -17790 27744 -17784
rect 27806 -17790 27852 -17784
rect 27698 -17796 27852 -17790
rect 27698 -18488 27704 -17796
rect 27738 -17800 27812 -17796
rect 27738 -18488 27812 -18480
rect 27846 -18488 27852 -17796
rect 27698 -18490 27852 -18488
rect 27698 -18500 27744 -18490
rect 27806 -18500 27852 -18490
rect 28334 -17796 28380 -17784
rect 28334 -18488 28340 -17796
rect 28374 -18488 28380 -17796
rect 28334 -18500 28380 -18488
rect 28770 -17796 28816 -17784
rect 28770 -18488 28776 -17796
rect 28810 -18488 28816 -17796
rect 28770 -18500 28816 -18488
rect 29298 -17790 29344 -17784
rect 29406 -17790 29452 -17784
rect 29298 -17796 29452 -17790
rect 29298 -18488 29304 -17796
rect 29338 -17800 29412 -17796
rect 29338 -18488 29412 -18480
rect 29446 -18488 29452 -17796
rect 29298 -18490 29452 -18488
rect 29298 -18500 29344 -18490
rect 29406 -18500 29452 -18490
rect 29934 -17796 29980 -17784
rect 29934 -18488 29940 -17796
rect 29974 -18488 29980 -17796
rect 29934 -18500 29980 -18488
rect 30370 -17796 30416 -17784
rect 30370 -18488 30376 -17796
rect 30410 -18488 30416 -17796
rect 30370 -18500 30416 -18488
rect 30898 -17790 30944 -17784
rect 31006 -17790 31052 -17784
rect 30898 -17796 31052 -17790
rect 30898 -18488 30904 -17796
rect 30938 -17800 31012 -17796
rect 30938 -18488 31012 -18480
rect 31046 -18488 31052 -17796
rect 30898 -18490 31052 -18488
rect 30898 -18500 30944 -18490
rect 31006 -18500 31052 -18490
rect 31534 -17796 31580 -17784
rect 31534 -18488 31540 -17796
rect 31574 -18488 31580 -17796
rect 31534 -18500 31580 -18488
rect 31970 -17796 32016 -17784
rect 31970 -18488 31976 -17796
rect 32010 -18488 32016 -17796
rect 31970 -18500 32016 -18488
rect 32498 -17790 32544 -17784
rect 32606 -17790 32652 -17784
rect 32498 -17796 32652 -17790
rect 32498 -18488 32504 -17796
rect 32538 -17800 32612 -17796
rect 32538 -18488 32612 -18480
rect 32646 -18488 32652 -17796
rect 32498 -18490 32652 -18488
rect 32498 -18500 32544 -18490
rect 32606 -18500 32652 -18490
rect 33134 -17796 33180 -17784
rect 33134 -18488 33140 -17796
rect 33174 -18488 33180 -17796
rect 33134 -18500 33180 -18488
rect 33570 -17796 33616 -17784
rect 33570 -18488 33576 -17796
rect 33610 -18488 33616 -17796
rect 33570 -18500 33616 -18488
rect 34098 -17790 34144 -17784
rect 34206 -17790 34252 -17784
rect 34098 -17796 34252 -17790
rect 34098 -18488 34104 -17796
rect 34138 -17800 34212 -17796
rect 34138 -18488 34212 -18480
rect 34246 -18488 34252 -17796
rect 34098 -18490 34252 -18488
rect 34098 -18500 34144 -18490
rect 34206 -18500 34252 -18490
rect 34734 -17796 34780 -17784
rect 34734 -18488 34740 -17796
rect 34774 -18488 34780 -17796
rect 34734 -18500 34780 -18488
rect 35170 -17796 35216 -17784
rect 35170 -18488 35176 -17796
rect 35210 -18488 35216 -17796
rect 35170 -18500 35216 -18488
rect 35698 -17790 35744 -17784
rect 35806 -17790 35852 -17784
rect 35698 -17796 35852 -17790
rect 35698 -18488 35704 -17796
rect 35738 -17800 35812 -17796
rect 35738 -18488 35812 -18480
rect 35846 -18488 35852 -17796
rect 35698 -18490 35852 -18488
rect 35698 -18500 35744 -18490
rect 35806 -18500 35852 -18490
rect 36334 -17796 36380 -17784
rect 36334 -18488 36340 -17796
rect 36374 -18488 36380 -17796
rect 36334 -18500 36380 -18488
rect 36770 -17796 36816 -17784
rect 36770 -18488 36776 -17796
rect 36810 -18488 36816 -17796
rect 36770 -18500 36816 -18488
rect 37298 -17796 37344 -17784
rect 37298 -18488 37304 -17796
rect 37338 -18488 37344 -17796
rect 37298 -18500 37344 -18488
rect 37406 -17796 37452 -17784
rect 37406 -18488 37412 -17796
rect 37446 -18488 37452 -17796
rect 37406 -18500 37452 -18488
rect 37934 -17796 37980 -17784
rect 37934 -18488 37940 -17796
rect 37974 -18488 37980 -17796
rect 37934 -18500 37980 -18488
rect 670 -18554 1093 -18548
rect 670 -18588 705 -18554
rect 1081 -18560 1093 -18554
rect 1657 -18554 2057 -18548
rect 1657 -18560 1669 -18554
rect 1081 -18588 1669 -18560
rect 2045 -18560 2057 -18554
rect 2293 -18554 2693 -18548
rect 2293 -18560 2305 -18554
rect 2045 -18588 2305 -18560
rect 2681 -18560 2693 -18554
rect 3257 -18554 3657 -18548
rect 3257 -18560 3269 -18554
rect 2681 -18588 3269 -18560
rect 3645 -18560 3657 -18554
rect 3893 -18554 4293 -18548
rect 3893 -18560 3905 -18554
rect 3645 -18588 3905 -18560
rect 4281 -18560 4293 -18554
rect 4857 -18554 5257 -18548
rect 4857 -18560 4869 -18554
rect 4281 -18588 4869 -18560
rect 5245 -18560 5257 -18554
rect 5493 -18554 5893 -18548
rect 5493 -18560 5505 -18554
rect 5245 -18588 5505 -18560
rect 5881 -18560 5893 -18554
rect 6457 -18554 6857 -18548
rect 6457 -18560 6469 -18554
rect 5881 -18588 6469 -18560
rect 6845 -18560 6857 -18554
rect 7093 -18554 7493 -18548
rect 7093 -18560 7105 -18554
rect 6845 -18588 7105 -18560
rect 7481 -18560 7493 -18554
rect 8057 -18554 8457 -18548
rect 8057 -18560 8069 -18554
rect 7481 -18588 8069 -18560
rect 8445 -18560 8457 -18554
rect 8693 -18554 9093 -18548
rect 8693 -18560 8705 -18554
rect 8445 -18588 8705 -18560
rect 9081 -18560 9093 -18554
rect 9657 -18554 10057 -18548
rect 9657 -18560 9669 -18554
rect 9081 -18588 9669 -18560
rect 10045 -18560 10057 -18554
rect 10293 -18554 10693 -18548
rect 10293 -18560 10305 -18554
rect 10045 -18588 10305 -18560
rect 10681 -18560 10693 -18554
rect 11257 -18554 11657 -18548
rect 11257 -18560 11269 -18554
rect 10681 -18588 11269 -18560
rect 11645 -18560 11657 -18554
rect 11893 -18554 12293 -18548
rect 11893 -18560 11905 -18554
rect 11645 -18588 11905 -18560
rect 12281 -18560 12293 -18554
rect 12857 -18554 13257 -18548
rect 12857 -18560 12869 -18554
rect 12281 -18588 12869 -18560
rect 13245 -18560 13257 -18554
rect 13493 -18554 13893 -18548
rect 13493 -18560 13505 -18554
rect 13245 -18588 13505 -18560
rect 13881 -18560 13893 -18554
rect 14457 -18554 14857 -18548
rect 14457 -18560 14469 -18554
rect 13881 -18588 14469 -18560
rect 14845 -18560 14857 -18554
rect 15093 -18554 15493 -18548
rect 15093 -18560 15105 -18554
rect 14845 -18588 15105 -18560
rect 15481 -18560 15493 -18554
rect 16057 -18554 16457 -18548
rect 16057 -18560 16069 -18554
rect 15481 -18588 16069 -18560
rect 16445 -18560 16457 -18554
rect 16693 -18554 17093 -18548
rect 16693 -18560 16705 -18554
rect 16445 -18588 16705 -18560
rect 17081 -18560 17093 -18554
rect 17657 -18554 18057 -18548
rect 17657 -18560 17669 -18554
rect 17081 -18588 17669 -18560
rect 18045 -18560 18057 -18554
rect 18293 -18554 18693 -18548
rect 18293 -18560 18305 -18554
rect 18045 -18588 18305 -18560
rect 18681 -18560 18693 -18554
rect 19257 -18554 19657 -18548
rect 19257 -18560 19269 -18554
rect 18681 -18588 19269 -18560
rect 19645 -18560 19657 -18554
rect 19893 -18554 20293 -18548
rect 19893 -18560 19905 -18554
rect 19645 -18588 19905 -18560
rect 20281 -18560 20293 -18554
rect 20857 -18554 21257 -18548
rect 20857 -18560 20869 -18554
rect 20281 -18588 20869 -18560
rect 21245 -18560 21257 -18554
rect 21493 -18554 21893 -18548
rect 21493 -18560 21505 -18554
rect 21245 -18588 21505 -18560
rect 21881 -18560 21893 -18554
rect 22457 -18554 22857 -18548
rect 22457 -18560 22469 -18554
rect 21881 -18588 22469 -18560
rect 22845 -18560 22857 -18554
rect 23093 -18554 23493 -18548
rect 23093 -18560 23105 -18554
rect 22845 -18588 23105 -18560
rect 23481 -18560 23493 -18554
rect 24057 -18554 24457 -18548
rect 24057 -18560 24069 -18554
rect 23481 -18588 24069 -18560
rect 24445 -18560 24457 -18554
rect 24693 -18554 25093 -18548
rect 24693 -18560 24705 -18554
rect 24445 -18588 24705 -18560
rect 25081 -18560 25093 -18554
rect 25657 -18554 26057 -18548
rect 25657 -18560 25669 -18554
rect 25081 -18588 25669 -18560
rect 26045 -18560 26057 -18554
rect 26293 -18554 26693 -18548
rect 26293 -18560 26305 -18554
rect 26045 -18588 26305 -18560
rect 26681 -18560 26693 -18554
rect 27257 -18554 27657 -18548
rect 27257 -18560 27269 -18554
rect 26681 -18588 27269 -18560
rect 27645 -18560 27657 -18554
rect 27893 -18554 28293 -18548
rect 27893 -18560 27905 -18554
rect 27645 -18588 27905 -18560
rect 28281 -18560 28293 -18554
rect 28857 -18554 29257 -18548
rect 28857 -18560 28869 -18554
rect 28281 -18588 28869 -18560
rect 29245 -18560 29257 -18554
rect 29493 -18554 29893 -18548
rect 29493 -18560 29505 -18554
rect 29245 -18588 29505 -18560
rect 29881 -18560 29893 -18554
rect 30457 -18554 30857 -18548
rect 30457 -18560 30469 -18554
rect 29881 -18588 30469 -18560
rect 30845 -18560 30857 -18554
rect 31093 -18554 31493 -18548
rect 31093 -18560 31105 -18554
rect 30845 -18588 31105 -18560
rect 31481 -18560 31493 -18554
rect 32057 -18554 32457 -18548
rect 32057 -18560 32069 -18554
rect 31481 -18588 32069 -18560
rect 32445 -18560 32457 -18554
rect 32693 -18554 33093 -18548
rect 32693 -18560 32705 -18554
rect 32445 -18588 32705 -18560
rect 33081 -18560 33093 -18554
rect 33657 -18554 34057 -18548
rect 33657 -18560 33669 -18554
rect 33081 -18588 33669 -18560
rect 34045 -18560 34057 -18554
rect 34293 -18554 34693 -18548
rect 34293 -18560 34305 -18554
rect 34045 -18588 34305 -18560
rect 34681 -18560 34693 -18554
rect 35257 -18554 35657 -18548
rect 35257 -18560 35269 -18554
rect 34681 -18588 35269 -18560
rect 35645 -18560 35657 -18554
rect 35893 -18554 36293 -18548
rect 35893 -18560 35905 -18554
rect 35645 -18588 35905 -18560
rect 36281 -18560 36293 -18554
rect 36857 -18554 37257 -18548
rect 36857 -18560 36869 -18554
rect 36281 -18588 36869 -18560
rect 37245 -18560 37257 -18554
rect 37493 -18554 37893 -18548
rect 37493 -18560 37505 -18554
rect 37245 -18588 37505 -18560
rect 37881 -18588 37893 -18554
rect 670 -18594 37893 -18588
rect 670 -18682 37880 -18594
rect 670 -18688 37949 -18682
rect 0 -18722 13 -18688
rect 1137 -18722 1613 -18688
rect 2737 -18722 3213 -18688
rect 4337 -18722 4813 -18688
rect 5937 -18722 6413 -18688
rect 7537 -18722 8013 -18688
rect 9137 -18722 9613 -18688
rect 10737 -18722 11213 -18688
rect 12337 -18722 12813 -18688
rect 13937 -18722 14413 -18688
rect 15537 -18722 16013 -18688
rect 17137 -18722 17613 -18688
rect 18737 -18722 19213 -18688
rect 20337 -18722 20813 -18688
rect 21937 -18722 22413 -18688
rect 23537 -18722 24013 -18688
rect 25137 -18722 25613 -18688
rect 26737 -18722 27213 -18688
rect 28337 -18722 28813 -18688
rect 29937 -18722 30413 -18688
rect 31537 -18722 32013 -18688
rect 33137 -18722 33613 -18688
rect 34737 -18722 35213 -18688
rect 36337 -18722 36813 -18688
rect 37937 -18722 37949 -18688
rect 0 -18820 490 -18722
rect 440 -18964 490 -18820
rect 57 -18970 490 -18964
rect 57 -19004 69 -18970
rect 445 -19004 490 -18970
rect 57 -19010 490 -19004
rect -30 -19057 16 -19045
rect -30 -19175 -24 -19057
rect 10 -19175 16 -19057
rect -30 -19187 16 -19175
rect 440 -19222 490 -19010
rect 670 -18728 37949 -18722
rect 670 -18820 37940 -18728
rect 670 -18964 720 -18820
rect 1200 -18870 1340 -18860
rect 670 -18970 1093 -18964
rect 670 -19004 705 -18970
rect 1081 -19004 1093 -18970
rect 1200 -18990 1210 -18870
rect 1330 -18880 1340 -18870
rect 2800 -18870 2940 -18860
rect 2800 -18880 2810 -18870
rect 1330 -18970 2810 -18880
rect 1330 -18980 1669 -18970
rect 1330 -18990 1340 -18980
rect 1200 -19000 1340 -18990
rect 670 -19010 1093 -19004
rect 1657 -19004 1669 -18980
rect 2045 -18980 2305 -18970
rect 2045 -19004 2057 -18980
rect 1657 -19010 2057 -19004
rect 2293 -19004 2305 -18980
rect 2681 -18980 2810 -18970
rect 2681 -19004 2693 -18980
rect 2800 -18990 2810 -18980
rect 2930 -18880 2940 -18870
rect 4400 -18870 4540 -18860
rect 4400 -18880 4410 -18870
rect 2930 -18970 4410 -18880
rect 2930 -18980 3269 -18970
rect 2930 -18990 2940 -18980
rect 2800 -19000 2940 -18990
rect 2293 -19010 2693 -19004
rect 3257 -19004 3269 -18980
rect 3645 -18980 3905 -18970
rect 3645 -19004 3657 -18980
rect 3257 -19010 3657 -19004
rect 3893 -19004 3905 -18980
rect 4281 -18980 4410 -18970
rect 4281 -19004 4293 -18980
rect 4400 -18990 4410 -18980
rect 4530 -18880 4540 -18870
rect 6000 -18870 6140 -18860
rect 6000 -18880 6010 -18870
rect 4530 -18970 6010 -18880
rect 4530 -18980 4869 -18970
rect 4530 -18990 4540 -18980
rect 4400 -19000 4540 -18990
rect 3893 -19010 4293 -19004
rect 4857 -19004 4869 -18980
rect 5245 -18980 5505 -18970
rect 5245 -19004 5257 -18980
rect 4857 -19010 5257 -19004
rect 5493 -19004 5505 -18980
rect 5881 -18980 6010 -18970
rect 5881 -19004 5893 -18980
rect 6000 -18990 6010 -18980
rect 6130 -18880 6140 -18870
rect 7600 -18870 7740 -18860
rect 7600 -18880 7610 -18870
rect 6130 -18970 7610 -18880
rect 6130 -18980 6469 -18970
rect 6130 -18990 6140 -18980
rect 6000 -19000 6140 -18990
rect 5493 -19010 5893 -19004
rect 6457 -19004 6469 -18980
rect 6845 -18980 7105 -18970
rect 6845 -19004 6857 -18980
rect 6457 -19010 6857 -19004
rect 7093 -19004 7105 -18980
rect 7481 -18980 7610 -18970
rect 7481 -19004 7493 -18980
rect 7600 -18990 7610 -18980
rect 7730 -18880 7740 -18870
rect 9200 -18870 9340 -18860
rect 15820 -18870 15960 -18860
rect 9200 -18880 9210 -18870
rect 7730 -18970 9210 -18880
rect 7730 -18980 8069 -18970
rect 7730 -18990 7740 -18980
rect 7600 -19000 7740 -18990
rect 7093 -19010 7493 -19004
rect 8057 -19004 8069 -18980
rect 8445 -18980 8705 -18970
rect 8445 -19004 8457 -18980
rect 8057 -19010 8457 -19004
rect 8693 -19004 8705 -18980
rect 9081 -18980 9210 -18970
rect 9081 -19004 9093 -18980
rect 9200 -18990 9210 -18980
rect 9330 -18880 9340 -18870
rect 12400 -18880 12540 -18870
rect 9330 -18970 10700 -18880
rect 9330 -18980 9669 -18970
rect 9330 -18990 9340 -18980
rect 9200 -19000 9340 -18990
rect 8693 -19010 9093 -19004
rect 9657 -19004 9669 -18980
rect 10045 -18980 10305 -18970
rect 10045 -19004 10057 -18980
rect 9657 -19010 10057 -19004
rect 10293 -19004 10305 -18980
rect 10681 -18980 10700 -18970
rect 11257 -18970 11657 -18964
rect 10681 -19004 10693 -18980
rect 10293 -19010 10693 -19004
rect 11257 -19004 11269 -18970
rect 11645 -19004 11657 -18970
rect 11257 -19010 11657 -19004
rect 11893 -18970 12293 -18964
rect 11893 -19004 11905 -18970
rect 12281 -19004 12293 -18970
rect 11893 -19010 12293 -19004
rect 12400 -19000 12410 -18880
rect 12530 -18910 12540 -18880
rect 12530 -18964 15490 -18910
rect 12530 -18970 15493 -18964
rect 12530 -19000 12869 -18970
rect 12400 -19010 12540 -19000
rect 12857 -19004 12869 -19000
rect 13245 -19000 13505 -18970
rect 13245 -19004 13257 -19000
rect 12857 -19010 13257 -19004
rect 13493 -19004 13505 -19000
rect 13881 -19000 14469 -18970
rect 13881 -19004 13893 -19000
rect 13493 -19010 13893 -19004
rect 14457 -19004 14469 -19000
rect 14845 -19000 15105 -18970
rect 14845 -19004 14857 -19000
rect 14457 -19010 14857 -19004
rect 15093 -19004 15105 -19000
rect 15481 -19004 15493 -18970
rect 15820 -18990 15830 -18870
rect 15950 -18900 15960 -18870
rect 17420 -18870 17560 -18860
rect 15950 -18964 17090 -18900
rect 15950 -18970 17093 -18964
rect 15950 -18990 16069 -18970
rect 15820 -19000 16069 -18990
rect 15093 -19010 15493 -19004
rect 16057 -19004 16069 -19000
rect 16445 -19000 16705 -18970
rect 16445 -19004 16457 -19000
rect 16057 -19010 16457 -19004
rect 16693 -19004 16705 -19000
rect 17081 -19004 17093 -18970
rect 17420 -18990 17430 -18870
rect 17550 -18900 17560 -18870
rect 19020 -18870 19160 -18860
rect 17550 -18964 18690 -18900
rect 17550 -18970 18693 -18964
rect 17550 -18990 17669 -18970
rect 17420 -19000 17669 -18990
rect 16693 -19010 17093 -19004
rect 17657 -19004 17669 -19000
rect 18045 -19000 18305 -18970
rect 18045 -19004 18057 -19000
rect 17657 -19010 18057 -19004
rect 18293 -19004 18305 -19000
rect 18681 -19004 18693 -18970
rect 19020 -18990 19030 -18870
rect 19150 -18900 19160 -18870
rect 20620 -18870 20760 -18860
rect 19150 -18964 20290 -18900
rect 19150 -18970 20293 -18964
rect 19150 -18990 19269 -18970
rect 19020 -19000 19269 -18990
rect 18293 -19010 18693 -19004
rect 19257 -19004 19269 -19000
rect 19645 -19000 19905 -18970
rect 19645 -19004 19657 -19000
rect 19257 -19010 19657 -19004
rect 19893 -19004 19905 -19000
rect 20281 -19004 20293 -18970
rect 20620 -18990 20630 -18870
rect 20750 -18900 20760 -18870
rect 22220 -18870 22360 -18860
rect 20750 -18964 21890 -18900
rect 20750 -18970 21893 -18964
rect 20750 -18990 20869 -18970
rect 20620 -19000 20869 -18990
rect 19893 -19010 20293 -19004
rect 20857 -19004 20869 -19000
rect 21245 -19000 21505 -18970
rect 21245 -19004 21257 -19000
rect 20857 -19010 21257 -19004
rect 21493 -19004 21505 -19000
rect 21881 -19004 21893 -18970
rect 22220 -18990 22230 -18870
rect 22350 -18900 22360 -18870
rect 23820 -18870 23960 -18860
rect 22350 -18964 23490 -18900
rect 22350 -18970 23493 -18964
rect 22350 -18990 22469 -18970
rect 22220 -19000 22469 -18990
rect 21493 -19010 21893 -19004
rect 22457 -19004 22469 -19000
rect 22845 -19000 23105 -18970
rect 22845 -19004 22857 -19000
rect 22457 -19010 22857 -19004
rect 23093 -19004 23105 -19000
rect 23481 -19004 23493 -18970
rect 23820 -18990 23830 -18870
rect 23950 -18900 23960 -18870
rect 27020 -18870 27160 -18860
rect 27020 -18900 27030 -18870
rect 23950 -18964 25090 -18900
rect 25660 -18964 27030 -18900
rect 23950 -18970 25093 -18964
rect 23950 -18990 24069 -18970
rect 23820 -19000 24069 -18990
rect 23093 -19010 23493 -19004
rect 24057 -19004 24069 -19000
rect 24445 -19000 24705 -18970
rect 24445 -19004 24457 -19000
rect 24057 -19010 24457 -19004
rect 24693 -19004 24705 -19000
rect 25081 -19004 25093 -18970
rect 24693 -19010 25093 -19004
rect 25657 -18970 27030 -18964
rect 25657 -19004 25669 -18970
rect 26045 -19000 26305 -18970
rect 26045 -19004 26057 -19000
rect 25657 -19010 26057 -19004
rect 26293 -19004 26305 -19000
rect 26681 -18990 27030 -18970
rect 27150 -18900 27160 -18870
rect 28620 -18870 28760 -18860
rect 27150 -18964 28290 -18900
rect 27150 -18970 28293 -18964
rect 27150 -18990 27269 -18970
rect 26681 -19000 27269 -18990
rect 26681 -19004 26693 -19000
rect 26293 -19010 26693 -19004
rect 27257 -19004 27269 -19000
rect 27645 -19000 27905 -18970
rect 27645 -19004 27657 -19000
rect 27257 -19010 27657 -19004
rect 27893 -19004 27905 -19000
rect 28281 -19004 28293 -18970
rect 28620 -18990 28630 -18870
rect 28750 -18900 28760 -18870
rect 31580 -18880 31720 -18870
rect 28750 -18964 31490 -18900
rect 28750 -18970 31493 -18964
rect 28750 -18990 28869 -18970
rect 28620 -19000 28869 -18990
rect 27893 -19010 28293 -19004
rect 28857 -19004 28869 -19000
rect 29245 -19000 29505 -18970
rect 29245 -19004 29257 -19000
rect 28857 -19010 29257 -19004
rect 29493 -19004 29505 -19000
rect 29881 -19000 30469 -18970
rect 29881 -19004 29893 -19000
rect 29493 -19010 29893 -19004
rect 30457 -19004 30469 -19000
rect 30845 -19000 31105 -18970
rect 30845 -19004 30857 -19000
rect 30457 -19010 30857 -19004
rect 31093 -19004 31105 -19000
rect 31481 -19004 31493 -18970
rect 31093 -19010 31493 -19004
rect 31580 -19000 31590 -18880
rect 31710 -18900 31720 -18880
rect 31710 -18964 36280 -18900
rect 31710 -18970 36293 -18964
rect 31710 -19000 32069 -18970
rect 31580 -19010 31720 -19000
rect 32057 -19004 32069 -19000
rect 32445 -19000 32705 -18970
rect 32445 -19004 32457 -19000
rect 32057 -19010 32457 -19004
rect 32693 -19004 32705 -19000
rect 33081 -19000 33669 -18970
rect 33081 -19004 33093 -19000
rect 32693 -19010 33093 -19004
rect 33657 -19004 33669 -19000
rect 34045 -19000 34305 -18970
rect 34045 -19004 34057 -19000
rect 33657 -19010 34057 -19004
rect 34293 -19004 34305 -19000
rect 34681 -19000 35269 -18970
rect 34681 -19004 34693 -19000
rect 34293 -19010 34693 -19004
rect 35257 -19004 35269 -19000
rect 35645 -19000 35905 -18970
rect 35645 -19004 35657 -19000
rect 35257 -19010 35657 -19004
rect 35893 -19004 35905 -19000
rect 36281 -19004 36293 -18970
rect 35893 -19010 36293 -19004
rect 36857 -18970 37257 -18964
rect 36857 -19004 36869 -18970
rect 37245 -19004 37257 -18970
rect 36857 -19010 37257 -19004
rect 37493 -18970 37893 -18964
rect 37493 -19004 37505 -18970
rect 37881 -19004 37893 -18970
rect 37493 -19010 37893 -19004
rect 57 -19228 490 -19222
rect 57 -19262 69 -19228
rect 445 -19262 490 -19228
rect 57 -19268 490 -19262
rect 440 -19490 490 -19268
rect 57 -19496 490 -19490
rect 57 -19530 69 -19496
rect 445 -19530 490 -19496
rect 57 -19536 490 -19530
rect -30 -19596 16 -19584
rect -30 -20288 -24 -19596
rect 10 -20288 16 -19596
rect -30 -20300 16 -20288
rect 440 -20348 490 -19536
rect 670 -19222 720 -19010
rect 1134 -19057 1180 -19045
rect 1134 -19175 1140 -19057
rect 1174 -19175 1180 -19057
rect 1570 -19057 1616 -19045
rect 1570 -19060 1576 -19057
rect 1134 -19187 1180 -19175
rect 1560 -19175 1576 -19060
rect 1610 -19060 1616 -19057
rect 2098 -19057 2144 -19045
rect 2098 -19060 2104 -19057
rect 1610 -19175 2104 -19060
rect 2138 -19060 2144 -19057
rect 2206 -19057 2252 -19045
rect 2206 -19060 2212 -19057
rect 2138 -19175 2212 -19060
rect 2246 -19060 2252 -19057
rect 2734 -19057 2780 -19045
rect 2734 -19060 2740 -19057
rect 2246 -19175 2740 -19060
rect 2774 -19060 2780 -19057
rect 3170 -19057 3216 -19045
rect 3170 -19060 3176 -19057
rect 2774 -19175 3176 -19060
rect 3210 -19060 3216 -19057
rect 3698 -19057 3744 -19045
rect 3698 -19060 3704 -19057
rect 3210 -19175 3704 -19060
rect 3738 -19060 3744 -19057
rect 3806 -19057 3852 -19045
rect 3806 -19060 3812 -19057
rect 3738 -19175 3812 -19060
rect 3846 -19060 3852 -19057
rect 4334 -19057 4380 -19045
rect 4334 -19060 4340 -19057
rect 3846 -19175 4340 -19060
rect 4374 -19060 4380 -19057
rect 4770 -19057 4816 -19045
rect 4770 -19060 4776 -19057
rect 4374 -19175 4776 -19060
rect 4810 -19060 4816 -19057
rect 5298 -19057 5344 -19045
rect 5298 -19060 5304 -19057
rect 4810 -19175 5304 -19060
rect 5338 -19060 5344 -19057
rect 5406 -19057 5452 -19045
rect 5406 -19060 5412 -19057
rect 5338 -19175 5412 -19060
rect 5446 -19060 5452 -19057
rect 5934 -19057 5980 -19045
rect 5934 -19060 5940 -19057
rect 5446 -19175 5940 -19060
rect 5974 -19060 5980 -19057
rect 6370 -19057 6416 -19045
rect 6370 -19060 6376 -19057
rect 5974 -19175 6376 -19060
rect 6410 -19060 6416 -19057
rect 6898 -19057 6944 -19045
rect 6898 -19060 6904 -19057
rect 6410 -19175 6904 -19060
rect 6938 -19060 6944 -19057
rect 7006 -19057 7052 -19045
rect 7006 -19060 7012 -19057
rect 6938 -19175 7012 -19060
rect 7046 -19060 7052 -19057
rect 7534 -19057 7580 -19045
rect 7534 -19060 7540 -19057
rect 7046 -19175 7540 -19060
rect 7574 -19060 7580 -19057
rect 7970 -19057 8016 -19045
rect 7970 -19060 7976 -19057
rect 7574 -19175 7976 -19060
rect 8010 -19060 8016 -19057
rect 8498 -19057 8544 -19045
rect 8498 -19060 8504 -19057
rect 8010 -19175 8504 -19060
rect 8538 -19060 8544 -19057
rect 8606 -19057 8652 -19045
rect 8606 -19060 8612 -19057
rect 8538 -19175 8612 -19060
rect 8646 -19060 8652 -19057
rect 9134 -19057 9180 -19045
rect 9134 -19060 9140 -19057
rect 8646 -19175 9140 -19060
rect 9174 -19060 9180 -19057
rect 9570 -19057 9616 -19045
rect 9570 -19060 9576 -19057
rect 9174 -19175 9576 -19060
rect 9610 -19060 9616 -19057
rect 10098 -19057 10144 -19045
rect 10098 -19060 10104 -19057
rect 9610 -19175 10104 -19060
rect 10138 -19060 10144 -19057
rect 10206 -19057 10252 -19045
rect 10206 -19060 10212 -19057
rect 10138 -19175 10212 -19060
rect 10246 -19060 10252 -19057
rect 10734 -19050 10780 -19045
rect 10734 -19057 10940 -19050
rect 10734 -19060 10740 -19057
rect 10246 -19175 10740 -19060
rect 10774 -19060 10940 -19057
rect 11170 -19057 11216 -19045
rect 11170 -19060 11176 -19057
rect 10774 -19175 10810 -19060
rect 1560 -19180 10810 -19175
rect 10930 -19175 11176 -19060
rect 11210 -19060 11216 -19057
rect 11400 -19060 11520 -19010
rect 11698 -19057 11744 -19045
rect 11698 -19060 11704 -19057
rect 11210 -19175 11704 -19060
rect 11738 -19060 11744 -19057
rect 11806 -19057 11852 -19045
rect 11806 -19060 11812 -19057
rect 11738 -19175 11812 -19060
rect 11846 -19060 11852 -19057
rect 12040 -19060 12160 -19010
rect 12334 -19057 12380 -19045
rect 12334 -19060 12340 -19057
rect 11846 -19175 12340 -19060
rect 12374 -19060 12380 -19057
rect 12770 -19057 12816 -19045
rect 12770 -19060 12776 -19057
rect 12374 -19175 12776 -19060
rect 12810 -19060 12816 -19057
rect 13298 -19057 13344 -19045
rect 13298 -19060 13304 -19057
rect 12810 -19175 13304 -19060
rect 13338 -19060 13344 -19057
rect 13406 -19057 13452 -19045
rect 13406 -19060 13412 -19057
rect 13338 -19175 13412 -19060
rect 13446 -19060 13452 -19057
rect 13934 -19057 13980 -19045
rect 13934 -19060 13940 -19057
rect 13446 -19175 13940 -19060
rect 13974 -19060 13980 -19057
rect 14370 -19057 14416 -19045
rect 14370 -19060 14376 -19057
rect 13974 -19175 14376 -19060
rect 14410 -19060 14416 -19057
rect 14898 -19057 14944 -19045
rect 14898 -19060 14904 -19057
rect 14410 -19175 14904 -19060
rect 14938 -19060 14944 -19057
rect 15006 -19057 15052 -19045
rect 15006 -19060 15012 -19057
rect 14938 -19175 15012 -19060
rect 15046 -19060 15052 -19057
rect 15534 -19057 15580 -19045
rect 15534 -19060 15540 -19057
rect 15046 -19175 15540 -19060
rect 15574 -19060 15580 -19057
rect 15970 -19057 16016 -19045
rect 15970 -19060 15976 -19057
rect 15574 -19175 15976 -19060
rect 16010 -19060 16016 -19057
rect 16498 -19057 16544 -19045
rect 16498 -19060 16504 -19057
rect 16010 -19175 16504 -19060
rect 16538 -19060 16544 -19057
rect 16606 -19057 16652 -19045
rect 16606 -19060 16612 -19057
rect 16538 -19175 16612 -19060
rect 16646 -19060 16652 -19057
rect 17134 -19057 17180 -19045
rect 17134 -19060 17140 -19057
rect 16646 -19175 17140 -19060
rect 17174 -19060 17180 -19057
rect 17570 -19057 17616 -19045
rect 17570 -19060 17576 -19057
rect 17174 -19175 17576 -19060
rect 17610 -19060 17616 -19057
rect 18098 -19057 18144 -19045
rect 18098 -19060 18104 -19057
rect 17610 -19175 18104 -19060
rect 18138 -19060 18144 -19057
rect 18206 -19057 18252 -19045
rect 18206 -19060 18212 -19057
rect 18138 -19175 18212 -19060
rect 18246 -19060 18252 -19057
rect 18734 -19057 18780 -19045
rect 18734 -19060 18740 -19057
rect 18246 -19175 18740 -19060
rect 18774 -19060 18780 -19057
rect 19170 -19057 19216 -19045
rect 19170 -19060 19176 -19057
rect 18774 -19175 19176 -19060
rect 19210 -19060 19216 -19057
rect 19698 -19057 19744 -19045
rect 19698 -19060 19704 -19057
rect 19210 -19175 19704 -19060
rect 19738 -19060 19744 -19057
rect 19806 -19057 19852 -19045
rect 19806 -19060 19812 -19057
rect 19738 -19175 19812 -19060
rect 19846 -19060 19852 -19057
rect 20334 -19057 20380 -19045
rect 20334 -19060 20340 -19057
rect 19846 -19175 20340 -19060
rect 20374 -19060 20380 -19057
rect 20770 -19057 20816 -19045
rect 20770 -19060 20776 -19057
rect 20374 -19175 20776 -19060
rect 20810 -19060 20816 -19057
rect 21298 -19057 21344 -19045
rect 21298 -19060 21304 -19057
rect 20810 -19175 21304 -19060
rect 21338 -19060 21344 -19057
rect 21406 -19057 21452 -19045
rect 21406 -19060 21412 -19057
rect 21338 -19175 21412 -19060
rect 21446 -19060 21452 -19057
rect 21934 -19057 21980 -19045
rect 21934 -19060 21940 -19057
rect 21446 -19175 21940 -19060
rect 21974 -19060 21980 -19057
rect 22370 -19057 22416 -19045
rect 22370 -19060 22376 -19057
rect 21974 -19175 22376 -19060
rect 22410 -19060 22416 -19057
rect 22898 -19057 22944 -19045
rect 22898 -19060 22904 -19057
rect 22410 -19175 22904 -19060
rect 22938 -19060 22944 -19057
rect 23006 -19057 23052 -19045
rect 23006 -19060 23012 -19057
rect 22938 -19175 23012 -19060
rect 23046 -19060 23052 -19057
rect 23534 -19057 23580 -19045
rect 23534 -19060 23540 -19057
rect 23046 -19175 23540 -19060
rect 23574 -19060 23580 -19057
rect 23970 -19057 24016 -19045
rect 23970 -19060 23976 -19057
rect 23574 -19175 23976 -19060
rect 24010 -19060 24016 -19057
rect 24498 -19057 24544 -19045
rect 24498 -19060 24504 -19057
rect 24010 -19175 24504 -19060
rect 24538 -19060 24544 -19057
rect 24606 -19057 24652 -19045
rect 24606 -19060 24612 -19057
rect 24538 -19175 24612 -19060
rect 24646 -19060 24652 -19057
rect 25134 -19057 25180 -19045
rect 25134 -19060 25140 -19057
rect 24646 -19175 25140 -19060
rect 25174 -19060 25180 -19057
rect 25570 -19057 25616 -19045
rect 25570 -19060 25576 -19057
rect 25174 -19175 25576 -19060
rect 25610 -19060 25616 -19057
rect 26098 -19057 26144 -19045
rect 26098 -19060 26104 -19057
rect 25610 -19175 26104 -19060
rect 26138 -19060 26144 -19057
rect 26206 -19057 26252 -19045
rect 26206 -19060 26212 -19057
rect 26138 -19175 26212 -19060
rect 26246 -19060 26252 -19057
rect 26734 -19057 26780 -19045
rect 26734 -19060 26740 -19057
rect 26246 -19175 26740 -19060
rect 26774 -19060 26780 -19057
rect 27170 -19057 27216 -19045
rect 27170 -19060 27176 -19057
rect 26774 -19175 27176 -19060
rect 27210 -19060 27216 -19057
rect 27698 -19057 27744 -19045
rect 27698 -19060 27704 -19057
rect 27210 -19175 27704 -19060
rect 27738 -19060 27744 -19057
rect 27806 -19057 27852 -19045
rect 27806 -19060 27812 -19057
rect 27738 -19175 27812 -19060
rect 27846 -19060 27852 -19057
rect 28334 -19057 28380 -19045
rect 28334 -19060 28340 -19057
rect 27846 -19175 28340 -19060
rect 28374 -19060 28380 -19057
rect 28770 -19057 28816 -19045
rect 28770 -19060 28776 -19057
rect 28374 -19175 28776 -19060
rect 28810 -19060 28816 -19057
rect 29298 -19057 29344 -19045
rect 29298 -19060 29304 -19057
rect 28810 -19175 29304 -19060
rect 29338 -19060 29344 -19057
rect 29406 -19057 29452 -19045
rect 29406 -19060 29412 -19057
rect 29338 -19175 29412 -19060
rect 29446 -19060 29452 -19057
rect 29934 -19057 29980 -19045
rect 29934 -19060 29940 -19057
rect 29446 -19175 29940 -19060
rect 29974 -19060 29980 -19057
rect 30370 -19057 30416 -19045
rect 30370 -19060 30376 -19057
rect 29974 -19175 30376 -19060
rect 30410 -19060 30416 -19057
rect 30898 -19057 30944 -19045
rect 30898 -19060 30904 -19057
rect 30410 -19175 30904 -19060
rect 30938 -19060 30944 -19057
rect 31006 -19057 31052 -19045
rect 31006 -19060 31012 -19057
rect 30938 -19175 31012 -19060
rect 31046 -19060 31052 -19057
rect 31534 -19057 31580 -19045
rect 31534 -19060 31540 -19057
rect 31046 -19175 31540 -19060
rect 31574 -19060 31580 -19057
rect 31970 -19057 32016 -19045
rect 31970 -19060 31976 -19057
rect 31574 -19175 31976 -19060
rect 32010 -19060 32016 -19057
rect 32498 -19057 32544 -19045
rect 32498 -19060 32504 -19057
rect 32010 -19175 32504 -19060
rect 32538 -19060 32544 -19057
rect 32606 -19057 32652 -19045
rect 32606 -19060 32612 -19057
rect 32538 -19175 32612 -19060
rect 32646 -19060 32652 -19057
rect 33134 -19057 33180 -19045
rect 33134 -19060 33140 -19057
rect 32646 -19175 33140 -19060
rect 33174 -19060 33180 -19057
rect 33570 -19057 33616 -19045
rect 33570 -19060 33576 -19057
rect 33174 -19175 33576 -19060
rect 33610 -19060 33616 -19057
rect 34098 -19057 34144 -19045
rect 34098 -19060 34104 -19057
rect 33610 -19175 34104 -19060
rect 34138 -19060 34144 -19057
rect 34206 -19057 34252 -19045
rect 34206 -19060 34212 -19057
rect 34138 -19175 34212 -19060
rect 34246 -19060 34252 -19057
rect 34734 -19057 34780 -19045
rect 34734 -19060 34740 -19057
rect 34246 -19175 34740 -19060
rect 34774 -19060 34780 -19057
rect 35170 -19057 35216 -19045
rect 35170 -19060 35176 -19057
rect 34774 -19175 35176 -19060
rect 35210 -19060 35216 -19057
rect 35698 -19057 35744 -19045
rect 35698 -19060 35704 -19057
rect 35210 -19175 35704 -19060
rect 35738 -19060 35744 -19057
rect 35806 -19057 35852 -19045
rect 35806 -19060 35812 -19057
rect 35738 -19175 35812 -19060
rect 35846 -19060 35852 -19057
rect 36334 -19057 36380 -19045
rect 36334 -19060 36340 -19057
rect 35846 -19175 36340 -19060
rect 36374 -19175 36380 -19057
rect 10930 -19180 36380 -19175
rect 1570 -19187 1616 -19180
rect 2098 -19187 2144 -19180
rect 2206 -19187 2252 -19180
rect 2734 -19187 2780 -19180
rect 3170 -19187 3216 -19180
rect 3698 -19187 3744 -19180
rect 3806 -19187 3852 -19180
rect 4334 -19187 4380 -19180
rect 4770 -19187 4816 -19180
rect 5298 -19187 5344 -19180
rect 5406 -19187 5452 -19180
rect 5934 -19187 5980 -19180
rect 6370 -19187 6416 -19180
rect 6898 -19187 6944 -19180
rect 7006 -19187 7052 -19180
rect 7534 -19187 7580 -19180
rect 7970 -19187 8016 -19180
rect 8498 -19187 8544 -19180
rect 8606 -19187 8652 -19180
rect 9134 -19187 9180 -19180
rect 9570 -19187 9616 -19180
rect 10098 -19187 10144 -19180
rect 10206 -19187 10252 -19180
rect 10734 -19187 10940 -19180
rect 11170 -19187 11216 -19180
rect 10750 -19190 10940 -19187
rect 11400 -19222 11520 -19180
rect 11698 -19187 11744 -19180
rect 11806 -19187 11852 -19180
rect 12040 -19222 12160 -19180
rect 12334 -19187 12380 -19180
rect 12770 -19187 12816 -19180
rect 13298 -19187 13344 -19180
rect 13406 -19187 13452 -19180
rect 13934 -19187 13980 -19180
rect 14370 -19187 14416 -19180
rect 14898 -19187 14944 -19180
rect 15006 -19187 15052 -19180
rect 15534 -19187 15580 -19180
rect 15970 -19187 16016 -19180
rect 16498 -19187 16544 -19180
rect 16606 -19187 16652 -19180
rect 17134 -19187 17180 -19180
rect 17570 -19187 17616 -19180
rect 18098 -19187 18144 -19180
rect 18206 -19187 18252 -19180
rect 18734 -19187 18780 -19180
rect 19170 -19187 19216 -19180
rect 19698 -19187 19744 -19180
rect 19806 -19187 19852 -19180
rect 20334 -19187 20380 -19180
rect 20770 -19187 20816 -19180
rect 21298 -19187 21344 -19180
rect 21406 -19187 21452 -19180
rect 21934 -19187 21980 -19180
rect 22370 -19187 22416 -19180
rect 22898 -19187 22944 -19180
rect 23006 -19187 23052 -19180
rect 23534 -19187 23580 -19180
rect 23970 -19187 24016 -19180
rect 24498 -19187 24544 -19180
rect 24606 -19187 24652 -19180
rect 25134 -19187 25180 -19180
rect 25570 -19187 25616 -19180
rect 26098 -19187 26144 -19180
rect 26206 -19187 26252 -19180
rect 26734 -19187 26780 -19180
rect 27170 -19187 27216 -19180
rect 27698 -19187 27744 -19180
rect 27806 -19187 27852 -19180
rect 28334 -19187 28380 -19180
rect 28770 -19187 28816 -19180
rect 29298 -19187 29344 -19180
rect 29406 -19187 29452 -19180
rect 29934 -19187 29980 -19180
rect 30370 -19187 30416 -19180
rect 30898 -19187 30944 -19180
rect 31006 -19187 31052 -19180
rect 31534 -19187 31580 -19180
rect 31970 -19187 32016 -19180
rect 32498 -19187 32544 -19180
rect 32606 -19187 32652 -19180
rect 33134 -19187 33180 -19180
rect 33570 -19187 33616 -19180
rect 34098 -19187 34144 -19180
rect 34206 -19187 34252 -19180
rect 34734 -19187 34780 -19180
rect 35170 -19187 35216 -19180
rect 35698 -19187 35744 -19180
rect 35806 -19187 35852 -19180
rect 36334 -19187 36380 -19180
rect 36770 -19057 36816 -19045
rect 36770 -19175 36776 -19057
rect 36810 -19175 36816 -19057
rect 36770 -19187 36816 -19175
rect 37298 -19057 37344 -19045
rect 37298 -19175 37304 -19057
rect 37338 -19175 37344 -19057
rect 37298 -19187 37344 -19175
rect 37406 -19057 37452 -19045
rect 37406 -19175 37412 -19057
rect 37446 -19175 37452 -19057
rect 37406 -19187 37452 -19175
rect 37934 -19057 37980 -19045
rect 37934 -19175 37940 -19057
rect 37974 -19175 37980 -19057
rect 37934 -19187 37980 -19175
rect 670 -19228 1093 -19222
rect 670 -19262 705 -19228
rect 1081 -19262 1093 -19228
rect 670 -19268 1093 -19262
rect 1657 -19228 2057 -19222
rect 1657 -19262 1669 -19228
rect 2045 -19230 2057 -19228
rect 2293 -19228 2693 -19222
rect 2293 -19230 2305 -19228
rect 2045 -19262 2060 -19230
rect 1657 -19268 2060 -19262
rect 670 -19490 720 -19268
rect 1420 -19310 1560 -19300
rect 1420 -19430 1430 -19310
rect 1550 -19320 1560 -19310
rect 1660 -19320 2060 -19268
rect 2290 -19262 2305 -19230
rect 2681 -19262 2693 -19228
rect 2290 -19268 2693 -19262
rect 3257 -19228 3657 -19222
rect 3257 -19262 3269 -19228
rect 3645 -19230 3657 -19228
rect 3893 -19228 4293 -19222
rect 3893 -19230 3905 -19228
rect 3645 -19262 3660 -19230
rect 3257 -19268 3660 -19262
rect 2290 -19320 2690 -19268
rect 3020 -19310 3160 -19300
rect 3020 -19320 3030 -19310
rect 1550 -19420 3030 -19320
rect 1550 -19430 1560 -19420
rect 1420 -19440 1560 -19430
rect 1660 -19440 2690 -19420
rect 3020 -19430 3030 -19420
rect 3150 -19320 3160 -19310
rect 3260 -19320 3660 -19268
rect 3890 -19262 3905 -19230
rect 4281 -19262 4293 -19228
rect 3890 -19268 4293 -19262
rect 4857 -19228 5257 -19222
rect 4857 -19262 4869 -19228
rect 5245 -19230 5257 -19228
rect 5493 -19228 5893 -19222
rect 5493 -19230 5505 -19228
rect 5245 -19262 5260 -19230
rect 4857 -19268 5260 -19262
rect 3890 -19320 4290 -19268
rect 4620 -19310 4760 -19300
rect 4620 -19320 4630 -19310
rect 3150 -19420 4630 -19320
rect 3150 -19430 3160 -19420
rect 3020 -19440 3160 -19430
rect 3260 -19440 4290 -19420
rect 4620 -19430 4630 -19420
rect 4750 -19320 4760 -19310
rect 4860 -19320 5260 -19268
rect 5490 -19262 5505 -19230
rect 5881 -19262 5893 -19228
rect 5490 -19268 5893 -19262
rect 6457 -19228 6857 -19222
rect 6457 -19262 6469 -19228
rect 6845 -19230 6857 -19228
rect 7093 -19228 7493 -19222
rect 7093 -19230 7105 -19228
rect 6845 -19262 6860 -19230
rect 6457 -19268 6860 -19262
rect 5490 -19320 5890 -19268
rect 6220 -19310 6360 -19300
rect 6220 -19320 6230 -19310
rect 4750 -19420 6230 -19320
rect 4750 -19430 4760 -19420
rect 4620 -19440 4760 -19430
rect 4860 -19440 5890 -19420
rect 6220 -19430 6230 -19420
rect 6350 -19320 6360 -19310
rect 6460 -19320 6860 -19268
rect 7090 -19262 7105 -19230
rect 7481 -19262 7493 -19228
rect 7090 -19268 7493 -19262
rect 8057 -19228 8457 -19222
rect 8057 -19262 8069 -19228
rect 8445 -19230 8457 -19228
rect 8693 -19228 9093 -19222
rect 8693 -19230 8705 -19228
rect 8445 -19262 8460 -19230
rect 8057 -19268 8460 -19262
rect 7090 -19320 7490 -19268
rect 7820 -19310 7960 -19300
rect 7820 -19320 7830 -19310
rect 6350 -19420 7830 -19320
rect 6350 -19430 6360 -19420
rect 6220 -19440 6360 -19430
rect 6460 -19440 7490 -19420
rect 7820 -19430 7830 -19420
rect 7950 -19320 7960 -19310
rect 8060 -19320 8460 -19268
rect 8690 -19262 8705 -19230
rect 9081 -19262 9093 -19228
rect 8690 -19268 9093 -19262
rect 9657 -19228 10057 -19222
rect 9657 -19262 9669 -19228
rect 10045 -19230 10057 -19228
rect 10293 -19228 10693 -19222
rect 10293 -19230 10305 -19228
rect 10045 -19262 10060 -19230
rect 9657 -19268 10060 -19262
rect 8690 -19320 9090 -19268
rect 9420 -19310 9560 -19300
rect 9420 -19320 9430 -19310
rect 7950 -19420 9430 -19320
rect 7950 -19430 7960 -19420
rect 7820 -19440 7960 -19430
rect 8060 -19440 9090 -19420
rect 9420 -19430 9430 -19420
rect 9550 -19320 9560 -19310
rect 9660 -19320 10060 -19268
rect 10290 -19262 10305 -19230
rect 10681 -19262 10693 -19228
rect 10290 -19268 10693 -19262
rect 11257 -19228 11657 -19222
rect 11257 -19262 11269 -19228
rect 11645 -19262 11657 -19228
rect 11257 -19268 11657 -19262
rect 11893 -19228 12293 -19222
rect 11893 -19262 11905 -19228
rect 12281 -19262 12293 -19228
rect 11893 -19268 12293 -19262
rect 12857 -19228 13257 -19222
rect 12857 -19262 12869 -19228
rect 13245 -19230 13257 -19228
rect 13493 -19228 13893 -19222
rect 13493 -19230 13505 -19228
rect 13245 -19262 13260 -19230
rect 12857 -19268 13260 -19262
rect 10290 -19320 10690 -19268
rect 9550 -19420 10690 -19320
rect 9550 -19430 9560 -19420
rect 9420 -19440 9560 -19430
rect 9660 -19440 10690 -19420
rect 1660 -19490 2060 -19440
rect 670 -19496 1093 -19490
rect 670 -19530 705 -19496
rect 1081 -19530 1093 -19496
rect 670 -19536 1093 -19530
rect 1657 -19496 2060 -19490
rect 1657 -19530 1669 -19496
rect 2045 -19530 2060 -19496
rect 2290 -19490 2690 -19440
rect 3260 -19490 3660 -19440
rect 2290 -19496 2693 -19490
rect 2290 -19530 2305 -19496
rect 2681 -19530 2693 -19496
rect 1657 -19536 2057 -19530
rect 2293 -19536 2693 -19530
rect 3257 -19496 3660 -19490
rect 3257 -19530 3269 -19496
rect 3645 -19530 3660 -19496
rect 3890 -19490 4290 -19440
rect 4860 -19490 5260 -19440
rect 3890 -19496 4293 -19490
rect 3890 -19530 3905 -19496
rect 4281 -19530 4293 -19496
rect 3257 -19536 3657 -19530
rect 3893 -19536 4293 -19530
rect 4857 -19496 5260 -19490
rect 4857 -19530 4869 -19496
rect 5245 -19530 5260 -19496
rect 5490 -19490 5890 -19440
rect 6460 -19490 6860 -19440
rect 5490 -19496 5893 -19490
rect 5490 -19530 5505 -19496
rect 5881 -19530 5893 -19496
rect 4857 -19536 5257 -19530
rect 5493 -19536 5893 -19530
rect 6457 -19496 6860 -19490
rect 6457 -19530 6469 -19496
rect 6845 -19530 6860 -19496
rect 7090 -19490 7490 -19440
rect 8060 -19490 8460 -19440
rect 7090 -19496 7493 -19490
rect 7090 -19530 7105 -19496
rect 7481 -19530 7493 -19496
rect 6457 -19536 6857 -19530
rect 7093 -19536 7493 -19530
rect 8057 -19496 8460 -19490
rect 8057 -19530 8069 -19496
rect 8445 -19530 8460 -19496
rect 8690 -19490 9090 -19440
rect 9660 -19490 10060 -19440
rect 8690 -19496 9093 -19490
rect 8690 -19530 8705 -19496
rect 9081 -19530 9093 -19496
rect 8057 -19536 8457 -19530
rect 8693 -19536 9093 -19530
rect 9657 -19496 10060 -19490
rect 9657 -19530 9669 -19496
rect 10045 -19530 10060 -19496
rect 10290 -19490 10690 -19440
rect 12860 -19320 13260 -19268
rect 13490 -19262 13505 -19230
rect 13881 -19262 13893 -19228
rect 13490 -19268 13893 -19262
rect 14457 -19228 14857 -19222
rect 14457 -19262 14469 -19228
rect 14845 -19230 14857 -19228
rect 15093 -19228 15493 -19222
rect 15093 -19230 15105 -19228
rect 14845 -19262 14860 -19230
rect 14457 -19268 14860 -19262
rect 13490 -19320 13890 -19268
rect 14460 -19320 14860 -19268
rect 15090 -19262 15105 -19230
rect 15481 -19262 15493 -19228
rect 15090 -19268 15493 -19262
rect 16057 -19228 16457 -19222
rect 16057 -19262 16069 -19228
rect 16445 -19262 16457 -19228
rect 16057 -19268 16457 -19262
rect 16693 -19228 17093 -19222
rect 16693 -19262 16705 -19228
rect 17081 -19262 17093 -19228
rect 16693 -19268 17093 -19262
rect 17657 -19228 18057 -19222
rect 17657 -19262 17669 -19228
rect 18045 -19262 18057 -19228
rect 17657 -19268 18057 -19262
rect 18293 -19228 18693 -19222
rect 18293 -19262 18305 -19228
rect 18681 -19262 18693 -19228
rect 18293 -19268 18693 -19262
rect 19257 -19228 19657 -19222
rect 19257 -19262 19269 -19228
rect 19645 -19262 19657 -19228
rect 19257 -19268 19657 -19262
rect 19893 -19228 20293 -19222
rect 19893 -19262 19905 -19228
rect 20281 -19262 20293 -19228
rect 19893 -19268 20293 -19262
rect 20857 -19228 21257 -19222
rect 20857 -19262 20869 -19228
rect 21245 -19262 21257 -19228
rect 20857 -19268 21257 -19262
rect 21493 -19228 21893 -19222
rect 21493 -19262 21505 -19228
rect 21881 -19262 21893 -19228
rect 21493 -19268 21893 -19262
rect 22457 -19228 22857 -19222
rect 22457 -19262 22469 -19228
rect 22845 -19262 22857 -19228
rect 22457 -19268 22857 -19262
rect 23093 -19228 23493 -19222
rect 23093 -19262 23105 -19228
rect 23481 -19262 23493 -19228
rect 23093 -19268 23493 -19262
rect 24057 -19228 24457 -19222
rect 24057 -19262 24069 -19228
rect 24445 -19262 24457 -19228
rect 24057 -19268 24457 -19262
rect 24693 -19228 25093 -19222
rect 24693 -19262 24705 -19228
rect 25081 -19262 25093 -19228
rect 24693 -19268 25093 -19262
rect 25657 -19228 26057 -19222
rect 25657 -19262 25669 -19228
rect 26045 -19262 26057 -19228
rect 25657 -19268 26057 -19262
rect 26293 -19228 26693 -19222
rect 26293 -19262 26305 -19228
rect 26681 -19262 26693 -19228
rect 26293 -19268 26693 -19262
rect 27257 -19228 27657 -19222
rect 27257 -19262 27269 -19228
rect 27645 -19262 27657 -19228
rect 27257 -19268 27657 -19262
rect 27893 -19228 28293 -19222
rect 27893 -19262 27905 -19228
rect 28281 -19262 28293 -19228
rect 27893 -19268 28293 -19262
rect 28857 -19228 29257 -19222
rect 28857 -19262 28869 -19228
rect 29245 -19262 29257 -19228
rect 28857 -19268 29257 -19262
rect 29493 -19228 29893 -19222
rect 29493 -19262 29505 -19228
rect 29881 -19262 29893 -19228
rect 29493 -19268 29893 -19262
rect 30457 -19228 30857 -19222
rect 30457 -19262 30469 -19228
rect 30845 -19262 30857 -19228
rect 30457 -19268 30857 -19262
rect 31093 -19228 31493 -19222
rect 31093 -19262 31105 -19228
rect 31481 -19262 31493 -19228
rect 32057 -19228 32457 -19222
rect 31093 -19268 31493 -19262
rect 31740 -19240 31820 -19230
rect 15090 -19320 15490 -19268
rect 12860 -19440 15490 -19320
rect 12860 -19490 13260 -19440
rect 10290 -19496 10693 -19490
rect 10290 -19530 10305 -19496
rect 10681 -19530 10693 -19496
rect 9657 -19536 10057 -19530
rect 10293 -19536 10693 -19530
rect 11257 -19496 11657 -19490
rect 11257 -19530 11269 -19496
rect 11645 -19530 11657 -19496
rect 11257 -19536 11657 -19530
rect 11893 -19496 12293 -19490
rect 11893 -19530 11905 -19496
rect 12281 -19530 12293 -19496
rect 11893 -19536 12293 -19530
rect 12857 -19496 13260 -19490
rect 12857 -19530 12869 -19496
rect 13245 -19530 13260 -19496
rect 13490 -19490 13890 -19440
rect 14460 -19490 14860 -19440
rect 13490 -19496 13893 -19490
rect 13490 -19530 13505 -19496
rect 13881 -19530 13893 -19496
rect 12857 -19536 13257 -19530
rect 13493 -19536 13893 -19530
rect 14457 -19496 14860 -19490
rect 14457 -19530 14469 -19496
rect 14845 -19530 14860 -19496
rect 15090 -19490 15490 -19440
rect 15600 -19320 15740 -19310
rect 15600 -19440 15610 -19320
rect 15730 -19330 15740 -19320
rect 16060 -19330 16450 -19268
rect 16700 -19330 17090 -19268
rect 15730 -19430 17090 -19330
rect 15730 -19440 15740 -19430
rect 15600 -19450 15740 -19440
rect 16060 -19490 16450 -19430
rect 16700 -19490 17090 -19430
rect 17200 -19320 17340 -19310
rect 17200 -19440 17210 -19320
rect 17330 -19330 17340 -19320
rect 17660 -19330 18050 -19268
rect 18300 -19330 18690 -19268
rect 17330 -19430 18690 -19330
rect 17330 -19440 17340 -19430
rect 17200 -19450 17340 -19440
rect 17660 -19490 18050 -19430
rect 18300 -19490 18690 -19430
rect 18800 -19320 18940 -19310
rect 18800 -19440 18810 -19320
rect 18930 -19330 18940 -19320
rect 19260 -19330 19650 -19268
rect 19900 -19330 20290 -19268
rect 18930 -19430 20290 -19330
rect 18930 -19440 18940 -19430
rect 18800 -19450 18940 -19440
rect 19260 -19490 19650 -19430
rect 19900 -19490 20290 -19430
rect 20400 -19320 20540 -19310
rect 20400 -19440 20410 -19320
rect 20530 -19330 20540 -19320
rect 20860 -19330 21250 -19268
rect 21500 -19330 21890 -19268
rect 20530 -19430 21890 -19330
rect 20530 -19440 20540 -19430
rect 20400 -19450 20540 -19440
rect 20860 -19490 21250 -19430
rect 21500 -19490 21890 -19430
rect 22000 -19320 22140 -19310
rect 22000 -19440 22010 -19320
rect 22130 -19330 22140 -19320
rect 22460 -19330 22850 -19268
rect 23100 -19330 23490 -19268
rect 22130 -19430 23490 -19330
rect 22130 -19440 22140 -19430
rect 22000 -19450 22140 -19440
rect 22460 -19490 22850 -19430
rect 23100 -19490 23490 -19430
rect 23600 -19320 23740 -19310
rect 23600 -19440 23610 -19320
rect 23730 -19330 23740 -19320
rect 24060 -19330 24450 -19268
rect 24700 -19330 25090 -19268
rect 23730 -19430 25090 -19330
rect 23730 -19440 23740 -19430
rect 23600 -19450 23740 -19440
rect 24060 -19490 24450 -19430
rect 24700 -19490 25090 -19430
rect 25660 -19330 26050 -19268
rect 26300 -19330 26690 -19268
rect 26800 -19320 26940 -19310
rect 26800 -19330 26810 -19320
rect 25660 -19430 26810 -19330
rect 25660 -19490 26050 -19430
rect 26300 -19490 26690 -19430
rect 26800 -19440 26810 -19430
rect 26930 -19330 26940 -19320
rect 27260 -19330 27650 -19268
rect 27900 -19330 28290 -19268
rect 26930 -19430 28290 -19330
rect 26930 -19440 26940 -19430
rect 26800 -19450 26940 -19440
rect 27260 -19490 27650 -19430
rect 27900 -19490 28290 -19430
rect 28400 -19320 28540 -19310
rect 28400 -19440 28410 -19320
rect 28530 -19330 28540 -19320
rect 28860 -19330 29250 -19268
rect 29500 -19330 29890 -19268
rect 30460 -19330 30850 -19268
rect 31100 -19330 31490 -19268
rect 28530 -19430 31490 -19330
rect 28530 -19440 28540 -19430
rect 28400 -19450 28540 -19440
rect 28860 -19490 29250 -19430
rect 29500 -19490 29890 -19430
rect 30460 -19490 30850 -19430
rect 31100 -19490 31490 -19430
rect 15090 -19496 15493 -19490
rect 15090 -19530 15105 -19496
rect 15481 -19530 15493 -19496
rect 14457 -19536 14857 -19530
rect 15093 -19536 15493 -19530
rect 16057 -19496 16457 -19490
rect 16057 -19530 16069 -19496
rect 16445 -19530 16457 -19496
rect 16057 -19536 16457 -19530
rect 16693 -19496 17093 -19490
rect 16693 -19530 16705 -19496
rect 17081 -19530 17093 -19496
rect 16693 -19536 17093 -19530
rect 17657 -19496 18057 -19490
rect 17657 -19530 17669 -19496
rect 18045 -19530 18057 -19496
rect 17657 -19536 18057 -19530
rect 18293 -19496 18693 -19490
rect 18293 -19530 18305 -19496
rect 18681 -19530 18693 -19496
rect 18293 -19536 18693 -19530
rect 19257 -19496 19657 -19490
rect 19257 -19530 19269 -19496
rect 19645 -19530 19657 -19496
rect 19257 -19536 19657 -19530
rect 19893 -19496 20293 -19490
rect 19893 -19530 19905 -19496
rect 20281 -19530 20293 -19496
rect 19893 -19536 20293 -19530
rect 20857 -19496 21257 -19490
rect 20857 -19530 20869 -19496
rect 21245 -19530 21257 -19496
rect 20857 -19536 21257 -19530
rect 21493 -19496 21893 -19490
rect 21493 -19530 21505 -19496
rect 21881 -19530 21893 -19496
rect 21493 -19536 21893 -19530
rect 22457 -19496 22857 -19490
rect 22457 -19530 22469 -19496
rect 22845 -19530 22857 -19496
rect 22457 -19536 22857 -19530
rect 23093 -19496 23493 -19490
rect 23093 -19530 23105 -19496
rect 23481 -19530 23493 -19496
rect 23093 -19536 23493 -19530
rect 24057 -19496 24457 -19490
rect 24057 -19530 24069 -19496
rect 24445 -19530 24457 -19496
rect 24057 -19536 24457 -19530
rect 24693 -19496 25093 -19490
rect 24693 -19530 24705 -19496
rect 25081 -19530 25093 -19496
rect 24693 -19536 25093 -19530
rect 25657 -19496 26057 -19490
rect 25657 -19530 25669 -19496
rect 26045 -19530 26057 -19496
rect 25657 -19536 26057 -19530
rect 26293 -19496 26693 -19490
rect 26293 -19530 26305 -19496
rect 26681 -19530 26693 -19496
rect 26293 -19536 26693 -19530
rect 27257 -19496 27657 -19490
rect 27257 -19530 27269 -19496
rect 27645 -19530 27657 -19496
rect 27257 -19536 27657 -19530
rect 27893 -19496 28293 -19490
rect 27893 -19530 27905 -19496
rect 28281 -19530 28293 -19496
rect 27893 -19536 28293 -19530
rect 28857 -19496 29257 -19490
rect 28857 -19530 28869 -19496
rect 29245 -19530 29257 -19496
rect 28857 -19536 29257 -19530
rect 29493 -19496 29893 -19490
rect 29493 -19530 29505 -19496
rect 29881 -19530 29893 -19496
rect 29493 -19536 29893 -19530
rect 30457 -19496 30857 -19490
rect 30457 -19530 30469 -19496
rect 30845 -19530 30857 -19496
rect 30457 -19536 30857 -19530
rect 31093 -19496 31493 -19490
rect 31093 -19530 31105 -19496
rect 31481 -19530 31493 -19496
rect 31740 -19520 31750 -19240
rect 31810 -19330 31820 -19240
rect 32057 -19262 32069 -19228
rect 32445 -19262 32457 -19228
rect 32057 -19268 32457 -19262
rect 32693 -19228 33093 -19222
rect 32693 -19262 32705 -19228
rect 33081 -19262 33093 -19228
rect 32693 -19268 33093 -19262
rect 33657 -19228 34057 -19222
rect 33657 -19262 33669 -19228
rect 34045 -19262 34057 -19228
rect 33657 -19268 34057 -19262
rect 34293 -19228 34693 -19222
rect 34293 -19262 34305 -19228
rect 34681 -19262 34693 -19228
rect 34293 -19268 34693 -19262
rect 35257 -19228 35657 -19222
rect 35257 -19262 35269 -19228
rect 35645 -19262 35657 -19228
rect 35257 -19268 35657 -19262
rect 35893 -19228 36293 -19222
rect 35893 -19262 35905 -19228
rect 36281 -19262 36293 -19228
rect 35893 -19268 36293 -19262
rect 36857 -19228 37257 -19222
rect 36857 -19262 36869 -19228
rect 37245 -19262 37257 -19228
rect 36857 -19268 37257 -19262
rect 37493 -19228 37893 -19222
rect 37493 -19262 37505 -19228
rect 37881 -19262 37893 -19228
rect 37493 -19268 37893 -19262
rect 32060 -19330 32450 -19268
rect 32700 -19330 33090 -19268
rect 33660 -19330 34050 -19268
rect 34300 -19330 34690 -19268
rect 35260 -19330 35650 -19268
rect 35900 -19330 36290 -19268
rect 31810 -19430 36290 -19330
rect 31810 -19520 31820 -19430
rect 32060 -19490 32450 -19430
rect 32700 -19490 33090 -19430
rect 33660 -19490 34050 -19430
rect 34300 -19490 34690 -19430
rect 35260 -19490 35650 -19430
rect 35900 -19490 36290 -19430
rect 31740 -19530 31820 -19520
rect 32057 -19496 32457 -19490
rect 32057 -19530 32069 -19496
rect 32445 -19530 32457 -19496
rect 31093 -19536 31493 -19530
rect 32057 -19536 32457 -19530
rect 32693 -19496 33093 -19490
rect 32693 -19530 32705 -19496
rect 33081 -19530 33093 -19496
rect 32693 -19536 33093 -19530
rect 33657 -19496 34057 -19490
rect 33657 -19530 33669 -19496
rect 34045 -19530 34057 -19496
rect 33657 -19536 34057 -19530
rect 34293 -19496 34693 -19490
rect 34293 -19530 34305 -19496
rect 34681 -19530 34693 -19496
rect 34293 -19536 34693 -19530
rect 35257 -19496 35657 -19490
rect 35257 -19530 35269 -19496
rect 35645 -19530 35657 -19496
rect 35257 -19536 35657 -19530
rect 35893 -19496 36293 -19490
rect 35893 -19530 35905 -19496
rect 36281 -19530 36293 -19496
rect 35893 -19536 36293 -19530
rect 36857 -19496 37257 -19490
rect 36857 -19530 36869 -19496
rect 37245 -19530 37257 -19496
rect 36857 -19536 37257 -19530
rect 37493 -19496 37893 -19490
rect 37493 -19530 37505 -19496
rect 37881 -19530 37893 -19496
rect 37493 -19536 37893 -19530
rect 57 -20354 490 -20348
rect 57 -20380 69 -20354
rect 0 -20388 69 -20380
rect 445 -20388 490 -20354
rect 0 -20488 490 -20388
rect 670 -20348 720 -19536
rect 1134 -19596 1180 -19584
rect 1134 -20288 1140 -19596
rect 1174 -20288 1180 -19596
rect 1134 -20300 1180 -20288
rect 1570 -19596 1616 -19584
rect 1570 -20288 1576 -19596
rect 1610 -20288 1616 -19596
rect 1570 -20300 1616 -20288
rect 2098 -19596 2144 -19584
rect 2098 -20288 2104 -19596
rect 2138 -19600 2144 -19596
rect 2206 -19596 2252 -19584
rect 2206 -19600 2212 -19596
rect 2138 -19610 2212 -19600
rect 2138 -20288 2144 -20270
rect 2098 -20300 2144 -20288
rect 2206 -20288 2212 -20270
rect 2246 -20288 2252 -19596
rect 2206 -20300 2252 -20288
rect 2734 -19596 2780 -19584
rect 2734 -20288 2740 -19596
rect 2774 -20288 2780 -19596
rect 2734 -20300 2780 -20288
rect 3170 -19596 3216 -19584
rect 3170 -20288 3176 -19596
rect 3210 -20288 3216 -19596
rect 3170 -20300 3216 -20288
rect 3698 -19596 3744 -19584
rect 3698 -20288 3704 -19596
rect 3738 -19600 3744 -19596
rect 3806 -19596 3852 -19584
rect 3806 -19600 3812 -19596
rect 3738 -19610 3812 -19600
rect 3738 -20288 3744 -20270
rect 3698 -20300 3744 -20288
rect 3806 -20288 3812 -20270
rect 3846 -20288 3852 -19596
rect 3806 -20300 3852 -20288
rect 4334 -19596 4380 -19584
rect 4334 -20288 4340 -19596
rect 4374 -20288 4380 -19596
rect 4334 -20300 4380 -20288
rect 4770 -19596 4816 -19584
rect 4770 -20288 4776 -19596
rect 4810 -20288 4816 -19596
rect 4770 -20300 4816 -20288
rect 5298 -19596 5344 -19584
rect 5298 -20288 5304 -19596
rect 5338 -19600 5344 -19596
rect 5406 -19596 5452 -19584
rect 5406 -19600 5412 -19596
rect 5338 -19610 5412 -19600
rect 5338 -20288 5344 -20270
rect 5298 -20300 5344 -20288
rect 5406 -20288 5412 -20270
rect 5446 -20288 5452 -19596
rect 5406 -20300 5452 -20288
rect 5934 -19596 5980 -19584
rect 5934 -20288 5940 -19596
rect 5974 -20288 5980 -19596
rect 5934 -20300 5980 -20288
rect 6370 -19596 6416 -19584
rect 6370 -20288 6376 -19596
rect 6410 -20288 6416 -19596
rect 6370 -20300 6416 -20288
rect 6898 -19596 6944 -19584
rect 6898 -20288 6904 -19596
rect 6938 -19600 6944 -19596
rect 7006 -19596 7052 -19584
rect 7006 -19600 7012 -19596
rect 6938 -19610 7012 -19600
rect 6938 -20288 6944 -20270
rect 6898 -20300 6944 -20288
rect 7006 -20288 7012 -20270
rect 7046 -20288 7052 -19596
rect 7006 -20300 7052 -20288
rect 7534 -19596 7580 -19584
rect 7534 -20288 7540 -19596
rect 7574 -20288 7580 -19596
rect 7534 -20300 7580 -20288
rect 7970 -19596 8016 -19584
rect 7970 -20288 7976 -19596
rect 8010 -20288 8016 -19596
rect 7970 -20300 8016 -20288
rect 8498 -19596 8544 -19584
rect 8498 -20288 8504 -19596
rect 8538 -19600 8544 -19596
rect 8606 -19596 8652 -19584
rect 8606 -19600 8612 -19596
rect 8538 -19610 8612 -19600
rect 8538 -20280 8612 -20270
rect 8538 -20288 8544 -20280
rect 8498 -20300 8544 -20288
rect 8606 -20288 8612 -20280
rect 8646 -20288 8652 -19596
rect 8606 -20300 8652 -20288
rect 9134 -19596 9180 -19584
rect 9134 -20288 9140 -19596
rect 9174 -20288 9180 -19596
rect 9134 -20300 9180 -20288
rect 9570 -19596 9616 -19584
rect 9570 -20288 9576 -19596
rect 9610 -20288 9616 -19596
rect 9570 -20300 9616 -20288
rect 10098 -19596 10144 -19584
rect 10098 -20288 10104 -19596
rect 10138 -19600 10144 -19596
rect 10206 -19596 10252 -19584
rect 10206 -19600 10212 -19596
rect 10138 -19610 10212 -19600
rect 10138 -20280 10212 -20270
rect 10138 -20288 10144 -20280
rect 10098 -20300 10144 -20288
rect 10206 -20288 10212 -20280
rect 10246 -20288 10252 -19596
rect 10206 -20300 10252 -20288
rect 10734 -19596 10780 -19584
rect 10734 -20288 10740 -19596
rect 10774 -20288 10780 -19596
rect 10734 -20300 10780 -20288
rect 11170 -19596 11216 -19584
rect 11170 -20288 11176 -19596
rect 11210 -19840 11216 -19596
rect 11370 -19840 11510 -19536
rect 11698 -19596 11744 -19584
rect 11698 -19840 11704 -19596
rect 11210 -20030 11704 -19840
rect 11210 -20288 11216 -20030
rect 11170 -20300 11216 -20288
rect 11370 -20348 11510 -20030
rect 11698 -20288 11704 -20030
rect 11738 -19840 11744 -19596
rect 11806 -19596 11852 -19584
rect 11806 -19840 11812 -19596
rect 11738 -20030 11812 -19840
rect 11738 -20288 11744 -20030
rect 11698 -20300 11744 -20288
rect 11806 -20288 11812 -20030
rect 11846 -19840 11852 -19596
rect 12030 -19840 12140 -19536
rect 12334 -19596 12380 -19584
rect 12334 -19840 12340 -19596
rect 11846 -20030 12340 -19840
rect 11846 -20288 11852 -20030
rect 11806 -20300 11852 -20288
rect 12030 -20348 12140 -20030
rect 12334 -20288 12340 -20030
rect 12374 -20288 12380 -19596
rect 12334 -20300 12380 -20288
rect 12770 -19596 12816 -19584
rect 12770 -20288 12776 -19596
rect 12810 -20288 12816 -19596
rect 12770 -20300 12816 -20288
rect 13298 -19596 13344 -19584
rect 13298 -20288 13304 -19596
rect 13338 -19600 13344 -19596
rect 13406 -19596 13452 -19584
rect 13406 -19600 13412 -19596
rect 13338 -19610 13412 -19600
rect 13338 -20280 13412 -20270
rect 13338 -20288 13344 -20280
rect 13298 -20300 13344 -20288
rect 13406 -20288 13412 -20280
rect 13446 -20288 13452 -19596
rect 13406 -20300 13452 -20288
rect 13934 -19596 13980 -19584
rect 13934 -20288 13940 -19596
rect 13974 -20288 13980 -19596
rect 13934 -20300 13980 -20288
rect 14370 -19596 14416 -19584
rect 14370 -20288 14376 -19596
rect 14410 -20288 14416 -19596
rect 14370 -20300 14416 -20288
rect 14898 -19596 14944 -19584
rect 14898 -20288 14904 -19596
rect 14938 -19600 14944 -19596
rect 15006 -19596 15052 -19584
rect 15006 -19600 15012 -19596
rect 14938 -19610 15012 -19600
rect 14938 -20280 15012 -20270
rect 14938 -20288 14944 -20280
rect 14898 -20300 14944 -20288
rect 15006 -20288 15012 -20280
rect 15046 -20288 15052 -19596
rect 15006 -20300 15052 -20288
rect 15534 -19596 15580 -19584
rect 15534 -20288 15540 -19596
rect 15574 -20288 15580 -19596
rect 15534 -20300 15580 -20288
rect 15970 -19596 16016 -19584
rect 15970 -20288 15976 -19596
rect 16010 -20288 16016 -19596
rect 15970 -20300 16016 -20288
rect 16498 -19590 16544 -19584
rect 16606 -19590 16652 -19584
rect 16498 -19596 16652 -19590
rect 16498 -20288 16504 -19596
rect 16538 -19600 16612 -19596
rect 16538 -20288 16612 -20280
rect 16646 -20288 16652 -19596
rect 16498 -20290 16652 -20288
rect 16498 -20300 16544 -20290
rect 16606 -20300 16652 -20290
rect 17134 -19596 17180 -19584
rect 17134 -20288 17140 -19596
rect 17174 -20288 17180 -19596
rect 17134 -20300 17180 -20288
rect 17570 -19596 17616 -19584
rect 17570 -20288 17576 -19596
rect 17610 -20288 17616 -19596
rect 17570 -20300 17616 -20288
rect 18098 -19590 18144 -19584
rect 18206 -19590 18252 -19584
rect 18098 -19596 18252 -19590
rect 18098 -20288 18104 -19596
rect 18138 -19600 18212 -19596
rect 18138 -20288 18212 -20280
rect 18246 -20288 18252 -19596
rect 18098 -20290 18252 -20288
rect 18098 -20300 18144 -20290
rect 18206 -20300 18252 -20290
rect 18734 -19596 18780 -19584
rect 18734 -20288 18740 -19596
rect 18774 -20288 18780 -19596
rect 18734 -20300 18780 -20288
rect 19170 -19596 19216 -19584
rect 19170 -20288 19176 -19596
rect 19210 -20288 19216 -19596
rect 19170 -20300 19216 -20288
rect 19698 -19590 19744 -19584
rect 19806 -19590 19852 -19584
rect 19698 -19596 19852 -19590
rect 19698 -20288 19704 -19596
rect 19738 -19600 19812 -19596
rect 19738 -20288 19812 -20280
rect 19846 -20288 19852 -19596
rect 19698 -20290 19852 -20288
rect 19698 -20300 19744 -20290
rect 19806 -20300 19852 -20290
rect 20334 -19596 20380 -19584
rect 20334 -20288 20340 -19596
rect 20374 -20288 20380 -19596
rect 20334 -20300 20380 -20288
rect 20770 -19596 20816 -19584
rect 20770 -20288 20776 -19596
rect 20810 -20288 20816 -19596
rect 20770 -20300 20816 -20288
rect 21298 -19590 21344 -19584
rect 21406 -19590 21452 -19584
rect 21298 -19596 21452 -19590
rect 21298 -20288 21304 -19596
rect 21338 -19600 21412 -19596
rect 21338 -20288 21412 -20280
rect 21446 -20288 21452 -19596
rect 21298 -20290 21452 -20288
rect 21298 -20300 21344 -20290
rect 21406 -20300 21452 -20290
rect 21934 -19596 21980 -19584
rect 21934 -20288 21940 -19596
rect 21974 -20288 21980 -19596
rect 21934 -20300 21980 -20288
rect 22370 -19596 22416 -19584
rect 22370 -20288 22376 -19596
rect 22410 -20288 22416 -19596
rect 22370 -20300 22416 -20288
rect 22898 -19590 22944 -19584
rect 23006 -19590 23052 -19584
rect 22898 -19596 23052 -19590
rect 22898 -20288 22904 -19596
rect 22938 -19600 23012 -19596
rect 22938 -20288 23012 -20280
rect 23046 -20288 23052 -19596
rect 22898 -20290 23052 -20288
rect 22898 -20300 22944 -20290
rect 23006 -20300 23052 -20290
rect 23534 -19596 23580 -19584
rect 23534 -20288 23540 -19596
rect 23574 -20288 23580 -19596
rect 23534 -20300 23580 -20288
rect 23970 -19596 24016 -19584
rect 23970 -20288 23976 -19596
rect 24010 -20288 24016 -19596
rect 23970 -20300 24016 -20288
rect 24498 -19590 24544 -19584
rect 24606 -19590 24652 -19584
rect 24498 -19596 24652 -19590
rect 24498 -20288 24504 -19596
rect 24538 -19600 24612 -19596
rect 24538 -20288 24612 -20280
rect 24646 -20288 24652 -19596
rect 24498 -20290 24652 -20288
rect 24498 -20300 24544 -20290
rect 24606 -20300 24652 -20290
rect 25134 -19596 25180 -19584
rect 25134 -20288 25140 -19596
rect 25174 -20288 25180 -19596
rect 25134 -20300 25180 -20288
rect 25570 -19596 25616 -19584
rect 25570 -20288 25576 -19596
rect 25610 -20288 25616 -19596
rect 25570 -20300 25616 -20288
rect 26098 -19590 26144 -19584
rect 26206 -19590 26252 -19584
rect 26098 -19596 26252 -19590
rect 26098 -20288 26104 -19596
rect 26138 -19600 26212 -19596
rect 26138 -20288 26212 -20280
rect 26246 -20288 26252 -19596
rect 26098 -20290 26252 -20288
rect 26098 -20300 26144 -20290
rect 26206 -20300 26252 -20290
rect 26734 -19596 26780 -19584
rect 26734 -20288 26740 -19596
rect 26774 -20288 26780 -19596
rect 26734 -20300 26780 -20288
rect 27170 -19596 27216 -19584
rect 27170 -20288 27176 -19596
rect 27210 -20288 27216 -19596
rect 27170 -20300 27216 -20288
rect 27698 -19590 27744 -19584
rect 27806 -19590 27852 -19584
rect 27698 -19596 27852 -19590
rect 27698 -20288 27704 -19596
rect 27738 -19600 27812 -19596
rect 27738 -20288 27812 -20280
rect 27846 -20288 27852 -19596
rect 27698 -20290 27852 -20288
rect 27698 -20300 27744 -20290
rect 27806 -20300 27852 -20290
rect 28334 -19596 28380 -19584
rect 28334 -20288 28340 -19596
rect 28374 -20288 28380 -19596
rect 28334 -20300 28380 -20288
rect 28770 -19596 28816 -19584
rect 28770 -20288 28776 -19596
rect 28810 -20288 28816 -19596
rect 28770 -20300 28816 -20288
rect 29298 -19590 29344 -19584
rect 29406 -19590 29452 -19584
rect 29298 -19596 29452 -19590
rect 29298 -20288 29304 -19596
rect 29338 -19600 29412 -19596
rect 29338 -20288 29412 -20280
rect 29446 -20288 29452 -19596
rect 29298 -20290 29452 -20288
rect 29298 -20300 29344 -20290
rect 29406 -20300 29452 -20290
rect 29934 -19596 29980 -19584
rect 29934 -20288 29940 -19596
rect 29974 -20288 29980 -19596
rect 29934 -20300 29980 -20288
rect 30370 -19596 30416 -19584
rect 30370 -20288 30376 -19596
rect 30410 -20288 30416 -19596
rect 30370 -20300 30416 -20288
rect 30898 -19590 30944 -19584
rect 31006 -19590 31052 -19584
rect 30898 -19596 31052 -19590
rect 30898 -20288 30904 -19596
rect 30938 -19600 31012 -19596
rect 30938 -20288 31012 -20280
rect 31046 -20288 31052 -19596
rect 30898 -20290 31052 -20288
rect 30898 -20300 30944 -20290
rect 31006 -20300 31052 -20290
rect 31534 -19596 31580 -19584
rect 31534 -20288 31540 -19596
rect 31574 -20288 31580 -19596
rect 31534 -20300 31580 -20288
rect 31970 -19596 32016 -19584
rect 31970 -20288 31976 -19596
rect 32010 -20288 32016 -19596
rect 31970 -20300 32016 -20288
rect 32498 -19590 32544 -19584
rect 32606 -19590 32652 -19584
rect 32498 -19596 32652 -19590
rect 32498 -20288 32504 -19596
rect 32538 -19600 32612 -19596
rect 32538 -20288 32612 -20280
rect 32646 -20288 32652 -19596
rect 32498 -20290 32652 -20288
rect 32498 -20300 32544 -20290
rect 32606 -20300 32652 -20290
rect 33134 -19596 33180 -19584
rect 33134 -20288 33140 -19596
rect 33174 -20288 33180 -19596
rect 33134 -20300 33180 -20288
rect 33570 -19596 33616 -19584
rect 33570 -20288 33576 -19596
rect 33610 -20288 33616 -19596
rect 33570 -20300 33616 -20288
rect 34098 -19590 34144 -19584
rect 34206 -19590 34252 -19584
rect 34098 -19596 34252 -19590
rect 34098 -20288 34104 -19596
rect 34138 -19600 34212 -19596
rect 34138 -20288 34212 -20280
rect 34246 -20288 34252 -19596
rect 34098 -20290 34252 -20288
rect 34098 -20300 34144 -20290
rect 34206 -20300 34252 -20290
rect 34734 -19596 34780 -19584
rect 34734 -20288 34740 -19596
rect 34774 -20288 34780 -19596
rect 34734 -20300 34780 -20288
rect 35170 -19596 35216 -19584
rect 35170 -20288 35176 -19596
rect 35210 -20288 35216 -19596
rect 35170 -20300 35216 -20288
rect 35698 -19590 35744 -19584
rect 35806 -19590 35852 -19584
rect 35698 -19596 35852 -19590
rect 35698 -20288 35704 -19596
rect 35738 -19600 35812 -19596
rect 35738 -20288 35812 -20280
rect 35846 -20288 35852 -19596
rect 35698 -20290 35852 -20288
rect 35698 -20300 35744 -20290
rect 35806 -20300 35852 -20290
rect 36334 -19596 36380 -19584
rect 36334 -20288 36340 -19596
rect 36374 -20288 36380 -19596
rect 36334 -20300 36380 -20288
rect 36770 -19596 36816 -19584
rect 36770 -20288 36776 -19596
rect 36810 -20288 36816 -19596
rect 36770 -20300 36816 -20288
rect 37298 -19596 37344 -19584
rect 37298 -20288 37304 -19596
rect 37338 -20288 37344 -19596
rect 37298 -20300 37344 -20288
rect 37406 -19596 37452 -19584
rect 37406 -20288 37412 -19596
rect 37446 -20288 37452 -19596
rect 37406 -20300 37452 -20288
rect 37934 -19596 37980 -19584
rect 37934 -20288 37940 -19596
rect 37974 -20288 37980 -19596
rect 37934 -20300 37980 -20288
rect 33180 -20340 33320 -20330
rect 670 -20354 1093 -20348
rect 670 -20388 705 -20354
rect 1081 -20380 1093 -20354
rect 1657 -20354 2057 -20348
rect 1657 -20380 1669 -20354
rect 1081 -20388 1669 -20380
rect 2045 -20380 2057 -20354
rect 2293 -20354 2693 -20348
rect 2293 -20380 2305 -20354
rect 2045 -20388 2305 -20380
rect 2681 -20380 2693 -20354
rect 3257 -20354 3657 -20348
rect 3257 -20380 3269 -20354
rect 2681 -20388 3269 -20380
rect 3645 -20380 3657 -20354
rect 3893 -20354 4293 -20348
rect 3893 -20380 3905 -20354
rect 3645 -20388 3905 -20380
rect 4281 -20380 4293 -20354
rect 4857 -20354 5257 -20348
rect 4857 -20380 4869 -20354
rect 4281 -20388 4869 -20380
rect 5245 -20380 5257 -20354
rect 5493 -20354 5893 -20348
rect 5493 -20380 5505 -20354
rect 5245 -20388 5505 -20380
rect 5881 -20380 5893 -20354
rect 6457 -20354 6857 -20348
rect 6457 -20380 6469 -20354
rect 5881 -20388 6469 -20380
rect 6845 -20380 6857 -20354
rect 7093 -20354 7493 -20348
rect 7093 -20380 7105 -20354
rect 6845 -20388 7105 -20380
rect 7481 -20380 7493 -20354
rect 8057 -20354 8457 -20348
rect 8057 -20380 8069 -20354
rect 7481 -20388 8069 -20380
rect 8445 -20380 8457 -20354
rect 8693 -20354 9093 -20348
rect 8693 -20380 8705 -20354
rect 8445 -20388 8705 -20380
rect 9081 -20380 9093 -20354
rect 9657 -20354 10057 -20348
rect 9657 -20380 9669 -20354
rect 9081 -20388 9669 -20380
rect 10045 -20380 10057 -20354
rect 10293 -20354 10693 -20348
rect 10293 -20380 10305 -20354
rect 10045 -20388 10305 -20380
rect 10681 -20380 10693 -20354
rect 11257 -20354 11657 -20348
rect 11257 -20380 11269 -20354
rect 10681 -20388 11269 -20380
rect 11645 -20380 11657 -20354
rect 11893 -20354 12293 -20348
rect 11893 -20380 11905 -20354
rect 11645 -20388 11905 -20380
rect 12281 -20380 12293 -20354
rect 12857 -20354 13257 -20348
rect 12857 -20380 12869 -20354
rect 12281 -20388 12869 -20380
rect 13245 -20380 13257 -20354
rect 13493 -20354 13893 -20348
rect 13493 -20380 13505 -20354
rect 13245 -20388 13505 -20380
rect 13881 -20380 13893 -20354
rect 14457 -20354 14857 -20348
rect 14457 -20380 14469 -20354
rect 13881 -20388 14469 -20380
rect 14845 -20380 14857 -20354
rect 15093 -20354 15493 -20348
rect 15093 -20380 15105 -20354
rect 14845 -20388 15105 -20380
rect 15481 -20380 15493 -20354
rect 16057 -20354 16457 -20348
rect 16057 -20380 16069 -20354
rect 15481 -20388 16069 -20380
rect 16445 -20380 16457 -20354
rect 16693 -20354 17093 -20348
rect 16693 -20380 16705 -20354
rect 16445 -20388 16705 -20380
rect 17081 -20380 17093 -20354
rect 17657 -20354 18057 -20348
rect 17657 -20380 17669 -20354
rect 17081 -20388 17669 -20380
rect 18045 -20380 18057 -20354
rect 18293 -20354 18693 -20348
rect 18293 -20380 18305 -20354
rect 18045 -20388 18305 -20380
rect 18681 -20380 18693 -20354
rect 19257 -20354 19657 -20348
rect 19257 -20380 19269 -20354
rect 18681 -20388 19269 -20380
rect 19645 -20380 19657 -20354
rect 19893 -20354 20293 -20348
rect 19893 -20380 19905 -20354
rect 19645 -20388 19905 -20380
rect 20281 -20380 20293 -20354
rect 20857 -20354 21257 -20348
rect 20857 -20380 20869 -20354
rect 20281 -20388 20869 -20380
rect 21245 -20380 21257 -20354
rect 21493 -20354 21893 -20348
rect 21493 -20380 21505 -20354
rect 21245 -20388 21505 -20380
rect 21881 -20380 21893 -20354
rect 22457 -20354 22857 -20348
rect 22457 -20380 22469 -20354
rect 21881 -20388 22469 -20380
rect 22845 -20380 22857 -20354
rect 23093 -20354 23493 -20348
rect 23093 -20380 23105 -20354
rect 22845 -20388 23105 -20380
rect 23481 -20380 23493 -20354
rect 24057 -20354 24457 -20348
rect 24057 -20380 24069 -20354
rect 23481 -20388 24069 -20380
rect 24445 -20380 24457 -20354
rect 24693 -20354 25093 -20348
rect 24693 -20380 24705 -20354
rect 24445 -20388 24705 -20380
rect 25081 -20380 25093 -20354
rect 25657 -20354 26057 -20348
rect 25657 -20380 25669 -20354
rect 25081 -20388 25669 -20380
rect 26045 -20380 26057 -20354
rect 26293 -20354 26693 -20348
rect 26293 -20380 26305 -20354
rect 26045 -20388 26305 -20380
rect 26681 -20380 26693 -20354
rect 27257 -20354 27657 -20348
rect 27257 -20380 27269 -20354
rect 26681 -20388 27269 -20380
rect 27645 -20380 27657 -20354
rect 27893 -20354 28293 -20348
rect 27893 -20380 27905 -20354
rect 27645 -20388 27905 -20380
rect 28281 -20380 28293 -20354
rect 28857 -20354 29257 -20348
rect 28857 -20380 28869 -20354
rect 28281 -20388 28869 -20380
rect 29245 -20380 29257 -20354
rect 29493 -20354 29893 -20348
rect 29493 -20380 29505 -20354
rect 29245 -20388 29505 -20380
rect 29881 -20380 29893 -20354
rect 30457 -20354 30857 -20348
rect 30457 -20380 30469 -20354
rect 29881 -20388 30469 -20380
rect 30845 -20380 30857 -20354
rect 31093 -20354 31493 -20348
rect 31093 -20380 31105 -20354
rect 30845 -20388 31105 -20380
rect 31481 -20388 31493 -20354
rect 670 -20394 31493 -20388
rect 32057 -20354 32457 -20348
rect 32057 -20388 32069 -20354
rect 32445 -20360 32457 -20354
rect 32693 -20354 33093 -20348
rect 32693 -20360 32705 -20354
rect 32445 -20388 32705 -20360
rect 33081 -20360 33093 -20354
rect 33180 -20360 33190 -20340
rect 33081 -20388 33190 -20360
rect 32057 -20394 33190 -20388
rect 670 -20482 31480 -20394
rect 32060 -20450 33190 -20394
rect 33180 -20460 33190 -20450
rect 33310 -20360 33320 -20340
rect 33657 -20354 34057 -20348
rect 33657 -20360 33669 -20354
rect 33310 -20388 33669 -20360
rect 34045 -20360 34057 -20354
rect 34293 -20354 34693 -20348
rect 34293 -20360 34305 -20354
rect 34045 -20388 34305 -20360
rect 34681 -20360 34693 -20354
rect 35257 -20354 35657 -20348
rect 35257 -20360 35269 -20354
rect 34681 -20388 35269 -20360
rect 35645 -20360 35657 -20354
rect 35893 -20354 36293 -20348
rect 35893 -20360 35905 -20354
rect 35645 -20388 35905 -20360
rect 36281 -20388 36293 -20354
rect 33310 -20394 36293 -20388
rect 36857 -20354 37257 -20348
rect 36857 -20388 36869 -20354
rect 37245 -20388 37257 -20354
rect 36857 -20394 37257 -20388
rect 37493 -20354 37893 -20348
rect 37493 -20388 37505 -20354
rect 37881 -20388 37893 -20354
rect 37493 -20394 37893 -20388
rect 33310 -20450 36280 -20394
rect 33310 -20460 33320 -20450
rect 33180 -20470 33320 -20460
rect 670 -20488 31549 -20482
rect 0 -20522 13 -20488
rect 1137 -20522 1613 -20488
rect 2737 -20522 3213 -20488
rect 4337 -20522 4813 -20488
rect 5937 -20522 6413 -20488
rect 7537 -20522 8013 -20488
rect 9137 -20522 9613 -20488
rect 10737 -20522 11213 -20488
rect 12337 -20522 12813 -20488
rect 13937 -20522 14413 -20488
rect 15537 -20522 16013 -20488
rect 17137 -20522 17613 -20488
rect 18737 -20522 19213 -20488
rect 20337 -20522 20813 -20488
rect 21937 -20522 22413 -20488
rect 23537 -20522 24013 -20488
rect 25137 -20522 25613 -20488
rect 26737 -20522 27213 -20488
rect 28337 -20522 28813 -20488
rect 29937 -20522 30413 -20488
rect 31537 -20500 31549 -20488
rect 32001 -20488 33149 -20482
rect 32001 -20500 32013 -20488
rect 31537 -20522 32013 -20500
rect 33137 -20500 33149 -20488
rect 33601 -20488 34749 -20482
rect 33601 -20500 33613 -20488
rect 33137 -20522 33613 -20500
rect 34737 -20500 34749 -20488
rect 35201 -20488 36349 -20482
rect 35201 -20500 35213 -20488
rect 34737 -20522 35213 -20500
rect 36337 -20500 36349 -20488
rect 36801 -20488 37949 -20482
rect 36801 -20500 36813 -20488
rect 36337 -20522 36813 -20500
rect 37937 -20522 37949 -20488
rect 0 -20620 490 -20522
rect 440 -20764 490 -20620
rect 57 -20770 490 -20764
rect 57 -20804 69 -20770
rect 445 -20804 490 -20770
rect 57 -20810 490 -20804
rect -30 -20857 16 -20845
rect -30 -20975 -24 -20857
rect 10 -20975 16 -20857
rect -30 -20987 16 -20975
rect 440 -21022 490 -20810
rect 670 -20528 37949 -20522
rect 670 -20620 37940 -20528
rect 670 -20764 720 -20620
rect 1200 -20670 1340 -20660
rect 670 -20770 1093 -20764
rect 670 -20804 705 -20770
rect 1081 -20804 1093 -20770
rect 1200 -20790 1210 -20670
rect 1330 -20680 1340 -20670
rect 2800 -20670 2940 -20660
rect 2800 -20680 2810 -20670
rect 1330 -20770 2810 -20680
rect 1330 -20780 1669 -20770
rect 1330 -20790 1340 -20780
rect 1200 -20800 1340 -20790
rect 670 -20810 1093 -20804
rect 1657 -20804 1669 -20780
rect 2045 -20780 2305 -20770
rect 2045 -20804 2057 -20780
rect 1657 -20810 2057 -20804
rect 2293 -20804 2305 -20780
rect 2681 -20780 2810 -20770
rect 2681 -20804 2693 -20780
rect 2800 -20790 2810 -20780
rect 2930 -20680 2940 -20670
rect 4400 -20670 4540 -20660
rect 4400 -20680 4410 -20670
rect 2930 -20770 4410 -20680
rect 2930 -20780 3269 -20770
rect 2930 -20790 2940 -20780
rect 2800 -20800 2940 -20790
rect 2293 -20810 2693 -20804
rect 3257 -20804 3269 -20780
rect 3645 -20780 3905 -20770
rect 3645 -20804 3657 -20780
rect 3257 -20810 3657 -20804
rect 3893 -20804 3905 -20780
rect 4281 -20780 4410 -20770
rect 4281 -20804 4293 -20780
rect 4400 -20790 4410 -20780
rect 4530 -20680 4540 -20670
rect 6000 -20670 6140 -20660
rect 6000 -20680 6010 -20670
rect 4530 -20770 6010 -20680
rect 4530 -20780 4869 -20770
rect 4530 -20790 4540 -20780
rect 4400 -20800 4540 -20790
rect 3893 -20810 4293 -20804
rect 4857 -20804 4869 -20780
rect 5245 -20780 5505 -20770
rect 5245 -20804 5257 -20780
rect 4857 -20810 5257 -20804
rect 5493 -20804 5505 -20780
rect 5881 -20780 6010 -20770
rect 5881 -20804 5893 -20780
rect 6000 -20790 6010 -20780
rect 6130 -20680 6140 -20670
rect 7600 -20670 7740 -20660
rect 7600 -20680 7610 -20670
rect 6130 -20770 7610 -20680
rect 6130 -20780 6469 -20770
rect 6130 -20790 6140 -20780
rect 6000 -20800 6140 -20790
rect 5493 -20810 5893 -20804
rect 6457 -20804 6469 -20780
rect 6845 -20780 7105 -20770
rect 6845 -20804 6857 -20780
rect 6457 -20810 6857 -20804
rect 7093 -20804 7105 -20780
rect 7481 -20780 7610 -20770
rect 7481 -20804 7493 -20780
rect 7600 -20790 7610 -20780
rect 7730 -20680 7740 -20670
rect 9200 -20670 9340 -20660
rect 15820 -20670 15960 -20660
rect 9200 -20680 9210 -20670
rect 7730 -20770 9210 -20680
rect 7730 -20780 8069 -20770
rect 7730 -20790 7740 -20780
rect 7600 -20800 7740 -20790
rect 7093 -20810 7493 -20804
rect 8057 -20804 8069 -20780
rect 8445 -20780 8705 -20770
rect 8445 -20804 8457 -20780
rect 8057 -20810 8457 -20804
rect 8693 -20804 8705 -20780
rect 9081 -20780 9210 -20770
rect 9081 -20804 9093 -20780
rect 9200 -20790 9210 -20780
rect 9330 -20680 9340 -20670
rect 12400 -20680 12540 -20670
rect 9330 -20770 10700 -20680
rect 12400 -20700 12410 -20680
rect 11260 -20764 12410 -20700
rect 9330 -20780 9669 -20770
rect 9330 -20790 9340 -20780
rect 9200 -20800 9340 -20790
rect 8693 -20810 9093 -20804
rect 9657 -20804 9669 -20780
rect 10045 -20780 10305 -20770
rect 10045 -20804 10057 -20780
rect 9657 -20810 10057 -20804
rect 10293 -20804 10305 -20780
rect 10681 -20780 10700 -20770
rect 11257 -20770 12410 -20764
rect 10681 -20804 10693 -20780
rect 10293 -20810 10693 -20804
rect 11257 -20804 11269 -20770
rect 11645 -20800 11905 -20770
rect 11645 -20804 11657 -20800
rect 11257 -20810 11657 -20804
rect 11893 -20804 11905 -20800
rect 12281 -20800 12410 -20770
rect 12530 -20800 12540 -20680
rect 12281 -20804 12293 -20800
rect 11893 -20810 12293 -20804
rect 12400 -20810 12540 -20800
rect 12857 -20770 13257 -20764
rect 12857 -20804 12869 -20770
rect 13245 -20804 13257 -20770
rect 12857 -20810 13257 -20804
rect 13493 -20770 13893 -20764
rect 13493 -20804 13505 -20770
rect 13881 -20804 13893 -20770
rect 13493 -20810 13893 -20804
rect 14457 -20770 14857 -20764
rect 14457 -20804 14469 -20770
rect 14845 -20804 14857 -20770
rect 14457 -20810 14857 -20804
rect 15093 -20770 15493 -20764
rect 15093 -20804 15105 -20770
rect 15481 -20804 15493 -20770
rect 15820 -20790 15830 -20670
rect 15950 -20700 15960 -20670
rect 17420 -20670 17560 -20660
rect 15950 -20764 17090 -20700
rect 15950 -20770 17093 -20764
rect 15950 -20790 16069 -20770
rect 15820 -20800 16069 -20790
rect 15093 -20810 15493 -20804
rect 16057 -20804 16069 -20800
rect 16445 -20800 16705 -20770
rect 16445 -20804 16457 -20800
rect 16057 -20810 16457 -20804
rect 16693 -20804 16705 -20800
rect 17081 -20804 17093 -20770
rect 17420 -20790 17430 -20670
rect 17550 -20700 17560 -20670
rect 19020 -20670 19160 -20660
rect 17550 -20764 18690 -20700
rect 17550 -20770 18693 -20764
rect 17550 -20790 17669 -20770
rect 17420 -20800 17669 -20790
rect 16693 -20810 17093 -20804
rect 17657 -20804 17669 -20800
rect 18045 -20800 18305 -20770
rect 18045 -20804 18057 -20800
rect 17657 -20810 18057 -20804
rect 18293 -20804 18305 -20800
rect 18681 -20804 18693 -20770
rect 19020 -20790 19030 -20670
rect 19150 -20700 19160 -20670
rect 20620 -20670 20760 -20660
rect 19150 -20764 20290 -20700
rect 19150 -20770 20293 -20764
rect 19150 -20790 19269 -20770
rect 19020 -20800 19269 -20790
rect 18293 -20810 18693 -20804
rect 19257 -20804 19269 -20800
rect 19645 -20800 19905 -20770
rect 19645 -20804 19657 -20800
rect 19257 -20810 19657 -20804
rect 19893 -20804 19905 -20800
rect 20281 -20804 20293 -20770
rect 20620 -20790 20630 -20670
rect 20750 -20700 20760 -20670
rect 22220 -20670 22360 -20660
rect 20750 -20764 21890 -20700
rect 20750 -20770 21893 -20764
rect 20750 -20790 20869 -20770
rect 20620 -20800 20869 -20790
rect 19893 -20810 20293 -20804
rect 20857 -20804 20869 -20800
rect 21245 -20800 21505 -20770
rect 21245 -20804 21257 -20800
rect 20857 -20810 21257 -20804
rect 21493 -20804 21505 -20800
rect 21881 -20804 21893 -20770
rect 22220 -20790 22230 -20670
rect 22350 -20700 22360 -20670
rect 23820 -20670 23960 -20660
rect 22350 -20764 23490 -20700
rect 22350 -20770 23493 -20764
rect 22350 -20790 22469 -20770
rect 22220 -20800 22469 -20790
rect 21493 -20810 21893 -20804
rect 22457 -20804 22469 -20800
rect 22845 -20800 23105 -20770
rect 22845 -20804 22857 -20800
rect 22457 -20810 22857 -20804
rect 23093 -20804 23105 -20800
rect 23481 -20804 23493 -20770
rect 23820 -20790 23830 -20670
rect 23950 -20700 23960 -20670
rect 27020 -20670 27160 -20660
rect 27020 -20700 27030 -20670
rect 23950 -20764 25090 -20700
rect 25660 -20764 27030 -20700
rect 23950 -20770 25093 -20764
rect 23950 -20790 24069 -20770
rect 23820 -20800 24069 -20790
rect 23093 -20810 23493 -20804
rect 24057 -20804 24069 -20800
rect 24445 -20800 24705 -20770
rect 24445 -20804 24457 -20800
rect 24057 -20810 24457 -20804
rect 24693 -20804 24705 -20800
rect 25081 -20804 25093 -20770
rect 24693 -20810 25093 -20804
rect 25657 -20770 27030 -20764
rect 25657 -20804 25669 -20770
rect 26045 -20800 26305 -20770
rect 26045 -20804 26057 -20800
rect 25657 -20810 26057 -20804
rect 26293 -20804 26305 -20800
rect 26681 -20790 27030 -20770
rect 27150 -20700 27160 -20670
rect 28620 -20670 28760 -20660
rect 27150 -20764 28290 -20700
rect 27150 -20770 28293 -20764
rect 27150 -20790 27269 -20770
rect 26681 -20800 27269 -20790
rect 26681 -20804 26693 -20800
rect 26293 -20810 26693 -20804
rect 27257 -20804 27269 -20800
rect 27645 -20800 27905 -20770
rect 27645 -20804 27657 -20800
rect 27257 -20810 27657 -20804
rect 27893 -20804 27905 -20800
rect 28281 -20804 28293 -20770
rect 28620 -20790 28630 -20670
rect 28750 -20700 28760 -20670
rect 31580 -20680 31720 -20670
rect 28750 -20764 31490 -20700
rect 28750 -20770 31493 -20764
rect 28750 -20790 28869 -20770
rect 28620 -20800 28869 -20790
rect 27893 -20810 28293 -20804
rect 28857 -20804 28869 -20800
rect 29245 -20800 29505 -20770
rect 29245 -20804 29257 -20800
rect 28857 -20810 29257 -20804
rect 29493 -20804 29505 -20800
rect 29881 -20800 30469 -20770
rect 29881 -20804 29893 -20800
rect 29493 -20810 29893 -20804
rect 30457 -20804 30469 -20800
rect 30845 -20800 31105 -20770
rect 30845 -20804 30857 -20800
rect 30457 -20810 30857 -20804
rect 31093 -20804 31105 -20800
rect 31481 -20804 31493 -20770
rect 31093 -20810 31493 -20804
rect 31580 -20800 31590 -20680
rect 31710 -20700 31720 -20680
rect 31710 -20764 36280 -20700
rect 31710 -20770 36293 -20764
rect 31710 -20800 32069 -20770
rect 31580 -20810 31720 -20800
rect 32057 -20804 32069 -20800
rect 32445 -20800 32705 -20770
rect 32445 -20804 32457 -20800
rect 32057 -20810 32457 -20804
rect 32693 -20804 32705 -20800
rect 33081 -20800 33669 -20770
rect 33081 -20804 33093 -20800
rect 32693 -20810 33093 -20804
rect 33657 -20804 33669 -20800
rect 34045 -20800 34305 -20770
rect 34045 -20804 34057 -20800
rect 33657 -20810 34057 -20804
rect 34293 -20804 34305 -20800
rect 34681 -20800 35269 -20770
rect 34681 -20804 34693 -20800
rect 34293 -20810 34693 -20804
rect 35257 -20804 35269 -20800
rect 35645 -20800 35905 -20770
rect 35645 -20804 35657 -20800
rect 35257 -20810 35657 -20804
rect 35893 -20804 35905 -20800
rect 36281 -20804 36293 -20770
rect 35893 -20810 36293 -20804
rect 36857 -20770 37257 -20764
rect 36857 -20804 36869 -20770
rect 37245 -20804 37257 -20770
rect 36857 -20810 37257 -20804
rect 37493 -20770 37893 -20764
rect 37493 -20804 37505 -20770
rect 37881 -20804 37893 -20770
rect 37493 -20810 37893 -20804
rect 57 -21028 490 -21022
rect 57 -21062 69 -21028
rect 445 -21062 490 -21028
rect 57 -21068 490 -21062
rect 440 -21290 490 -21068
rect 57 -21296 490 -21290
rect 57 -21330 69 -21296
rect 445 -21330 490 -21296
rect 57 -21336 490 -21330
rect -30 -21396 16 -21384
rect -30 -22088 -24 -21396
rect 10 -22088 16 -21396
rect -30 -22100 16 -22088
rect 440 -22148 490 -21336
rect 670 -21022 720 -20810
rect 1134 -20857 1180 -20845
rect 1134 -20975 1140 -20857
rect 1174 -20975 1180 -20857
rect 1570 -20857 1616 -20845
rect 1570 -20860 1576 -20857
rect 1134 -20987 1180 -20975
rect 1560 -20975 1576 -20860
rect 1610 -20860 1616 -20857
rect 2098 -20857 2144 -20845
rect 2098 -20860 2104 -20857
rect 1610 -20975 2104 -20860
rect 2138 -20860 2144 -20857
rect 2206 -20857 2252 -20845
rect 2206 -20860 2212 -20857
rect 2138 -20975 2212 -20860
rect 2246 -20860 2252 -20857
rect 2734 -20857 2780 -20845
rect 2734 -20860 2740 -20857
rect 2246 -20975 2740 -20860
rect 2774 -20860 2780 -20857
rect 3170 -20857 3216 -20845
rect 3170 -20860 3176 -20857
rect 2774 -20975 3176 -20860
rect 3210 -20860 3216 -20857
rect 3698 -20857 3744 -20845
rect 3698 -20860 3704 -20857
rect 3210 -20975 3704 -20860
rect 3738 -20860 3744 -20857
rect 3806 -20857 3852 -20845
rect 3806 -20860 3812 -20857
rect 3738 -20975 3812 -20860
rect 3846 -20860 3852 -20857
rect 4334 -20857 4380 -20845
rect 4334 -20860 4340 -20857
rect 3846 -20975 4340 -20860
rect 4374 -20860 4380 -20857
rect 4770 -20857 4816 -20845
rect 4770 -20860 4776 -20857
rect 4374 -20975 4776 -20860
rect 4810 -20860 4816 -20857
rect 5298 -20857 5344 -20845
rect 5298 -20860 5304 -20857
rect 4810 -20975 5304 -20860
rect 5338 -20860 5344 -20857
rect 5406 -20857 5452 -20845
rect 5406 -20860 5412 -20857
rect 5338 -20975 5412 -20860
rect 5446 -20860 5452 -20857
rect 5934 -20857 5980 -20845
rect 5934 -20860 5940 -20857
rect 5446 -20975 5940 -20860
rect 5974 -20860 5980 -20857
rect 6370 -20857 6416 -20845
rect 6370 -20860 6376 -20857
rect 5974 -20975 6376 -20860
rect 6410 -20860 6416 -20857
rect 6898 -20857 6944 -20845
rect 6898 -20860 6904 -20857
rect 6410 -20975 6904 -20860
rect 6938 -20860 6944 -20857
rect 7006 -20857 7052 -20845
rect 7006 -20860 7012 -20857
rect 6938 -20975 7012 -20860
rect 7046 -20860 7052 -20857
rect 7534 -20857 7580 -20845
rect 7534 -20860 7540 -20857
rect 7046 -20975 7540 -20860
rect 7574 -20860 7580 -20857
rect 7970 -20857 8016 -20845
rect 7970 -20860 7976 -20857
rect 7574 -20975 7976 -20860
rect 8010 -20860 8016 -20857
rect 8498 -20857 8544 -20845
rect 8498 -20860 8504 -20857
rect 8010 -20975 8504 -20860
rect 8538 -20860 8544 -20857
rect 8606 -20857 8652 -20845
rect 8606 -20860 8612 -20857
rect 8538 -20975 8612 -20860
rect 8646 -20860 8652 -20857
rect 9134 -20857 9180 -20845
rect 9134 -20860 9140 -20857
rect 8646 -20975 9140 -20860
rect 9174 -20860 9180 -20857
rect 9570 -20857 9616 -20845
rect 9570 -20860 9576 -20857
rect 9174 -20975 9576 -20860
rect 9610 -20860 9616 -20857
rect 10098 -20857 10144 -20845
rect 10098 -20860 10104 -20857
rect 9610 -20975 10104 -20860
rect 10138 -20860 10144 -20857
rect 10206 -20857 10252 -20845
rect 10206 -20860 10212 -20857
rect 10138 -20975 10212 -20860
rect 10246 -20860 10252 -20857
rect 10734 -20850 10780 -20845
rect 10734 -20857 10940 -20850
rect 10734 -20860 10740 -20857
rect 10246 -20975 10740 -20860
rect 10774 -20860 10940 -20857
rect 11170 -20857 11216 -20845
rect 11170 -20860 11176 -20857
rect 10774 -20975 10810 -20860
rect 1560 -20980 10810 -20975
rect 10930 -20975 11176 -20860
rect 11210 -20860 11216 -20857
rect 11698 -20857 11744 -20845
rect 11698 -20860 11704 -20857
rect 11210 -20975 11704 -20860
rect 11738 -20860 11744 -20857
rect 11806 -20857 11852 -20845
rect 11806 -20860 11812 -20857
rect 11738 -20975 11812 -20860
rect 11846 -20860 11852 -20857
rect 12334 -20857 12380 -20845
rect 12334 -20860 12340 -20857
rect 11846 -20975 12340 -20860
rect 12374 -20860 12380 -20857
rect 12770 -20857 12816 -20845
rect 12770 -20860 12776 -20857
rect 12374 -20975 12776 -20860
rect 12810 -20860 12816 -20857
rect 13000 -20860 13120 -20810
rect 13298 -20857 13344 -20845
rect 13298 -20860 13304 -20857
rect 12810 -20975 13304 -20860
rect 13338 -20860 13344 -20857
rect 13406 -20857 13452 -20845
rect 13406 -20860 13412 -20857
rect 13338 -20975 13412 -20860
rect 13446 -20860 13452 -20857
rect 13640 -20860 13760 -20810
rect 13934 -20857 13980 -20845
rect 13934 -20860 13940 -20857
rect 13446 -20975 13940 -20860
rect 13974 -20860 13980 -20857
rect 14370 -20857 14416 -20845
rect 14370 -20860 14376 -20857
rect 13974 -20975 14376 -20860
rect 14410 -20860 14416 -20857
rect 14600 -20860 14720 -20810
rect 14898 -20857 14944 -20845
rect 14898 -20860 14904 -20857
rect 14410 -20975 14904 -20860
rect 14938 -20860 14944 -20857
rect 15006 -20857 15052 -20845
rect 15006 -20860 15012 -20857
rect 14938 -20975 15012 -20860
rect 15046 -20860 15052 -20857
rect 15240 -20860 15360 -20810
rect 15534 -20857 15580 -20845
rect 15534 -20860 15540 -20857
rect 15046 -20975 15540 -20860
rect 15574 -20860 15580 -20857
rect 15970 -20857 16016 -20845
rect 15970 -20860 15976 -20857
rect 15574 -20975 15976 -20860
rect 16010 -20860 16016 -20857
rect 16498 -20857 16544 -20845
rect 16498 -20860 16504 -20857
rect 16010 -20975 16504 -20860
rect 16538 -20860 16544 -20857
rect 16606 -20857 16652 -20845
rect 16606 -20860 16612 -20857
rect 16538 -20975 16612 -20860
rect 16646 -20860 16652 -20857
rect 17134 -20857 17180 -20845
rect 17134 -20860 17140 -20857
rect 16646 -20975 17140 -20860
rect 17174 -20860 17180 -20857
rect 17570 -20857 17616 -20845
rect 17570 -20860 17576 -20857
rect 17174 -20975 17576 -20860
rect 17610 -20860 17616 -20857
rect 18098 -20857 18144 -20845
rect 18098 -20860 18104 -20857
rect 17610 -20975 18104 -20860
rect 18138 -20860 18144 -20857
rect 18206 -20857 18252 -20845
rect 18206 -20860 18212 -20857
rect 18138 -20975 18212 -20860
rect 18246 -20860 18252 -20857
rect 18734 -20857 18780 -20845
rect 18734 -20860 18740 -20857
rect 18246 -20975 18740 -20860
rect 18774 -20860 18780 -20857
rect 19170 -20857 19216 -20845
rect 19170 -20860 19176 -20857
rect 18774 -20975 19176 -20860
rect 19210 -20860 19216 -20857
rect 19698 -20857 19744 -20845
rect 19698 -20860 19704 -20857
rect 19210 -20975 19704 -20860
rect 19738 -20860 19744 -20857
rect 19806 -20857 19852 -20845
rect 19806 -20860 19812 -20857
rect 19738 -20975 19812 -20860
rect 19846 -20860 19852 -20857
rect 20334 -20857 20380 -20845
rect 20334 -20860 20340 -20857
rect 19846 -20975 20340 -20860
rect 20374 -20860 20380 -20857
rect 20770 -20857 20816 -20845
rect 20770 -20860 20776 -20857
rect 20374 -20975 20776 -20860
rect 20810 -20860 20816 -20857
rect 21298 -20857 21344 -20845
rect 21298 -20860 21304 -20857
rect 20810 -20975 21304 -20860
rect 21338 -20860 21344 -20857
rect 21406 -20857 21452 -20845
rect 21406 -20860 21412 -20857
rect 21338 -20975 21412 -20860
rect 21446 -20860 21452 -20857
rect 21934 -20857 21980 -20845
rect 21934 -20860 21940 -20857
rect 21446 -20975 21940 -20860
rect 21974 -20860 21980 -20857
rect 22370 -20857 22416 -20845
rect 22370 -20860 22376 -20857
rect 21974 -20975 22376 -20860
rect 22410 -20860 22416 -20857
rect 22898 -20857 22944 -20845
rect 22898 -20860 22904 -20857
rect 22410 -20975 22904 -20860
rect 22938 -20860 22944 -20857
rect 23006 -20857 23052 -20845
rect 23006 -20860 23012 -20857
rect 22938 -20975 23012 -20860
rect 23046 -20860 23052 -20857
rect 23534 -20857 23580 -20845
rect 23534 -20860 23540 -20857
rect 23046 -20975 23540 -20860
rect 23574 -20860 23580 -20857
rect 23970 -20857 24016 -20845
rect 23970 -20860 23976 -20857
rect 23574 -20975 23976 -20860
rect 24010 -20860 24016 -20857
rect 24498 -20857 24544 -20845
rect 24498 -20860 24504 -20857
rect 24010 -20975 24504 -20860
rect 24538 -20860 24544 -20857
rect 24606 -20857 24652 -20845
rect 24606 -20860 24612 -20857
rect 24538 -20975 24612 -20860
rect 24646 -20860 24652 -20857
rect 25134 -20857 25180 -20845
rect 25134 -20860 25140 -20857
rect 24646 -20975 25140 -20860
rect 25174 -20860 25180 -20857
rect 25570 -20857 25616 -20845
rect 25570 -20860 25576 -20857
rect 25174 -20975 25576 -20860
rect 25610 -20860 25616 -20857
rect 26098 -20857 26144 -20845
rect 26098 -20860 26104 -20857
rect 25610 -20975 26104 -20860
rect 26138 -20860 26144 -20857
rect 26206 -20857 26252 -20845
rect 26206 -20860 26212 -20857
rect 26138 -20975 26212 -20860
rect 26246 -20860 26252 -20857
rect 26734 -20857 26780 -20845
rect 26734 -20860 26740 -20857
rect 26246 -20975 26740 -20860
rect 26774 -20860 26780 -20857
rect 27170 -20857 27216 -20845
rect 27170 -20860 27176 -20857
rect 26774 -20975 27176 -20860
rect 27210 -20860 27216 -20857
rect 27698 -20857 27744 -20845
rect 27698 -20860 27704 -20857
rect 27210 -20975 27704 -20860
rect 27738 -20860 27744 -20857
rect 27806 -20857 27852 -20845
rect 27806 -20860 27812 -20857
rect 27738 -20975 27812 -20860
rect 27846 -20860 27852 -20857
rect 28334 -20857 28380 -20845
rect 28334 -20860 28340 -20857
rect 27846 -20975 28340 -20860
rect 28374 -20860 28380 -20857
rect 28770 -20857 28816 -20845
rect 28770 -20860 28776 -20857
rect 28374 -20975 28776 -20860
rect 28810 -20860 28816 -20857
rect 29298 -20857 29344 -20845
rect 29298 -20860 29304 -20857
rect 28810 -20975 29304 -20860
rect 29338 -20860 29344 -20857
rect 29406 -20857 29452 -20845
rect 29406 -20860 29412 -20857
rect 29338 -20975 29412 -20860
rect 29446 -20860 29452 -20857
rect 29934 -20857 29980 -20845
rect 29934 -20860 29940 -20857
rect 29446 -20975 29940 -20860
rect 29974 -20860 29980 -20857
rect 30370 -20857 30416 -20845
rect 30370 -20860 30376 -20857
rect 29974 -20975 30376 -20860
rect 30410 -20860 30416 -20857
rect 30898 -20857 30944 -20845
rect 30898 -20860 30904 -20857
rect 30410 -20975 30904 -20860
rect 30938 -20860 30944 -20857
rect 31006 -20857 31052 -20845
rect 31006 -20860 31012 -20857
rect 30938 -20975 31012 -20860
rect 31046 -20860 31052 -20857
rect 31534 -20857 31580 -20845
rect 31534 -20860 31540 -20857
rect 31046 -20975 31540 -20860
rect 31574 -20860 31580 -20857
rect 31970 -20857 32016 -20845
rect 31970 -20860 31976 -20857
rect 31574 -20975 31976 -20860
rect 32010 -20860 32016 -20857
rect 32498 -20857 32544 -20845
rect 32498 -20860 32504 -20857
rect 32010 -20975 32504 -20860
rect 32538 -20860 32544 -20857
rect 32606 -20857 32652 -20845
rect 32606 -20860 32612 -20857
rect 32538 -20975 32612 -20860
rect 32646 -20860 32652 -20857
rect 33134 -20857 33180 -20845
rect 33134 -20860 33140 -20857
rect 32646 -20975 33140 -20860
rect 33174 -20860 33180 -20857
rect 33570 -20857 33616 -20845
rect 33570 -20860 33576 -20857
rect 33174 -20975 33576 -20860
rect 33610 -20860 33616 -20857
rect 34098 -20857 34144 -20845
rect 34098 -20860 34104 -20857
rect 33610 -20975 34104 -20860
rect 34138 -20860 34144 -20857
rect 34206 -20857 34252 -20845
rect 34206 -20860 34212 -20857
rect 34138 -20975 34212 -20860
rect 34246 -20860 34252 -20857
rect 34734 -20857 34780 -20845
rect 34734 -20860 34740 -20857
rect 34246 -20975 34740 -20860
rect 34774 -20860 34780 -20857
rect 35170 -20857 35216 -20845
rect 35170 -20860 35176 -20857
rect 34774 -20975 35176 -20860
rect 35210 -20860 35216 -20857
rect 35698 -20857 35744 -20845
rect 35698 -20860 35704 -20857
rect 35210 -20975 35704 -20860
rect 35738 -20860 35744 -20857
rect 35806 -20857 35852 -20845
rect 35806 -20860 35812 -20857
rect 35738 -20975 35812 -20860
rect 35846 -20860 35852 -20857
rect 36334 -20857 36380 -20845
rect 36334 -20860 36340 -20857
rect 35846 -20975 36340 -20860
rect 36374 -20975 36380 -20857
rect 10930 -20980 36380 -20975
rect 1570 -20987 1616 -20980
rect 2098 -20987 2144 -20980
rect 2206 -20987 2252 -20980
rect 2734 -20987 2780 -20980
rect 3170 -20987 3216 -20980
rect 3698 -20987 3744 -20980
rect 3806 -20987 3852 -20980
rect 4334 -20987 4380 -20980
rect 4770 -20987 4816 -20980
rect 5298 -20987 5344 -20980
rect 5406 -20987 5452 -20980
rect 5934 -20987 5980 -20980
rect 6370 -20987 6416 -20980
rect 6898 -20987 6944 -20980
rect 7006 -20987 7052 -20980
rect 7534 -20987 7580 -20980
rect 7970 -20987 8016 -20980
rect 8498 -20987 8544 -20980
rect 8606 -20987 8652 -20980
rect 9134 -20987 9180 -20980
rect 9570 -20987 9616 -20980
rect 10098 -20987 10144 -20980
rect 10206 -20987 10252 -20980
rect 10734 -20987 10940 -20980
rect 11170 -20987 11216 -20980
rect 11698 -20987 11744 -20980
rect 11806 -20987 11852 -20980
rect 12334 -20987 12380 -20980
rect 12770 -20987 12816 -20980
rect 10750 -20990 10940 -20987
rect 13000 -21022 13120 -20980
rect 13298 -20987 13344 -20980
rect 13406 -20987 13452 -20980
rect 13640 -21022 13760 -20980
rect 13934 -20987 13980 -20980
rect 14370 -20987 14416 -20980
rect 14600 -21022 14720 -20980
rect 14898 -20987 14944 -20980
rect 15006 -20987 15052 -20980
rect 15240 -21022 15360 -20980
rect 15534 -20987 15580 -20980
rect 15970 -20987 16016 -20980
rect 16498 -20987 16544 -20980
rect 16606 -20987 16652 -20980
rect 17134 -20987 17180 -20980
rect 17570 -20987 17616 -20980
rect 18098 -20987 18144 -20980
rect 18206 -20987 18252 -20980
rect 18734 -20987 18780 -20980
rect 19170 -20987 19216 -20980
rect 19698 -20987 19744 -20980
rect 19806 -20987 19852 -20980
rect 20334 -20987 20380 -20980
rect 20770 -20987 20816 -20980
rect 21298 -20987 21344 -20980
rect 21406 -20987 21452 -20980
rect 21934 -20987 21980 -20980
rect 22370 -20987 22416 -20980
rect 22898 -20987 22944 -20980
rect 23006 -20987 23052 -20980
rect 23534 -20987 23580 -20980
rect 23970 -20987 24016 -20980
rect 24498 -20987 24544 -20980
rect 24606 -20987 24652 -20980
rect 25134 -20987 25180 -20980
rect 25570 -20987 25616 -20980
rect 26098 -20987 26144 -20980
rect 26206 -20987 26252 -20980
rect 26734 -20987 26780 -20980
rect 27170 -20987 27216 -20980
rect 27698 -20987 27744 -20980
rect 27806 -20987 27852 -20980
rect 28334 -20987 28380 -20980
rect 28770 -20987 28816 -20980
rect 29298 -20987 29344 -20980
rect 29406 -20987 29452 -20980
rect 29934 -20987 29980 -20980
rect 30370 -20987 30416 -20980
rect 30898 -20987 30944 -20980
rect 31006 -20987 31052 -20980
rect 31534 -20987 31580 -20980
rect 31970 -20987 32016 -20980
rect 32498 -20987 32544 -20980
rect 32606 -20987 32652 -20980
rect 33134 -20987 33180 -20980
rect 33570 -20987 33616 -20980
rect 34098 -20987 34144 -20980
rect 34206 -20987 34252 -20980
rect 34734 -20987 34780 -20980
rect 35170 -20987 35216 -20980
rect 35698 -20987 35744 -20980
rect 35806 -20987 35852 -20980
rect 36334 -20987 36380 -20980
rect 36770 -20857 36816 -20845
rect 36770 -20975 36776 -20857
rect 36810 -20975 36816 -20857
rect 36770 -20987 36816 -20975
rect 37298 -20857 37344 -20845
rect 37298 -20975 37304 -20857
rect 37338 -20975 37344 -20857
rect 37298 -20987 37344 -20975
rect 37406 -20857 37452 -20845
rect 37406 -20975 37412 -20857
rect 37446 -20975 37452 -20857
rect 37406 -20987 37452 -20975
rect 37934 -20857 37980 -20845
rect 37934 -20975 37940 -20857
rect 37974 -20975 37980 -20857
rect 37934 -20987 37980 -20975
rect 670 -21028 1093 -21022
rect 670 -21062 705 -21028
rect 1081 -21062 1093 -21028
rect 670 -21068 1093 -21062
rect 1657 -21028 2057 -21022
rect 1657 -21062 1669 -21028
rect 2045 -21030 2057 -21028
rect 2293 -21028 2693 -21022
rect 2293 -21030 2305 -21028
rect 2045 -21062 2060 -21030
rect 1657 -21068 2060 -21062
rect 670 -21290 720 -21068
rect 1420 -21110 1560 -21100
rect 1420 -21230 1430 -21110
rect 1550 -21120 1560 -21110
rect 1660 -21120 2060 -21068
rect 2290 -21062 2305 -21030
rect 2681 -21062 2693 -21028
rect 2290 -21068 2693 -21062
rect 3257 -21028 3657 -21022
rect 3257 -21062 3269 -21028
rect 3645 -21030 3657 -21028
rect 3893 -21028 4293 -21022
rect 3893 -21030 3905 -21028
rect 3645 -21062 3660 -21030
rect 3257 -21068 3660 -21062
rect 2290 -21120 2690 -21068
rect 3020 -21110 3160 -21100
rect 3020 -21120 3030 -21110
rect 1550 -21220 3030 -21120
rect 1550 -21230 1560 -21220
rect 1420 -21240 1560 -21230
rect 1660 -21240 2690 -21220
rect 3020 -21230 3030 -21220
rect 3150 -21120 3160 -21110
rect 3260 -21120 3660 -21068
rect 3890 -21062 3905 -21030
rect 4281 -21062 4293 -21028
rect 3890 -21068 4293 -21062
rect 4857 -21028 5257 -21022
rect 4857 -21062 4869 -21028
rect 5245 -21030 5257 -21028
rect 5493 -21028 5893 -21022
rect 5493 -21030 5505 -21028
rect 5245 -21062 5260 -21030
rect 4857 -21068 5260 -21062
rect 3890 -21120 4290 -21068
rect 4620 -21110 4760 -21100
rect 4620 -21120 4630 -21110
rect 3150 -21220 4630 -21120
rect 3150 -21230 3160 -21220
rect 3020 -21240 3160 -21230
rect 3260 -21240 4290 -21220
rect 4620 -21230 4630 -21220
rect 4750 -21120 4760 -21110
rect 4860 -21120 5260 -21068
rect 5490 -21062 5505 -21030
rect 5881 -21062 5893 -21028
rect 5490 -21068 5893 -21062
rect 6457 -21028 6857 -21022
rect 6457 -21062 6469 -21028
rect 6845 -21030 6857 -21028
rect 7093 -21028 7493 -21022
rect 7093 -21030 7105 -21028
rect 6845 -21062 6860 -21030
rect 6457 -21068 6860 -21062
rect 5490 -21120 5890 -21068
rect 6220 -21110 6360 -21100
rect 6220 -21120 6230 -21110
rect 4750 -21220 6230 -21120
rect 4750 -21230 4760 -21220
rect 4620 -21240 4760 -21230
rect 4860 -21240 5890 -21220
rect 6220 -21230 6230 -21220
rect 6350 -21120 6360 -21110
rect 6460 -21120 6860 -21068
rect 7090 -21062 7105 -21030
rect 7481 -21062 7493 -21028
rect 7090 -21068 7493 -21062
rect 8057 -21028 8457 -21022
rect 8057 -21062 8069 -21028
rect 8445 -21030 8457 -21028
rect 8693 -21028 9093 -21022
rect 8693 -21030 8705 -21028
rect 8445 -21062 8460 -21030
rect 8057 -21068 8460 -21062
rect 7090 -21120 7490 -21068
rect 7820 -21110 7960 -21100
rect 7820 -21120 7830 -21110
rect 6350 -21220 7830 -21120
rect 6350 -21230 6360 -21220
rect 6220 -21240 6360 -21230
rect 6460 -21240 7490 -21220
rect 7820 -21230 7830 -21220
rect 7950 -21120 7960 -21110
rect 8060 -21120 8460 -21068
rect 8690 -21062 8705 -21030
rect 9081 -21062 9093 -21028
rect 8690 -21068 9093 -21062
rect 9657 -21028 10057 -21022
rect 9657 -21062 9669 -21028
rect 10045 -21030 10057 -21028
rect 10293 -21028 10693 -21022
rect 10293 -21030 10305 -21028
rect 10045 -21062 10060 -21030
rect 9657 -21068 10060 -21062
rect 8690 -21120 9090 -21068
rect 9420 -21110 9560 -21100
rect 9420 -21120 9430 -21110
rect 7950 -21220 9430 -21120
rect 7950 -21230 7960 -21220
rect 7820 -21240 7960 -21230
rect 8060 -21240 9090 -21220
rect 9420 -21230 9430 -21220
rect 9550 -21120 9560 -21110
rect 9660 -21120 10060 -21068
rect 10290 -21062 10305 -21030
rect 10681 -21062 10693 -21028
rect 10290 -21068 10693 -21062
rect 11257 -21028 11657 -21022
rect 11257 -21062 11269 -21028
rect 11645 -21030 11657 -21028
rect 11893 -21028 12293 -21022
rect 11893 -21030 11905 -21028
rect 11645 -21062 11660 -21030
rect 11257 -21068 11660 -21062
rect 10290 -21120 10690 -21068
rect 9550 -21220 10690 -21120
rect 9550 -21230 9560 -21220
rect 9420 -21240 9560 -21230
rect 9660 -21240 10690 -21220
rect 1660 -21290 2060 -21240
rect 670 -21296 1093 -21290
rect 670 -21330 705 -21296
rect 1081 -21330 1093 -21296
rect 670 -21336 1093 -21330
rect 1657 -21296 2060 -21290
rect 1657 -21330 1669 -21296
rect 2045 -21330 2060 -21296
rect 2290 -21290 2690 -21240
rect 3260 -21290 3660 -21240
rect 2290 -21296 2693 -21290
rect 2290 -21330 2305 -21296
rect 2681 -21330 2693 -21296
rect 1657 -21336 2057 -21330
rect 2293 -21336 2693 -21330
rect 3257 -21296 3660 -21290
rect 3257 -21330 3269 -21296
rect 3645 -21330 3660 -21296
rect 3890 -21290 4290 -21240
rect 4860 -21290 5260 -21240
rect 3890 -21296 4293 -21290
rect 3890 -21330 3905 -21296
rect 4281 -21330 4293 -21296
rect 3257 -21336 3657 -21330
rect 3893 -21336 4293 -21330
rect 4857 -21296 5260 -21290
rect 4857 -21330 4869 -21296
rect 5245 -21330 5260 -21296
rect 5490 -21290 5890 -21240
rect 6460 -21290 6860 -21240
rect 5490 -21296 5893 -21290
rect 5490 -21330 5505 -21296
rect 5881 -21330 5893 -21296
rect 4857 -21336 5257 -21330
rect 5493 -21336 5893 -21330
rect 6457 -21296 6860 -21290
rect 6457 -21330 6469 -21296
rect 6845 -21330 6860 -21296
rect 7090 -21290 7490 -21240
rect 8060 -21290 8460 -21240
rect 7090 -21296 7493 -21290
rect 7090 -21330 7105 -21296
rect 7481 -21330 7493 -21296
rect 6457 -21336 6857 -21330
rect 7093 -21336 7493 -21330
rect 8057 -21296 8460 -21290
rect 8057 -21330 8069 -21296
rect 8445 -21330 8460 -21296
rect 8690 -21290 9090 -21240
rect 9660 -21290 10060 -21240
rect 8690 -21296 9093 -21290
rect 8690 -21330 8705 -21296
rect 9081 -21330 9093 -21296
rect 8057 -21336 8457 -21330
rect 8693 -21336 9093 -21330
rect 9657 -21296 10060 -21290
rect 9657 -21330 9669 -21296
rect 10045 -21330 10060 -21296
rect 10290 -21290 10690 -21240
rect 11260 -21120 11660 -21068
rect 11890 -21062 11905 -21030
rect 12281 -21062 12293 -21028
rect 11890 -21068 12293 -21062
rect 12857 -21028 13257 -21022
rect 12857 -21062 12869 -21028
rect 13245 -21062 13257 -21028
rect 12857 -21068 13257 -21062
rect 13493 -21028 13893 -21022
rect 13493 -21062 13505 -21028
rect 13881 -21062 13893 -21028
rect 13493 -21068 13893 -21062
rect 14457 -21028 14857 -21022
rect 14457 -21062 14469 -21028
rect 14845 -21062 14857 -21028
rect 14457 -21068 14857 -21062
rect 15093 -21028 15493 -21022
rect 15093 -21062 15105 -21028
rect 15481 -21062 15493 -21028
rect 15093 -21068 15493 -21062
rect 16057 -21028 16457 -21022
rect 16057 -21062 16069 -21028
rect 16445 -21062 16457 -21028
rect 16057 -21068 16457 -21062
rect 16693 -21028 17093 -21022
rect 16693 -21062 16705 -21028
rect 17081 -21062 17093 -21028
rect 16693 -21068 17093 -21062
rect 17657 -21028 18057 -21022
rect 17657 -21062 17669 -21028
rect 18045 -21062 18057 -21028
rect 17657 -21068 18057 -21062
rect 18293 -21028 18693 -21022
rect 18293 -21062 18305 -21028
rect 18681 -21062 18693 -21028
rect 18293 -21068 18693 -21062
rect 19257 -21028 19657 -21022
rect 19257 -21062 19269 -21028
rect 19645 -21062 19657 -21028
rect 19257 -21068 19657 -21062
rect 19893 -21028 20293 -21022
rect 19893 -21062 19905 -21028
rect 20281 -21062 20293 -21028
rect 19893 -21068 20293 -21062
rect 20857 -21028 21257 -21022
rect 20857 -21062 20869 -21028
rect 21245 -21062 21257 -21028
rect 20857 -21068 21257 -21062
rect 21493 -21028 21893 -21022
rect 21493 -21062 21505 -21028
rect 21881 -21062 21893 -21028
rect 21493 -21068 21893 -21062
rect 22457 -21028 22857 -21022
rect 22457 -21062 22469 -21028
rect 22845 -21062 22857 -21028
rect 22457 -21068 22857 -21062
rect 23093 -21028 23493 -21022
rect 23093 -21062 23105 -21028
rect 23481 -21062 23493 -21028
rect 23093 -21068 23493 -21062
rect 24057 -21028 24457 -21022
rect 24057 -21062 24069 -21028
rect 24445 -21062 24457 -21028
rect 24057 -21068 24457 -21062
rect 24693 -21028 25093 -21022
rect 24693 -21062 24705 -21028
rect 25081 -21062 25093 -21028
rect 24693 -21068 25093 -21062
rect 25657 -21028 26057 -21022
rect 25657 -21062 25669 -21028
rect 26045 -21062 26057 -21028
rect 25657 -21068 26057 -21062
rect 26293 -21028 26693 -21022
rect 26293 -21062 26305 -21028
rect 26681 -21062 26693 -21028
rect 26293 -21068 26693 -21062
rect 27257 -21028 27657 -21022
rect 27257 -21062 27269 -21028
rect 27645 -21062 27657 -21028
rect 27257 -21068 27657 -21062
rect 27893 -21028 28293 -21022
rect 27893 -21062 27905 -21028
rect 28281 -21062 28293 -21028
rect 27893 -21068 28293 -21062
rect 28857 -21028 29257 -21022
rect 28857 -21062 28869 -21028
rect 29245 -21062 29257 -21028
rect 28857 -21068 29257 -21062
rect 29493 -21028 29893 -21022
rect 29493 -21062 29505 -21028
rect 29881 -21062 29893 -21028
rect 29493 -21068 29893 -21062
rect 30457 -21028 30857 -21022
rect 30457 -21062 30469 -21028
rect 30845 -21062 30857 -21028
rect 30457 -21068 30857 -21062
rect 31093 -21028 31493 -21022
rect 31093 -21062 31105 -21028
rect 31481 -21062 31493 -21028
rect 32057 -21028 32457 -21022
rect 31093 -21068 31493 -21062
rect 31740 -21040 31820 -21030
rect 11890 -21120 12290 -21068
rect 11260 -21240 12290 -21120
rect 11260 -21290 11660 -21240
rect 10290 -21296 10693 -21290
rect 10290 -21330 10305 -21296
rect 10681 -21330 10693 -21296
rect 9657 -21336 10057 -21330
rect 10293 -21336 10693 -21330
rect 11257 -21296 11660 -21290
rect 11257 -21330 11269 -21296
rect 11645 -21330 11660 -21296
rect 11890 -21290 12290 -21240
rect 15600 -21120 15740 -21110
rect 15600 -21240 15610 -21120
rect 15730 -21130 15740 -21120
rect 16060 -21130 16450 -21068
rect 16700 -21130 17090 -21068
rect 15730 -21230 17090 -21130
rect 15730 -21240 15740 -21230
rect 15600 -21250 15740 -21240
rect 16060 -21290 16450 -21230
rect 16700 -21290 17090 -21230
rect 17200 -21120 17340 -21110
rect 17200 -21240 17210 -21120
rect 17330 -21130 17340 -21120
rect 17660 -21130 18050 -21068
rect 18300 -21130 18690 -21068
rect 17330 -21230 18690 -21130
rect 17330 -21240 17340 -21230
rect 17200 -21250 17340 -21240
rect 17660 -21290 18050 -21230
rect 18300 -21290 18690 -21230
rect 18800 -21120 18940 -21110
rect 18800 -21240 18810 -21120
rect 18930 -21130 18940 -21120
rect 19260 -21130 19650 -21068
rect 19900 -21130 20290 -21068
rect 18930 -21230 20290 -21130
rect 18930 -21240 18940 -21230
rect 18800 -21250 18940 -21240
rect 19260 -21290 19650 -21230
rect 19900 -21290 20290 -21230
rect 20400 -21120 20540 -21110
rect 20400 -21240 20410 -21120
rect 20530 -21130 20540 -21120
rect 20860 -21130 21250 -21068
rect 21500 -21130 21890 -21068
rect 20530 -21230 21890 -21130
rect 20530 -21240 20540 -21230
rect 20400 -21250 20540 -21240
rect 20860 -21290 21250 -21230
rect 21500 -21290 21890 -21230
rect 22000 -21120 22140 -21110
rect 22000 -21240 22010 -21120
rect 22130 -21130 22140 -21120
rect 22460 -21130 22850 -21068
rect 23100 -21130 23490 -21068
rect 22130 -21230 23490 -21130
rect 22130 -21240 22140 -21230
rect 22000 -21250 22140 -21240
rect 22460 -21290 22850 -21230
rect 23100 -21290 23490 -21230
rect 23600 -21120 23740 -21110
rect 23600 -21240 23610 -21120
rect 23730 -21130 23740 -21120
rect 24060 -21130 24450 -21068
rect 24700 -21130 25090 -21068
rect 23730 -21230 25090 -21130
rect 23730 -21240 23740 -21230
rect 23600 -21250 23740 -21240
rect 24060 -21290 24450 -21230
rect 24700 -21290 25090 -21230
rect 25660 -21130 26050 -21068
rect 26300 -21130 26690 -21068
rect 26800 -21120 26940 -21110
rect 26800 -21130 26810 -21120
rect 25660 -21230 26810 -21130
rect 25660 -21290 26050 -21230
rect 26300 -21290 26690 -21230
rect 26800 -21240 26810 -21230
rect 26930 -21130 26940 -21120
rect 27260 -21130 27650 -21068
rect 27900 -21130 28290 -21068
rect 26930 -21230 28290 -21130
rect 26930 -21240 26940 -21230
rect 26800 -21250 26940 -21240
rect 27260 -21290 27650 -21230
rect 27900 -21290 28290 -21230
rect 28400 -21120 28540 -21110
rect 28400 -21240 28410 -21120
rect 28530 -21130 28540 -21120
rect 28860 -21130 29250 -21068
rect 29500 -21130 29890 -21068
rect 30460 -21130 30850 -21068
rect 31100 -21130 31490 -21068
rect 28530 -21230 31490 -21130
rect 28530 -21240 28540 -21230
rect 28400 -21250 28540 -21240
rect 28860 -21290 29250 -21230
rect 29500 -21290 29890 -21230
rect 30460 -21290 30850 -21230
rect 31100 -21290 31490 -21230
rect 11890 -21296 12293 -21290
rect 11890 -21330 11905 -21296
rect 12281 -21330 12293 -21296
rect 11257 -21336 11657 -21330
rect 11893 -21336 12293 -21330
rect 12857 -21296 13257 -21290
rect 12857 -21330 12869 -21296
rect 13245 -21330 13257 -21296
rect 12857 -21336 13257 -21330
rect 13493 -21296 13893 -21290
rect 13493 -21330 13505 -21296
rect 13881 -21330 13893 -21296
rect 13493 -21336 13893 -21330
rect 14457 -21296 14857 -21290
rect 14457 -21330 14469 -21296
rect 14845 -21330 14857 -21296
rect 14457 -21336 14857 -21330
rect 15093 -21296 15493 -21290
rect 15093 -21330 15105 -21296
rect 15481 -21330 15493 -21296
rect 15093 -21336 15493 -21330
rect 16057 -21296 16457 -21290
rect 16057 -21330 16069 -21296
rect 16445 -21330 16457 -21296
rect 16057 -21336 16457 -21330
rect 16693 -21296 17093 -21290
rect 16693 -21330 16705 -21296
rect 17081 -21330 17093 -21296
rect 16693 -21336 17093 -21330
rect 17657 -21296 18057 -21290
rect 17657 -21330 17669 -21296
rect 18045 -21330 18057 -21296
rect 17657 -21336 18057 -21330
rect 18293 -21296 18693 -21290
rect 18293 -21330 18305 -21296
rect 18681 -21330 18693 -21296
rect 18293 -21336 18693 -21330
rect 19257 -21296 19657 -21290
rect 19257 -21330 19269 -21296
rect 19645 -21330 19657 -21296
rect 19257 -21336 19657 -21330
rect 19893 -21296 20293 -21290
rect 19893 -21330 19905 -21296
rect 20281 -21330 20293 -21296
rect 19893 -21336 20293 -21330
rect 20857 -21296 21257 -21290
rect 20857 -21330 20869 -21296
rect 21245 -21330 21257 -21296
rect 20857 -21336 21257 -21330
rect 21493 -21296 21893 -21290
rect 21493 -21330 21505 -21296
rect 21881 -21330 21893 -21296
rect 21493 -21336 21893 -21330
rect 22457 -21296 22857 -21290
rect 22457 -21330 22469 -21296
rect 22845 -21330 22857 -21296
rect 22457 -21336 22857 -21330
rect 23093 -21296 23493 -21290
rect 23093 -21330 23105 -21296
rect 23481 -21330 23493 -21296
rect 23093 -21336 23493 -21330
rect 24057 -21296 24457 -21290
rect 24057 -21330 24069 -21296
rect 24445 -21330 24457 -21296
rect 24057 -21336 24457 -21330
rect 24693 -21296 25093 -21290
rect 24693 -21330 24705 -21296
rect 25081 -21330 25093 -21296
rect 24693 -21336 25093 -21330
rect 25657 -21296 26057 -21290
rect 25657 -21330 25669 -21296
rect 26045 -21330 26057 -21296
rect 25657 -21336 26057 -21330
rect 26293 -21296 26693 -21290
rect 26293 -21330 26305 -21296
rect 26681 -21330 26693 -21296
rect 26293 -21336 26693 -21330
rect 27257 -21296 27657 -21290
rect 27257 -21330 27269 -21296
rect 27645 -21330 27657 -21296
rect 27257 -21336 27657 -21330
rect 27893 -21296 28293 -21290
rect 27893 -21330 27905 -21296
rect 28281 -21330 28293 -21296
rect 27893 -21336 28293 -21330
rect 28857 -21296 29257 -21290
rect 28857 -21330 28869 -21296
rect 29245 -21330 29257 -21296
rect 28857 -21336 29257 -21330
rect 29493 -21296 29893 -21290
rect 29493 -21330 29505 -21296
rect 29881 -21330 29893 -21296
rect 29493 -21336 29893 -21330
rect 30457 -21296 30857 -21290
rect 30457 -21330 30469 -21296
rect 30845 -21330 30857 -21296
rect 30457 -21336 30857 -21330
rect 31093 -21296 31493 -21290
rect 31093 -21330 31105 -21296
rect 31481 -21330 31493 -21296
rect 31740 -21320 31750 -21040
rect 31810 -21130 31820 -21040
rect 32057 -21062 32069 -21028
rect 32445 -21062 32457 -21028
rect 32057 -21068 32457 -21062
rect 32693 -21028 33093 -21022
rect 32693 -21062 32705 -21028
rect 33081 -21062 33093 -21028
rect 32693 -21068 33093 -21062
rect 33657 -21028 34057 -21022
rect 33657 -21062 33669 -21028
rect 34045 -21062 34057 -21028
rect 33657 -21068 34057 -21062
rect 34293 -21028 34693 -21022
rect 34293 -21062 34305 -21028
rect 34681 -21062 34693 -21028
rect 34293 -21068 34693 -21062
rect 35257 -21028 35657 -21022
rect 35257 -21062 35269 -21028
rect 35645 -21062 35657 -21028
rect 35257 -21068 35657 -21062
rect 35893 -21028 36293 -21022
rect 35893 -21062 35905 -21028
rect 36281 -21062 36293 -21028
rect 35893 -21068 36293 -21062
rect 36857 -21028 37257 -21022
rect 36857 -21062 36869 -21028
rect 37245 -21062 37257 -21028
rect 36857 -21068 37257 -21062
rect 37493 -21028 37893 -21022
rect 37493 -21062 37505 -21028
rect 37881 -21062 37893 -21028
rect 37493 -21068 37893 -21062
rect 32060 -21130 32450 -21068
rect 32700 -21130 33090 -21068
rect 31810 -21230 33090 -21130
rect 31810 -21320 31820 -21230
rect 32060 -21290 32450 -21230
rect 32700 -21290 33090 -21230
rect 33660 -21130 34050 -21068
rect 34300 -21130 34690 -21068
rect 35260 -21130 35650 -21068
rect 35900 -21130 36290 -21068
rect 33660 -21230 36290 -21130
rect 33660 -21290 34050 -21230
rect 34300 -21290 34690 -21230
rect 35260 -21290 35650 -21230
rect 35900 -21290 36290 -21230
rect 31740 -21330 31820 -21320
rect 32057 -21296 32457 -21290
rect 32057 -21330 32069 -21296
rect 32445 -21330 32457 -21296
rect 31093 -21336 31493 -21330
rect 32057 -21336 32457 -21330
rect 32693 -21296 33093 -21290
rect 32693 -21330 32705 -21296
rect 33081 -21330 33093 -21296
rect 32693 -21336 33093 -21330
rect 33657 -21296 34057 -21290
rect 33657 -21330 33669 -21296
rect 34045 -21330 34057 -21296
rect 33657 -21336 34057 -21330
rect 34293 -21296 34693 -21290
rect 34293 -21330 34305 -21296
rect 34681 -21330 34693 -21296
rect 34293 -21336 34693 -21330
rect 35257 -21296 35657 -21290
rect 35257 -21330 35269 -21296
rect 35645 -21330 35657 -21296
rect 35257 -21336 35657 -21330
rect 35893 -21296 36293 -21290
rect 35893 -21330 35905 -21296
rect 36281 -21330 36293 -21296
rect 35893 -21336 36293 -21330
rect 36857 -21296 37257 -21290
rect 36857 -21330 36869 -21296
rect 37245 -21330 37257 -21296
rect 36857 -21336 37257 -21330
rect 37493 -21296 37893 -21290
rect 37493 -21330 37505 -21296
rect 37881 -21330 37893 -21296
rect 37493 -21336 37893 -21330
rect 57 -22154 490 -22148
rect 57 -22160 69 -22154
rect 0 -22188 69 -22160
rect 445 -22188 490 -22154
rect 0 -22288 490 -22188
rect 670 -22148 720 -21336
rect 1134 -21396 1180 -21384
rect 1134 -22088 1140 -21396
rect 1174 -22088 1180 -21396
rect 1134 -22100 1180 -22088
rect 1570 -21396 1616 -21384
rect 1570 -22088 1576 -21396
rect 1610 -22088 1616 -21396
rect 1570 -22100 1616 -22088
rect 2098 -21396 2144 -21384
rect 2098 -22088 2104 -21396
rect 2138 -21400 2144 -21396
rect 2206 -21396 2252 -21384
rect 2206 -21400 2212 -21396
rect 2138 -21410 2212 -21400
rect 2138 -22080 2212 -22070
rect 2138 -22088 2144 -22080
rect 2098 -22100 2144 -22088
rect 2206 -22088 2212 -22080
rect 2246 -22088 2252 -21396
rect 2206 -22100 2252 -22088
rect 2734 -21396 2780 -21384
rect 2734 -22088 2740 -21396
rect 2774 -22088 2780 -21396
rect 2734 -22100 2780 -22088
rect 3170 -21396 3216 -21384
rect 3170 -22088 3176 -21396
rect 3210 -22088 3216 -21396
rect 3170 -22100 3216 -22088
rect 3698 -21396 3744 -21384
rect 3698 -22088 3704 -21396
rect 3738 -21400 3744 -21396
rect 3806 -21396 3852 -21384
rect 3806 -21400 3812 -21396
rect 3738 -21410 3812 -21400
rect 3738 -22080 3812 -22070
rect 3738 -22088 3744 -22080
rect 3698 -22100 3744 -22088
rect 3806 -22088 3812 -22080
rect 3846 -22088 3852 -21396
rect 3806 -22100 3852 -22088
rect 4334 -21396 4380 -21384
rect 4334 -22088 4340 -21396
rect 4374 -22088 4380 -21396
rect 4334 -22100 4380 -22088
rect 4770 -21396 4816 -21384
rect 4770 -22088 4776 -21396
rect 4810 -22088 4816 -21396
rect 4770 -22100 4816 -22088
rect 5298 -21396 5344 -21384
rect 5298 -22088 5304 -21396
rect 5338 -21400 5344 -21396
rect 5406 -21396 5452 -21384
rect 5406 -21400 5412 -21396
rect 5338 -21410 5412 -21400
rect 5338 -22080 5412 -22070
rect 5338 -22088 5344 -22080
rect 5298 -22100 5344 -22088
rect 5406 -22088 5412 -22080
rect 5446 -22088 5452 -21396
rect 5406 -22100 5452 -22088
rect 5934 -21396 5980 -21384
rect 5934 -22088 5940 -21396
rect 5974 -22088 5980 -21396
rect 5934 -22100 5980 -22088
rect 6370 -21396 6416 -21384
rect 6370 -22088 6376 -21396
rect 6410 -22088 6416 -21396
rect 6370 -22100 6416 -22088
rect 6898 -21396 6944 -21384
rect 6898 -22088 6904 -21396
rect 6938 -21400 6944 -21396
rect 7006 -21396 7052 -21384
rect 7006 -21400 7012 -21396
rect 6938 -21410 7012 -21400
rect 6938 -22080 7012 -22070
rect 6938 -22088 6944 -22080
rect 6898 -22100 6944 -22088
rect 7006 -22088 7012 -22080
rect 7046 -22088 7052 -21396
rect 7006 -22100 7052 -22088
rect 7534 -21396 7580 -21384
rect 7534 -22088 7540 -21396
rect 7574 -22088 7580 -21396
rect 7534 -22100 7580 -22088
rect 7970 -21396 8016 -21384
rect 7970 -22088 7976 -21396
rect 8010 -22088 8016 -21396
rect 7970 -22100 8016 -22088
rect 8498 -21396 8544 -21384
rect 8498 -22088 8504 -21396
rect 8538 -21400 8544 -21396
rect 8606 -21396 8652 -21384
rect 8606 -21400 8612 -21396
rect 8538 -21410 8612 -21400
rect 8538 -22080 8612 -22070
rect 8538 -22088 8544 -22080
rect 8498 -22100 8544 -22088
rect 8606 -22088 8612 -22080
rect 8646 -22088 8652 -21396
rect 8606 -22100 8652 -22088
rect 9134 -21396 9180 -21384
rect 9134 -22088 9140 -21396
rect 9174 -22088 9180 -21396
rect 9134 -22100 9180 -22088
rect 9570 -21396 9616 -21384
rect 9570 -22088 9576 -21396
rect 9610 -22088 9616 -21396
rect 9570 -22100 9616 -22088
rect 10098 -21396 10144 -21384
rect 10098 -22088 10104 -21396
rect 10138 -21400 10144 -21396
rect 10206 -21396 10252 -21384
rect 10206 -21400 10212 -21396
rect 10138 -21410 10212 -21400
rect 10138 -22080 10212 -22070
rect 10138 -22088 10144 -22080
rect 10098 -22100 10144 -22088
rect 10206 -22088 10212 -22080
rect 10246 -22088 10252 -21396
rect 10206 -22100 10252 -22088
rect 10734 -21396 10780 -21384
rect 10734 -22088 10740 -21396
rect 10774 -22088 10780 -21396
rect 10734 -22100 10780 -22088
rect 11170 -21396 11216 -21384
rect 11170 -22088 11176 -21396
rect 11210 -22088 11216 -21396
rect 11170 -22100 11216 -22088
rect 11698 -21390 11744 -21384
rect 11806 -21390 11852 -21384
rect 11698 -21396 11852 -21390
rect 11698 -22088 11704 -21396
rect 11738 -21400 11812 -21396
rect 11738 -22088 11812 -22080
rect 11846 -22088 11852 -21396
rect 11698 -22090 11852 -22088
rect 11698 -22100 11744 -22090
rect 11806 -22100 11852 -22090
rect 12334 -21396 12380 -21384
rect 12334 -22088 12340 -21396
rect 12374 -22088 12380 -21396
rect 12334 -22100 12380 -22088
rect 12770 -21396 12816 -21384
rect 12770 -22088 12776 -21396
rect 12810 -21650 12816 -21396
rect 13010 -21650 13110 -21336
rect 13298 -21396 13344 -21384
rect 13298 -21650 13304 -21396
rect 12810 -21810 13304 -21650
rect 12810 -22088 12816 -21810
rect 12770 -22100 12816 -22088
rect 13010 -22148 13110 -21810
rect 13298 -22088 13304 -21810
rect 13338 -21650 13344 -21396
rect 13406 -21396 13452 -21384
rect 13406 -21650 13412 -21396
rect 13338 -21810 13412 -21650
rect 13338 -22088 13344 -21810
rect 13298 -22100 13344 -22088
rect 13406 -22088 13412 -21810
rect 13446 -21650 13452 -21396
rect 13640 -21650 13740 -21336
rect 13934 -21396 13980 -21384
rect 13934 -21650 13940 -21396
rect 13446 -21810 13940 -21650
rect 13446 -22088 13452 -21810
rect 13406 -22100 13452 -22088
rect 13640 -22148 13740 -21810
rect 13934 -22088 13940 -21810
rect 13974 -22088 13980 -21396
rect 13934 -22100 13980 -22088
rect 14370 -21396 14416 -21384
rect 14370 -22088 14376 -21396
rect 14410 -21640 14416 -21396
rect 14630 -21640 14700 -21336
rect 14898 -21396 14944 -21384
rect 14898 -21640 14904 -21396
rect 14410 -21780 14904 -21640
rect 14410 -22088 14416 -21780
rect 14370 -22100 14416 -22088
rect 14630 -22148 14700 -21780
rect 14898 -22088 14904 -21780
rect 14938 -21640 14944 -21396
rect 15006 -21396 15052 -21384
rect 15006 -21640 15012 -21396
rect 14938 -21780 15012 -21640
rect 14938 -22088 14944 -21780
rect 14898 -22100 14944 -22088
rect 15006 -22088 15012 -21780
rect 15046 -21640 15052 -21396
rect 15260 -21640 15330 -21336
rect 15534 -21396 15580 -21384
rect 15534 -21640 15540 -21396
rect 15046 -21780 15540 -21640
rect 15046 -22088 15052 -21780
rect 15006 -22100 15052 -22088
rect 15260 -22148 15330 -21780
rect 15534 -22088 15540 -21780
rect 15574 -22088 15580 -21396
rect 15534 -22100 15580 -22088
rect 15970 -21396 16016 -21384
rect 15970 -22088 15976 -21396
rect 16010 -22088 16016 -21396
rect 15970 -22100 16016 -22088
rect 16498 -21390 16544 -21384
rect 16606 -21390 16652 -21384
rect 16498 -21396 16652 -21390
rect 16498 -22088 16504 -21396
rect 16538 -21400 16612 -21396
rect 16538 -22088 16612 -22080
rect 16646 -22088 16652 -21396
rect 16498 -22090 16652 -22088
rect 16498 -22100 16544 -22090
rect 16606 -22100 16652 -22090
rect 17134 -21396 17180 -21384
rect 17134 -22088 17140 -21396
rect 17174 -22088 17180 -21396
rect 17134 -22100 17180 -22088
rect 17570 -21396 17616 -21384
rect 17570 -22088 17576 -21396
rect 17610 -22088 17616 -21396
rect 17570 -22100 17616 -22088
rect 18098 -21390 18144 -21384
rect 18206 -21390 18252 -21384
rect 18098 -21396 18252 -21390
rect 18098 -22088 18104 -21396
rect 18138 -21400 18212 -21396
rect 18138 -22088 18212 -22080
rect 18246 -22088 18252 -21396
rect 18098 -22090 18252 -22088
rect 18098 -22100 18144 -22090
rect 18206 -22100 18252 -22090
rect 18734 -21396 18780 -21384
rect 18734 -22088 18740 -21396
rect 18774 -22088 18780 -21396
rect 18734 -22100 18780 -22088
rect 19170 -21396 19216 -21384
rect 19170 -22088 19176 -21396
rect 19210 -22088 19216 -21396
rect 19170 -22100 19216 -22088
rect 19698 -21390 19744 -21384
rect 19806 -21390 19852 -21384
rect 19698 -21396 19852 -21390
rect 19698 -22088 19704 -21396
rect 19738 -21400 19812 -21396
rect 19738 -22088 19812 -22080
rect 19846 -22088 19852 -21396
rect 19698 -22090 19852 -22088
rect 19698 -22100 19744 -22090
rect 19806 -22100 19852 -22090
rect 20334 -21396 20380 -21384
rect 20334 -22088 20340 -21396
rect 20374 -22088 20380 -21396
rect 20334 -22100 20380 -22088
rect 20770 -21396 20816 -21384
rect 20770 -22088 20776 -21396
rect 20810 -22088 20816 -21396
rect 20770 -22100 20816 -22088
rect 21298 -21390 21344 -21384
rect 21406 -21390 21452 -21384
rect 21298 -21396 21452 -21390
rect 21298 -22088 21304 -21396
rect 21338 -21400 21412 -21396
rect 21338 -22088 21412 -22080
rect 21446 -22088 21452 -21396
rect 21298 -22090 21452 -22088
rect 21298 -22100 21344 -22090
rect 21406 -22100 21452 -22090
rect 21934 -21396 21980 -21384
rect 21934 -22088 21940 -21396
rect 21974 -22088 21980 -21396
rect 21934 -22100 21980 -22088
rect 22370 -21396 22416 -21384
rect 22370 -22088 22376 -21396
rect 22410 -22088 22416 -21396
rect 22370 -22100 22416 -22088
rect 22898 -21390 22944 -21384
rect 23006 -21390 23052 -21384
rect 22898 -21396 23052 -21390
rect 22898 -22088 22904 -21396
rect 22938 -21400 23012 -21396
rect 22938 -22088 23012 -22080
rect 23046 -22088 23052 -21396
rect 22898 -22090 23052 -22088
rect 22898 -22100 22944 -22090
rect 23006 -22100 23052 -22090
rect 23534 -21396 23580 -21384
rect 23534 -22088 23540 -21396
rect 23574 -22088 23580 -21396
rect 23534 -22100 23580 -22088
rect 23970 -21396 24016 -21384
rect 23970 -22088 23976 -21396
rect 24010 -22088 24016 -21396
rect 23970 -22100 24016 -22088
rect 24498 -21390 24544 -21384
rect 24606 -21390 24652 -21384
rect 24498 -21396 24652 -21390
rect 24498 -22088 24504 -21396
rect 24538 -21400 24612 -21396
rect 24538 -22088 24612 -22080
rect 24646 -22088 24652 -21396
rect 24498 -22090 24652 -22088
rect 24498 -22100 24544 -22090
rect 24606 -22100 24652 -22090
rect 25134 -21396 25180 -21384
rect 25134 -22088 25140 -21396
rect 25174 -22088 25180 -21396
rect 25134 -22100 25180 -22088
rect 25570 -21396 25616 -21384
rect 25570 -22088 25576 -21396
rect 25610 -22088 25616 -21396
rect 25570 -22100 25616 -22088
rect 26098 -21390 26144 -21384
rect 26206 -21390 26252 -21384
rect 26098 -21396 26252 -21390
rect 26098 -22088 26104 -21396
rect 26138 -21400 26212 -21396
rect 26138 -22088 26212 -22080
rect 26246 -22088 26252 -21396
rect 26098 -22090 26252 -22088
rect 26098 -22100 26144 -22090
rect 26206 -22100 26252 -22090
rect 26734 -21396 26780 -21384
rect 26734 -22088 26740 -21396
rect 26774 -22088 26780 -21396
rect 26734 -22100 26780 -22088
rect 27170 -21396 27216 -21384
rect 27170 -22088 27176 -21396
rect 27210 -22088 27216 -21396
rect 27170 -22100 27216 -22088
rect 27698 -21390 27744 -21384
rect 27806 -21390 27852 -21384
rect 27698 -21396 27852 -21390
rect 27698 -22088 27704 -21396
rect 27738 -21400 27812 -21396
rect 27738 -22088 27812 -22080
rect 27846 -22088 27852 -21396
rect 27698 -22090 27852 -22088
rect 27698 -22100 27744 -22090
rect 27806 -22100 27852 -22090
rect 28334 -21396 28380 -21384
rect 28334 -22088 28340 -21396
rect 28374 -22088 28380 -21396
rect 28334 -22100 28380 -22088
rect 28770 -21396 28816 -21384
rect 28770 -22088 28776 -21396
rect 28810 -22088 28816 -21396
rect 28770 -22100 28816 -22088
rect 29298 -21390 29344 -21384
rect 29406 -21390 29452 -21384
rect 29298 -21396 29452 -21390
rect 29298 -22088 29304 -21396
rect 29338 -21400 29412 -21396
rect 29338 -22088 29412 -22080
rect 29446 -22088 29452 -21396
rect 29298 -22090 29452 -22088
rect 29298 -22100 29344 -22090
rect 29406 -22100 29452 -22090
rect 29934 -21396 29980 -21384
rect 29934 -22088 29940 -21396
rect 29974 -22088 29980 -21396
rect 29934 -22100 29980 -22088
rect 30370 -21396 30416 -21384
rect 30370 -22088 30376 -21396
rect 30410 -22088 30416 -21396
rect 30370 -22100 30416 -22088
rect 30898 -21390 30944 -21384
rect 31006 -21390 31052 -21384
rect 30898 -21396 31052 -21390
rect 30898 -22088 30904 -21396
rect 30938 -21400 31012 -21396
rect 30938 -22088 31012 -22080
rect 31046 -22088 31052 -21396
rect 30898 -22090 31052 -22088
rect 30898 -22100 30944 -22090
rect 31006 -22100 31052 -22090
rect 31534 -21396 31580 -21384
rect 31534 -22088 31540 -21396
rect 31574 -22088 31580 -21396
rect 31534 -22100 31580 -22088
rect 31970 -21396 32016 -21384
rect 31970 -22088 31976 -21396
rect 32010 -22088 32016 -21396
rect 31970 -22100 32016 -22088
rect 32498 -21390 32544 -21384
rect 32606 -21390 32652 -21384
rect 32498 -21396 32652 -21390
rect 32498 -22088 32504 -21396
rect 32538 -21400 32612 -21396
rect 32538 -22088 32612 -22080
rect 32646 -22088 32652 -21396
rect 32498 -22090 32652 -22088
rect 32498 -22100 32544 -22090
rect 32606 -22100 32652 -22090
rect 33134 -21396 33180 -21384
rect 33134 -22088 33140 -21396
rect 33174 -22088 33180 -21396
rect 33134 -22100 33180 -22088
rect 33570 -21396 33616 -21384
rect 33570 -22088 33576 -21396
rect 33610 -22088 33616 -21396
rect 33570 -22100 33616 -22088
rect 34098 -21390 34144 -21384
rect 34206 -21390 34252 -21384
rect 34098 -21396 34252 -21390
rect 34098 -22088 34104 -21396
rect 34138 -21400 34212 -21396
rect 34138 -22088 34212 -22080
rect 34246 -22088 34252 -21396
rect 34098 -22090 34252 -22088
rect 34098 -22100 34144 -22090
rect 34206 -22100 34252 -22090
rect 34734 -21396 34780 -21384
rect 34734 -22088 34740 -21396
rect 34774 -22088 34780 -21396
rect 34734 -22100 34780 -22088
rect 35170 -21396 35216 -21384
rect 35170 -22088 35176 -21396
rect 35210 -22088 35216 -21396
rect 35170 -22100 35216 -22088
rect 35698 -21390 35744 -21384
rect 35806 -21390 35852 -21384
rect 35698 -21396 35852 -21390
rect 35698 -22088 35704 -21396
rect 35738 -21400 35812 -21396
rect 35738 -22088 35812 -22080
rect 35846 -22088 35852 -21396
rect 35698 -22090 35852 -22088
rect 35698 -22100 35744 -22090
rect 35806 -22100 35852 -22090
rect 36334 -21396 36380 -21384
rect 36334 -22088 36340 -21396
rect 36374 -22088 36380 -21396
rect 36334 -22100 36380 -22088
rect 36770 -21396 36816 -21384
rect 36770 -22088 36776 -21396
rect 36810 -22088 36816 -21396
rect 36770 -22100 36816 -22088
rect 37298 -21396 37344 -21384
rect 37298 -22088 37304 -21396
rect 37338 -22088 37344 -21396
rect 37298 -22100 37344 -22088
rect 37406 -21396 37452 -21384
rect 37406 -22088 37412 -21396
rect 37446 -22088 37452 -21396
rect 37406 -22100 37452 -22088
rect 37934 -21396 37980 -21384
rect 37934 -22088 37940 -21396
rect 37974 -22088 37980 -21396
rect 37934 -22100 37980 -22088
rect 33200 -22140 33300 -22130
rect 670 -22154 1093 -22148
rect 670 -22188 705 -22154
rect 1081 -22160 1093 -22154
rect 1657 -22154 2057 -22148
rect 1657 -22160 1669 -22154
rect 1081 -22188 1669 -22160
rect 2045 -22160 2057 -22154
rect 2293 -22154 2693 -22148
rect 2293 -22160 2305 -22154
rect 2045 -22188 2305 -22160
rect 2681 -22160 2693 -22154
rect 3257 -22154 3657 -22148
rect 3257 -22160 3269 -22154
rect 2681 -22188 3269 -22160
rect 3645 -22160 3657 -22154
rect 3893 -22154 4293 -22148
rect 3893 -22160 3905 -22154
rect 3645 -22188 3905 -22160
rect 4281 -22160 4293 -22154
rect 4857 -22154 5257 -22148
rect 4857 -22160 4869 -22154
rect 4281 -22188 4869 -22160
rect 5245 -22160 5257 -22154
rect 5493 -22154 5893 -22148
rect 5493 -22160 5505 -22154
rect 5245 -22188 5505 -22160
rect 5881 -22160 5893 -22154
rect 6457 -22154 6857 -22148
rect 6457 -22160 6469 -22154
rect 5881 -22188 6469 -22160
rect 6845 -22160 6857 -22154
rect 7093 -22154 7493 -22148
rect 7093 -22160 7105 -22154
rect 6845 -22188 7105 -22160
rect 7481 -22160 7493 -22154
rect 8057 -22154 8457 -22148
rect 8057 -22160 8069 -22154
rect 7481 -22188 8069 -22160
rect 8445 -22160 8457 -22154
rect 8693 -22154 9093 -22148
rect 8693 -22160 8705 -22154
rect 8445 -22188 8705 -22160
rect 9081 -22160 9093 -22154
rect 9657 -22154 10057 -22148
rect 9657 -22160 9669 -22154
rect 9081 -22188 9669 -22160
rect 10045 -22160 10057 -22154
rect 10293 -22154 10693 -22148
rect 10293 -22160 10305 -22154
rect 10045 -22188 10305 -22160
rect 10681 -22160 10693 -22154
rect 11257 -22154 11657 -22148
rect 11257 -22160 11269 -22154
rect 10681 -22188 11269 -22160
rect 11645 -22160 11657 -22154
rect 11893 -22154 12293 -22148
rect 11893 -22160 11905 -22154
rect 11645 -22188 11905 -22160
rect 12281 -22160 12293 -22154
rect 12857 -22154 13257 -22148
rect 12857 -22160 12869 -22154
rect 12281 -22188 12869 -22160
rect 13245 -22160 13257 -22154
rect 13493 -22154 13893 -22148
rect 13493 -22160 13505 -22154
rect 13245 -22188 13505 -22160
rect 13881 -22160 13893 -22154
rect 14457 -22154 14857 -22148
rect 14457 -22160 14469 -22154
rect 13881 -22188 14469 -22160
rect 14845 -22160 14857 -22154
rect 15093 -22154 15493 -22148
rect 15093 -22160 15105 -22154
rect 14845 -22188 15105 -22160
rect 15481 -22160 15493 -22154
rect 16057 -22154 16457 -22148
rect 16057 -22160 16069 -22154
rect 15481 -22188 16069 -22160
rect 16445 -22160 16457 -22154
rect 16693 -22154 17093 -22148
rect 16693 -22160 16705 -22154
rect 16445 -22188 16705 -22160
rect 17081 -22160 17093 -22154
rect 17657 -22154 18057 -22148
rect 17657 -22160 17669 -22154
rect 17081 -22188 17669 -22160
rect 18045 -22160 18057 -22154
rect 18293 -22154 18693 -22148
rect 18293 -22160 18305 -22154
rect 18045 -22188 18305 -22160
rect 18681 -22160 18693 -22154
rect 19257 -22154 19657 -22148
rect 19257 -22160 19269 -22154
rect 18681 -22188 19269 -22160
rect 19645 -22160 19657 -22154
rect 19893 -22154 20293 -22148
rect 19893 -22160 19905 -22154
rect 19645 -22188 19905 -22160
rect 20281 -22160 20293 -22154
rect 20857 -22154 21257 -22148
rect 20857 -22160 20869 -22154
rect 20281 -22188 20869 -22160
rect 21245 -22160 21257 -22154
rect 21493 -22154 21893 -22148
rect 21493 -22160 21505 -22154
rect 21245 -22188 21505 -22160
rect 21881 -22160 21893 -22154
rect 22457 -22154 22857 -22148
rect 22457 -22160 22469 -22154
rect 21881 -22188 22469 -22160
rect 22845 -22160 22857 -22154
rect 23093 -22154 23493 -22148
rect 23093 -22160 23105 -22154
rect 22845 -22188 23105 -22160
rect 23481 -22160 23493 -22154
rect 24057 -22154 24457 -22148
rect 24057 -22160 24069 -22154
rect 23481 -22188 24069 -22160
rect 24445 -22160 24457 -22154
rect 24693 -22154 25093 -22148
rect 24693 -22160 24705 -22154
rect 24445 -22188 24705 -22160
rect 25081 -22160 25093 -22154
rect 25657 -22154 26057 -22148
rect 25657 -22160 25669 -22154
rect 25081 -22188 25669 -22160
rect 26045 -22160 26057 -22154
rect 26293 -22154 26693 -22148
rect 26293 -22160 26305 -22154
rect 26045 -22188 26305 -22160
rect 26681 -22160 26693 -22154
rect 27257 -22154 27657 -22148
rect 27257 -22160 27269 -22154
rect 26681 -22188 27269 -22160
rect 27645 -22160 27657 -22154
rect 27893 -22154 28293 -22148
rect 27893 -22160 27905 -22154
rect 27645 -22188 27905 -22160
rect 28281 -22160 28293 -22154
rect 28857 -22154 29257 -22148
rect 28857 -22160 28869 -22154
rect 28281 -22188 28869 -22160
rect 29245 -22160 29257 -22154
rect 29493 -22154 29893 -22148
rect 29493 -22160 29505 -22154
rect 29245 -22188 29505 -22160
rect 29881 -22160 29893 -22154
rect 30457 -22154 30857 -22148
rect 30457 -22160 30469 -22154
rect 29881 -22188 30469 -22160
rect 30845 -22160 30857 -22154
rect 31093 -22154 31493 -22148
rect 31093 -22160 31105 -22154
rect 30845 -22188 31105 -22160
rect 31481 -22188 31493 -22154
rect 670 -22194 31493 -22188
rect 32057 -22154 32457 -22148
rect 32057 -22188 32069 -22154
rect 32445 -22160 32457 -22154
rect 32693 -22150 33093 -22148
rect 33200 -22150 33210 -22140
rect 32693 -22154 33210 -22150
rect 32693 -22160 32705 -22154
rect 32445 -22188 32705 -22160
rect 33081 -22188 33210 -22154
rect 32057 -22194 33210 -22188
rect 670 -22282 31480 -22194
rect 32060 -22240 33210 -22194
rect 33290 -22240 33300 -22140
rect 33657 -22154 34057 -22148
rect 33657 -22188 33669 -22154
rect 34045 -22160 34057 -22154
rect 34293 -22154 34693 -22148
rect 34293 -22160 34305 -22154
rect 34045 -22170 34305 -22160
rect 34681 -22160 34693 -22154
rect 35257 -22154 35657 -22148
rect 35257 -22160 35269 -22154
rect 34681 -22188 35269 -22160
rect 35645 -22160 35657 -22154
rect 35893 -22154 36293 -22148
rect 35893 -22160 35905 -22154
rect 35645 -22188 35905 -22160
rect 36281 -22188 36293 -22154
rect 33657 -22194 34020 -22188
rect 32060 -22250 33300 -22240
rect 33660 -22240 34020 -22194
rect 34360 -22194 36293 -22188
rect 36857 -22154 37257 -22148
rect 36857 -22188 36869 -22154
rect 37245 -22188 37257 -22154
rect 36857 -22194 37257 -22188
rect 37493 -22154 37893 -22148
rect 37493 -22188 37505 -22154
rect 37881 -22188 37893 -22154
rect 37493 -22194 37893 -22188
rect 34360 -22240 36290 -22194
rect 33660 -22250 34000 -22240
rect 34320 -22250 36290 -22240
rect 670 -22288 31549 -22282
rect 0 -22322 13 -22288
rect 1137 -22322 1613 -22288
rect 2737 -22322 3213 -22288
rect 4337 -22322 4813 -22288
rect 5937 -22322 6413 -22288
rect 7537 -22322 8013 -22288
rect 9137 -22322 9613 -22288
rect 10737 -22322 11213 -22288
rect 12337 -22322 12813 -22288
rect 13937 -22322 14413 -22288
rect 15537 -22322 16013 -22288
rect 17137 -22322 17613 -22288
rect 18737 -22322 19213 -22288
rect 20337 -22322 20813 -22288
rect 21937 -22322 22413 -22288
rect 23537 -22322 24013 -22288
rect 25137 -22322 25613 -22288
rect 26737 -22322 27213 -22288
rect 28337 -22322 28813 -22288
rect 29937 -22322 30413 -22288
rect 31537 -22300 31549 -22288
rect 32001 -22288 33149 -22282
rect 32001 -22300 32013 -22288
rect 31537 -22322 32013 -22300
rect 33137 -22300 33149 -22288
rect 33601 -22288 34749 -22282
rect 33601 -22300 33613 -22288
rect 33137 -22322 33613 -22300
rect 34737 -22300 34749 -22288
rect 35201 -22288 36349 -22282
rect 35201 -22300 35213 -22288
rect 34737 -22322 35213 -22300
rect 36337 -22300 36349 -22288
rect 36801 -22288 37949 -22282
rect 36801 -22300 36813 -22288
rect 36337 -22322 36813 -22300
rect 37937 -22322 37949 -22288
rect 0 -22380 490 -22322
rect 670 -22328 37949 -22322
rect 670 -22380 37940 -22328
rect 0 -22390 37940 -22380
rect 0 -22420 32490 -22390
rect 36180 -22420 37940 -22390
rect 28500 -22672 28540 -22420
rect 28820 -22672 28860 -22420
rect 28346 -22684 28392 -22672
rect 28346 -22720 28352 -22684
rect 28140 -22730 28352 -22720
rect 28140 -22870 28150 -22730
rect 28140 -22880 28352 -22870
rect 28346 -23460 28352 -22880
rect 28386 -23460 28392 -22684
rect 28500 -22684 28550 -22672
rect 28500 -22760 28510 -22684
rect 28346 -23472 28392 -23460
rect 28504 -23460 28510 -22760
rect 28544 -23460 28550 -22684
rect 28662 -22684 28708 -22672
rect 28662 -22730 28668 -22684
rect 28620 -22740 28668 -22730
rect 28702 -22730 28708 -22684
rect 28820 -22684 28866 -22672
rect 28702 -22740 28750 -22730
rect 28620 -22870 28630 -22740
rect 28740 -22870 28750 -22740
rect 28620 -22880 28668 -22870
rect 28504 -23472 28550 -23460
rect 28662 -23460 28668 -22880
rect 28702 -22880 28750 -22870
rect 28702 -23460 28708 -22880
rect 28662 -23472 28708 -23460
rect 28820 -23460 28826 -22684
rect 28860 -23460 28866 -22684
rect 28820 -23472 28866 -23460
rect 28978 -22684 29024 -22672
rect 28978 -23460 28984 -22684
rect 29018 -22720 29024 -22684
rect 29018 -22730 29230 -22720
rect 29220 -22870 29230 -22730
rect 29018 -22880 29230 -22870
rect 29018 -23460 29024 -22880
rect 31890 -23240 32390 -22420
rect 32620 -22430 33310 -22420
rect 32620 -22490 32630 -22430
rect 33300 -22490 33310 -22430
rect 32620 -22500 33310 -22490
rect 34030 -22430 34320 -22420
rect 34030 -22490 34040 -22430
rect 34310 -22490 34320 -22430
rect 34030 -22500 34320 -22490
rect 32492 -22515 32538 -22503
rect 32492 -23131 32498 -22515
rect 32532 -23131 32538 -22515
rect 32699 -22542 32757 -22536
rect 32699 -22576 32711 -22542
rect 32745 -22576 32757 -22542
rect 32699 -22582 32757 -22576
rect 32626 -22635 32672 -22623
rect 32626 -22840 32632 -22635
rect 32492 -23143 32538 -23131
rect 32620 -23011 32632 -22840
rect 32666 -23011 32672 -22635
rect 32620 -23023 32672 -23011
rect 32620 -23202 32660 -23023
rect 32710 -23060 32750 -22582
rect 32790 -22623 32820 -22500
rect 32857 -22542 32915 -22536
rect 32857 -22576 32869 -22542
rect 32903 -22576 32915 -22542
rect 32857 -22582 32915 -22576
rect 33015 -22542 33073 -22536
rect 33015 -22576 33027 -22542
rect 33061 -22576 33073 -22542
rect 33015 -22582 33073 -22576
rect 32784 -22635 32830 -22623
rect 32784 -23011 32790 -22635
rect 32824 -23011 32830 -22635
rect 32784 -23023 32830 -23011
rect 32870 -23060 32910 -22582
rect 32942 -22635 32988 -22623
rect 32942 -23011 32948 -22635
rect 32982 -23011 32988 -22635
rect 32942 -23023 32988 -23011
rect 32690 -23070 32920 -23060
rect 32690 -23150 32700 -23070
rect 32910 -23150 32920 -23070
rect 32690 -23160 32920 -23150
rect 32950 -23202 32980 -23023
rect 33030 -23060 33070 -22582
rect 33110 -22623 33140 -22500
rect 33392 -22515 33438 -22503
rect 33173 -22542 33231 -22536
rect 33173 -22576 33185 -22542
rect 33219 -22576 33231 -22542
rect 33173 -22582 33231 -22576
rect 33100 -22635 33146 -22623
rect 33100 -23011 33106 -22635
rect 33140 -23011 33146 -22635
rect 33100 -23023 33146 -23011
rect 33180 -23060 33220 -22582
rect 33258 -22630 33304 -22623
rect 33258 -22635 33330 -22630
rect 33258 -23011 33264 -22635
rect 33298 -23011 33330 -22635
rect 33258 -23023 33330 -23011
rect 33010 -23070 33240 -23060
rect 33010 -23150 33020 -23070
rect 33230 -23150 33240 -23070
rect 33010 -23160 33240 -23150
rect 33290 -23202 33330 -23023
rect 33392 -23131 33398 -22515
rect 33432 -23131 33438 -22515
rect 33392 -23143 33438 -23131
rect 33862 -22535 33908 -22523
rect 33862 -23151 33868 -22535
rect 33902 -23151 33908 -22535
rect 34069 -22562 34127 -22556
rect 34069 -22596 34081 -22562
rect 34115 -22596 34127 -22562
rect 34069 -22602 34127 -22596
rect 33996 -22655 34042 -22643
rect 33996 -23031 34002 -22655
rect 34036 -23031 34042 -22655
rect 33996 -23043 34042 -23031
rect 33862 -23163 33908 -23151
rect 32607 -23208 33330 -23202
rect 32607 -23240 32619 -23208
rect 31890 -23242 32619 -23240
rect 33311 -23240 33330 -23208
rect 34000 -23222 34030 -23043
rect 34080 -23084 34120 -22602
rect 34160 -22643 34190 -22500
rect 34446 -22535 34492 -22523
rect 34227 -22562 34285 -22556
rect 34227 -22596 34239 -22562
rect 34273 -22596 34285 -22562
rect 34227 -22602 34285 -22596
rect 34154 -22655 34200 -22643
rect 34154 -23031 34160 -22655
rect 34194 -23031 34200 -22655
rect 34154 -23043 34200 -23031
rect 34240 -23084 34280 -22602
rect 34312 -22655 34358 -22643
rect 34312 -23031 34318 -22655
rect 34352 -22960 34358 -22655
rect 34352 -23031 34380 -22960
rect 34312 -23043 34380 -23031
rect 34069 -23090 34127 -23084
rect 34227 -23090 34285 -23084
rect 34060 -23100 34081 -23090
rect 34115 -23100 34239 -23090
rect 34273 -23100 34310 -23090
rect 34060 -23160 34070 -23100
rect 34300 -23160 34310 -23100
rect 34060 -23170 34310 -23160
rect 34350 -23222 34380 -23043
rect 34446 -23151 34452 -22535
rect 34486 -23151 34492 -22535
rect 34446 -23163 34492 -23151
rect 33945 -23228 34409 -23222
rect 33945 -23240 33957 -23228
rect 33311 -23242 33957 -23240
rect 31890 -23262 33957 -23242
rect 34397 -23240 34409 -23228
rect 34397 -23262 34480 -23240
rect 31890 -23370 34480 -23262
rect 32300 -23460 34480 -23370
rect 28978 -23472 29024 -23460
rect 28402 -23519 28494 -23513
rect 28402 -23520 28414 -23519
rect 28370 -23553 28414 -23520
rect 28482 -23520 28494 -23519
rect 28560 -23519 28652 -23513
rect 28560 -23520 28572 -23519
rect 28482 -23553 28572 -23520
rect 28640 -23520 28652 -23519
rect 28718 -23519 28810 -23513
rect 28718 -23520 28730 -23519
rect 28640 -23553 28730 -23520
rect 28798 -23520 28810 -23519
rect 28876 -23519 28968 -23513
rect 28876 -23520 28888 -23519
rect 28798 -23553 28888 -23520
rect 28956 -23520 28968 -23519
rect 29740 -23520 29890 -23510
rect 28956 -23553 29750 -23520
rect 28370 -23590 29750 -23553
rect 29880 -23590 29890 -23520
rect 29740 -23600 29890 -23590
rect 32540 -23645 33040 -23460
rect 33400 -23560 33920 -23550
rect 33400 -23590 33410 -23560
rect 33170 -23620 33410 -23590
rect 33910 -23590 33920 -23560
rect 34620 -23560 37030 -23550
rect 33910 -23620 34150 -23590
rect 33170 -23630 34150 -23620
rect 34620 -23620 35000 -23560
rect 37020 -23620 37030 -23560
rect 34620 -23630 35180 -23620
rect 35210 -23630 37030 -23620
rect 32540 -23657 33076 -23645
rect 32540 -24273 33036 -23657
rect 33070 -24273 33076 -23657
rect 33170 -23765 33200 -23630
rect 33237 -23684 33295 -23678
rect 33237 -23718 33249 -23684
rect 33283 -23718 33295 -23684
rect 33237 -23724 33295 -23718
rect 33395 -23684 33453 -23678
rect 33395 -23718 33407 -23684
rect 33441 -23718 33453 -23684
rect 33395 -23724 33453 -23718
rect 33164 -23777 33210 -23765
rect 33164 -24153 33170 -23777
rect 33204 -24153 33210 -23777
rect 33164 -24165 33210 -24153
rect 33250 -24206 33290 -23724
rect 33322 -23777 33368 -23765
rect 33322 -24153 33328 -23777
rect 33362 -24153 33368 -23777
rect 33322 -24165 33368 -24153
rect 33237 -24210 33295 -24206
rect 32540 -24285 33076 -24273
rect 33160 -24212 33295 -24210
rect 33160 -24220 33249 -24212
rect 33160 -24280 33170 -24220
rect 33283 -24246 33295 -24212
rect 33280 -24252 33295 -24246
rect 33280 -24280 33290 -24252
rect 32540 -24360 33040 -24285
rect 33160 -24290 33290 -24280
rect 33330 -24344 33360 -24165
rect 33410 -24206 33440 -23724
rect 33490 -23765 33520 -23630
rect 33553 -23684 33611 -23678
rect 33553 -23718 33565 -23684
rect 33599 -23718 33611 -23684
rect 33553 -23724 33611 -23718
rect 33711 -23684 33769 -23678
rect 33711 -23718 33723 -23684
rect 33757 -23718 33769 -23684
rect 33711 -23724 33769 -23718
rect 33480 -23777 33526 -23765
rect 33480 -24153 33486 -23777
rect 33520 -24153 33526 -23777
rect 33480 -24165 33526 -24153
rect 33570 -24206 33600 -23724
rect 33638 -23777 33684 -23765
rect 33638 -24153 33644 -23777
rect 33678 -24153 33684 -23777
rect 33638 -24165 33684 -24153
rect 33395 -24210 33453 -24206
rect 33553 -24210 33611 -24206
rect 33395 -24212 33611 -24210
rect 33395 -24246 33407 -24212
rect 33441 -24220 33565 -24212
rect 33599 -24220 33611 -24212
rect 33395 -24252 33410 -24246
rect 33400 -24280 33410 -24252
rect 33600 -24252 33611 -24220
rect 33600 -24280 33610 -24252
rect 33400 -24290 33610 -24280
rect 33650 -24344 33680 -24165
rect 33730 -24206 33760 -23724
rect 33810 -23765 33840 -23630
rect 33869 -23684 33927 -23678
rect 33869 -23718 33881 -23684
rect 33915 -23718 33927 -23684
rect 33869 -23724 33927 -23718
rect 34027 -23684 34085 -23678
rect 34027 -23718 34039 -23684
rect 34073 -23718 34085 -23684
rect 34027 -23724 34085 -23718
rect 33796 -23777 33842 -23765
rect 33796 -24153 33802 -23777
rect 33836 -24153 33842 -23777
rect 33796 -24165 33842 -24153
rect 33890 -24206 33920 -23724
rect 33954 -23777 34000 -23765
rect 33954 -24153 33960 -23777
rect 33994 -24153 34000 -23777
rect 33954 -24165 34000 -24153
rect 33711 -24210 33769 -24206
rect 33869 -24210 33927 -24206
rect 33711 -24212 33930 -24210
rect 33711 -24246 33723 -24212
rect 33757 -24220 33881 -24212
rect 33915 -24220 33930 -24212
rect 33711 -24252 33730 -24246
rect 33720 -24280 33730 -24252
rect 33920 -24280 33930 -24220
rect 33720 -24290 33930 -24280
rect 33960 -24344 33990 -24165
rect 34040 -24206 34080 -23724
rect 34120 -23765 34150 -23630
rect 34246 -23657 34292 -23645
rect 34112 -23777 34158 -23765
rect 34112 -24153 34118 -23777
rect 34152 -24153 34158 -23777
rect 34112 -24165 34158 -24153
rect 34027 -24210 34085 -24206
rect 34027 -24212 34150 -24210
rect 34027 -24246 34039 -24212
rect 34073 -24220 34150 -24212
rect 34027 -24252 34040 -24246
rect 34030 -24280 34040 -24252
rect 34140 -24280 34150 -24220
rect 34030 -24290 34150 -24280
rect 34246 -24273 34252 -23657
rect 34286 -24273 34292 -23657
rect 34246 -24285 34292 -24273
rect 34402 -23655 34448 -23643
rect 34402 -24271 34408 -23655
rect 34442 -24271 34448 -23655
rect 34609 -23682 34667 -23676
rect 34609 -23716 34621 -23682
rect 34655 -23716 34667 -23682
rect 34609 -23722 34667 -23716
rect 34536 -23775 34582 -23763
rect 34536 -24151 34542 -23775
rect 34576 -24151 34582 -23775
rect 34536 -24163 34582 -24151
rect 34402 -24283 34448 -24271
rect 33176 -24350 34146 -24344
rect 33176 -24360 33188 -24350
rect 32540 -24384 33188 -24360
rect 34134 -24360 34146 -24350
rect 34540 -24360 34570 -24163
rect 34620 -24204 34650 -23722
rect 34700 -23763 34730 -23630
rect 34767 -23682 34825 -23676
rect 34767 -23716 34779 -23682
rect 34813 -23716 34825 -23682
rect 34767 -23722 34825 -23716
rect 34925 -23682 34983 -23676
rect 34925 -23716 34937 -23682
rect 34971 -23716 34983 -23682
rect 34925 -23722 34983 -23716
rect 34694 -23775 34740 -23763
rect 34694 -24151 34700 -23775
rect 34734 -24151 34740 -23775
rect 34694 -24163 34740 -24151
rect 34780 -24204 34810 -23722
rect 34852 -23775 34898 -23763
rect 34852 -24151 34858 -23775
rect 34892 -24151 34898 -23775
rect 34852 -24163 34898 -24151
rect 34609 -24210 34667 -24204
rect 34767 -24210 34825 -24204
rect 34609 -24220 34621 -24210
rect 34655 -24220 34779 -24210
rect 34609 -24250 34620 -24220
rect 34770 -24244 34779 -24220
rect 34813 -24244 34825 -24210
rect 34610 -24280 34620 -24250
rect 34770 -24250 34825 -24244
rect 34770 -24280 34820 -24250
rect 34610 -24290 34820 -24280
rect 34860 -24342 34890 -24163
rect 34940 -24204 34970 -23722
rect 35020 -23763 35050 -23630
rect 35083 -23682 35141 -23676
rect 35083 -23716 35095 -23682
rect 35129 -23716 35141 -23682
rect 35083 -23722 35141 -23716
rect 35241 -23682 35299 -23676
rect 35241 -23716 35253 -23682
rect 35287 -23716 35299 -23682
rect 35241 -23722 35299 -23716
rect 35010 -23775 35056 -23763
rect 35010 -24151 35016 -23775
rect 35050 -24151 35056 -23775
rect 35010 -24163 35056 -24151
rect 35100 -24204 35130 -23722
rect 35168 -23775 35214 -23763
rect 35168 -24151 35174 -23775
rect 35208 -24151 35214 -23775
rect 35168 -24163 35214 -24151
rect 34925 -24210 34983 -24204
rect 35083 -24210 35141 -24204
rect 34925 -24244 34937 -24210
rect 34971 -24220 35095 -24210
rect 35129 -24220 35141 -24210
rect 34971 -24244 34990 -24220
rect 34925 -24250 34990 -24244
rect 34930 -24280 34990 -24250
rect 35130 -24250 35141 -24220
rect 35130 -24280 35140 -24250
rect 34930 -24290 35140 -24280
rect 35180 -24342 35210 -24163
rect 35250 -24204 35280 -23722
rect 35330 -23763 35360 -23630
rect 35399 -23682 35457 -23676
rect 35399 -23716 35411 -23682
rect 35445 -23716 35457 -23682
rect 35399 -23722 35457 -23716
rect 35557 -23682 35615 -23676
rect 35557 -23716 35569 -23682
rect 35603 -23716 35615 -23682
rect 35557 -23722 35615 -23716
rect 35326 -23775 35372 -23763
rect 35326 -24151 35332 -23775
rect 35366 -24151 35372 -23775
rect 35326 -24163 35372 -24151
rect 35410 -24204 35440 -23722
rect 35484 -23775 35530 -23763
rect 35484 -24151 35490 -23775
rect 35524 -24151 35530 -23775
rect 35484 -24163 35530 -24151
rect 35241 -24210 35299 -24204
rect 35399 -24210 35457 -24204
rect 35241 -24244 35253 -24210
rect 35287 -24220 35411 -24210
rect 35445 -24220 35460 -24210
rect 35241 -24250 35260 -24244
rect 35250 -24280 35260 -24250
rect 35450 -24280 35460 -24220
rect 35250 -24290 35460 -24280
rect 35490 -24342 35520 -24163
rect 35570 -24204 35600 -23722
rect 35650 -23763 35680 -23630
rect 35715 -23682 35773 -23676
rect 35715 -23716 35727 -23682
rect 35761 -23716 35773 -23682
rect 35715 -23722 35773 -23716
rect 35873 -23682 35931 -23676
rect 35873 -23716 35885 -23682
rect 35919 -23716 35931 -23682
rect 35873 -23722 35931 -23716
rect 35642 -23775 35688 -23763
rect 35642 -24151 35648 -23775
rect 35682 -24151 35688 -23775
rect 35642 -24163 35688 -24151
rect 35730 -24204 35760 -23722
rect 35800 -23775 35846 -23763
rect 35800 -24151 35806 -23775
rect 35840 -24151 35846 -23775
rect 35800 -24163 35846 -24151
rect 35557 -24210 35615 -24204
rect 35715 -24210 35773 -24204
rect 35557 -24244 35569 -24210
rect 35603 -24220 35727 -24210
rect 35761 -24244 35773 -24210
rect 35557 -24250 35570 -24244
rect 35560 -24280 35570 -24250
rect 35760 -24250 35773 -24244
rect 35760 -24280 35770 -24250
rect 35560 -24290 35770 -24280
rect 35810 -24342 35840 -24163
rect 35890 -24204 35920 -23722
rect 35970 -23763 36000 -23630
rect 36031 -23682 36089 -23676
rect 36031 -23716 36043 -23682
rect 36077 -23716 36089 -23682
rect 36031 -23722 36089 -23716
rect 36189 -23682 36247 -23676
rect 36189 -23716 36201 -23682
rect 36235 -23716 36247 -23682
rect 36189 -23722 36247 -23716
rect 35958 -23775 36004 -23763
rect 35958 -24151 35964 -23775
rect 35998 -24151 36004 -23775
rect 35958 -24163 36004 -24151
rect 36050 -24204 36080 -23722
rect 36116 -23775 36162 -23763
rect 36116 -24151 36122 -23775
rect 36156 -24151 36162 -23775
rect 36116 -24163 36162 -24151
rect 35873 -24210 35931 -24204
rect 36031 -24210 36089 -24204
rect 35873 -24244 35885 -24210
rect 35919 -24220 36043 -24210
rect 36077 -24220 36090 -24210
rect 35873 -24250 35890 -24244
rect 35880 -24280 35890 -24250
rect 36080 -24280 36090 -24220
rect 35880 -24290 36090 -24280
rect 36120 -24342 36150 -24163
rect 36200 -24204 36230 -23722
rect 36280 -23763 36310 -23630
rect 36347 -23682 36405 -23676
rect 36347 -23716 36359 -23682
rect 36393 -23716 36405 -23682
rect 36347 -23722 36405 -23716
rect 36505 -23682 36563 -23676
rect 36505 -23716 36517 -23682
rect 36551 -23716 36563 -23682
rect 36505 -23722 36563 -23716
rect 36274 -23775 36320 -23763
rect 36274 -24151 36280 -23775
rect 36314 -24151 36320 -23775
rect 36274 -24163 36320 -24151
rect 36360 -24204 36390 -23722
rect 36432 -23775 36478 -23763
rect 36432 -24151 36438 -23775
rect 36472 -24151 36478 -23775
rect 36432 -24163 36478 -24151
rect 36189 -24210 36247 -24204
rect 36347 -24210 36405 -24204
rect 36189 -24220 36201 -24210
rect 36235 -24220 36359 -24210
rect 36189 -24250 36200 -24220
rect 36393 -24244 36405 -24210
rect 36190 -24280 36200 -24250
rect 36390 -24250 36405 -24244
rect 36390 -24280 36400 -24250
rect 36190 -24290 36400 -24280
rect 36440 -24342 36470 -24163
rect 36520 -24204 36550 -23722
rect 36600 -23763 36630 -23630
rect 36663 -23682 36721 -23676
rect 36663 -23716 36675 -23682
rect 36709 -23716 36721 -23682
rect 36663 -23722 36721 -23716
rect 36821 -23682 36879 -23676
rect 36821 -23716 36833 -23682
rect 36867 -23716 36879 -23682
rect 36821 -23722 36879 -23716
rect 36590 -23775 36636 -23763
rect 36590 -24151 36596 -23775
rect 36630 -24151 36636 -23775
rect 36590 -24163 36636 -24151
rect 36680 -24204 36710 -23722
rect 36748 -23775 36794 -23763
rect 36748 -24151 36754 -23775
rect 36788 -24151 36794 -23775
rect 36748 -24163 36794 -24151
rect 36505 -24210 36563 -24204
rect 36663 -24210 36721 -24204
rect 36505 -24244 36517 -24210
rect 36551 -24220 36675 -24210
rect 36709 -24220 36721 -24210
rect 36505 -24250 36520 -24244
rect 36510 -24280 36520 -24250
rect 36710 -24250 36721 -24220
rect 36710 -24280 36720 -24250
rect 36510 -24290 36720 -24280
rect 36750 -24342 36780 -24163
rect 36830 -24204 36860 -23722
rect 36910 -23763 36940 -23630
rect 37198 -23655 37244 -23643
rect 36979 -23682 37037 -23676
rect 36979 -23716 36991 -23682
rect 37025 -23716 37037 -23682
rect 36979 -23722 37037 -23716
rect 36906 -23775 36952 -23763
rect 36906 -24151 36912 -23775
rect 36946 -24151 36952 -23775
rect 36906 -24163 36952 -24151
rect 36990 -24204 37020 -23722
rect 37064 -23775 37110 -23763
rect 37064 -24151 37070 -23775
rect 37104 -24151 37110 -23775
rect 37064 -24163 37110 -24151
rect 36821 -24210 36879 -24204
rect 36979 -24210 37037 -24204
rect 36820 -24220 36833 -24210
rect 36867 -24220 36991 -24210
rect 36820 -24280 36830 -24220
rect 37025 -24244 37037 -24210
rect 37020 -24250 37037 -24244
rect 37020 -24280 37030 -24250
rect 36820 -24290 37030 -24280
rect 34706 -24348 36940 -24342
rect 34706 -24360 34718 -24348
rect 34134 -24382 34718 -24360
rect 36928 -24360 36940 -24348
rect 37070 -24360 37100 -24163
rect 37198 -24271 37204 -23655
rect 37238 -24271 37244 -23655
rect 37198 -24283 37244 -24271
rect 36928 -24382 37260 -24360
rect 34134 -24384 37260 -24382
rect 27940 -24496 29990 -24390
rect 32540 -24410 37260 -24384
rect 32980 -24420 37260 -24410
rect 27919 -24502 29990 -24496
rect 22458 -24514 26802 -24508
rect 22458 -24548 22470 -24514
rect 26790 -24548 26802 -24514
rect 27919 -24536 27931 -24502
rect 28805 -24520 29990 -24502
rect 28805 -24536 28817 -24520
rect 27919 -24542 28817 -24536
rect 22458 -24554 26802 -24548
rect 28908 -24611 28954 -24599
rect 27870 -24634 28760 -24630
rect 27870 -24640 28764 -24634
rect 27870 -24674 27984 -24640
rect 28752 -24674 28764 -24640
rect 22351 -24683 22913 -24677
rect 22190 -24922 22236 -24910
rect 2500 -25070 4020 -25060
rect 2500 -25100 2510 -25070
rect 2467 -25106 2510 -25100
rect 4010 -25100 4020 -25070
rect 4700 -25070 6220 -25060
rect 4700 -25100 4710 -25070
rect 4010 -25106 4067 -25100
rect 2467 -25140 2479 -25106
rect 4055 -25140 4067 -25106
rect 2467 -25146 4067 -25140
rect 4667 -25106 4710 -25100
rect 6210 -25100 6220 -25070
rect 6900 -25070 8420 -25060
rect 6900 -25100 6910 -25070
rect 6210 -25106 6267 -25100
rect 4667 -25140 4679 -25106
rect 6255 -25140 6267 -25106
rect 4667 -25146 6267 -25140
rect 6867 -25106 6910 -25100
rect 8410 -25100 8420 -25070
rect 9100 -25070 10620 -25060
rect 9100 -25100 9110 -25070
rect 8410 -25106 8467 -25100
rect 6867 -25140 6879 -25106
rect 8455 -25140 8467 -25106
rect 6867 -25146 8467 -25140
rect 9067 -25106 9110 -25100
rect 10610 -25100 10620 -25070
rect 11300 -25070 12820 -25060
rect 11300 -25100 11310 -25070
rect 10610 -25106 10667 -25100
rect 9067 -25140 9079 -25106
rect 10655 -25140 10667 -25106
rect 9067 -25146 10667 -25140
rect 11267 -25106 11310 -25100
rect 12810 -25100 12820 -25070
rect 13500 -25070 15020 -25060
rect 13500 -25100 13510 -25070
rect 12810 -25106 12867 -25100
rect 11267 -25140 11279 -25106
rect 12855 -25140 12867 -25106
rect 11267 -25146 12867 -25140
rect 13467 -25106 13510 -25100
rect 15010 -25100 15020 -25070
rect 15700 -25070 17220 -25060
rect 15700 -25100 15710 -25070
rect 15010 -25106 15067 -25100
rect 13467 -25140 13479 -25106
rect 15055 -25140 15067 -25106
rect 13467 -25146 15067 -25140
rect 15667 -25106 15710 -25100
rect 17210 -25100 17220 -25070
rect 17900 -25070 19420 -25060
rect 17900 -25100 17910 -25070
rect 17210 -25106 17267 -25100
rect 15667 -25140 15679 -25106
rect 17255 -25140 17267 -25106
rect 15667 -25146 17267 -25140
rect 17867 -25106 17910 -25100
rect 19410 -25100 19420 -25070
rect 19410 -25106 19467 -25100
rect 17867 -25140 17879 -25106
rect 19455 -25140 19467 -25106
rect 17867 -25146 19467 -25140
rect 2380 -25168 2426 -25156
rect 2380 -25260 2386 -25168
rect 2010 -25320 2240 -25260
rect 2300 -25320 2386 -25260
rect 2380 -25436 2386 -25320
rect 2420 -25436 2426 -25168
rect 4108 -25168 4154 -25156
rect 4108 -25170 4114 -25168
rect 4100 -25230 4114 -25170
rect 2380 -25448 2426 -25436
rect 4108 -25436 4114 -25230
rect 4148 -25170 4154 -25168
rect 4580 -25168 4626 -25156
rect 4148 -25230 4440 -25170
rect 4500 -25230 4510 -25170
rect 4148 -25436 4154 -25230
rect 4580 -25280 4586 -25168
rect 4210 -25340 4440 -25280
rect 4500 -25340 4586 -25280
rect 4108 -25448 4154 -25436
rect 4580 -25436 4586 -25340
rect 4620 -25436 4626 -25168
rect 6308 -25168 6354 -25156
rect 6308 -25170 6314 -25168
rect 6300 -25230 6314 -25170
rect 4580 -25448 4626 -25436
rect 6308 -25436 6314 -25230
rect 6348 -25170 6354 -25168
rect 6780 -25168 6826 -25156
rect 6348 -25230 6640 -25170
rect 6700 -25230 6710 -25170
rect 6348 -25436 6354 -25230
rect 6780 -25280 6786 -25168
rect 6410 -25340 6420 -25280
rect 6480 -25340 6786 -25280
rect 6308 -25448 6354 -25436
rect 6780 -25436 6786 -25340
rect 6820 -25436 6826 -25168
rect 8508 -25168 8554 -25156
rect 8508 -25170 8514 -25168
rect 8500 -25230 8514 -25170
rect 6780 -25448 6826 -25436
rect 8508 -25436 8514 -25230
rect 8548 -25170 8554 -25168
rect 8980 -25168 9026 -25156
rect 8548 -25230 8620 -25170
rect 8680 -25230 8910 -25170
rect 8548 -25436 8554 -25230
rect 8980 -25280 8986 -25168
rect 8610 -25340 8620 -25280
rect 8680 -25340 8986 -25280
rect 8508 -25448 8554 -25436
rect 8980 -25436 8986 -25340
rect 9020 -25436 9026 -25168
rect 10708 -25168 10754 -25156
rect 10708 -25170 10714 -25168
rect 10700 -25230 10714 -25170
rect 8980 -25448 9026 -25436
rect 10708 -25436 10714 -25230
rect 10748 -25170 10754 -25168
rect 11180 -25168 11226 -25156
rect 10748 -25230 10820 -25170
rect 10880 -25230 11110 -25170
rect 10748 -25436 10754 -25230
rect 11180 -25280 11186 -25168
rect 10810 -25340 10820 -25280
rect 10880 -25340 11186 -25280
rect 10708 -25448 10754 -25436
rect 11180 -25436 11186 -25340
rect 11220 -25436 11226 -25168
rect 12908 -25168 12954 -25156
rect 12908 -25170 12914 -25168
rect 12900 -25230 12914 -25170
rect 11180 -25448 11226 -25436
rect 12908 -25436 12914 -25230
rect 12948 -25170 12954 -25168
rect 13380 -25168 13426 -25156
rect 12948 -25230 13020 -25170
rect 13080 -25230 13310 -25170
rect 12948 -25436 12954 -25230
rect 13380 -25280 13386 -25168
rect 13010 -25340 13020 -25280
rect 13080 -25340 13386 -25280
rect 12908 -25448 12954 -25436
rect 13380 -25436 13386 -25340
rect 13420 -25436 13426 -25168
rect 15108 -25168 15154 -25156
rect 15108 -25170 15114 -25168
rect 15100 -25230 15114 -25170
rect 13380 -25448 13426 -25436
rect 15108 -25436 15114 -25230
rect 15148 -25170 15154 -25168
rect 15580 -25168 15626 -25156
rect 15148 -25230 15220 -25170
rect 15280 -25230 15510 -25170
rect 15148 -25436 15154 -25230
rect 15580 -25280 15586 -25168
rect 15210 -25340 15440 -25280
rect 15500 -25340 15586 -25280
rect 15108 -25448 15154 -25436
rect 15580 -25436 15586 -25340
rect 15620 -25436 15626 -25168
rect 17308 -25168 17354 -25156
rect 17308 -25170 17314 -25168
rect 17300 -25230 17314 -25170
rect 15580 -25448 15626 -25436
rect 17308 -25436 17314 -25230
rect 17348 -25170 17354 -25168
rect 17780 -25168 17826 -25156
rect 17348 -25230 17640 -25170
rect 17700 -25230 17710 -25170
rect 17348 -25436 17354 -25230
rect 17780 -25280 17786 -25168
rect 17410 -25340 17640 -25280
rect 17700 -25340 17786 -25280
rect 17308 -25448 17354 -25436
rect 17780 -25436 17786 -25340
rect 17820 -25436 17826 -25168
rect 19508 -25168 19554 -25156
rect 19508 -25170 19514 -25168
rect 19500 -25230 19514 -25170
rect 17780 -25448 17826 -25436
rect 19508 -25436 19514 -25230
rect 19548 -25170 19554 -25168
rect 19548 -25230 19840 -25170
rect 19900 -25230 19910 -25170
rect 19548 -25436 19554 -25230
rect 19508 -25448 19554 -25436
rect 2467 -25464 4067 -25458
rect 2467 -25498 2479 -25464
rect 4055 -25498 4067 -25464
rect 2467 -25504 4067 -25498
rect 4667 -25464 6267 -25458
rect 4667 -25498 4679 -25464
rect 6255 -25498 6267 -25464
rect 4667 -25504 6267 -25498
rect 6867 -25464 8467 -25458
rect 6867 -25498 6879 -25464
rect 8455 -25498 8467 -25464
rect 6867 -25504 8467 -25498
rect 9067 -25464 10667 -25458
rect 9067 -25498 9079 -25464
rect 10655 -25498 10667 -25464
rect 9067 -25504 10667 -25498
rect 11267 -25464 12867 -25458
rect 11267 -25498 11279 -25464
rect 12855 -25498 12867 -25464
rect 11267 -25504 12867 -25498
rect 13467 -25464 15067 -25458
rect 13467 -25498 13479 -25464
rect 15055 -25498 15067 -25464
rect 13467 -25504 15067 -25498
rect 15667 -25464 17267 -25458
rect 15667 -25498 15679 -25464
rect 17255 -25498 17267 -25464
rect 15667 -25504 17267 -25498
rect 17867 -25464 19467 -25458
rect 17867 -25498 17879 -25464
rect 19455 -25498 19467 -25464
rect 17867 -25504 19467 -25498
rect 2500 -25700 2700 -25504
rect 2500 -25760 2510 -25700
rect 2690 -25760 2700 -25700
rect 3160 -25700 3360 -25504
rect 3160 -25760 3170 -25700
rect 3350 -25760 3360 -25700
rect 3820 -25700 4020 -25504
rect 3820 -25760 3830 -25700
rect 4010 -25760 4020 -25700
rect 4700 -25700 4900 -25504
rect 4700 -25760 4710 -25700
rect 4890 -25760 4900 -25700
rect 5360 -25700 5560 -25504
rect 5360 -25760 5370 -25700
rect 5550 -25760 5560 -25700
rect 6020 -25700 6220 -25504
rect 6020 -25760 6030 -25700
rect 6210 -25760 6220 -25700
rect 6900 -25560 7100 -25504
rect 6900 -25620 6910 -25560
rect 7090 -25620 7100 -25560
rect 6900 -25760 7100 -25620
rect 7560 -25560 7760 -25504
rect 7560 -25620 7570 -25560
rect 7750 -25620 7760 -25560
rect 7560 -25760 7760 -25620
rect 8220 -25560 8420 -25504
rect 8220 -25620 8230 -25560
rect 8410 -25620 8420 -25560
rect 8220 -25760 8420 -25620
rect 9100 -25560 9300 -25504
rect 9100 -25620 9110 -25560
rect 9290 -25620 9300 -25560
rect 9100 -25760 9300 -25620
rect 9760 -25560 9960 -25504
rect 9760 -25620 9770 -25560
rect 9950 -25620 9960 -25560
rect 9760 -25760 9960 -25620
rect 10420 -25560 10620 -25504
rect 10420 -25620 10430 -25560
rect 10610 -25620 10620 -25560
rect 10420 -25760 10620 -25620
rect 11300 -25560 11500 -25504
rect 11300 -25620 11310 -25560
rect 11490 -25620 11500 -25560
rect 11300 -25760 11500 -25620
rect 11960 -25560 12160 -25504
rect 11960 -25620 11970 -25560
rect 12150 -25620 12160 -25560
rect 11960 -25760 12160 -25620
rect 12620 -25560 12820 -25504
rect 12620 -25620 12630 -25560
rect 12810 -25620 12820 -25560
rect 12620 -25760 12820 -25620
rect 13500 -25560 13700 -25504
rect 13500 -25620 13510 -25560
rect 13690 -25620 13700 -25560
rect 13500 -25760 13700 -25620
rect 14160 -25560 14360 -25504
rect 14160 -25620 14170 -25560
rect 14350 -25620 14360 -25560
rect 14160 -25760 14360 -25620
rect 14820 -25560 15020 -25504
rect 14820 -25620 14830 -25560
rect 15010 -25620 15020 -25560
rect 14820 -25760 15020 -25620
rect 15700 -25700 15900 -25504
rect 15700 -25760 15710 -25700
rect 15890 -25760 15900 -25700
rect 16360 -25700 16560 -25504
rect 16360 -25760 16370 -25700
rect 16550 -25760 16560 -25700
rect 17020 -25700 17220 -25504
rect 17020 -25760 17030 -25700
rect 17210 -25760 17220 -25700
rect 17900 -25700 18100 -25504
rect 17900 -25760 17910 -25700
rect 18090 -25760 18100 -25700
rect 18560 -25700 18760 -25504
rect 18560 -25760 18570 -25700
rect 18750 -25760 18760 -25700
rect 19220 -25700 19420 -25504
rect 19220 -25760 19230 -25700
rect 19410 -25760 19420 -25700
rect 2500 -25870 4020 -25860
rect 2500 -25900 2510 -25870
rect 2467 -25906 2510 -25900
rect 4010 -25900 4020 -25870
rect 4700 -25870 6220 -25860
rect 4700 -25900 4710 -25870
rect 4010 -25906 4067 -25900
rect 2467 -25940 2479 -25906
rect 4055 -25940 4067 -25906
rect 2467 -25946 4067 -25940
rect 4667 -25906 4710 -25900
rect 6210 -25900 6220 -25870
rect 6900 -25870 8420 -25860
rect 6900 -25900 6910 -25870
rect 6210 -25906 6267 -25900
rect 4667 -25940 4679 -25906
rect 6255 -25940 6267 -25906
rect 4667 -25946 6267 -25940
rect 6867 -25906 6910 -25900
rect 8410 -25900 8420 -25870
rect 9100 -25870 10620 -25860
rect 9100 -25900 9110 -25870
rect 8410 -25906 8467 -25900
rect 6867 -25940 6879 -25906
rect 8455 -25940 8467 -25906
rect 6867 -25946 8467 -25940
rect 9067 -25906 9110 -25900
rect 10610 -25900 10620 -25870
rect 11300 -25870 12820 -25860
rect 11300 -25900 11310 -25870
rect 10610 -25906 10667 -25900
rect 9067 -25940 9079 -25906
rect 10655 -25940 10667 -25906
rect 9067 -25946 10667 -25940
rect 11267 -25906 11310 -25900
rect 12810 -25900 12820 -25870
rect 13500 -25870 15020 -25860
rect 13500 -25900 13510 -25870
rect 12810 -25906 12867 -25900
rect 11267 -25940 11279 -25906
rect 12855 -25940 12867 -25906
rect 11267 -25946 12867 -25940
rect 13467 -25906 13510 -25900
rect 15010 -25900 15020 -25870
rect 15700 -25870 17220 -25860
rect 15700 -25900 15710 -25870
rect 15010 -25906 15067 -25900
rect 13467 -25940 13479 -25906
rect 15055 -25940 15067 -25906
rect 13467 -25946 15067 -25940
rect 15667 -25906 15710 -25900
rect 17210 -25900 17220 -25870
rect 17900 -25870 19420 -25860
rect 17900 -25900 17910 -25870
rect 17210 -25906 17267 -25900
rect 15667 -25940 15679 -25906
rect 17255 -25940 17267 -25906
rect 15667 -25946 17267 -25940
rect 17867 -25906 17910 -25900
rect 19410 -25900 19420 -25870
rect 19410 -25906 19467 -25900
rect 17867 -25940 17879 -25906
rect 19455 -25940 19467 -25906
rect 17867 -25946 19467 -25940
rect 2380 -25968 2426 -25956
rect 2380 -26060 2386 -25968
rect 2010 -26120 2020 -26060
rect 2080 -26120 2386 -26060
rect 2380 -26236 2386 -26120
rect 2420 -26236 2426 -25968
rect 4108 -25968 4154 -25956
rect 4108 -25970 4114 -25968
rect 4100 -26030 4114 -25970
rect 2380 -26248 2426 -26236
rect 4108 -26236 4114 -26030
rect 4148 -25970 4154 -25968
rect 4580 -25968 4626 -25956
rect 4148 -26030 4220 -25970
rect 4280 -26030 4510 -25970
rect 4148 -26236 4154 -26030
rect 4580 -26080 4586 -25968
rect 4210 -26140 4220 -26080
rect 4280 -26140 4586 -26080
rect 4108 -26248 4154 -26236
rect 4580 -26236 4586 -26140
rect 4620 -26236 4626 -25968
rect 6308 -25968 6354 -25956
rect 6308 -25970 6314 -25968
rect 6300 -26030 6314 -25970
rect 4580 -26248 4626 -26236
rect 6308 -26236 6314 -26030
rect 6348 -25970 6354 -25968
rect 6780 -25968 6826 -25956
rect 6348 -26030 6420 -25970
rect 6480 -26030 6710 -25970
rect 6348 -26236 6354 -26030
rect 6780 -26080 6786 -25968
rect 6410 -26140 6640 -26080
rect 6700 -26140 6786 -26080
rect 6308 -26248 6354 -26236
rect 6780 -26236 6786 -26140
rect 6820 -26236 6826 -25968
rect 8508 -25968 8554 -25956
rect 8508 -25970 8514 -25968
rect 8500 -26030 8514 -25970
rect 6780 -26248 6826 -26236
rect 8508 -26236 8514 -26030
rect 8548 -25970 8554 -25968
rect 8980 -25968 9026 -25956
rect 8548 -26030 8840 -25970
rect 8900 -26030 8910 -25970
rect 8548 -26236 8554 -26030
rect 8980 -26080 8986 -25968
rect 8610 -26140 8840 -26080
rect 8900 -26140 8986 -26080
rect 8508 -26248 8554 -26236
rect 8980 -26236 8986 -26140
rect 9020 -26236 9026 -25968
rect 10708 -25968 10754 -25956
rect 10708 -25970 10714 -25968
rect 10700 -26030 10714 -25970
rect 8980 -26248 9026 -26236
rect 10708 -26236 10714 -26030
rect 10748 -25970 10754 -25968
rect 11180 -25968 11226 -25956
rect 10748 -26030 11040 -25970
rect 11100 -26030 11110 -25970
rect 10748 -26236 10754 -26030
rect 11180 -26080 11186 -25968
rect 10810 -26140 11040 -26080
rect 11100 -26140 11186 -26080
rect 10708 -26248 10754 -26236
rect 11180 -26236 11186 -26140
rect 11220 -26236 11226 -25968
rect 12908 -25968 12954 -25956
rect 12908 -25970 12914 -25968
rect 12900 -26030 12914 -25970
rect 11180 -26248 11226 -26236
rect 12908 -26236 12914 -26030
rect 12948 -25970 12954 -25968
rect 13380 -25968 13426 -25956
rect 12948 -26030 13240 -25970
rect 13300 -26030 13310 -25970
rect 12948 -26236 12954 -26030
rect 13380 -26080 13386 -25968
rect 13010 -26140 13240 -26080
rect 13300 -26140 13386 -26080
rect 12908 -26248 12954 -26236
rect 13380 -26236 13386 -26140
rect 13420 -26236 13426 -25968
rect 15108 -25968 15154 -25956
rect 15108 -25970 15114 -25968
rect 15100 -26030 15114 -25970
rect 13380 -26248 13426 -26236
rect 15108 -26236 15114 -26030
rect 15148 -25970 15154 -25968
rect 15580 -25968 15626 -25956
rect 15148 -26030 15440 -25970
rect 15500 -26030 15510 -25970
rect 15148 -26236 15154 -26030
rect 15580 -26080 15586 -25968
rect 15210 -26140 15220 -26080
rect 15280 -26140 15586 -26080
rect 15108 -26248 15154 -26236
rect 15580 -26236 15586 -26140
rect 15620 -26236 15626 -25968
rect 17308 -25968 17354 -25956
rect 17308 -25970 17314 -25968
rect 17300 -26030 17314 -25970
rect 15580 -26248 15626 -26236
rect 17308 -26236 17314 -26030
rect 17348 -25970 17354 -25968
rect 17780 -25968 17826 -25956
rect 17348 -26030 17420 -25970
rect 17480 -26030 17710 -25970
rect 17348 -26236 17354 -26030
rect 17780 -26080 17786 -25968
rect 17410 -26140 17420 -26080
rect 17480 -26140 17786 -26080
rect 17308 -26248 17354 -26236
rect 17780 -26236 17786 -26140
rect 17820 -26236 17826 -25968
rect 19508 -25968 19554 -25956
rect 19508 -25970 19514 -25968
rect 19500 -26030 19514 -25970
rect 17780 -26248 17826 -26236
rect 19508 -26236 19514 -26030
rect 19548 -25970 19554 -25968
rect 19548 -26030 19620 -25970
rect 19680 -26030 19910 -25970
rect 19548 -26236 19554 -26030
rect 19508 -26248 19554 -26236
rect 2467 -26264 4067 -26258
rect 2467 -26298 2479 -26264
rect 4055 -26298 4067 -26264
rect 2467 -26304 4067 -26298
rect 4667 -26264 6267 -26258
rect 4667 -26298 4679 -26264
rect 6255 -26298 6267 -26264
rect 4667 -26304 6267 -26298
rect 6867 -26264 8467 -26258
rect 6867 -26298 6879 -26264
rect 8455 -26298 8467 -26264
rect 6867 -26304 8467 -26298
rect 9067 -26264 10667 -26258
rect 9067 -26298 9079 -26264
rect 10655 -26298 10667 -26264
rect 9067 -26304 10667 -26298
rect 11267 -26264 12867 -26258
rect 11267 -26298 11279 -26264
rect 12855 -26298 12867 -26264
rect 11267 -26304 12867 -26298
rect 13467 -26264 15067 -26258
rect 13467 -26298 13479 -26264
rect 15055 -26298 15067 -26264
rect 13467 -26304 15067 -26298
rect 15667 -26264 17267 -26258
rect 15667 -26298 15679 -26264
rect 17255 -26298 17267 -26264
rect 15667 -26304 17267 -26298
rect 17867 -26264 19467 -26258
rect 17867 -26298 17879 -26264
rect 19455 -26298 19467 -26264
rect 17867 -26304 19467 -26298
rect 2500 -26360 2700 -26304
rect 2500 -26420 2510 -26360
rect 2690 -26420 2700 -26360
rect 2500 -26560 2700 -26420
rect 3160 -26360 3360 -26304
rect 3160 -26420 3170 -26360
rect 3350 -26420 3360 -26360
rect 3160 -26560 3360 -26420
rect 3820 -26360 4020 -26304
rect 3820 -26420 3830 -26360
rect 4010 -26420 4020 -26360
rect 3820 -26560 4020 -26420
rect 4700 -26360 4900 -26304
rect 4700 -26420 4710 -26360
rect 4890 -26420 4900 -26360
rect 4700 -26560 4900 -26420
rect 5360 -26360 5560 -26304
rect 5360 -26420 5370 -26360
rect 5550 -26420 5560 -26360
rect 5360 -26560 5560 -26420
rect 6020 -26360 6220 -26304
rect 6020 -26420 6030 -26360
rect 6210 -26420 6220 -26360
rect 6020 -26560 6220 -26420
rect 6900 -26500 7100 -26304
rect 6900 -26560 6910 -26500
rect 7090 -26560 7100 -26500
rect 7560 -26500 7760 -26304
rect 7560 -26560 7570 -26500
rect 7750 -26560 7760 -26500
rect 8220 -26500 8420 -26304
rect 8220 -26560 8230 -26500
rect 8410 -26560 8420 -26500
rect 9100 -26500 9300 -26304
rect 9100 -26560 9110 -26500
rect 9290 -26560 9300 -26500
rect 9760 -26500 9960 -26304
rect 9760 -26560 9770 -26500
rect 9950 -26560 9960 -26500
rect 10420 -26500 10620 -26304
rect 10420 -26560 10430 -26500
rect 10610 -26560 10620 -26500
rect 11300 -26500 11500 -26304
rect 11300 -26560 11310 -26500
rect 11490 -26560 11500 -26500
rect 11960 -26500 12160 -26304
rect 11960 -26560 11970 -26500
rect 12150 -26560 12160 -26500
rect 12620 -26500 12820 -26304
rect 12620 -26560 12630 -26500
rect 12810 -26560 12820 -26500
rect 13500 -26500 13700 -26304
rect 13500 -26560 13510 -26500
rect 13690 -26560 13700 -26500
rect 14160 -26500 14360 -26304
rect 14160 -26560 14170 -26500
rect 14350 -26560 14360 -26500
rect 14820 -26500 15020 -26304
rect 14820 -26560 14830 -26500
rect 15010 -26560 15020 -26500
rect 15700 -26360 15900 -26304
rect 15700 -26420 15710 -26360
rect 15890 -26420 15900 -26360
rect 15700 -26560 15900 -26420
rect 16360 -26360 16560 -26304
rect 16360 -26420 16370 -26360
rect 16550 -26420 16560 -26360
rect 16360 -26560 16560 -26420
rect 17020 -26360 17220 -26304
rect 17020 -26420 17030 -26360
rect 17210 -26420 17220 -26360
rect 17020 -26560 17220 -26420
rect 17900 -26360 18100 -26304
rect 17900 -26420 17910 -26360
rect 18090 -26420 18100 -26360
rect 17900 -26560 18100 -26420
rect 18560 -26360 18760 -26304
rect 18560 -26420 18570 -26360
rect 18750 -26420 18760 -26360
rect 18560 -26560 18760 -26420
rect 19220 -26360 19420 -26304
rect 19220 -26420 19230 -26360
rect 19410 -26420 19420 -26360
rect 19220 -26560 19420 -26420
rect 420 -26630 620 -26620
rect 420 -26710 430 -26630
rect 610 -26640 620 -26630
rect 21300 -26630 21500 -26620
rect 21300 -26640 21310 -26630
rect 610 -26700 4040 -26640
rect 4700 -26670 6220 -26660
rect 4700 -26700 4710 -26670
rect 610 -26710 620 -26700
rect 420 -26720 620 -26710
rect 2467 -26706 4067 -26700
rect 2467 -26740 2479 -26706
rect 4055 -26740 4067 -26706
rect 2467 -26746 4067 -26740
rect 4667 -26706 4710 -26700
rect 6210 -26700 6220 -26670
rect 6900 -26670 8420 -26660
rect 6900 -26700 6910 -26670
rect 6210 -26706 6267 -26700
rect 4667 -26740 4679 -26706
rect 6255 -26740 6267 -26706
rect 4667 -26746 6267 -26740
rect 6867 -26706 6910 -26700
rect 8410 -26700 8420 -26670
rect 9100 -26670 10620 -26660
rect 9100 -26700 9110 -26670
rect 8410 -26706 8467 -26700
rect 6867 -26740 6879 -26706
rect 8455 -26740 8467 -26706
rect 6867 -26746 8467 -26740
rect 9067 -26706 9110 -26700
rect 10610 -26700 10620 -26670
rect 11300 -26670 12820 -26660
rect 11300 -26700 11310 -26670
rect 10610 -26706 10667 -26700
rect 9067 -26740 9079 -26706
rect 10655 -26740 10667 -26706
rect 9067 -26746 10667 -26740
rect 11267 -26706 11310 -26700
rect 12810 -26700 12820 -26670
rect 13500 -26670 15020 -26660
rect 13500 -26700 13510 -26670
rect 12810 -26706 12867 -26700
rect 11267 -26740 11279 -26706
rect 12855 -26740 12867 -26706
rect 11267 -26746 12867 -26740
rect 13467 -26706 13510 -26700
rect 15010 -26700 15020 -26670
rect 15700 -26670 17220 -26660
rect 15700 -26700 15710 -26670
rect 15010 -26706 15067 -26700
rect 13467 -26740 13479 -26706
rect 15055 -26740 15067 -26706
rect 13467 -26746 15067 -26740
rect 15667 -26706 15710 -26700
rect 17210 -26700 17220 -26670
rect 17880 -26700 21310 -26640
rect 17210 -26706 17267 -26700
rect 15667 -26740 15679 -26706
rect 17255 -26740 17267 -26706
rect 15667 -26746 17267 -26740
rect 17867 -26706 19467 -26700
rect 17867 -26740 17879 -26706
rect 19455 -26740 19467 -26706
rect 21300 -26710 21310 -26700
rect 21490 -26710 21500 -26630
rect 21300 -26720 21500 -26710
rect 17867 -26746 19467 -26740
rect 2380 -26768 2426 -26756
rect 2380 -26860 2386 -26768
rect 1410 -26870 2386 -26860
rect 1410 -27020 1420 -26870
rect 1480 -26920 2386 -26870
rect 1480 -27020 1490 -26920
rect 1410 -27030 1490 -27020
rect 2380 -27036 2386 -26920
rect 2420 -27036 2426 -26768
rect 4108 -26768 4154 -26756
rect 4108 -26770 4114 -26768
rect 4100 -26830 4114 -26770
rect 2380 -27048 2426 -27036
rect 4108 -27036 4114 -26830
rect 4148 -26770 4154 -26768
rect 4580 -26768 4626 -26756
rect 4148 -26830 4510 -26770
rect 4148 -27036 4154 -26830
rect 4580 -26880 4586 -26768
rect 4210 -26940 4440 -26880
rect 4500 -26940 4586 -26880
rect 4108 -27048 4154 -27036
rect 4580 -27036 4586 -26940
rect 4620 -27036 4626 -26768
rect 6308 -26768 6354 -26756
rect 6308 -26770 6314 -26768
rect 6300 -26830 6314 -26770
rect 4580 -27048 4626 -27036
rect 6308 -27036 6314 -26830
rect 6348 -26770 6354 -26768
rect 6780 -26768 6826 -26756
rect 6348 -26830 6640 -26770
rect 6700 -26830 6710 -26770
rect 6348 -27036 6354 -26830
rect 6780 -26880 6786 -26768
rect 6410 -26940 6420 -26880
rect 6480 -26940 6786 -26880
rect 6308 -27048 6354 -27036
rect 6780 -27036 6786 -26940
rect 6820 -27036 6826 -26768
rect 8508 -26768 8554 -26756
rect 8508 -26770 8514 -26768
rect 8500 -26830 8514 -26770
rect 6780 -27048 6826 -27036
rect 8508 -27036 8514 -26830
rect 8548 -26770 8554 -26768
rect 8980 -26768 9026 -26756
rect 8548 -26830 8620 -26770
rect 8680 -26830 8910 -26770
rect 8548 -27036 8554 -26830
rect 8980 -26880 8986 -26768
rect 8610 -26940 8620 -26880
rect 8680 -26940 8986 -26880
rect 8508 -27048 8554 -27036
rect 8980 -27036 8986 -26940
rect 9020 -27036 9026 -26768
rect 10708 -26768 10754 -26756
rect 10708 -26770 10714 -26768
rect 10700 -26830 10714 -26770
rect 8980 -27048 9026 -27036
rect 10708 -27036 10714 -26830
rect 10748 -26770 10754 -26768
rect 11180 -26768 11226 -26756
rect 10748 -26830 10820 -26770
rect 10880 -26830 11110 -26770
rect 10748 -27036 10754 -26830
rect 11180 -26880 11186 -26768
rect 10810 -26940 10820 -26880
rect 10880 -26940 11186 -26880
rect 10708 -27048 10754 -27036
rect 11180 -27036 11186 -26940
rect 11220 -27036 11226 -26768
rect 12908 -26768 12954 -26756
rect 12908 -26770 12914 -26768
rect 12900 -26830 12914 -26770
rect 11180 -27048 11226 -27036
rect 12908 -27036 12914 -26830
rect 12948 -26770 12954 -26768
rect 13380 -26768 13426 -26756
rect 12948 -26830 13020 -26770
rect 13080 -26830 13310 -26770
rect 12948 -27036 12954 -26830
rect 13380 -26880 13386 -26768
rect 13010 -26940 13020 -26880
rect 13080 -26940 13386 -26880
rect 12908 -27048 12954 -27036
rect 13380 -27036 13386 -26940
rect 13420 -27036 13426 -26768
rect 15108 -26768 15154 -26756
rect 15108 -26770 15114 -26768
rect 15100 -26830 15114 -26770
rect 13380 -27048 13426 -27036
rect 15108 -27036 15114 -26830
rect 15148 -26770 15154 -26768
rect 15580 -26768 15626 -26756
rect 15148 -26830 15220 -26770
rect 15280 -26830 15510 -26770
rect 15148 -27036 15154 -26830
rect 15580 -26880 15586 -26768
rect 15210 -26940 15440 -26880
rect 15500 -26940 15586 -26880
rect 15108 -27048 15154 -27036
rect 15580 -27036 15586 -26940
rect 15620 -27036 15626 -26768
rect 17308 -26768 17354 -26756
rect 17308 -26770 17314 -26768
rect 17300 -26830 17314 -26770
rect 15580 -27048 15626 -27036
rect 17308 -27036 17314 -26830
rect 17348 -26770 17354 -26768
rect 17780 -26768 17826 -26756
rect 17348 -26830 17640 -26770
rect 17700 -26830 17710 -26770
rect 17348 -27036 17354 -26830
rect 17780 -26880 17786 -26768
rect 17410 -26940 17786 -26880
rect 17308 -27048 17354 -27036
rect 17780 -27036 17786 -26940
rect 17820 -27036 17826 -26768
rect 19508 -26768 19554 -26756
rect 19508 -26770 19514 -26768
rect 19500 -26830 19514 -26770
rect 17780 -27048 17826 -27036
rect 19508 -27036 19514 -26830
rect 19548 -26770 19554 -26768
rect 19548 -26780 20310 -26770
rect 19548 -26830 20240 -26780
rect 19548 -27036 19554 -26830
rect 20230 -26930 20240 -26830
rect 20300 -26930 20310 -26780
rect 20230 -26940 20310 -26930
rect 19508 -27048 19554 -27036
rect 2467 -27064 4067 -27058
rect 2467 -27098 2479 -27064
rect 4055 -27098 4067 -27064
rect 2467 -27104 4067 -27098
rect 4667 -27064 6267 -27058
rect 4667 -27098 4679 -27064
rect 6255 -27098 6267 -27064
rect 4667 -27104 6267 -27098
rect 6867 -27064 8467 -27058
rect 6867 -27098 6879 -27064
rect 8455 -27098 8467 -27064
rect 6867 -27104 8467 -27098
rect 9067 -27064 10667 -27058
rect 9067 -27098 9079 -27064
rect 10655 -27098 10667 -27064
rect 9067 -27104 10667 -27098
rect 11267 -27064 12867 -27058
rect 11267 -27098 11279 -27064
rect 12855 -27098 12867 -27064
rect 11267 -27104 12867 -27098
rect 13467 -27064 15067 -27058
rect 13467 -27098 13479 -27064
rect 15055 -27098 15067 -27064
rect 13467 -27104 15067 -27098
rect 15667 -27064 17267 -27058
rect 15667 -27098 15679 -27064
rect 17255 -27098 17267 -27064
rect 15667 -27104 17267 -27098
rect 17867 -27064 19467 -27058
rect 17867 -27098 17879 -27064
rect 19455 -27098 19467 -27064
rect 17867 -27104 19467 -27098
rect 2500 -27300 2700 -27104
rect 2500 -27360 2510 -27300
rect 2690 -27360 2700 -27300
rect 3160 -27300 3360 -27104
rect 3160 -27360 3170 -27300
rect 3350 -27360 3360 -27300
rect 3820 -27300 4020 -27104
rect 3820 -27360 3830 -27300
rect 4010 -27360 4020 -27300
rect 4700 -27300 4900 -27104
rect 4700 -27360 4710 -27300
rect 4890 -27360 4900 -27300
rect 5360 -27300 5560 -27104
rect 5360 -27360 5370 -27300
rect 5550 -27360 5560 -27300
rect 6020 -27300 6220 -27104
rect 6020 -27360 6030 -27300
rect 6210 -27360 6220 -27300
rect 6900 -27160 7100 -27104
rect 6900 -27220 6910 -27160
rect 7090 -27220 7100 -27160
rect 6900 -27360 7100 -27220
rect 7560 -27160 7760 -27104
rect 7560 -27220 7570 -27160
rect 7750 -27220 7760 -27160
rect 7560 -27360 7760 -27220
rect 8220 -27160 8420 -27104
rect 8220 -27220 8230 -27160
rect 8410 -27220 8420 -27160
rect 8220 -27360 8420 -27220
rect 9100 -27160 9300 -27104
rect 9100 -27220 9110 -27160
rect 9290 -27220 9300 -27160
rect 9100 -27360 9300 -27220
rect 9760 -27160 9960 -27104
rect 9760 -27220 9770 -27160
rect 9950 -27220 9960 -27160
rect 9760 -27360 9960 -27220
rect 10420 -27160 10620 -27104
rect 10420 -27220 10430 -27160
rect 10610 -27220 10620 -27160
rect 10420 -27360 10620 -27220
rect 11300 -27160 11500 -27104
rect 11300 -27220 11310 -27160
rect 11490 -27220 11500 -27160
rect 11300 -27360 11500 -27220
rect 11960 -27160 12160 -27104
rect 11960 -27220 11970 -27160
rect 12150 -27220 12160 -27160
rect 11960 -27360 12160 -27220
rect 12620 -27160 12820 -27104
rect 12620 -27220 12630 -27160
rect 12810 -27220 12820 -27160
rect 12620 -27360 12820 -27220
rect 13500 -27160 13700 -27104
rect 13500 -27220 13510 -27160
rect 13690 -27220 13700 -27160
rect 13500 -27360 13700 -27220
rect 14160 -27160 14360 -27104
rect 14160 -27220 14170 -27160
rect 14350 -27220 14360 -27160
rect 14160 -27360 14360 -27220
rect 14820 -27160 15020 -27104
rect 14820 -27220 14830 -27160
rect 15010 -27220 15020 -27160
rect 14820 -27360 15020 -27220
rect 15700 -27300 15900 -27104
rect 15700 -27360 15710 -27300
rect 15890 -27360 15900 -27300
rect 16360 -27300 16560 -27104
rect 16360 -27360 16370 -27300
rect 16550 -27360 16560 -27300
rect 17020 -27300 17220 -27104
rect 17020 -27360 17030 -27300
rect 17210 -27360 17220 -27300
rect 17900 -27300 18100 -27104
rect 17900 -27360 17910 -27300
rect 18090 -27360 18100 -27300
rect 18560 -27300 18760 -27104
rect 18560 -27360 18570 -27300
rect 18750 -27360 18760 -27300
rect 19220 -27300 19420 -27104
rect 19220 -27360 19230 -27300
rect 19410 -27360 19420 -27300
rect 420 -27430 620 -27420
rect 420 -27510 430 -27430
rect 610 -27440 620 -27430
rect 21300 -27430 21500 -27420
rect 21300 -27440 21310 -27430
rect 610 -27500 4040 -27440
rect 4700 -27470 6220 -27460
rect 4700 -27500 4710 -27470
rect 610 -27510 620 -27500
rect 420 -27520 620 -27510
rect 2467 -27506 4067 -27500
rect 2467 -27540 2479 -27506
rect 4055 -27540 4067 -27506
rect 2467 -27546 4067 -27540
rect 4667 -27506 4710 -27500
rect 6210 -27500 6220 -27470
rect 6900 -27470 8420 -27460
rect 6900 -27500 6910 -27470
rect 6210 -27506 6267 -27500
rect 4667 -27540 4679 -27506
rect 6255 -27540 6267 -27506
rect 4667 -27546 6267 -27540
rect 6867 -27506 6910 -27500
rect 8410 -27500 8420 -27470
rect 9100 -27470 10620 -27460
rect 9100 -27500 9110 -27470
rect 8410 -27506 8467 -27500
rect 6867 -27540 6879 -27506
rect 8455 -27540 8467 -27506
rect 6867 -27546 8467 -27540
rect 9067 -27506 9110 -27500
rect 10610 -27500 10620 -27470
rect 11300 -27470 12820 -27460
rect 11300 -27500 11310 -27470
rect 10610 -27506 10667 -27500
rect 9067 -27540 9079 -27506
rect 10655 -27540 10667 -27506
rect 9067 -27546 10667 -27540
rect 11267 -27506 11310 -27500
rect 12810 -27500 12820 -27470
rect 13500 -27470 15020 -27460
rect 13500 -27500 13510 -27470
rect 12810 -27506 12867 -27500
rect 11267 -27540 11279 -27506
rect 12855 -27540 12867 -27506
rect 11267 -27546 12867 -27540
rect 13467 -27506 13510 -27500
rect 15010 -27500 15020 -27470
rect 15700 -27470 17220 -27460
rect 15700 -27500 15710 -27470
rect 15010 -27506 15067 -27500
rect 13467 -27540 13479 -27506
rect 15055 -27540 15067 -27506
rect 13467 -27546 15067 -27540
rect 15667 -27506 15710 -27500
rect 17210 -27500 17220 -27470
rect 17880 -27500 21310 -27440
rect 17210 -27506 17267 -27500
rect 15667 -27540 15679 -27506
rect 17255 -27540 17267 -27506
rect 15667 -27546 17267 -27540
rect 17867 -27506 19467 -27500
rect 17867 -27540 17879 -27506
rect 19455 -27540 19467 -27506
rect 21300 -27510 21310 -27500
rect 21490 -27510 21500 -27430
rect 21300 -27520 21500 -27510
rect 17867 -27546 19467 -27540
rect 2380 -27568 2426 -27556
rect 2380 -27660 2386 -27568
rect 1610 -27670 2386 -27660
rect 1610 -27820 1620 -27670
rect 1680 -27720 2386 -27670
rect 1680 -27820 1690 -27720
rect 1610 -27830 1690 -27820
rect 2380 -27836 2386 -27720
rect 2420 -27836 2426 -27568
rect 4108 -27568 4154 -27556
rect 4108 -27570 4114 -27568
rect 4100 -27630 4114 -27570
rect 2380 -27848 2426 -27836
rect 4108 -27836 4114 -27630
rect 4148 -27570 4154 -27568
rect 4580 -27568 4626 -27556
rect 4148 -27630 4510 -27570
rect 4148 -27836 4154 -27630
rect 4580 -27680 4586 -27568
rect 4210 -27740 4220 -27680
rect 4280 -27740 4586 -27680
rect 4108 -27848 4154 -27836
rect 4580 -27836 4586 -27740
rect 4620 -27836 4626 -27568
rect 6308 -27568 6354 -27556
rect 6308 -27570 6314 -27568
rect 6300 -27630 6314 -27570
rect 4580 -27848 4626 -27836
rect 6308 -27836 6314 -27630
rect 6348 -27570 6354 -27568
rect 6780 -27568 6826 -27556
rect 6348 -27630 6420 -27570
rect 6480 -27630 6710 -27570
rect 6348 -27836 6354 -27630
rect 6780 -27680 6786 -27568
rect 6410 -27740 6640 -27680
rect 6700 -27740 6786 -27680
rect 6308 -27848 6354 -27836
rect 6780 -27836 6786 -27740
rect 6820 -27836 6826 -27568
rect 8508 -27568 8554 -27556
rect 8508 -27570 8514 -27568
rect 8500 -27630 8514 -27570
rect 6780 -27848 6826 -27836
rect 8508 -27836 8514 -27630
rect 8548 -27570 8554 -27568
rect 8980 -27568 9026 -27556
rect 8548 -27630 8840 -27570
rect 8900 -27630 8910 -27570
rect 8548 -27836 8554 -27630
rect 8980 -27680 8986 -27568
rect 8610 -27740 8840 -27680
rect 8900 -27740 8986 -27680
rect 8508 -27848 8554 -27836
rect 8980 -27836 8986 -27740
rect 9020 -27836 9026 -27568
rect 10708 -27568 10754 -27556
rect 10708 -27570 10714 -27568
rect 10700 -27630 10714 -27570
rect 8980 -27848 9026 -27836
rect 10708 -27836 10714 -27630
rect 10748 -27570 10754 -27568
rect 11180 -27568 11226 -27556
rect 10748 -27630 11040 -27570
rect 11100 -27630 11110 -27570
rect 10748 -27836 10754 -27630
rect 11180 -27680 11186 -27568
rect 10810 -27740 11040 -27680
rect 11100 -27740 11186 -27680
rect 10708 -27848 10754 -27836
rect 11180 -27836 11186 -27740
rect 11220 -27836 11226 -27568
rect 12908 -27568 12954 -27556
rect 12908 -27570 12914 -27568
rect 12900 -27630 12914 -27570
rect 11180 -27848 11226 -27836
rect 12908 -27836 12914 -27630
rect 12948 -27570 12954 -27568
rect 13380 -27568 13426 -27556
rect 12948 -27630 13240 -27570
rect 13300 -27630 13310 -27570
rect 12948 -27836 12954 -27630
rect 13380 -27680 13386 -27568
rect 13010 -27740 13240 -27680
rect 13300 -27740 13386 -27680
rect 12908 -27848 12954 -27836
rect 13380 -27836 13386 -27740
rect 13420 -27836 13426 -27568
rect 15108 -27568 15154 -27556
rect 15108 -27570 15114 -27568
rect 15100 -27630 15114 -27570
rect 13380 -27848 13426 -27836
rect 15108 -27836 15114 -27630
rect 15148 -27570 15154 -27568
rect 15580 -27568 15626 -27556
rect 15148 -27630 15440 -27570
rect 15500 -27630 15510 -27570
rect 15148 -27836 15154 -27630
rect 15580 -27680 15586 -27568
rect 15210 -27740 15220 -27680
rect 15280 -27740 15586 -27680
rect 15108 -27848 15154 -27836
rect 15580 -27836 15586 -27740
rect 15620 -27836 15626 -27568
rect 17308 -27568 17354 -27556
rect 17308 -27570 17314 -27568
rect 17300 -27630 17314 -27570
rect 15580 -27848 15626 -27836
rect 17308 -27836 17314 -27630
rect 17348 -27570 17354 -27568
rect 17780 -27568 17826 -27556
rect 17348 -27630 17420 -27570
rect 17480 -27630 17710 -27570
rect 17348 -27836 17354 -27630
rect 17780 -27680 17786 -27568
rect 17410 -27740 17786 -27680
rect 17308 -27848 17354 -27836
rect 17780 -27836 17786 -27740
rect 17820 -27836 17826 -27568
rect 19508 -27568 19554 -27556
rect 19508 -27570 19514 -27568
rect 19500 -27630 19514 -27570
rect 17780 -27848 17826 -27836
rect 19508 -27836 19514 -27630
rect 19548 -27570 19554 -27568
rect 19548 -27580 20510 -27570
rect 19548 -27630 20440 -27580
rect 19548 -27836 19554 -27630
rect 20430 -27730 20440 -27630
rect 20500 -27730 20510 -27580
rect 20430 -27740 20510 -27730
rect 19508 -27848 19554 -27836
rect 2467 -27864 4067 -27858
rect 2467 -27898 2479 -27864
rect 4055 -27898 4067 -27864
rect 2467 -27904 4067 -27898
rect 4667 -27864 6267 -27858
rect 4667 -27898 4679 -27864
rect 6255 -27898 6267 -27864
rect 4667 -27904 6267 -27898
rect 6867 -27864 8467 -27858
rect 6867 -27898 6879 -27864
rect 8455 -27898 8467 -27864
rect 6867 -27904 8467 -27898
rect 9067 -27864 10667 -27858
rect 9067 -27898 9079 -27864
rect 10655 -27898 10667 -27864
rect 9067 -27904 10667 -27898
rect 11267 -27864 12867 -27858
rect 11267 -27898 11279 -27864
rect 12855 -27898 12867 -27864
rect 11267 -27904 12867 -27898
rect 13467 -27864 15067 -27858
rect 13467 -27898 13479 -27864
rect 15055 -27898 15067 -27864
rect 13467 -27904 15067 -27898
rect 15667 -27864 17267 -27858
rect 15667 -27898 15679 -27864
rect 17255 -27898 17267 -27864
rect 15667 -27904 17267 -27898
rect 17867 -27864 19467 -27858
rect 17867 -27898 17879 -27864
rect 19455 -27898 19467 -27864
rect 17867 -27904 19467 -27898
rect 2500 -27960 2700 -27904
rect 2500 -28020 2510 -27960
rect 2690 -28020 2700 -27960
rect 2500 -28160 2700 -28020
rect 3160 -27960 3360 -27904
rect 3160 -28020 3170 -27960
rect 3350 -28020 3360 -27960
rect 3160 -28160 3360 -28020
rect 3820 -27960 4020 -27904
rect 3820 -28020 3830 -27960
rect 4010 -28020 4020 -27960
rect 3820 -28160 4020 -28020
rect 4700 -27960 4900 -27904
rect 4700 -28020 4710 -27960
rect 4890 -28020 4900 -27960
rect 4700 -28160 4900 -28020
rect 5360 -27960 5560 -27904
rect 5360 -28020 5370 -27960
rect 5550 -28020 5560 -27960
rect 5360 -28160 5560 -28020
rect 6020 -27960 6220 -27904
rect 6020 -28020 6030 -27960
rect 6210 -28020 6220 -27960
rect 6020 -28160 6220 -28020
rect 6900 -28100 7100 -27904
rect 6900 -28160 6910 -28100
rect 7090 -28160 7100 -28100
rect 7560 -28100 7760 -27904
rect 7560 -28160 7570 -28100
rect 7750 -28160 7760 -28100
rect 8220 -28100 8420 -27904
rect 8220 -28160 8230 -28100
rect 8410 -28160 8420 -28100
rect 9100 -28100 9300 -27904
rect 9100 -28160 9110 -28100
rect 9290 -28160 9300 -28100
rect 9760 -28100 9960 -27904
rect 9760 -28160 9770 -28100
rect 9950 -28160 9960 -28100
rect 10420 -28100 10620 -27904
rect 10420 -28160 10430 -28100
rect 10610 -28160 10620 -28100
rect 11300 -28100 11500 -27904
rect 11300 -28160 11310 -28100
rect 11490 -28160 11500 -28100
rect 11960 -28100 12160 -27904
rect 11960 -28160 11970 -28100
rect 12150 -28160 12160 -28100
rect 12620 -28100 12820 -27904
rect 12620 -28160 12630 -28100
rect 12810 -28160 12820 -28100
rect 13500 -28100 13700 -27904
rect 13500 -28160 13510 -28100
rect 13690 -28160 13700 -28100
rect 14160 -28100 14360 -27904
rect 14160 -28160 14170 -28100
rect 14350 -28160 14360 -28100
rect 14820 -28100 15020 -27904
rect 14820 -28160 14830 -28100
rect 15010 -28160 15020 -28100
rect 15700 -27960 15900 -27904
rect 15700 -28020 15710 -27960
rect 15890 -28020 15900 -27960
rect 15700 -28160 15900 -28020
rect 16360 -27960 16560 -27904
rect 16360 -28020 16370 -27960
rect 16550 -28020 16560 -27960
rect 16360 -28160 16560 -28020
rect 17020 -27960 17220 -27904
rect 17020 -28020 17030 -27960
rect 17210 -28020 17220 -27960
rect 17020 -28160 17220 -28020
rect 17900 -27960 18100 -27904
rect 17900 -28020 17910 -27960
rect 18090 -28020 18100 -27960
rect 17900 -28160 18100 -28020
rect 18560 -27960 18760 -27904
rect 18560 -28020 18570 -27960
rect 18750 -28020 18760 -27960
rect 18560 -28160 18760 -28020
rect 19220 -27960 19420 -27904
rect 19220 -28020 19230 -27960
rect 19410 -28020 19420 -27960
rect 19220 -28160 19420 -28020
rect 420 -28230 620 -28220
rect 420 -28310 430 -28230
rect 610 -28240 620 -28230
rect 21300 -28230 21500 -28220
rect 21300 -28240 21310 -28230
rect 610 -28300 4040 -28240
rect 4700 -28270 6220 -28260
rect 4700 -28300 4710 -28270
rect 610 -28310 620 -28300
rect 420 -28320 620 -28310
rect 2467 -28306 4067 -28300
rect 2467 -28340 2479 -28306
rect 4055 -28340 4067 -28306
rect 2467 -28346 4067 -28340
rect 4667 -28306 4710 -28300
rect 6210 -28300 6220 -28270
rect 6900 -28270 8420 -28260
rect 6900 -28300 6910 -28270
rect 6210 -28306 6267 -28300
rect 4667 -28340 4679 -28306
rect 6255 -28340 6267 -28306
rect 4667 -28346 6267 -28340
rect 6867 -28306 6910 -28300
rect 8410 -28300 8420 -28270
rect 9100 -28270 10620 -28260
rect 9100 -28300 9110 -28270
rect 8410 -28306 8467 -28300
rect 6867 -28340 6879 -28306
rect 8455 -28340 8467 -28306
rect 6867 -28346 8467 -28340
rect 9067 -28306 9110 -28300
rect 10610 -28300 10620 -28270
rect 11300 -28270 12820 -28260
rect 11300 -28300 11310 -28270
rect 10610 -28306 10667 -28300
rect 9067 -28340 9079 -28306
rect 10655 -28340 10667 -28306
rect 9067 -28346 10667 -28340
rect 11267 -28306 11310 -28300
rect 12810 -28300 12820 -28270
rect 13500 -28270 15020 -28260
rect 13500 -28300 13510 -28270
rect 12810 -28306 12867 -28300
rect 11267 -28340 11279 -28306
rect 12855 -28340 12867 -28306
rect 11267 -28346 12867 -28340
rect 13467 -28306 13510 -28300
rect 15010 -28300 15020 -28270
rect 15700 -28270 17220 -28260
rect 15700 -28300 15710 -28270
rect 15010 -28306 15067 -28300
rect 13467 -28340 13479 -28306
rect 15055 -28340 15067 -28306
rect 13467 -28346 15067 -28340
rect 15667 -28306 15710 -28300
rect 17210 -28300 17220 -28270
rect 17880 -28300 21310 -28240
rect 17210 -28306 17267 -28300
rect 15667 -28340 15679 -28306
rect 17255 -28340 17267 -28306
rect 15667 -28346 17267 -28340
rect 17867 -28306 19467 -28300
rect 17867 -28340 17879 -28306
rect 19455 -28340 19467 -28306
rect 21300 -28310 21310 -28300
rect 21490 -28310 21500 -28230
rect 21300 -28320 21500 -28310
rect 17867 -28346 19467 -28340
rect 2380 -28368 2426 -28356
rect 2380 -28460 2386 -28368
rect 1610 -28470 2386 -28460
rect 1610 -28620 1620 -28470
rect 1680 -28520 2386 -28470
rect 1680 -28620 1690 -28520
rect 1610 -28630 1690 -28620
rect 2380 -28636 2386 -28520
rect 2420 -28636 2426 -28368
rect 4108 -28368 4154 -28356
rect 4108 -28370 4114 -28368
rect 4100 -28430 4114 -28370
rect 2380 -28648 2426 -28636
rect 4108 -28636 4114 -28430
rect 4148 -28370 4154 -28368
rect 4580 -28368 4626 -28356
rect 4148 -28430 4510 -28370
rect 4148 -28636 4154 -28430
rect 4580 -28480 4586 -28368
rect 4210 -28540 4220 -28480
rect 4280 -28540 4586 -28480
rect 4108 -28648 4154 -28636
rect 4580 -28636 4586 -28540
rect 4620 -28636 4626 -28368
rect 6308 -28368 6354 -28356
rect 6308 -28370 6314 -28368
rect 6300 -28430 6314 -28370
rect 4580 -28648 4626 -28636
rect 6308 -28636 6314 -28430
rect 6348 -28370 6354 -28368
rect 6780 -28368 6826 -28356
rect 6348 -28430 6420 -28370
rect 6480 -28430 6710 -28370
rect 6348 -28636 6354 -28430
rect 6780 -28480 6786 -28368
rect 6410 -28540 6640 -28480
rect 6700 -28540 6786 -28480
rect 6308 -28648 6354 -28636
rect 6780 -28636 6786 -28540
rect 6820 -28636 6826 -28368
rect 8508 -28368 8554 -28356
rect 8508 -28370 8514 -28368
rect 8500 -28430 8514 -28370
rect 6780 -28648 6826 -28636
rect 8508 -28636 8514 -28430
rect 8548 -28370 8554 -28368
rect 8980 -28368 9026 -28356
rect 8548 -28430 8840 -28370
rect 8900 -28430 8910 -28370
rect 8548 -28636 8554 -28430
rect 8980 -28480 8986 -28368
rect 8610 -28540 8840 -28480
rect 8900 -28540 8986 -28480
rect 8508 -28648 8554 -28636
rect 8980 -28636 8986 -28540
rect 9020 -28636 9026 -28368
rect 10708 -28368 10754 -28356
rect 10708 -28370 10714 -28368
rect 10700 -28430 10714 -28370
rect 8980 -28648 9026 -28636
rect 10708 -28636 10714 -28430
rect 10748 -28370 10754 -28368
rect 11180 -28368 11226 -28356
rect 10748 -28430 11040 -28370
rect 11100 -28430 11110 -28370
rect 10748 -28636 10754 -28430
rect 11180 -28480 11186 -28368
rect 10810 -28540 11040 -28480
rect 11100 -28540 11186 -28480
rect 10708 -28648 10754 -28636
rect 11180 -28636 11186 -28540
rect 11220 -28636 11226 -28368
rect 12908 -28368 12954 -28356
rect 12908 -28370 12914 -28368
rect 12900 -28430 12914 -28370
rect 11180 -28648 11226 -28636
rect 12908 -28636 12914 -28430
rect 12948 -28370 12954 -28368
rect 13380 -28368 13426 -28356
rect 12948 -28430 13240 -28370
rect 13300 -28430 13310 -28370
rect 12948 -28636 12954 -28430
rect 13380 -28480 13386 -28368
rect 13010 -28540 13240 -28480
rect 13300 -28540 13386 -28480
rect 12908 -28648 12954 -28636
rect 13380 -28636 13386 -28540
rect 13420 -28636 13426 -28368
rect 15108 -28368 15154 -28356
rect 15108 -28370 15114 -28368
rect 15100 -28430 15114 -28370
rect 13380 -28648 13426 -28636
rect 15108 -28636 15114 -28430
rect 15148 -28370 15154 -28368
rect 15580 -28368 15626 -28356
rect 15148 -28430 15440 -28370
rect 15500 -28430 15510 -28370
rect 15148 -28636 15154 -28430
rect 15580 -28480 15586 -28368
rect 15210 -28540 15220 -28480
rect 15280 -28540 15586 -28480
rect 15108 -28648 15154 -28636
rect 15580 -28636 15586 -28540
rect 15620 -28636 15626 -28368
rect 17308 -28368 17354 -28356
rect 17308 -28370 17314 -28368
rect 17300 -28430 17314 -28370
rect 15580 -28648 15626 -28636
rect 17308 -28636 17314 -28430
rect 17348 -28370 17354 -28368
rect 17780 -28368 17826 -28356
rect 17348 -28430 17420 -28370
rect 17480 -28430 17710 -28370
rect 17348 -28636 17354 -28430
rect 17780 -28480 17786 -28368
rect 17410 -28540 17786 -28480
rect 17308 -28648 17354 -28636
rect 17780 -28636 17786 -28540
rect 17820 -28636 17826 -28368
rect 19508 -28368 19554 -28356
rect 19508 -28370 19514 -28368
rect 19500 -28430 19514 -28370
rect 17780 -28648 17826 -28636
rect 19508 -28636 19514 -28430
rect 19548 -28370 19554 -28368
rect 19548 -28380 20510 -28370
rect 19548 -28430 20440 -28380
rect 19548 -28636 19554 -28430
rect 20430 -28530 20440 -28430
rect 20500 -28530 20510 -28380
rect 20430 -28540 20510 -28530
rect 19508 -28648 19554 -28636
rect 2467 -28664 4067 -28658
rect 2467 -28698 2479 -28664
rect 4055 -28698 4067 -28664
rect 2467 -28704 4067 -28698
rect 4667 -28664 6267 -28658
rect 4667 -28698 4679 -28664
rect 6255 -28698 6267 -28664
rect 4667 -28704 6267 -28698
rect 6867 -28664 8467 -28658
rect 6867 -28698 6879 -28664
rect 8455 -28698 8467 -28664
rect 6867 -28704 8467 -28698
rect 9067 -28664 10667 -28658
rect 9067 -28698 9079 -28664
rect 10655 -28698 10667 -28664
rect 9067 -28704 10667 -28698
rect 11267 -28664 12867 -28658
rect 11267 -28698 11279 -28664
rect 12855 -28698 12867 -28664
rect 11267 -28704 12867 -28698
rect 13467 -28664 15067 -28658
rect 13467 -28698 13479 -28664
rect 15055 -28698 15067 -28664
rect 13467 -28704 15067 -28698
rect 15667 -28664 17267 -28658
rect 15667 -28698 15679 -28664
rect 17255 -28698 17267 -28664
rect 15667 -28704 17267 -28698
rect 17867 -28664 19467 -28658
rect 17867 -28698 17879 -28664
rect 19455 -28698 19467 -28664
rect 17867 -28704 19467 -28698
rect 2500 -28760 2700 -28704
rect 2500 -28820 2510 -28760
rect 2690 -28820 2700 -28760
rect 2500 -28960 2700 -28820
rect 3160 -28760 3360 -28704
rect 3160 -28820 3170 -28760
rect 3350 -28820 3360 -28760
rect 3160 -28960 3360 -28820
rect 3820 -28760 4020 -28704
rect 3820 -28820 3830 -28760
rect 4010 -28820 4020 -28760
rect 3820 -28960 4020 -28820
rect 4700 -28760 4900 -28704
rect 4700 -28820 4710 -28760
rect 4890 -28820 4900 -28760
rect 4700 -28960 4900 -28820
rect 5360 -28760 5560 -28704
rect 5360 -28820 5370 -28760
rect 5550 -28820 5560 -28760
rect 5360 -28960 5560 -28820
rect 6020 -28760 6220 -28704
rect 6020 -28820 6030 -28760
rect 6210 -28820 6220 -28760
rect 6020 -28960 6220 -28820
rect 6900 -28900 7100 -28704
rect 6900 -28960 6910 -28900
rect 7090 -28960 7100 -28900
rect 7560 -28900 7760 -28704
rect 7560 -28960 7570 -28900
rect 7750 -28960 7760 -28900
rect 8220 -28900 8420 -28704
rect 8220 -28960 8230 -28900
rect 8410 -28960 8420 -28900
rect 9100 -28900 9300 -28704
rect 9100 -28960 9110 -28900
rect 9290 -28960 9300 -28900
rect 9760 -28900 9960 -28704
rect 9760 -28960 9770 -28900
rect 9950 -28960 9960 -28900
rect 10420 -28900 10620 -28704
rect 10420 -28960 10430 -28900
rect 10610 -28960 10620 -28900
rect 11300 -28900 11500 -28704
rect 11300 -28960 11310 -28900
rect 11490 -28960 11500 -28900
rect 11960 -28900 12160 -28704
rect 11960 -28960 11970 -28900
rect 12150 -28960 12160 -28900
rect 12620 -28900 12820 -28704
rect 12620 -28960 12630 -28900
rect 12810 -28960 12820 -28900
rect 13500 -28900 13700 -28704
rect 13500 -28960 13510 -28900
rect 13690 -28960 13700 -28900
rect 14160 -28900 14360 -28704
rect 14160 -28960 14170 -28900
rect 14350 -28960 14360 -28900
rect 14820 -28900 15020 -28704
rect 14820 -28960 14830 -28900
rect 15010 -28960 15020 -28900
rect 15700 -28760 15900 -28704
rect 15700 -28820 15710 -28760
rect 15890 -28820 15900 -28760
rect 15700 -28960 15900 -28820
rect 16360 -28760 16560 -28704
rect 16360 -28820 16370 -28760
rect 16550 -28820 16560 -28760
rect 16360 -28960 16560 -28820
rect 17020 -28760 17220 -28704
rect 17020 -28820 17030 -28760
rect 17210 -28820 17220 -28760
rect 17020 -28960 17220 -28820
rect 17900 -28760 18100 -28704
rect 17900 -28820 17910 -28760
rect 18090 -28820 18100 -28760
rect 17900 -28960 18100 -28820
rect 18560 -28760 18760 -28704
rect 18560 -28820 18570 -28760
rect 18750 -28820 18760 -28760
rect 18560 -28960 18760 -28820
rect 19220 -28760 19420 -28704
rect 19220 -28820 19230 -28760
rect 19410 -28820 19420 -28760
rect 19220 -28960 19420 -28820
rect 420 -29030 620 -29020
rect 420 -29110 430 -29030
rect 610 -29040 620 -29030
rect 21300 -29030 21500 -29020
rect 21300 -29040 21310 -29030
rect 610 -29100 4040 -29040
rect 4700 -29070 6220 -29060
rect 4700 -29100 4710 -29070
rect 610 -29110 620 -29100
rect 420 -29120 620 -29110
rect 2467 -29106 4067 -29100
rect 2467 -29140 2479 -29106
rect 4055 -29140 4067 -29106
rect 2467 -29146 4067 -29140
rect 4667 -29106 4710 -29100
rect 6210 -29100 6220 -29070
rect 6900 -29070 8420 -29060
rect 6900 -29100 6910 -29070
rect 6210 -29106 6267 -29100
rect 4667 -29140 4679 -29106
rect 6255 -29140 6267 -29106
rect 4667 -29146 6267 -29140
rect 6867 -29106 6910 -29100
rect 8410 -29100 8420 -29070
rect 9100 -29070 10620 -29060
rect 9100 -29100 9110 -29070
rect 8410 -29106 8467 -29100
rect 6867 -29140 6879 -29106
rect 8455 -29140 8467 -29106
rect 6867 -29146 8467 -29140
rect 9067 -29106 9110 -29100
rect 10610 -29100 10620 -29070
rect 11300 -29070 12820 -29060
rect 11300 -29100 11310 -29070
rect 10610 -29106 10667 -29100
rect 9067 -29140 9079 -29106
rect 10655 -29140 10667 -29106
rect 9067 -29146 10667 -29140
rect 11267 -29106 11310 -29100
rect 12810 -29100 12820 -29070
rect 13500 -29070 15020 -29060
rect 13500 -29100 13510 -29070
rect 12810 -29106 12867 -29100
rect 11267 -29140 11279 -29106
rect 12855 -29140 12867 -29106
rect 11267 -29146 12867 -29140
rect 13467 -29106 13510 -29100
rect 15010 -29100 15020 -29070
rect 15700 -29070 17220 -29060
rect 15700 -29100 15710 -29070
rect 15010 -29106 15067 -29100
rect 13467 -29140 13479 -29106
rect 15055 -29140 15067 -29106
rect 13467 -29146 15067 -29140
rect 15667 -29106 15710 -29100
rect 17210 -29100 17220 -29070
rect 17880 -29100 21310 -29040
rect 17210 -29106 17267 -29100
rect 15667 -29140 15679 -29106
rect 17255 -29140 17267 -29106
rect 15667 -29146 17267 -29140
rect 17867 -29106 19467 -29100
rect 17867 -29140 17879 -29106
rect 19455 -29140 19467 -29106
rect 21300 -29110 21310 -29100
rect 21490 -29110 21500 -29030
rect 21300 -29120 21500 -29110
rect 17867 -29146 19467 -29140
rect 2380 -29168 2426 -29156
rect 2380 -29260 2386 -29168
rect 1410 -29270 2386 -29260
rect 1410 -29420 1420 -29270
rect 1480 -29320 2386 -29270
rect 1480 -29420 1490 -29320
rect 1410 -29430 1490 -29420
rect 2380 -29436 2386 -29320
rect 2420 -29436 2426 -29168
rect 4108 -29168 4154 -29156
rect 4108 -29170 4114 -29168
rect 4100 -29230 4114 -29170
rect 2380 -29448 2426 -29436
rect 4108 -29436 4114 -29230
rect 4148 -29170 4154 -29168
rect 4580 -29168 4626 -29156
rect 4148 -29230 4510 -29170
rect 4148 -29436 4154 -29230
rect 4580 -29280 4586 -29168
rect 4210 -29340 4440 -29280
rect 4500 -29340 4586 -29280
rect 4108 -29448 4154 -29436
rect 4580 -29436 4586 -29340
rect 4620 -29436 4626 -29168
rect 6308 -29168 6354 -29156
rect 6308 -29170 6314 -29168
rect 6300 -29230 6314 -29170
rect 4580 -29448 4626 -29436
rect 6308 -29436 6314 -29230
rect 6348 -29170 6354 -29168
rect 6780 -29168 6826 -29156
rect 6348 -29230 6640 -29170
rect 6700 -29230 6710 -29170
rect 6348 -29436 6354 -29230
rect 6780 -29280 6786 -29168
rect 6410 -29340 6420 -29280
rect 6480 -29340 6786 -29280
rect 6308 -29448 6354 -29436
rect 6780 -29436 6786 -29340
rect 6820 -29436 6826 -29168
rect 8508 -29168 8554 -29156
rect 8508 -29170 8514 -29168
rect 8500 -29230 8514 -29170
rect 6780 -29448 6826 -29436
rect 8508 -29436 8514 -29230
rect 8548 -29170 8554 -29168
rect 8980 -29168 9026 -29156
rect 8548 -29230 8620 -29170
rect 8680 -29230 8910 -29170
rect 8548 -29436 8554 -29230
rect 8980 -29280 8986 -29168
rect 8610 -29340 8620 -29280
rect 8680 -29340 8986 -29280
rect 8508 -29448 8554 -29436
rect 8980 -29436 8986 -29340
rect 9020 -29436 9026 -29168
rect 10708 -29168 10754 -29156
rect 10708 -29170 10714 -29168
rect 10700 -29230 10714 -29170
rect 8980 -29448 9026 -29436
rect 10708 -29436 10714 -29230
rect 10748 -29170 10754 -29168
rect 11180 -29168 11226 -29156
rect 10748 -29230 10820 -29170
rect 10880 -29230 11110 -29170
rect 10748 -29436 10754 -29230
rect 11180 -29280 11186 -29168
rect 10810 -29340 10820 -29280
rect 10880 -29340 11186 -29280
rect 10708 -29448 10754 -29436
rect 11180 -29436 11186 -29340
rect 11220 -29436 11226 -29168
rect 12908 -29168 12954 -29156
rect 12908 -29170 12914 -29168
rect 12900 -29230 12914 -29170
rect 11180 -29448 11226 -29436
rect 12908 -29436 12914 -29230
rect 12948 -29170 12954 -29168
rect 13380 -29168 13426 -29156
rect 12948 -29230 13020 -29170
rect 13080 -29230 13310 -29170
rect 12948 -29436 12954 -29230
rect 13380 -29280 13386 -29168
rect 13010 -29340 13020 -29280
rect 13080 -29340 13386 -29280
rect 12908 -29448 12954 -29436
rect 13380 -29436 13386 -29340
rect 13420 -29436 13426 -29168
rect 15108 -29168 15154 -29156
rect 15108 -29170 15114 -29168
rect 15100 -29230 15114 -29170
rect 13380 -29448 13426 -29436
rect 15108 -29436 15114 -29230
rect 15148 -29170 15154 -29168
rect 15580 -29168 15626 -29156
rect 15148 -29230 15220 -29170
rect 15280 -29230 15510 -29170
rect 15148 -29436 15154 -29230
rect 15580 -29280 15586 -29168
rect 15210 -29340 15440 -29280
rect 15500 -29340 15586 -29280
rect 15108 -29448 15154 -29436
rect 15580 -29436 15586 -29340
rect 15620 -29436 15626 -29168
rect 17308 -29168 17354 -29156
rect 17308 -29170 17314 -29168
rect 17300 -29230 17314 -29170
rect 15580 -29448 15626 -29436
rect 17308 -29436 17314 -29230
rect 17348 -29170 17354 -29168
rect 17780 -29168 17826 -29156
rect 17348 -29230 17640 -29170
rect 17700 -29230 17710 -29170
rect 17348 -29436 17354 -29230
rect 17780 -29280 17786 -29168
rect 17410 -29340 17786 -29280
rect 17308 -29448 17354 -29436
rect 17780 -29436 17786 -29340
rect 17820 -29436 17826 -29168
rect 19508 -29168 19554 -29156
rect 19508 -29170 19514 -29168
rect 19500 -29230 19514 -29170
rect 17780 -29448 17826 -29436
rect 19508 -29436 19514 -29230
rect 19548 -29170 19554 -29168
rect 19548 -29180 20310 -29170
rect 19548 -29230 20240 -29180
rect 19548 -29436 19554 -29230
rect 20230 -29330 20240 -29230
rect 20300 -29330 20310 -29180
rect 20230 -29340 20310 -29330
rect 19508 -29448 19554 -29436
rect 2467 -29464 4067 -29458
rect 2467 -29498 2479 -29464
rect 4055 -29498 4067 -29464
rect 2467 -29504 4067 -29498
rect 4667 -29464 6267 -29458
rect 4667 -29498 4679 -29464
rect 6255 -29498 6267 -29464
rect 4667 -29504 6267 -29498
rect 6867 -29464 8467 -29458
rect 6867 -29498 6879 -29464
rect 8455 -29498 8467 -29464
rect 6867 -29504 8467 -29498
rect 9067 -29464 10667 -29458
rect 9067 -29498 9079 -29464
rect 10655 -29498 10667 -29464
rect 9067 -29504 10667 -29498
rect 11267 -29464 12867 -29458
rect 11267 -29498 11279 -29464
rect 12855 -29498 12867 -29464
rect 11267 -29504 12867 -29498
rect 13467 -29464 15067 -29458
rect 13467 -29498 13479 -29464
rect 15055 -29498 15067 -29464
rect 13467 -29504 15067 -29498
rect 15667 -29464 17267 -29458
rect 15667 -29498 15679 -29464
rect 17255 -29498 17267 -29464
rect 15667 -29504 17267 -29498
rect 17867 -29464 19467 -29458
rect 17867 -29498 17879 -29464
rect 19455 -29498 19467 -29464
rect 17867 -29504 19467 -29498
rect 2500 -29700 2700 -29504
rect 2500 -29760 2510 -29700
rect 2690 -29760 2700 -29700
rect 3160 -29700 3360 -29504
rect 3160 -29760 3170 -29700
rect 3350 -29760 3360 -29700
rect 3820 -29700 4020 -29504
rect 3820 -29760 3830 -29700
rect 4010 -29760 4020 -29700
rect 4700 -29700 4900 -29504
rect 4700 -29760 4710 -29700
rect 4890 -29760 4900 -29700
rect 5360 -29700 5560 -29504
rect 5360 -29760 5370 -29700
rect 5550 -29760 5560 -29700
rect 6020 -29700 6220 -29504
rect 6020 -29760 6030 -29700
rect 6210 -29760 6220 -29700
rect 6900 -29560 7100 -29504
rect 6900 -29620 6910 -29560
rect 7090 -29620 7100 -29560
rect 6900 -29760 7100 -29620
rect 7560 -29560 7760 -29504
rect 7560 -29620 7570 -29560
rect 7750 -29620 7760 -29560
rect 7560 -29760 7760 -29620
rect 8220 -29560 8420 -29504
rect 8220 -29620 8230 -29560
rect 8410 -29620 8420 -29560
rect 8220 -29760 8420 -29620
rect 9100 -29560 9300 -29504
rect 9100 -29620 9110 -29560
rect 9290 -29620 9300 -29560
rect 9100 -29760 9300 -29620
rect 9760 -29560 9960 -29504
rect 9760 -29620 9770 -29560
rect 9950 -29620 9960 -29560
rect 9760 -29760 9960 -29620
rect 10420 -29560 10620 -29504
rect 10420 -29620 10430 -29560
rect 10610 -29620 10620 -29560
rect 10420 -29760 10620 -29620
rect 11300 -29560 11500 -29504
rect 11300 -29620 11310 -29560
rect 11490 -29620 11500 -29560
rect 11300 -29760 11500 -29620
rect 11960 -29560 12160 -29504
rect 11960 -29620 11970 -29560
rect 12150 -29620 12160 -29560
rect 11960 -29760 12160 -29620
rect 12620 -29560 12820 -29504
rect 12620 -29620 12630 -29560
rect 12810 -29620 12820 -29560
rect 12620 -29760 12820 -29620
rect 13500 -29560 13700 -29504
rect 13500 -29620 13510 -29560
rect 13690 -29620 13700 -29560
rect 13500 -29760 13700 -29620
rect 14160 -29560 14360 -29504
rect 14160 -29620 14170 -29560
rect 14350 -29620 14360 -29560
rect 14160 -29760 14360 -29620
rect 14820 -29560 15020 -29504
rect 14820 -29620 14830 -29560
rect 15010 -29620 15020 -29560
rect 14820 -29760 15020 -29620
rect 15700 -29700 15900 -29504
rect 15700 -29760 15710 -29700
rect 15890 -29760 15900 -29700
rect 16360 -29700 16560 -29504
rect 16360 -29760 16370 -29700
rect 16550 -29760 16560 -29700
rect 17020 -29700 17220 -29504
rect 17020 -29760 17030 -29700
rect 17210 -29760 17220 -29700
rect 17900 -29700 18100 -29504
rect 17900 -29760 17910 -29700
rect 18090 -29760 18100 -29700
rect 18560 -29700 18760 -29504
rect 18560 -29760 18570 -29700
rect 18750 -29760 18760 -29700
rect 19220 -29700 19420 -29504
rect 19220 -29760 19230 -29700
rect 19410 -29760 19420 -29700
rect 2500 -29870 4020 -29860
rect 2500 -29900 2510 -29870
rect 2467 -29906 2510 -29900
rect 4010 -29900 4020 -29870
rect 4700 -29870 6220 -29860
rect 4700 -29900 4710 -29870
rect 4010 -29906 4067 -29900
rect 2467 -29940 2479 -29906
rect 4055 -29940 4067 -29906
rect 2467 -29946 4067 -29940
rect 4667 -29906 4710 -29900
rect 6210 -29900 6220 -29870
rect 6900 -29870 8420 -29860
rect 6900 -29900 6910 -29870
rect 6210 -29906 6267 -29900
rect 4667 -29940 4679 -29906
rect 6255 -29940 6267 -29906
rect 4667 -29946 6267 -29940
rect 6867 -29906 6910 -29900
rect 8410 -29900 8420 -29870
rect 9100 -29870 10620 -29860
rect 9100 -29900 9110 -29870
rect 8410 -29906 8467 -29900
rect 6867 -29940 6879 -29906
rect 8455 -29940 8467 -29906
rect 6867 -29946 8467 -29940
rect 9067 -29906 9110 -29900
rect 10610 -29900 10620 -29870
rect 11300 -29870 12820 -29860
rect 11300 -29900 11310 -29870
rect 10610 -29906 10667 -29900
rect 9067 -29940 9079 -29906
rect 10655 -29940 10667 -29906
rect 9067 -29946 10667 -29940
rect 11267 -29906 11310 -29900
rect 12810 -29900 12820 -29870
rect 13500 -29870 15020 -29860
rect 13500 -29900 13510 -29870
rect 12810 -29906 12867 -29900
rect 11267 -29940 11279 -29906
rect 12855 -29940 12867 -29906
rect 11267 -29946 12867 -29940
rect 13467 -29906 13510 -29900
rect 15010 -29900 15020 -29870
rect 15700 -29870 17220 -29860
rect 15700 -29900 15710 -29870
rect 15010 -29906 15067 -29900
rect 13467 -29940 13479 -29906
rect 15055 -29940 15067 -29906
rect 13467 -29946 15067 -29940
rect 15667 -29906 15710 -29900
rect 17210 -29900 17220 -29870
rect 17900 -29870 19420 -29860
rect 17900 -29900 17910 -29870
rect 17210 -29906 17267 -29900
rect 15667 -29940 15679 -29906
rect 17255 -29940 17267 -29906
rect 15667 -29946 17267 -29940
rect 17867 -29906 17910 -29900
rect 19410 -29900 19420 -29870
rect 19410 -29906 19467 -29900
rect 17867 -29940 17879 -29906
rect 19455 -29940 19467 -29906
rect 17867 -29946 19467 -29940
rect 2380 -29968 2426 -29956
rect 2380 -30060 2386 -29968
rect 2010 -30120 2020 -30060
rect 2080 -30120 2386 -30060
rect 2380 -30236 2386 -30120
rect 2420 -30236 2426 -29968
rect 4108 -29968 4154 -29956
rect 4108 -29970 4114 -29968
rect 4100 -30030 4114 -29970
rect 2380 -30248 2426 -30236
rect 4108 -30236 4114 -30030
rect 4148 -29970 4154 -29968
rect 4580 -29968 4626 -29956
rect 4148 -30030 4220 -29970
rect 4280 -30030 4510 -29970
rect 4148 -30236 4154 -30030
rect 4580 -30080 4586 -29968
rect 4210 -30140 4220 -30080
rect 4280 -30140 4586 -30080
rect 4108 -30248 4154 -30236
rect 4580 -30236 4586 -30140
rect 4620 -30236 4626 -29968
rect 6308 -29968 6354 -29956
rect 6308 -29970 6314 -29968
rect 6300 -30030 6314 -29970
rect 4580 -30248 4626 -30236
rect 6308 -30236 6314 -30030
rect 6348 -29970 6354 -29968
rect 6780 -29968 6826 -29956
rect 6348 -30030 6420 -29970
rect 6480 -30030 6710 -29970
rect 6348 -30236 6354 -30030
rect 6780 -30080 6786 -29968
rect 6410 -30140 6640 -30080
rect 6700 -30140 6786 -30080
rect 6308 -30248 6354 -30236
rect 6780 -30236 6786 -30140
rect 6820 -30236 6826 -29968
rect 8508 -29968 8554 -29956
rect 8508 -29970 8514 -29968
rect 8500 -30030 8514 -29970
rect 6780 -30248 6826 -30236
rect 8508 -30236 8514 -30030
rect 8548 -29970 8554 -29968
rect 8980 -29968 9026 -29956
rect 8548 -30030 8840 -29970
rect 8900 -30030 8910 -29970
rect 8548 -30236 8554 -30030
rect 8980 -30080 8986 -29968
rect 8610 -30140 8840 -30080
rect 8900 -30140 8986 -30080
rect 8508 -30248 8554 -30236
rect 8980 -30236 8986 -30140
rect 9020 -30236 9026 -29968
rect 10708 -29968 10754 -29956
rect 10708 -29970 10714 -29968
rect 10700 -30030 10714 -29970
rect 8980 -30248 9026 -30236
rect 10708 -30236 10714 -30030
rect 10748 -29970 10754 -29968
rect 11180 -29968 11226 -29956
rect 10748 -30030 11040 -29970
rect 11100 -30030 11110 -29970
rect 10748 -30236 10754 -30030
rect 11180 -30080 11186 -29968
rect 10810 -30140 11040 -30080
rect 11100 -30140 11186 -30080
rect 10708 -30248 10754 -30236
rect 11180 -30236 11186 -30140
rect 11220 -30236 11226 -29968
rect 12908 -29968 12954 -29956
rect 12908 -29970 12914 -29968
rect 12900 -30030 12914 -29970
rect 11180 -30248 11226 -30236
rect 12908 -30236 12914 -30030
rect 12948 -29970 12954 -29968
rect 13380 -29968 13426 -29956
rect 12948 -30030 13240 -29970
rect 13300 -30030 13310 -29970
rect 12948 -30236 12954 -30030
rect 13380 -30080 13386 -29968
rect 13010 -30140 13240 -30080
rect 13300 -30140 13386 -30080
rect 12908 -30248 12954 -30236
rect 13380 -30236 13386 -30140
rect 13420 -30236 13426 -29968
rect 15108 -29968 15154 -29956
rect 15108 -29970 15114 -29968
rect 15100 -30030 15114 -29970
rect 13380 -30248 13426 -30236
rect 15108 -30236 15114 -30030
rect 15148 -29970 15154 -29968
rect 15580 -29968 15626 -29956
rect 15148 -30030 15440 -29970
rect 15500 -30030 15510 -29970
rect 15148 -30236 15154 -30030
rect 15580 -30080 15586 -29968
rect 15210 -30140 15220 -30080
rect 15280 -30140 15586 -30080
rect 15108 -30248 15154 -30236
rect 15580 -30236 15586 -30140
rect 15620 -30236 15626 -29968
rect 17308 -29968 17354 -29956
rect 17308 -29970 17314 -29968
rect 17300 -30030 17314 -29970
rect 15580 -30248 15626 -30236
rect 17308 -30236 17314 -30030
rect 17348 -29970 17354 -29968
rect 17780 -29968 17826 -29956
rect 17348 -30030 17420 -29970
rect 17480 -30030 17710 -29970
rect 17348 -30236 17354 -30030
rect 17780 -30080 17786 -29968
rect 17410 -30140 17420 -30080
rect 17480 -30140 17786 -30080
rect 17308 -30248 17354 -30236
rect 17780 -30236 17786 -30140
rect 17820 -30236 17826 -29968
rect 19508 -29968 19554 -29956
rect 19508 -29970 19514 -29968
rect 19500 -30030 19514 -29970
rect 17780 -30248 17826 -30236
rect 19508 -30236 19514 -30030
rect 19548 -29970 19554 -29968
rect 19548 -30030 19620 -29970
rect 19680 -30030 19910 -29970
rect 19548 -30236 19554 -30030
rect 19508 -30248 19554 -30236
rect 2467 -30264 4067 -30258
rect 2467 -30298 2479 -30264
rect 4055 -30298 4067 -30264
rect 2467 -30304 4067 -30298
rect 4667 -30264 6267 -30258
rect 4667 -30298 4679 -30264
rect 6255 -30298 6267 -30264
rect 4667 -30304 6267 -30298
rect 6867 -30264 8467 -30258
rect 6867 -30298 6879 -30264
rect 8455 -30298 8467 -30264
rect 6867 -30304 8467 -30298
rect 9067 -30264 10667 -30258
rect 9067 -30298 9079 -30264
rect 10655 -30298 10667 -30264
rect 9067 -30304 10667 -30298
rect 11267 -30264 12867 -30258
rect 11267 -30298 11279 -30264
rect 12855 -30298 12867 -30264
rect 11267 -30304 12867 -30298
rect 13467 -30264 15067 -30258
rect 13467 -30298 13479 -30264
rect 15055 -30298 15067 -30264
rect 13467 -30304 15067 -30298
rect 15667 -30264 17267 -30258
rect 15667 -30298 15679 -30264
rect 17255 -30298 17267 -30264
rect 15667 -30304 17267 -30298
rect 17867 -30264 19467 -30258
rect 17867 -30298 17879 -30264
rect 19455 -30298 19467 -30264
rect 17867 -30304 19467 -30298
rect 2500 -30360 2700 -30304
rect 2500 -30420 2510 -30360
rect 2690 -30420 2700 -30360
rect 2500 -30560 2700 -30420
rect 3160 -30360 3360 -30304
rect 3160 -30420 3170 -30360
rect 3350 -30420 3360 -30360
rect 3160 -30560 3360 -30420
rect 3820 -30360 4020 -30304
rect 3820 -30420 3830 -30360
rect 4010 -30420 4020 -30360
rect 3820 -30560 4020 -30420
rect 4700 -30360 4900 -30304
rect 4700 -30420 4710 -30360
rect 4890 -30420 4900 -30360
rect 4700 -30560 4900 -30420
rect 5360 -30360 5560 -30304
rect 5360 -30420 5370 -30360
rect 5550 -30420 5560 -30360
rect 5360 -30560 5560 -30420
rect 6020 -30360 6220 -30304
rect 6020 -30420 6030 -30360
rect 6210 -30420 6220 -30360
rect 6020 -30560 6220 -30420
rect 6900 -30500 7100 -30304
rect 6900 -30560 6910 -30500
rect 7090 -30560 7100 -30500
rect 7560 -30500 7760 -30304
rect 7560 -30560 7570 -30500
rect 7750 -30560 7760 -30500
rect 8220 -30500 8420 -30304
rect 8220 -30560 8230 -30500
rect 8410 -30560 8420 -30500
rect 9100 -30500 9300 -30304
rect 9100 -30560 9110 -30500
rect 9290 -30560 9300 -30500
rect 9760 -30500 9960 -30304
rect 9760 -30560 9770 -30500
rect 9950 -30560 9960 -30500
rect 10420 -30500 10620 -30304
rect 10420 -30560 10430 -30500
rect 10610 -30560 10620 -30500
rect 11300 -30500 11500 -30304
rect 11300 -30560 11310 -30500
rect 11490 -30560 11500 -30500
rect 11960 -30500 12160 -30304
rect 11960 -30560 11970 -30500
rect 12150 -30560 12160 -30500
rect 12620 -30500 12820 -30304
rect 12620 -30560 12630 -30500
rect 12810 -30560 12820 -30500
rect 13500 -30500 13700 -30304
rect 13500 -30560 13510 -30500
rect 13690 -30560 13700 -30500
rect 14160 -30500 14360 -30304
rect 14160 -30560 14170 -30500
rect 14350 -30560 14360 -30500
rect 14820 -30500 15020 -30304
rect 14820 -30560 14830 -30500
rect 15010 -30560 15020 -30500
rect 15700 -30360 15900 -30304
rect 15700 -30420 15710 -30360
rect 15890 -30420 15900 -30360
rect 15700 -30560 15900 -30420
rect 16360 -30360 16560 -30304
rect 16360 -30420 16370 -30360
rect 16550 -30420 16560 -30360
rect 16360 -30560 16560 -30420
rect 17020 -30360 17220 -30304
rect 17020 -30420 17030 -30360
rect 17210 -30420 17220 -30360
rect 17020 -30560 17220 -30420
rect 17900 -30360 18100 -30304
rect 17900 -30420 17910 -30360
rect 18090 -30420 18100 -30360
rect 17900 -30560 18100 -30420
rect 18560 -30360 18760 -30304
rect 18560 -30420 18570 -30360
rect 18750 -30420 18760 -30360
rect 18560 -30560 18760 -30420
rect 19220 -30360 19420 -30304
rect 19220 -30420 19230 -30360
rect 19410 -30420 19420 -30360
rect 19220 -30560 19420 -30420
rect 2500 -30670 4020 -30660
rect 2500 -30700 2510 -30670
rect 2467 -30706 2510 -30700
rect 4010 -30700 4020 -30670
rect 4700 -30670 6220 -30660
rect 4700 -30700 4710 -30670
rect 4010 -30706 4067 -30700
rect 2467 -30740 2479 -30706
rect 4055 -30740 4067 -30706
rect 2467 -30746 4067 -30740
rect 4667 -30706 4710 -30700
rect 6210 -30700 6220 -30670
rect 6900 -30670 8420 -30660
rect 6900 -30700 6910 -30670
rect 6210 -30706 6267 -30700
rect 4667 -30740 4679 -30706
rect 6255 -30740 6267 -30706
rect 4667 -30746 6267 -30740
rect 6867 -30706 6910 -30700
rect 8410 -30700 8420 -30670
rect 9100 -30670 10620 -30660
rect 9100 -30700 9110 -30670
rect 8410 -30706 8467 -30700
rect 6867 -30740 6879 -30706
rect 8455 -30740 8467 -30706
rect 6867 -30746 8467 -30740
rect 9067 -30706 9110 -30700
rect 10610 -30700 10620 -30670
rect 11300 -30670 12820 -30660
rect 11300 -30700 11310 -30670
rect 10610 -30706 10667 -30700
rect 9067 -30740 9079 -30706
rect 10655 -30740 10667 -30706
rect 9067 -30746 10667 -30740
rect 11267 -30706 11310 -30700
rect 12810 -30700 12820 -30670
rect 13500 -30670 15020 -30660
rect 13500 -30700 13510 -30670
rect 12810 -30706 12867 -30700
rect 11267 -30740 11279 -30706
rect 12855 -30740 12867 -30706
rect 11267 -30746 12867 -30740
rect 13467 -30706 13510 -30700
rect 15010 -30700 15020 -30670
rect 15700 -30670 17220 -30660
rect 15700 -30700 15710 -30670
rect 15010 -30706 15067 -30700
rect 13467 -30740 13479 -30706
rect 15055 -30740 15067 -30706
rect 13467 -30746 15067 -30740
rect 15667 -30706 15710 -30700
rect 17210 -30700 17220 -30670
rect 17900 -30670 19420 -30660
rect 17900 -30700 17910 -30670
rect 17210 -30706 17267 -30700
rect 15667 -30740 15679 -30706
rect 17255 -30740 17267 -30706
rect 15667 -30746 17267 -30740
rect 17867 -30706 17910 -30700
rect 19410 -30700 19420 -30670
rect 19410 -30706 19467 -30700
rect 17867 -30740 17879 -30706
rect 19455 -30740 19467 -30706
rect 17867 -30746 19467 -30740
rect 2380 -30768 2426 -30756
rect 2380 -30860 2386 -30768
rect 2010 -30920 2240 -30860
rect 2300 -30920 2386 -30860
rect 2380 -31036 2386 -30920
rect 2420 -31036 2426 -30768
rect 4108 -30768 4154 -30756
rect 4108 -30770 4114 -30768
rect 4100 -30830 4114 -30770
rect 2380 -31048 2426 -31036
rect 4108 -31036 4114 -30830
rect 4148 -30770 4154 -30768
rect 4580 -30768 4626 -30756
rect 4148 -30830 4440 -30770
rect 4500 -30830 4510 -30770
rect 4148 -31036 4154 -30830
rect 4580 -30880 4586 -30768
rect 4210 -30940 4440 -30880
rect 4500 -30940 4586 -30880
rect 4108 -31048 4154 -31036
rect 4580 -31036 4586 -30940
rect 4620 -31036 4626 -30768
rect 6308 -30768 6354 -30756
rect 6308 -30770 6314 -30768
rect 6300 -30830 6314 -30770
rect 4580 -31048 4626 -31036
rect 6308 -31036 6314 -30830
rect 6348 -30770 6354 -30768
rect 6780 -30768 6826 -30756
rect 6348 -30830 6640 -30770
rect 6700 -30830 6710 -30770
rect 6348 -31036 6354 -30830
rect 6780 -30880 6786 -30768
rect 6410 -30940 6420 -30880
rect 6480 -30940 6786 -30880
rect 6308 -31048 6354 -31036
rect 6780 -31036 6786 -30940
rect 6820 -31036 6826 -30768
rect 8508 -30768 8554 -30756
rect 8508 -30770 8514 -30768
rect 8500 -30830 8514 -30770
rect 6780 -31048 6826 -31036
rect 8508 -31036 8514 -30830
rect 8548 -30770 8554 -30768
rect 8980 -30768 9026 -30756
rect 8548 -30830 8620 -30770
rect 8680 -30830 8910 -30770
rect 8548 -31036 8554 -30830
rect 8980 -30880 8986 -30768
rect 8610 -30940 8620 -30880
rect 8680 -30940 8986 -30880
rect 8508 -31048 8554 -31036
rect 8980 -31036 8986 -30940
rect 9020 -31036 9026 -30768
rect 10708 -30768 10754 -30756
rect 10708 -30770 10714 -30768
rect 10700 -30830 10714 -30770
rect 8980 -31048 9026 -31036
rect 10708 -31036 10714 -30830
rect 10748 -30770 10754 -30768
rect 11180 -30768 11226 -30756
rect 10748 -30830 10820 -30770
rect 10880 -30830 11110 -30770
rect 10748 -31036 10754 -30830
rect 11180 -30880 11186 -30768
rect 10810 -30940 10820 -30880
rect 10880 -30940 11186 -30880
rect 10708 -31048 10754 -31036
rect 11180 -31036 11186 -30940
rect 11220 -31036 11226 -30768
rect 12908 -30768 12954 -30756
rect 12908 -30770 12914 -30768
rect 12900 -30830 12914 -30770
rect 11180 -31048 11226 -31036
rect 12908 -31036 12914 -30830
rect 12948 -30770 12954 -30768
rect 13380 -30768 13426 -30756
rect 12948 -30830 13020 -30770
rect 13080 -30830 13310 -30770
rect 12948 -31036 12954 -30830
rect 13380 -30880 13386 -30768
rect 13010 -30940 13020 -30880
rect 13080 -30940 13386 -30880
rect 12908 -31048 12954 -31036
rect 13380 -31036 13386 -30940
rect 13420 -31036 13426 -30768
rect 15108 -30768 15154 -30756
rect 15108 -30770 15114 -30768
rect 15100 -30830 15114 -30770
rect 13380 -31048 13426 -31036
rect 15108 -31036 15114 -30830
rect 15148 -30770 15154 -30768
rect 15580 -30768 15626 -30756
rect 15148 -30830 15220 -30770
rect 15280 -30830 15510 -30770
rect 15148 -31036 15154 -30830
rect 15580 -30880 15586 -30768
rect 15210 -30940 15440 -30880
rect 15500 -30940 15586 -30880
rect 15108 -31048 15154 -31036
rect 15580 -31036 15586 -30940
rect 15620 -31036 15626 -30768
rect 17308 -30768 17354 -30756
rect 17308 -30770 17314 -30768
rect 17300 -30830 17314 -30770
rect 15580 -31048 15626 -31036
rect 17308 -31036 17314 -30830
rect 17348 -30770 17354 -30768
rect 17780 -30768 17826 -30756
rect 17348 -30830 17640 -30770
rect 17700 -30830 17710 -30770
rect 17348 -31036 17354 -30830
rect 17780 -30880 17786 -30768
rect 17410 -30940 17640 -30880
rect 17700 -30940 17786 -30880
rect 17308 -31048 17354 -31036
rect 17780 -31036 17786 -30940
rect 17820 -31036 17826 -30768
rect 19508 -30768 19554 -30756
rect 19508 -30770 19514 -30768
rect 19500 -30830 19514 -30770
rect 17780 -31048 17826 -31036
rect 19508 -31036 19514 -30830
rect 19548 -30770 19554 -30768
rect 19548 -30830 19840 -30770
rect 19900 -30830 19910 -30770
rect 19548 -31036 19554 -30830
rect 19508 -31048 19554 -31036
rect 2467 -31064 4067 -31058
rect 2467 -31098 2479 -31064
rect 4055 -31098 4067 -31064
rect 2467 -31104 4067 -31098
rect 4667 -31064 6267 -31058
rect 4667 -31098 4679 -31064
rect 6255 -31098 6267 -31064
rect 4667 -31104 6267 -31098
rect 6867 -31064 8467 -31058
rect 6867 -31098 6879 -31064
rect 8455 -31098 8467 -31064
rect 6867 -31104 8467 -31098
rect 9067 -31064 10667 -31058
rect 9067 -31098 9079 -31064
rect 10655 -31098 10667 -31064
rect 9067 -31104 10667 -31098
rect 11267 -31064 12867 -31058
rect 11267 -31098 11279 -31064
rect 12855 -31098 12867 -31064
rect 11267 -31104 12867 -31098
rect 13467 -31064 15067 -31058
rect 13467 -31098 13479 -31064
rect 15055 -31098 15067 -31064
rect 13467 -31104 15067 -31098
rect 15667 -31064 17267 -31058
rect 15667 -31098 15679 -31064
rect 17255 -31098 17267 -31064
rect 15667 -31104 17267 -31098
rect 17867 -31064 19467 -31058
rect 17867 -31098 17879 -31064
rect 19455 -31098 19467 -31064
rect 17867 -31104 19467 -31098
rect 2500 -31300 2700 -31104
rect 2500 -31360 2510 -31300
rect 2690 -31360 2700 -31300
rect 3160 -31300 3360 -31104
rect 3160 -31360 3170 -31300
rect 3350 -31360 3360 -31300
rect 3820 -31300 4020 -31104
rect 3820 -31360 3830 -31300
rect 4010 -31360 4020 -31300
rect 4700 -31300 4900 -31104
rect 4700 -31360 4710 -31300
rect 4890 -31360 4900 -31300
rect 5360 -31300 5560 -31104
rect 5360 -31360 5370 -31300
rect 5550 -31360 5560 -31300
rect 6020 -31300 6220 -31104
rect 6020 -31360 6030 -31300
rect 6210 -31360 6220 -31300
rect 6900 -31160 7100 -31104
rect 6900 -31220 6910 -31160
rect 7090 -31220 7100 -31160
rect 6900 -31360 7100 -31220
rect 7560 -31160 7760 -31104
rect 7560 -31220 7570 -31160
rect 7750 -31220 7760 -31160
rect 7560 -31360 7760 -31220
rect 8220 -31160 8420 -31104
rect 8220 -31220 8230 -31160
rect 8410 -31220 8420 -31160
rect 8220 -31360 8420 -31220
rect 9100 -31160 9300 -31104
rect 9100 -31220 9110 -31160
rect 9290 -31220 9300 -31160
rect 9100 -31360 9300 -31220
rect 9760 -31160 9960 -31104
rect 9760 -31220 9770 -31160
rect 9950 -31220 9960 -31160
rect 9760 -31360 9960 -31220
rect 10420 -31160 10620 -31104
rect 10420 -31220 10430 -31160
rect 10610 -31220 10620 -31160
rect 10420 -31360 10620 -31220
rect 11300 -31160 11500 -31104
rect 11300 -31220 11310 -31160
rect 11490 -31220 11500 -31160
rect 11300 -31360 11500 -31220
rect 11960 -31160 12160 -31104
rect 11960 -31220 11970 -31160
rect 12150 -31220 12160 -31160
rect 11960 -31360 12160 -31220
rect 12620 -31160 12820 -31104
rect 12620 -31220 12630 -31160
rect 12810 -31220 12820 -31160
rect 12620 -31360 12820 -31220
rect 13500 -31160 13700 -31104
rect 13500 -31220 13510 -31160
rect 13690 -31220 13700 -31160
rect 13500 -31360 13700 -31220
rect 14160 -31160 14360 -31104
rect 14160 -31220 14170 -31160
rect 14350 -31220 14360 -31160
rect 14160 -31360 14360 -31220
rect 14820 -31160 15020 -31104
rect 14820 -31220 14830 -31160
rect 15010 -31220 15020 -31160
rect 14820 -31360 15020 -31220
rect 15700 -31300 15900 -31104
rect 15700 -31360 15710 -31300
rect 15890 -31360 15900 -31300
rect 16360 -31300 16560 -31104
rect 16360 -31360 16370 -31300
rect 16550 -31360 16560 -31300
rect 17020 -31300 17220 -31104
rect 17020 -31360 17030 -31300
rect 17210 -31360 17220 -31300
rect 17900 -31300 18100 -31104
rect 17900 -31360 17910 -31300
rect 18090 -31360 18100 -31300
rect 18560 -31300 18760 -31104
rect 18560 -31360 18570 -31300
rect 18750 -31360 18760 -31300
rect 19220 -31300 19420 -31104
rect 19220 -31360 19230 -31300
rect 19410 -31360 19420 -31300
rect 22190 -31656 22196 -24922
rect 22230 -31656 22236 -24922
rect 22351 -25080 22363 -24683
rect 22901 -25080 22913 -24683
rect 22351 -25086 22913 -25080
rect 23017 -24683 23579 -24677
rect 23017 -25080 23029 -24683
rect 23567 -25080 23579 -24683
rect 23017 -25086 23579 -25080
rect 23683 -24680 24245 -24677
rect 24349 -24680 24911 -24677
rect 23683 -24683 24911 -24680
rect 23683 -25080 23695 -24683
rect 24233 -25080 24361 -24683
rect 24899 -25080 24911 -24683
rect 23683 -25086 24245 -25080
rect 24349 -25086 24911 -25080
rect 25015 -24680 25577 -24677
rect 25681 -24680 26243 -24677
rect 25015 -24683 26243 -24680
rect 25015 -25080 25027 -24683
rect 25565 -25080 25693 -24683
rect 26231 -25080 26243 -24683
rect 25015 -25086 25577 -25080
rect 25681 -25086 26243 -25080
rect 26347 -24683 26909 -24677
rect 26347 -25080 26359 -24683
rect 26897 -25080 26909 -24683
rect 27870 -24680 28764 -24674
rect 27870 -24720 27970 -24680
rect 28774 -24720 28820 -24712
rect 28908 -24720 28914 -24611
rect 27870 -24724 27962 -24720
rect 27870 -24810 27922 -24724
rect 27250 -24910 27922 -24810
rect 26347 -25086 26909 -25080
rect 27024 -24922 27070 -24910
rect 22190 -31668 22236 -31656
rect 22351 -31498 22913 -31492
rect 22351 -31895 22363 -31498
rect 22901 -31895 22913 -31498
rect 22351 -31901 22913 -31895
rect 23017 -31498 23579 -31492
rect 23017 -31895 23029 -31498
rect 23567 -31500 23579 -31498
rect 23683 -31498 24245 -31492
rect 23683 -31500 23695 -31498
rect 23567 -31895 23695 -31500
rect 24233 -31895 24245 -31498
rect 23017 -31900 24245 -31895
rect 23017 -31901 23579 -31900
rect 23683 -31901 24245 -31900
rect 24349 -31498 24911 -31492
rect 24349 -31895 24361 -31498
rect 24899 -31500 24911 -31498
rect 25015 -31498 25577 -31492
rect 25015 -31500 25027 -31498
rect 24899 -31895 25027 -31500
rect 25565 -31895 25577 -31498
rect 24349 -31900 25577 -31895
rect 24349 -31901 24911 -31900
rect 25015 -31901 25577 -31900
rect 25681 -31498 26243 -31492
rect 25681 -31895 25693 -31498
rect 26231 -31895 26243 -31498
rect 25681 -31901 26243 -31895
rect 26347 -31498 26909 -31492
rect 26347 -31895 26359 -31498
rect 26897 -31895 26909 -31498
rect 27024 -31656 27030 -24922
rect 27064 -31656 27070 -24922
rect 27250 -25510 27330 -24910
rect 27870 -25100 27922 -24910
rect 27956 -25100 27962 -24724
rect 27870 -25110 27962 -25100
rect 28774 -24724 28914 -24720
rect 28774 -25100 28780 -24724
rect 28814 -25100 28914 -24724
rect 28774 -25110 28914 -25100
rect 27870 -25144 27990 -25110
rect 28774 -25112 28820 -25110
rect 27870 -25150 28764 -25144
rect 27870 -25184 27984 -25150
rect 28752 -25184 28764 -25150
rect 27870 -25190 28764 -25184
rect 27870 -25200 28760 -25190
rect 28908 -25213 28914 -25110
rect 28948 -25213 28954 -24611
rect 28908 -25225 28954 -25213
rect 27919 -25288 28817 -25282
rect 27919 -25322 27931 -25288
rect 28805 -25300 28817 -25288
rect 29790 -25300 29990 -24520
rect 34800 -24490 34940 -24480
rect 35960 -24490 36140 -24460
rect 34800 -24610 34810 -24490
rect 34930 -24610 36140 -24490
rect 34800 -24620 34940 -24610
rect 28805 -25322 29990 -25300
rect 27919 -25328 29990 -25322
rect 27930 -25402 29990 -25328
rect 27910 -25408 29990 -25402
rect 27910 -25442 27931 -25408
rect 28803 -25430 29990 -25408
rect 28803 -25442 28815 -25430
rect 27910 -25448 28815 -25442
rect 27250 -25600 27260 -25510
rect 27320 -25536 27330 -25510
rect 27320 -25542 28736 -25536
rect 27320 -25576 27948 -25542
rect 28724 -25576 28736 -25542
rect 27320 -25582 28736 -25576
rect 27320 -25600 27330 -25582
rect 27250 -25610 27330 -25600
rect 28767 -25611 28814 -25599
rect 27730 -25670 27810 -25660
rect 27730 -25694 27740 -25670
rect 27260 -25740 27740 -25694
rect 27730 -25760 27740 -25740
rect 27800 -25694 27810 -25670
rect 28767 -25665 28774 -25611
rect 28808 -25665 28814 -25611
rect 28767 -25677 28814 -25665
rect 27800 -25700 28736 -25694
rect 27800 -25734 27948 -25700
rect 28724 -25734 28736 -25700
rect 27800 -25740 28736 -25734
rect 27800 -25760 27810 -25740
rect 28770 -25757 28810 -25677
rect 27730 -25770 27810 -25760
rect 28767 -25769 28814 -25757
rect 27250 -25830 27330 -25820
rect 27250 -25920 27260 -25830
rect 27320 -25852 27330 -25830
rect 28767 -25823 28774 -25769
rect 28808 -25823 28814 -25769
rect 28767 -25830 28814 -25823
rect 29370 -25770 29450 -25760
rect 29370 -25830 29380 -25770
rect 28767 -25835 29380 -25830
rect 27320 -25858 28736 -25852
rect 27320 -25892 27948 -25858
rect 28724 -25892 28736 -25858
rect 27320 -25898 28736 -25892
rect 27320 -25920 27330 -25898
rect 28770 -25915 29380 -25835
rect 27250 -25930 27330 -25920
rect 28767 -25920 29380 -25915
rect 28767 -25927 28814 -25920
rect 27730 -25985 27810 -25975
rect 27730 -26010 27740 -25985
rect 27260 -26056 27740 -26010
rect 27730 -26075 27740 -26056
rect 27800 -26010 27810 -25985
rect 28767 -25981 28774 -25927
rect 28808 -25981 28814 -25927
rect 29370 -25970 29380 -25920
rect 29440 -25970 29450 -25770
rect 29370 -25980 29450 -25970
rect 28767 -25993 28814 -25981
rect 27800 -26016 28736 -26010
rect 27800 -26050 27948 -26016
rect 28724 -26050 28736 -26016
rect 27800 -26056 28736 -26050
rect 27800 -26075 27810 -26056
rect 28770 -26073 28810 -25993
rect 27730 -26085 27810 -26075
rect 28767 -26085 28814 -26073
rect 27250 -26145 27330 -26135
rect 27250 -26235 27260 -26145
rect 27320 -26168 27330 -26145
rect 28767 -26139 28774 -26085
rect 28808 -26139 28814 -26085
rect 28767 -26151 28814 -26139
rect 27320 -26174 28736 -26168
rect 27320 -26208 27948 -26174
rect 28724 -26208 28736 -26174
rect 27320 -26214 28736 -26208
rect 27320 -26235 27330 -26214
rect 27250 -26245 27330 -26235
rect 27910 -26308 28815 -26302
rect 27910 -26342 27931 -26308
rect 28803 -26330 28815 -26308
rect 29790 -26330 29990 -25430
rect 28803 -26342 29990 -26330
rect 27910 -26348 29990 -26342
rect 27930 -26442 29990 -26348
rect 27910 -26448 29990 -26442
rect 27910 -26482 27931 -26448
rect 28803 -26460 29990 -26448
rect 28803 -26482 28815 -26460
rect 27910 -26488 28815 -26482
rect 27730 -26550 27810 -26540
rect 27730 -26576 27740 -26550
rect 27260 -26622 27740 -26576
rect 27730 -26640 27740 -26622
rect 27800 -26576 27810 -26550
rect 27800 -26582 28736 -26576
rect 27800 -26616 27948 -26582
rect 28724 -26616 28736 -26582
rect 27800 -26622 28736 -26616
rect 27800 -26640 27810 -26622
rect 27730 -26650 27810 -26640
rect 28767 -26651 28814 -26639
rect 27370 -26710 27450 -26700
rect 27370 -26734 27380 -26710
rect 27260 -26780 27380 -26734
rect 27370 -26800 27380 -26780
rect 27440 -26734 27450 -26710
rect 28767 -26705 28774 -26651
rect 28808 -26705 28814 -26651
rect 28767 -26717 28814 -26705
rect 27440 -26740 28736 -26734
rect 27440 -26774 27948 -26740
rect 28724 -26774 28736 -26740
rect 27440 -26780 28736 -26774
rect 27440 -26800 27450 -26780
rect 28770 -26797 28810 -26717
rect 27370 -26810 27450 -26800
rect 28767 -26809 28814 -26797
rect 27730 -26870 27810 -26860
rect 27730 -26892 27740 -26870
rect 27260 -26938 27740 -26892
rect 27730 -26960 27740 -26938
rect 27800 -26892 27810 -26870
rect 28767 -26863 28774 -26809
rect 28808 -26863 28814 -26809
rect 28767 -26870 28814 -26863
rect 29520 -26810 29600 -26800
rect 29520 -26870 29530 -26810
rect 28767 -26875 29530 -26870
rect 27800 -26898 28736 -26892
rect 27800 -26932 27948 -26898
rect 28724 -26932 28736 -26898
rect 27800 -26938 28736 -26932
rect 27800 -26960 27810 -26938
rect 28770 -26955 29530 -26875
rect 27730 -26970 27810 -26960
rect 28767 -26960 29530 -26955
rect 28767 -26967 28814 -26960
rect 27370 -27025 27450 -27015
rect 27370 -27050 27380 -27025
rect 27260 -27096 27380 -27050
rect 27370 -27115 27380 -27096
rect 27440 -27050 27450 -27025
rect 28767 -27021 28774 -26967
rect 28808 -27021 28814 -26967
rect 29520 -27010 29530 -26960
rect 29590 -27010 29600 -26810
rect 29520 -27020 29600 -27010
rect 28767 -27033 28814 -27021
rect 27440 -27056 28736 -27050
rect 27440 -27090 27948 -27056
rect 28724 -27090 28736 -27056
rect 27440 -27096 28736 -27090
rect 27440 -27115 27450 -27096
rect 28770 -27113 28810 -27033
rect 27370 -27125 27450 -27115
rect 28767 -27125 28814 -27113
rect 27730 -27185 27810 -27175
rect 27730 -27208 27740 -27185
rect 27260 -27254 27740 -27208
rect 27730 -27275 27740 -27254
rect 27800 -27208 27810 -27185
rect 28767 -27179 28774 -27125
rect 28808 -27179 28814 -27125
rect 28767 -27191 28814 -27179
rect 27800 -27214 28736 -27208
rect 27800 -27248 27948 -27214
rect 28724 -27248 28736 -27214
rect 27800 -27254 28736 -27248
rect 27800 -27275 27810 -27254
rect 27730 -27285 27810 -27275
rect 27910 -27348 28815 -27342
rect 27910 -27382 27931 -27348
rect 28803 -27370 28815 -27348
rect 29790 -27370 29990 -26460
rect 34630 -24830 34730 -24700
rect 34977 -24830 35777 -24824
rect 34630 -24860 34989 -24830
rect 34630 -25350 34730 -24860
rect 34977 -24864 34989 -24860
rect 35765 -24864 35777 -24830
rect 34977 -24870 35777 -24864
rect 34890 -24909 34936 -24897
rect 34890 -24930 34896 -24909
rect 34800 -24940 34896 -24930
rect 34930 -24930 34936 -24909
rect 35818 -24909 35864 -24897
rect 35818 -24930 35824 -24909
rect 34800 -25010 34810 -24940
rect 34800 -25043 34896 -25010
rect 34930 -25020 35824 -24930
rect 34930 -25043 34936 -25020
rect 34800 -25055 34936 -25043
rect 35818 -25043 35824 -25020
rect 35858 -25043 35864 -24909
rect 35818 -25055 35864 -25043
rect 34800 -25155 34900 -25055
rect 34977 -25088 35777 -25082
rect 34977 -25122 34989 -25088
rect 35765 -25090 35777 -25088
rect 35960 -25090 36140 -24610
rect 36317 -24830 37117 -24824
rect 37330 -24830 37430 -24710
rect 36317 -24864 36329 -24830
rect 37105 -24860 37430 -24830
rect 37105 -24864 37117 -24860
rect 36317 -24870 37117 -24864
rect 36230 -24909 36276 -24897
rect 36230 -25043 36236 -24909
rect 36270 -24930 36276 -24909
rect 37158 -24909 37204 -24897
rect 37158 -24930 37164 -24909
rect 36270 -25020 37164 -24930
rect 37198 -24930 37204 -24909
rect 37198 -24940 37290 -24930
rect 37280 -25010 37290 -24940
rect 36270 -25043 36276 -25020
rect 36230 -25055 36276 -25043
rect 37158 -25043 37164 -25020
rect 37198 -25043 37290 -25010
rect 37158 -25055 37290 -25043
rect 36317 -25088 37117 -25082
rect 36317 -25090 36329 -25088
rect 35765 -25120 36329 -25090
rect 35765 -25122 35777 -25120
rect 34977 -25128 35777 -25122
rect 34800 -25167 34936 -25155
rect 34800 -25200 34896 -25167
rect 34930 -25190 34936 -25167
rect 35818 -25167 35864 -25155
rect 35818 -25190 35824 -25167
rect 34800 -25270 34810 -25200
rect 34800 -25280 34896 -25270
rect 34890 -25301 34896 -25280
rect 34930 -25280 35824 -25190
rect 34930 -25301 34936 -25280
rect 34890 -25313 34936 -25301
rect 35818 -25301 35824 -25280
rect 35858 -25301 35864 -25167
rect 35818 -25313 35864 -25301
rect 34977 -25346 35777 -25340
rect 34977 -25350 34989 -25346
rect 34630 -25380 34989 -25350
rect 35765 -25380 35777 -25346
rect 34630 -25860 34730 -25380
rect 34977 -25386 35777 -25380
rect 34890 -25425 34936 -25413
rect 34890 -25450 34896 -25425
rect 34800 -25460 34896 -25450
rect 34930 -25450 34936 -25425
rect 35818 -25425 35864 -25413
rect 35818 -25450 35824 -25425
rect 34800 -25530 34810 -25460
rect 34800 -25559 34896 -25530
rect 34930 -25540 35824 -25450
rect 34930 -25559 34936 -25540
rect 34800 -25571 34936 -25559
rect 35818 -25559 35824 -25540
rect 35858 -25559 35864 -25425
rect 35818 -25571 35864 -25559
rect 34800 -25671 34900 -25571
rect 34977 -25604 35777 -25598
rect 34977 -25638 34989 -25604
rect 35765 -25610 35777 -25604
rect 35960 -25610 36140 -25120
rect 36317 -25122 36329 -25120
rect 37105 -25122 37117 -25088
rect 36317 -25128 37117 -25122
rect 37180 -25155 37290 -25055
rect 36230 -25167 36276 -25155
rect 36230 -25301 36236 -25167
rect 36270 -25190 36276 -25167
rect 37158 -25167 37290 -25155
rect 37158 -25190 37164 -25167
rect 36270 -25280 37164 -25190
rect 37198 -25200 37290 -25167
rect 37280 -25270 37290 -25200
rect 36270 -25301 36276 -25280
rect 36230 -25313 36276 -25301
rect 37158 -25301 37164 -25280
rect 37198 -25280 37290 -25270
rect 37198 -25301 37204 -25280
rect 37158 -25313 37204 -25301
rect 36317 -25346 37117 -25340
rect 36317 -25380 36329 -25346
rect 37105 -25350 37117 -25346
rect 37330 -25350 37430 -24860
rect 37105 -25380 37430 -25350
rect 36317 -25386 37117 -25380
rect 36230 -25425 36276 -25413
rect 36230 -25559 36236 -25425
rect 36270 -25450 36276 -25425
rect 37158 -25425 37204 -25413
rect 37158 -25450 37164 -25425
rect 36270 -25540 37164 -25450
rect 37198 -25450 37204 -25425
rect 37198 -25460 37290 -25450
rect 37280 -25530 37290 -25460
rect 36270 -25559 36276 -25540
rect 36230 -25571 36276 -25559
rect 37158 -25559 37164 -25540
rect 37198 -25559 37290 -25530
rect 37158 -25571 37290 -25559
rect 36317 -25604 37117 -25598
rect 36317 -25610 36329 -25604
rect 35765 -25638 36329 -25610
rect 37105 -25638 37117 -25604
rect 34977 -25640 37117 -25638
rect 34977 -25644 35777 -25640
rect 34800 -25683 34936 -25671
rect 34800 -25720 34896 -25683
rect 34930 -25710 34936 -25683
rect 35818 -25683 35864 -25671
rect 35818 -25710 35824 -25683
rect 34800 -25790 34810 -25720
rect 34800 -25800 34896 -25790
rect 34890 -25817 34896 -25800
rect 34930 -25800 35824 -25710
rect 34930 -25817 34936 -25800
rect 34890 -25829 34936 -25817
rect 35818 -25817 35824 -25800
rect 35858 -25817 35864 -25683
rect 35818 -25829 35864 -25817
rect 34977 -25860 35777 -25856
rect 34630 -25862 35777 -25860
rect 34630 -25890 34989 -25862
rect 34630 -26380 34730 -25890
rect 34977 -25896 34989 -25890
rect 35765 -25896 35777 -25862
rect 34977 -25902 35777 -25896
rect 34890 -25941 34936 -25929
rect 34890 -25970 34896 -25941
rect 34800 -25980 34896 -25970
rect 34930 -25970 34936 -25941
rect 35818 -25941 35864 -25929
rect 35818 -25970 35824 -25941
rect 34800 -26050 34810 -25980
rect 34800 -26075 34896 -26050
rect 34930 -26060 35824 -25970
rect 34930 -26075 34936 -26060
rect 34800 -26087 34936 -26075
rect 35818 -26075 35824 -26060
rect 35858 -26075 35864 -25941
rect 35818 -26087 35864 -26075
rect 34800 -26187 34900 -26087
rect 34977 -26120 35777 -26114
rect 35960 -26120 36140 -25640
rect 36317 -25644 37117 -25640
rect 37180 -25671 37290 -25571
rect 36230 -25683 36276 -25671
rect 36230 -25817 36236 -25683
rect 36270 -25710 36276 -25683
rect 37158 -25683 37290 -25671
rect 37158 -25710 37164 -25683
rect 36270 -25800 37164 -25710
rect 37198 -25720 37290 -25683
rect 37280 -25790 37290 -25720
rect 36270 -25817 36276 -25800
rect 36230 -25829 36276 -25817
rect 37158 -25817 37164 -25800
rect 37198 -25800 37290 -25790
rect 37198 -25817 37204 -25800
rect 37158 -25829 37204 -25817
rect 36317 -25860 37117 -25856
rect 37330 -25860 37430 -25380
rect 36317 -25862 37430 -25860
rect 36317 -25896 36329 -25862
rect 37105 -25890 37430 -25862
rect 37105 -25896 37117 -25890
rect 36317 -25902 37117 -25896
rect 36230 -25941 36276 -25929
rect 36230 -26075 36236 -25941
rect 36270 -25970 36276 -25941
rect 37158 -25941 37204 -25929
rect 37158 -25970 37164 -25941
rect 36270 -26060 37164 -25970
rect 37198 -25970 37204 -25941
rect 37198 -25980 37290 -25970
rect 37280 -26050 37290 -25980
rect 36270 -26075 36276 -26060
rect 36230 -26087 36276 -26075
rect 37158 -26075 37164 -26060
rect 37198 -26075 37290 -26050
rect 37158 -26087 37290 -26075
rect 36317 -26120 37117 -26114
rect 34977 -26154 34989 -26120
rect 35765 -26150 36329 -26120
rect 35765 -26154 35777 -26150
rect 34977 -26160 35777 -26154
rect 34800 -26199 34936 -26187
rect 34800 -26240 34896 -26199
rect 34930 -26230 34936 -26199
rect 35818 -26199 35864 -26187
rect 35818 -26230 35824 -26199
rect 34800 -26310 34810 -26240
rect 34800 -26320 34896 -26310
rect 34890 -26333 34896 -26320
rect 34930 -26320 35824 -26230
rect 34930 -26333 34936 -26320
rect 34890 -26345 34936 -26333
rect 35818 -26333 35824 -26320
rect 35858 -26333 35864 -26199
rect 35818 -26345 35864 -26333
rect 34977 -26378 35777 -26372
rect 34977 -26380 34989 -26378
rect 34630 -26410 34989 -26380
rect 34630 -26900 34730 -26410
rect 34977 -26412 34989 -26410
rect 35765 -26412 35777 -26378
rect 34977 -26418 35777 -26412
rect 34890 -26457 34936 -26445
rect 34890 -26490 34896 -26457
rect 34800 -26500 34896 -26490
rect 34930 -26490 34936 -26457
rect 35818 -26457 35864 -26445
rect 35818 -26490 35824 -26457
rect 34800 -26570 34810 -26500
rect 34800 -26591 34896 -26570
rect 34930 -26580 35824 -26490
rect 34930 -26591 34936 -26580
rect 34800 -26603 34936 -26591
rect 35818 -26591 35824 -26580
rect 35858 -26591 35864 -26457
rect 35818 -26603 35864 -26591
rect 34800 -26703 34900 -26603
rect 34977 -26636 35777 -26630
rect 34977 -26670 34989 -26636
rect 35765 -26640 35777 -26636
rect 35960 -26640 36140 -26150
rect 36317 -26154 36329 -26150
rect 37105 -26154 37117 -26120
rect 36317 -26160 37117 -26154
rect 37180 -26187 37290 -26087
rect 36230 -26199 36276 -26187
rect 36230 -26333 36236 -26199
rect 36270 -26230 36276 -26199
rect 37158 -26199 37290 -26187
rect 37158 -26230 37164 -26199
rect 36270 -26320 37164 -26230
rect 37198 -26240 37290 -26199
rect 37280 -26310 37290 -26240
rect 36270 -26333 36276 -26320
rect 36230 -26345 36276 -26333
rect 37158 -26333 37164 -26320
rect 37198 -26320 37290 -26310
rect 37198 -26333 37204 -26320
rect 37158 -26345 37204 -26333
rect 36317 -26378 37117 -26372
rect 36317 -26412 36329 -26378
rect 37105 -26380 37117 -26378
rect 37330 -26380 37430 -25890
rect 37105 -26410 37430 -26380
rect 37105 -26412 37117 -26410
rect 36317 -26418 37117 -26412
rect 36230 -26457 36276 -26445
rect 36230 -26591 36236 -26457
rect 36270 -26490 36276 -26457
rect 37158 -26457 37204 -26445
rect 37158 -26490 37164 -26457
rect 36270 -26580 37164 -26490
rect 37198 -26490 37204 -26457
rect 37198 -26500 37290 -26490
rect 37280 -26570 37290 -26500
rect 36270 -26591 36276 -26580
rect 36230 -26603 36276 -26591
rect 37158 -26591 37164 -26580
rect 37198 -26591 37290 -26570
rect 37158 -26603 37290 -26591
rect 36317 -26636 37117 -26630
rect 36317 -26640 36329 -26636
rect 35765 -26670 36329 -26640
rect 37105 -26670 37117 -26636
rect 34977 -26676 35777 -26670
rect 34800 -26715 34936 -26703
rect 34800 -26760 34896 -26715
rect 34930 -26750 34936 -26715
rect 35818 -26715 35864 -26703
rect 35818 -26750 35824 -26715
rect 34800 -26830 34810 -26760
rect 34800 -26840 34896 -26830
rect 34890 -26849 34896 -26840
rect 34930 -26840 35824 -26750
rect 34930 -26849 34936 -26840
rect 34890 -26861 34936 -26849
rect 35818 -26849 35824 -26840
rect 35858 -26849 35864 -26715
rect 35818 -26861 35864 -26849
rect 34977 -26894 35777 -26888
rect 34977 -26900 34989 -26894
rect 34630 -26928 34989 -26900
rect 35765 -26928 35777 -26894
rect 35960 -26910 36140 -26670
rect 36317 -26676 37117 -26670
rect 37180 -26703 37290 -26603
rect 36230 -26715 36276 -26703
rect 36230 -26849 36236 -26715
rect 36270 -26750 36276 -26715
rect 37158 -26715 37290 -26703
rect 37158 -26750 37164 -26715
rect 36270 -26840 37164 -26750
rect 37198 -26760 37290 -26715
rect 37280 -26830 37290 -26760
rect 36270 -26849 36276 -26840
rect 36230 -26861 36276 -26849
rect 37158 -26849 37164 -26840
rect 37198 -26840 37290 -26830
rect 37198 -26849 37204 -26840
rect 37158 -26861 37204 -26849
rect 36317 -26894 37117 -26888
rect 34630 -26930 35777 -26928
rect 34630 -27020 34730 -26930
rect 34977 -26934 35777 -26930
rect 36317 -26928 36329 -26894
rect 37105 -26900 37117 -26894
rect 37330 -26900 37430 -26410
rect 37105 -26928 37430 -26900
rect 36317 -26930 37430 -26928
rect 36317 -26934 37117 -26930
rect 36020 -27010 36420 -27000
rect 36020 -27020 36030 -27010
rect 34630 -27130 36030 -27020
rect 36020 -27140 36030 -27130
rect 36410 -27140 36420 -27010
rect 36020 -27150 36420 -27140
rect 36520 -27010 36920 -27000
rect 36520 -27140 36530 -27010
rect 36910 -27020 36920 -27010
rect 37330 -27020 37430 -26930
rect 36910 -27130 37430 -27020
rect 36910 -27140 36920 -27130
rect 36520 -27150 36920 -27140
rect 28803 -27382 29990 -27370
rect 27910 -27388 29990 -27382
rect 27930 -27482 29990 -27388
rect 27910 -27488 29990 -27482
rect 27910 -27522 27931 -27488
rect 28803 -27500 29990 -27488
rect 28803 -27522 28815 -27500
rect 27910 -27528 28815 -27522
rect 27250 -27595 27330 -27585
rect 27250 -27685 27260 -27595
rect 27320 -27616 27330 -27595
rect 27320 -27622 28736 -27616
rect 27320 -27656 27948 -27622
rect 28724 -27656 28736 -27622
rect 27320 -27662 28736 -27656
rect 27320 -27685 27330 -27662
rect 27250 -27695 27330 -27685
rect 28767 -27691 28814 -27679
rect 27490 -27750 27570 -27740
rect 27490 -27774 27500 -27750
rect 27260 -27820 27500 -27774
rect 27490 -27840 27500 -27820
rect 27560 -27774 27570 -27750
rect 28767 -27745 28774 -27691
rect 28808 -27745 28814 -27691
rect 28767 -27757 28814 -27745
rect 27560 -27780 28736 -27774
rect 27560 -27814 27948 -27780
rect 28724 -27814 28736 -27780
rect 27560 -27820 28736 -27814
rect 27560 -27840 27570 -27820
rect 28770 -27837 28810 -27757
rect 27490 -27850 27570 -27840
rect 28767 -27849 28814 -27837
rect 27250 -27910 27330 -27900
rect 27250 -28000 27260 -27910
rect 27320 -27932 27330 -27910
rect 28767 -27903 28774 -27849
rect 28808 -27903 28814 -27849
rect 28767 -27910 28814 -27903
rect 29070 -27850 29150 -27840
rect 29070 -27910 29080 -27850
rect 28767 -27915 29080 -27910
rect 27320 -27938 28736 -27932
rect 27320 -27972 27948 -27938
rect 28724 -27972 28736 -27938
rect 27320 -27978 28736 -27972
rect 27320 -28000 27330 -27978
rect 28770 -27995 29080 -27915
rect 27250 -28010 27330 -28000
rect 28767 -28000 29080 -27995
rect 28767 -28007 28814 -28000
rect 27490 -28065 27570 -28055
rect 27490 -28090 27500 -28065
rect 27260 -28136 27500 -28090
rect 27490 -28155 27500 -28136
rect 27560 -28090 27570 -28065
rect 28767 -28061 28774 -28007
rect 28808 -28061 28814 -28007
rect 29070 -28050 29080 -28000
rect 29140 -28050 29150 -27850
rect 29070 -28060 29150 -28050
rect 28767 -28073 28814 -28061
rect 27560 -28096 28736 -28090
rect 27560 -28130 27948 -28096
rect 28724 -28130 28736 -28096
rect 27560 -28136 28736 -28130
rect 27560 -28155 27570 -28136
rect 28770 -28153 28810 -28073
rect 27490 -28165 27570 -28155
rect 28767 -28165 28814 -28153
rect 27250 -28225 27330 -28215
rect 27250 -28315 27260 -28225
rect 27320 -28248 27330 -28225
rect 28767 -28219 28774 -28165
rect 28808 -28219 28814 -28165
rect 28767 -28231 28814 -28219
rect 27320 -28254 28736 -28248
rect 27320 -28288 27948 -28254
rect 28724 -28288 28736 -28254
rect 27320 -28294 28736 -28288
rect 27320 -28315 27330 -28294
rect 27250 -28325 27330 -28315
rect 27910 -28388 28815 -28382
rect 27910 -28422 27931 -28388
rect 28803 -28410 28815 -28388
rect 29790 -28410 29990 -27500
rect 31630 -28050 38160 -28020
rect 31630 -28290 31820 -28050
rect 33160 -28290 38160 -28050
rect 31630 -28302 38160 -28290
rect 31630 -28336 31712 -28302
rect 32104 -28336 32152 -28302
rect 32544 -28336 32592 -28302
rect 32984 -28320 33912 -28302
rect 32984 -28336 33710 -28320
rect 31630 -28360 33710 -28336
rect 33830 -28336 33912 -28320
rect 34304 -28336 34352 -28302
rect 34744 -28336 34792 -28302
rect 35184 -28320 36112 -28302
rect 35184 -28336 35910 -28320
rect 33830 -28360 35910 -28336
rect 36030 -28336 36112 -28320
rect 36504 -28336 36552 -28302
rect 36944 -28336 36992 -28302
rect 37384 -28320 38160 -28302
rect 37384 -28336 38110 -28320
rect 36030 -28360 38110 -28336
rect 28803 -28422 29990 -28410
rect 27910 -28428 29990 -28422
rect 27930 -28522 29990 -28428
rect 27910 -28528 29990 -28522
rect 27910 -28562 27931 -28528
rect 28803 -28540 29990 -28528
rect 28803 -28562 28815 -28540
rect 27910 -28568 28815 -28562
rect 27250 -28630 27330 -28620
rect 27250 -28720 27260 -28630
rect 27320 -28656 27330 -28630
rect 27320 -28662 28736 -28656
rect 27320 -28696 27948 -28662
rect 28724 -28696 28736 -28662
rect 27320 -28702 28736 -28696
rect 27320 -28720 27330 -28702
rect 27250 -28730 27330 -28720
rect 28767 -28731 28814 -28719
rect 27610 -28790 27690 -28780
rect 27610 -28814 27620 -28790
rect 27260 -28860 27620 -28814
rect 27610 -28880 27620 -28860
rect 27680 -28814 27690 -28790
rect 28767 -28785 28774 -28731
rect 28808 -28785 28814 -28731
rect 28767 -28797 28814 -28785
rect 27680 -28820 28736 -28814
rect 27680 -28854 27948 -28820
rect 28724 -28854 28736 -28820
rect 27680 -28860 28736 -28854
rect 27680 -28880 27690 -28860
rect 28770 -28877 28810 -28797
rect 27610 -28890 27690 -28880
rect 28767 -28889 28814 -28877
rect 27250 -28950 27330 -28940
rect 27250 -29040 27260 -28950
rect 27320 -28972 27330 -28950
rect 28767 -28943 28774 -28889
rect 28808 -28943 28814 -28889
rect 28767 -28950 28814 -28943
rect 29220 -28890 29300 -28880
rect 29220 -28950 29230 -28890
rect 28767 -28955 29230 -28950
rect 27320 -28978 28736 -28972
rect 27320 -29012 27948 -28978
rect 28724 -29012 28736 -28978
rect 27320 -29018 28736 -29012
rect 27320 -29040 27330 -29018
rect 28770 -29035 29230 -28955
rect 27250 -29050 27330 -29040
rect 28767 -29040 29230 -29035
rect 28767 -29047 28814 -29040
rect 27610 -29110 27690 -29100
rect 27610 -29130 27620 -29110
rect 27260 -29176 27620 -29130
rect 27610 -29200 27620 -29176
rect 27680 -29130 27690 -29110
rect 28767 -29101 28774 -29047
rect 28808 -29101 28814 -29047
rect 29220 -29090 29230 -29040
rect 29290 -29090 29300 -28890
rect 29220 -29100 29300 -29090
rect 28767 -29113 28814 -29101
rect 27680 -29136 28736 -29130
rect 27680 -29170 27948 -29136
rect 28724 -29170 28736 -29136
rect 27680 -29176 28736 -29170
rect 27680 -29200 27690 -29176
rect 28770 -29193 28810 -29113
rect 27610 -29210 27690 -29200
rect 28767 -29205 28814 -29193
rect 27250 -29260 27330 -29250
rect 27250 -29350 27260 -29260
rect 27320 -29288 27330 -29260
rect 28767 -29259 28774 -29205
rect 28808 -29259 28814 -29205
rect 28767 -29271 28814 -29259
rect 27320 -29294 28736 -29288
rect 27320 -29328 27948 -29294
rect 28724 -29328 28736 -29294
rect 27320 -29334 28736 -29328
rect 27320 -29350 27330 -29334
rect 27250 -29360 27330 -29350
rect 27910 -29428 28815 -29422
rect 27910 -29462 27931 -29428
rect 28803 -29450 28815 -29428
rect 29790 -29450 29990 -28540
rect 31784 -28521 31828 -28360
rect 31876 -28440 32152 -28434
rect 31876 -28474 31888 -28440
rect 31928 -28474 32152 -28440
rect 31876 -28480 32152 -28474
rect 32316 -28440 32380 -28434
rect 32316 -28474 32328 -28440
rect 32368 -28474 32380 -28440
rect 32316 -28480 32380 -28474
rect 31784 -28533 31852 -28521
rect 31784 -28909 31812 -28533
rect 31846 -28909 31852 -28533
rect 31784 -28920 31852 -28909
rect 31806 -28921 31852 -28920
rect 31888 -28962 31928 -28480
rect 31964 -28522 32010 -28521
rect 31964 -28528 32058 -28522
rect 31964 -28533 31994 -28528
rect 31964 -28909 31970 -28533
rect 32052 -28874 32058 -28528
rect 32104 -28524 32152 -28480
rect 32246 -28522 32292 -28521
rect 32200 -28524 32292 -28522
rect 32104 -28528 32292 -28524
rect 32104 -28570 32206 -28528
rect 32264 -28533 32292 -28528
rect 31964 -28914 31994 -28909
rect 32052 -28914 32152 -28874
rect 31964 -28920 32152 -28914
rect 32200 -28914 32206 -28570
rect 32286 -28909 32292 -28533
rect 32264 -28914 32292 -28909
rect 32200 -28920 32292 -28914
rect 31964 -28921 32010 -28920
rect 32104 -28962 32152 -28920
rect 32246 -28921 32292 -28920
rect 32328 -28962 32368 -28480
rect 32428 -28521 32472 -28360
rect 32756 -28440 32820 -28434
rect 32756 -28474 32768 -28440
rect 32808 -28474 32820 -28440
rect 32756 -28480 32820 -28474
rect 32404 -28533 32472 -28521
rect 32686 -28522 32732 -28521
rect 32404 -28909 32410 -28533
rect 32444 -28909 32472 -28533
rect 32404 -28920 32472 -28909
rect 32664 -28533 32732 -28522
rect 32664 -28909 32692 -28533
rect 32726 -28909 32732 -28533
rect 32404 -28921 32450 -28920
rect 32664 -28921 32732 -28909
rect 31876 -28968 31940 -28962
rect 31876 -29002 31888 -28968
rect 31928 -29002 31940 -28968
rect 31876 -29008 31940 -29002
rect 32104 -28968 32380 -28962
rect 32104 -29002 32328 -28968
rect 32368 -29002 32380 -28968
rect 32104 -29008 32380 -29002
rect 31888 -29020 31928 -29008
rect 32328 -29020 32368 -29008
rect 32664 -29152 32708 -28921
rect 32768 -28962 32808 -28480
rect 32866 -28521 32910 -28360
rect 32844 -28533 32910 -28521
rect 32844 -28909 32850 -28533
rect 32884 -28909 32910 -28533
rect 32994 -28602 33710 -28360
rect 32994 -28608 33075 -28602
rect 32844 -28920 32910 -28909
rect 32966 -28636 33075 -28608
rect 33629 -28636 33710 -28602
rect 32966 -28642 33710 -28636
rect 33984 -28521 34028 -28360
rect 34076 -28440 34352 -28434
rect 34076 -28474 34088 -28440
rect 34128 -28474 34352 -28440
rect 34076 -28480 34352 -28474
rect 34516 -28440 34580 -28434
rect 34516 -28474 34528 -28440
rect 34568 -28474 34580 -28440
rect 34516 -28480 34580 -28474
rect 33984 -28533 34052 -28521
rect 32966 -28683 33012 -28642
rect 32844 -28921 32890 -28920
rect 32756 -28968 32820 -28962
rect 32756 -29002 32768 -28968
rect 32808 -29002 32820 -28968
rect 32756 -29008 32820 -29002
rect 28803 -29462 29990 -29450
rect 27910 -29468 29990 -29462
rect 31888 -29212 32708 -29152
rect 31888 -29463 31928 -29212
rect 32328 -29276 32478 -29270
rect 32328 -29334 32334 -29276
rect 32472 -29334 32478 -29276
rect 32328 -29340 32478 -29334
rect 32102 -29420 32160 -29408
rect 27920 -29562 29990 -29468
rect 31863 -29469 31955 -29463
rect 31863 -29503 31875 -29469
rect 31943 -29503 31955 -29469
rect 31863 -29509 31955 -29503
rect 27910 -29568 29990 -29562
rect 27910 -29602 27931 -29568
rect 28803 -29580 29990 -29568
rect 28803 -29602 28815 -29580
rect 27910 -29608 28815 -29602
rect 27370 -29670 27450 -29660
rect 27370 -29696 27380 -29670
rect 27260 -29742 27380 -29696
rect 27370 -29760 27380 -29742
rect 27440 -29696 27450 -29670
rect 27440 -29702 28736 -29696
rect 27440 -29736 27948 -29702
rect 28724 -29736 28736 -29702
rect 27440 -29742 28736 -29736
rect 27440 -29760 27450 -29742
rect 27370 -29770 27450 -29760
rect 28767 -29771 28814 -29759
rect 27610 -29830 27690 -29820
rect 27610 -29854 27620 -29830
rect 27260 -29900 27620 -29854
rect 27610 -29920 27620 -29900
rect 27680 -29854 27690 -29830
rect 28767 -29825 28774 -29771
rect 28808 -29825 28814 -29771
rect 28767 -29837 28814 -29825
rect 27680 -29860 28736 -29854
rect 27680 -29894 27948 -29860
rect 28724 -29894 28736 -29860
rect 27680 -29900 28736 -29894
rect 27680 -29920 27690 -29900
rect 28770 -29917 28810 -29837
rect 29790 -29900 29990 -29580
rect 31786 -29541 31830 -29538
rect 31786 -29553 31853 -29541
rect 31786 -29729 31813 -29553
rect 31847 -29729 31853 -29553
rect 31786 -29741 31853 -29729
rect 31786 -29900 31830 -29741
rect 31888 -29773 31928 -29509
rect 31965 -29542 32011 -29541
rect 31965 -29548 32058 -29542
rect 31965 -29553 31994 -29548
rect 31965 -29729 31971 -29553
rect 31965 -29734 31994 -29729
rect 32052 -29734 32058 -29548
rect 31965 -29740 32058 -29734
rect 31965 -29741 32011 -29740
rect 31863 -29779 31955 -29773
rect 31863 -29813 31875 -29779
rect 31943 -29813 31955 -29779
rect 31863 -29819 31955 -29813
rect 31888 -29820 31928 -29819
rect 32102 -29862 32119 -29420
rect 32153 -29862 32160 -29420
rect 32328 -29463 32368 -29340
rect 32303 -29469 32395 -29463
rect 32303 -29503 32315 -29469
rect 32383 -29503 32395 -29469
rect 32303 -29509 32395 -29503
rect 32247 -29542 32293 -29541
rect 32226 -29544 32293 -29542
rect 32200 -29550 32293 -29544
rect 32200 -29736 32206 -29550
rect 32264 -29553 32293 -29550
rect 32287 -29729 32293 -29553
rect 32264 -29736 32293 -29729
rect 32200 -29741 32293 -29736
rect 32200 -29742 32270 -29741
rect 32328 -29773 32368 -29509
rect 32428 -29541 32472 -29538
rect 32405 -29553 32472 -29541
rect 32405 -29729 32411 -29553
rect 32445 -29729 32472 -29553
rect 32405 -29741 32472 -29729
rect 32303 -29779 32395 -29773
rect 32303 -29813 32315 -29779
rect 32383 -29813 32395 -29779
rect 32303 -29819 32395 -29813
rect 32328 -29820 32368 -29819
rect 32102 -29900 32160 -29862
rect 32428 -29900 32472 -29741
rect 32664 -29541 32708 -29212
rect 32768 -29152 32808 -29008
rect 32966 -29059 32972 -28683
rect 33006 -29059 33012 -28683
rect 33230 -28740 33474 -28734
rect 33230 -28774 33242 -28740
rect 33462 -28774 33474 -28740
rect 33100 -28822 33146 -28821
rect 32966 -29118 33012 -29059
rect 33078 -28833 33146 -28822
rect 33078 -28909 33106 -28833
rect 33140 -28909 33146 -28833
rect 33078 -28921 33146 -28909
rect 33078 -29152 33122 -28921
rect 33230 -28968 33474 -28774
rect 33558 -28833 33604 -28642
rect 33558 -28909 33564 -28833
rect 33598 -28909 33604 -28833
rect 33558 -28921 33604 -28909
rect 33984 -28909 34012 -28533
rect 34046 -28909 34052 -28533
rect 33984 -28920 34052 -28909
rect 34006 -28921 34052 -28920
rect 34088 -28962 34128 -28480
rect 34164 -28522 34210 -28521
rect 34164 -28528 34258 -28522
rect 34164 -28533 34194 -28528
rect 34164 -28909 34170 -28533
rect 34252 -28874 34258 -28528
rect 34304 -28524 34352 -28480
rect 34446 -28522 34492 -28521
rect 34400 -28524 34492 -28522
rect 34304 -28528 34492 -28524
rect 34304 -28570 34406 -28528
rect 34464 -28533 34492 -28528
rect 34164 -28914 34194 -28909
rect 34252 -28914 34352 -28874
rect 34164 -28920 34352 -28914
rect 34400 -28914 34406 -28570
rect 34486 -28909 34492 -28533
rect 34464 -28914 34492 -28909
rect 34400 -28920 34492 -28914
rect 34164 -28921 34210 -28920
rect 34304 -28962 34352 -28920
rect 34446 -28921 34492 -28920
rect 34528 -28962 34568 -28480
rect 34628 -28521 34672 -28360
rect 34956 -28440 35020 -28434
rect 34956 -28474 34968 -28440
rect 35008 -28474 35020 -28440
rect 34956 -28480 35020 -28474
rect 34604 -28533 34672 -28521
rect 34886 -28522 34932 -28521
rect 34604 -28909 34610 -28533
rect 34644 -28909 34672 -28533
rect 34604 -28920 34672 -28909
rect 34864 -28533 34932 -28522
rect 34864 -28909 34892 -28533
rect 34926 -28909 34932 -28533
rect 34604 -28921 34650 -28920
rect 34864 -28921 34932 -28909
rect 33230 -29002 33242 -28968
rect 33462 -29002 33474 -28968
rect 33230 -29008 33474 -29002
rect 34076 -28968 34140 -28962
rect 34076 -29002 34088 -28968
rect 34128 -29002 34140 -28968
rect 34076 -29008 34140 -29002
rect 34304 -28968 34580 -28962
rect 34304 -29002 34528 -28968
rect 34568 -29002 34580 -28968
rect 34304 -29008 34580 -29002
rect 32768 -29212 33148 -29152
rect 33366 -29200 33406 -29008
rect 34088 -29020 34128 -29008
rect 34528 -29020 34568 -29008
rect 34864 -29152 34908 -28921
rect 34968 -28962 35008 -28480
rect 35066 -28521 35110 -28360
rect 35044 -28533 35110 -28521
rect 35044 -28909 35050 -28533
rect 35084 -28909 35110 -28533
rect 35194 -28602 35910 -28360
rect 35194 -28608 35275 -28602
rect 35044 -28920 35110 -28909
rect 35166 -28636 35275 -28608
rect 35829 -28636 35910 -28602
rect 35166 -28642 35910 -28636
rect 36184 -28521 36228 -28360
rect 36276 -28440 36552 -28434
rect 36276 -28474 36288 -28440
rect 36328 -28474 36552 -28440
rect 36276 -28480 36552 -28474
rect 36716 -28440 36780 -28434
rect 36716 -28474 36728 -28440
rect 36768 -28474 36780 -28440
rect 36716 -28480 36780 -28474
rect 36184 -28533 36252 -28521
rect 35166 -28683 35212 -28642
rect 35044 -28921 35090 -28920
rect 34956 -28968 35020 -28962
rect 34956 -29002 34968 -28968
rect 35008 -29002 35020 -28968
rect 34956 -29008 35020 -29002
rect 32768 -29463 32808 -29212
rect 33104 -29270 33148 -29212
rect 32998 -29276 33148 -29270
rect 32998 -29334 33004 -29276
rect 33142 -29334 33148 -29276
rect 33350 -29210 33570 -29200
rect 33350 -29290 33360 -29210
rect 33560 -29290 33570 -29210
rect 33350 -29300 33570 -29290
rect 34088 -29212 34908 -29152
rect 32998 -29340 33148 -29334
rect 32986 -29420 33038 -29408
rect 32757 -29469 32821 -29463
rect 32757 -29503 32769 -29469
rect 32809 -29503 32821 -29469
rect 32757 -29509 32821 -29503
rect 32664 -29553 32733 -29541
rect 32664 -29729 32693 -29553
rect 32727 -29729 32733 -29553
rect 32664 -29741 32733 -29729
rect 32664 -29742 32708 -29741
rect 32768 -29773 32808 -29509
rect 32868 -29541 32912 -29538
rect 32845 -29553 32912 -29541
rect 32845 -29729 32851 -29553
rect 32885 -29729 32912 -29553
rect 32845 -29741 32912 -29729
rect 32757 -29779 32821 -29773
rect 32757 -29813 32769 -29779
rect 32809 -29813 32821 -29779
rect 32757 -29819 32821 -29813
rect 32768 -29820 32808 -29819
rect 32868 -29900 32912 -29741
rect 32986 -29862 32998 -29420
rect 33032 -29862 33038 -29420
rect 33104 -29540 33148 -29340
rect 33208 -29463 33248 -29446
rect 33366 -29463 33406 -29300
rect 33448 -29378 33594 -29376
rect 33448 -29430 33454 -29378
rect 33588 -29430 33594 -29378
rect 33448 -29432 33594 -29430
rect 33196 -29464 33260 -29463
rect 33354 -29464 33418 -29463
rect 33196 -29469 33418 -29464
rect 33196 -29503 33208 -29469
rect 33248 -29503 33366 -29469
rect 33406 -29503 33418 -29469
rect 33196 -29508 33418 -29503
rect 33196 -29509 33260 -29508
rect 33354 -29509 33418 -29508
rect 33072 -29546 33172 -29540
rect 33072 -29736 33078 -29546
rect 33166 -29736 33172 -29546
rect 33072 -29742 33172 -29736
rect 33208 -29773 33248 -29509
rect 33284 -29553 33330 -29541
rect 33284 -29729 33290 -29553
rect 33324 -29729 33330 -29553
rect 33284 -29741 33330 -29729
rect 33196 -29779 33260 -29773
rect 33196 -29813 33208 -29779
rect 33248 -29813 33260 -29779
rect 33196 -29819 33260 -29813
rect 32986 -29900 33038 -29862
rect 33288 -29900 33326 -29741
rect 33366 -29773 33406 -29509
rect 33448 -29541 33482 -29432
rect 33524 -29463 33564 -29462
rect 34088 -29463 34128 -29212
rect 34528 -29276 34678 -29270
rect 34528 -29334 34534 -29276
rect 34672 -29334 34678 -29276
rect 34528 -29340 34678 -29334
rect 34302 -29420 34360 -29408
rect 33512 -29469 33576 -29463
rect 33512 -29503 33524 -29469
rect 33564 -29503 33576 -29469
rect 33512 -29509 33576 -29503
rect 34063 -29469 34155 -29463
rect 34063 -29503 34075 -29469
rect 34143 -29503 34155 -29469
rect 34063 -29509 34155 -29503
rect 33442 -29553 33488 -29541
rect 33442 -29729 33448 -29553
rect 33482 -29729 33488 -29553
rect 33442 -29741 33488 -29729
rect 33524 -29773 33564 -29509
rect 33986 -29541 34030 -29538
rect 33600 -29542 33646 -29541
rect 33600 -29553 33658 -29542
rect 33600 -29729 33606 -29553
rect 33640 -29729 33658 -29553
rect 33600 -29741 33658 -29729
rect 33354 -29774 33418 -29773
rect 33512 -29774 33576 -29773
rect 33354 -29779 33576 -29774
rect 33354 -29813 33366 -29779
rect 33406 -29813 33524 -29779
rect 33564 -29813 33576 -29779
rect 33354 -29814 33576 -29813
rect 33354 -29819 33418 -29814
rect 33512 -29819 33576 -29814
rect 33612 -29900 33658 -29741
rect 33986 -29553 34053 -29541
rect 33986 -29729 34013 -29553
rect 34047 -29729 34053 -29553
rect 33986 -29741 34053 -29729
rect 33986 -29900 34030 -29741
rect 34088 -29773 34128 -29509
rect 34165 -29542 34211 -29541
rect 34165 -29548 34258 -29542
rect 34165 -29553 34194 -29548
rect 34165 -29729 34171 -29553
rect 34165 -29734 34194 -29729
rect 34252 -29734 34258 -29548
rect 34165 -29740 34258 -29734
rect 34165 -29741 34211 -29740
rect 34063 -29779 34155 -29773
rect 34063 -29813 34075 -29779
rect 34143 -29813 34155 -29779
rect 34063 -29819 34155 -29813
rect 34088 -29820 34128 -29819
rect 34302 -29862 34319 -29420
rect 34353 -29862 34360 -29420
rect 34528 -29463 34568 -29340
rect 34503 -29469 34595 -29463
rect 34503 -29503 34515 -29469
rect 34583 -29503 34595 -29469
rect 34503 -29509 34595 -29503
rect 34447 -29542 34493 -29541
rect 34426 -29544 34493 -29542
rect 34400 -29550 34493 -29544
rect 34400 -29736 34406 -29550
rect 34464 -29553 34493 -29550
rect 34487 -29729 34493 -29553
rect 34464 -29736 34493 -29729
rect 34400 -29741 34493 -29736
rect 34400 -29742 34470 -29741
rect 34528 -29773 34568 -29509
rect 34628 -29541 34672 -29538
rect 34605 -29553 34672 -29541
rect 34605 -29729 34611 -29553
rect 34645 -29729 34672 -29553
rect 34605 -29741 34672 -29729
rect 34503 -29779 34595 -29773
rect 34503 -29813 34515 -29779
rect 34583 -29813 34595 -29779
rect 34503 -29819 34595 -29813
rect 34528 -29820 34568 -29819
rect 34302 -29900 34360 -29862
rect 34628 -29900 34672 -29741
rect 34864 -29541 34908 -29212
rect 34968 -29152 35008 -29008
rect 35166 -29059 35172 -28683
rect 35206 -29059 35212 -28683
rect 35430 -28740 35674 -28734
rect 35430 -28774 35442 -28740
rect 35662 -28774 35674 -28740
rect 35300 -28822 35346 -28821
rect 35166 -29118 35212 -29059
rect 35278 -28833 35346 -28822
rect 35278 -28909 35306 -28833
rect 35340 -28909 35346 -28833
rect 35278 -28921 35346 -28909
rect 35278 -29152 35322 -28921
rect 35430 -28968 35674 -28774
rect 35758 -28833 35804 -28642
rect 35758 -28909 35764 -28833
rect 35798 -28909 35804 -28833
rect 35758 -28921 35804 -28909
rect 36184 -28909 36212 -28533
rect 36246 -28909 36252 -28533
rect 36184 -28920 36252 -28909
rect 36206 -28921 36252 -28920
rect 36288 -28962 36328 -28480
rect 36364 -28522 36410 -28521
rect 36364 -28528 36458 -28522
rect 36364 -28533 36394 -28528
rect 36364 -28909 36370 -28533
rect 36452 -28874 36458 -28528
rect 36504 -28524 36552 -28480
rect 36646 -28522 36692 -28521
rect 36600 -28524 36692 -28522
rect 36504 -28528 36692 -28524
rect 36504 -28570 36606 -28528
rect 36664 -28533 36692 -28528
rect 36364 -28914 36394 -28909
rect 36452 -28914 36552 -28874
rect 36364 -28920 36552 -28914
rect 36600 -28914 36606 -28570
rect 36686 -28909 36692 -28533
rect 36664 -28914 36692 -28909
rect 36600 -28920 36692 -28914
rect 36364 -28921 36410 -28920
rect 36504 -28962 36552 -28920
rect 36646 -28921 36692 -28920
rect 36728 -28962 36768 -28480
rect 36828 -28521 36872 -28360
rect 37156 -28440 37220 -28434
rect 37156 -28474 37168 -28440
rect 37208 -28474 37220 -28440
rect 37156 -28480 37220 -28474
rect 36804 -28533 36872 -28521
rect 37086 -28522 37132 -28521
rect 36804 -28909 36810 -28533
rect 36844 -28909 36872 -28533
rect 36804 -28920 36872 -28909
rect 37064 -28533 37132 -28522
rect 37064 -28909 37092 -28533
rect 37126 -28909 37132 -28533
rect 36804 -28921 36850 -28920
rect 37064 -28921 37132 -28909
rect 35430 -29002 35442 -28968
rect 35662 -29002 35674 -28968
rect 35430 -29008 35674 -29002
rect 36276 -28968 36340 -28962
rect 36276 -29002 36288 -28968
rect 36328 -29002 36340 -28968
rect 36276 -29008 36340 -29002
rect 36504 -28968 36780 -28962
rect 36504 -29002 36728 -28968
rect 36768 -29002 36780 -28968
rect 36504 -29008 36780 -29002
rect 34968 -29212 35348 -29152
rect 35566 -29200 35606 -29008
rect 36288 -29020 36328 -29008
rect 36728 -29020 36768 -29008
rect 37064 -29152 37108 -28921
rect 37168 -28962 37208 -28480
rect 37266 -28521 37310 -28360
rect 37244 -28533 37310 -28521
rect 37244 -28909 37250 -28533
rect 37284 -28909 37310 -28533
rect 37394 -28602 38110 -28360
rect 37394 -28608 37475 -28602
rect 37244 -28920 37310 -28909
rect 37366 -28636 37475 -28608
rect 38029 -28636 38110 -28602
rect 37366 -28642 38110 -28636
rect 37366 -28683 37412 -28642
rect 37244 -28921 37290 -28920
rect 37156 -28968 37220 -28962
rect 37156 -29002 37168 -28968
rect 37208 -29002 37220 -28968
rect 37156 -29008 37220 -29002
rect 34968 -29463 35008 -29212
rect 35304 -29270 35348 -29212
rect 35198 -29276 35348 -29270
rect 35198 -29334 35204 -29276
rect 35342 -29334 35348 -29276
rect 35550 -29210 35770 -29200
rect 35550 -29290 35560 -29210
rect 35760 -29290 35770 -29210
rect 35550 -29300 35770 -29290
rect 36288 -29212 37108 -29152
rect 35198 -29340 35348 -29334
rect 35186 -29420 35238 -29408
rect 34957 -29469 35021 -29463
rect 34957 -29503 34969 -29469
rect 35009 -29503 35021 -29469
rect 34957 -29509 35021 -29503
rect 34864 -29553 34933 -29541
rect 34864 -29729 34893 -29553
rect 34927 -29729 34933 -29553
rect 34864 -29741 34933 -29729
rect 34864 -29742 34908 -29741
rect 34968 -29773 35008 -29509
rect 35068 -29541 35112 -29538
rect 35045 -29553 35112 -29541
rect 35045 -29729 35051 -29553
rect 35085 -29729 35112 -29553
rect 35045 -29741 35112 -29729
rect 34957 -29779 35021 -29773
rect 34957 -29813 34969 -29779
rect 35009 -29813 35021 -29779
rect 34957 -29819 35021 -29813
rect 34968 -29820 35008 -29819
rect 35068 -29900 35112 -29741
rect 35186 -29862 35198 -29420
rect 35232 -29862 35238 -29420
rect 35304 -29540 35348 -29340
rect 35408 -29463 35448 -29446
rect 35566 -29463 35606 -29300
rect 35648 -29378 35794 -29376
rect 35648 -29430 35654 -29378
rect 35788 -29430 35794 -29378
rect 35648 -29432 35794 -29430
rect 35396 -29464 35460 -29463
rect 35554 -29464 35618 -29463
rect 35396 -29469 35618 -29464
rect 35396 -29503 35408 -29469
rect 35448 -29503 35566 -29469
rect 35606 -29503 35618 -29469
rect 35396 -29508 35618 -29503
rect 35396 -29509 35460 -29508
rect 35554 -29509 35618 -29508
rect 35272 -29546 35372 -29540
rect 35272 -29736 35278 -29546
rect 35366 -29736 35372 -29546
rect 35272 -29742 35372 -29736
rect 35408 -29773 35448 -29509
rect 35484 -29553 35530 -29541
rect 35484 -29729 35490 -29553
rect 35524 -29729 35530 -29553
rect 35484 -29741 35530 -29729
rect 35396 -29779 35460 -29773
rect 35396 -29813 35408 -29779
rect 35448 -29813 35460 -29779
rect 35396 -29819 35460 -29813
rect 35186 -29900 35238 -29862
rect 35488 -29900 35526 -29741
rect 35566 -29773 35606 -29509
rect 35648 -29541 35682 -29432
rect 35724 -29463 35764 -29462
rect 36288 -29463 36328 -29212
rect 36728 -29276 36878 -29270
rect 36728 -29334 36734 -29276
rect 36872 -29334 36878 -29276
rect 36728 -29340 36878 -29334
rect 36502 -29420 36560 -29408
rect 35712 -29469 35776 -29463
rect 35712 -29503 35724 -29469
rect 35764 -29503 35776 -29469
rect 35712 -29509 35776 -29503
rect 36263 -29469 36355 -29463
rect 36263 -29503 36275 -29469
rect 36343 -29503 36355 -29469
rect 36263 -29509 36355 -29503
rect 35642 -29553 35688 -29541
rect 35642 -29729 35648 -29553
rect 35682 -29729 35688 -29553
rect 35642 -29741 35688 -29729
rect 35724 -29773 35764 -29509
rect 36186 -29541 36230 -29538
rect 35800 -29542 35846 -29541
rect 35800 -29553 35858 -29542
rect 35800 -29729 35806 -29553
rect 35840 -29729 35858 -29553
rect 35800 -29741 35858 -29729
rect 35554 -29774 35618 -29773
rect 35712 -29774 35776 -29773
rect 35554 -29779 35776 -29774
rect 35554 -29813 35566 -29779
rect 35606 -29813 35724 -29779
rect 35764 -29813 35776 -29779
rect 35554 -29814 35776 -29813
rect 35554 -29819 35618 -29814
rect 35712 -29819 35776 -29814
rect 35812 -29900 35858 -29741
rect 36186 -29553 36253 -29541
rect 36186 -29729 36213 -29553
rect 36247 -29729 36253 -29553
rect 36186 -29741 36253 -29729
rect 36186 -29900 36230 -29741
rect 36288 -29773 36328 -29509
rect 36365 -29542 36411 -29541
rect 36365 -29548 36458 -29542
rect 36365 -29553 36394 -29548
rect 36365 -29729 36371 -29553
rect 36365 -29734 36394 -29729
rect 36452 -29734 36458 -29548
rect 36365 -29740 36458 -29734
rect 36365 -29741 36411 -29740
rect 36263 -29779 36355 -29773
rect 36263 -29813 36275 -29779
rect 36343 -29813 36355 -29779
rect 36263 -29819 36355 -29813
rect 36288 -29820 36328 -29819
rect 36502 -29862 36519 -29420
rect 36553 -29862 36560 -29420
rect 36728 -29463 36768 -29340
rect 36703 -29469 36795 -29463
rect 36703 -29503 36715 -29469
rect 36783 -29503 36795 -29469
rect 36703 -29509 36795 -29503
rect 36647 -29542 36693 -29541
rect 36626 -29544 36693 -29542
rect 36600 -29550 36693 -29544
rect 36600 -29736 36606 -29550
rect 36664 -29553 36693 -29550
rect 36687 -29729 36693 -29553
rect 36664 -29736 36693 -29729
rect 36600 -29741 36693 -29736
rect 36600 -29742 36670 -29741
rect 36728 -29773 36768 -29509
rect 36828 -29541 36872 -29538
rect 36805 -29553 36872 -29541
rect 36805 -29729 36811 -29553
rect 36845 -29729 36872 -29553
rect 36805 -29741 36872 -29729
rect 36703 -29779 36795 -29773
rect 36703 -29813 36715 -29779
rect 36783 -29813 36795 -29779
rect 36703 -29819 36795 -29813
rect 36728 -29820 36768 -29819
rect 36502 -29900 36560 -29862
rect 36828 -29900 36872 -29741
rect 37064 -29541 37108 -29212
rect 37168 -29152 37208 -29008
rect 37366 -29059 37372 -28683
rect 37406 -29059 37412 -28683
rect 37630 -28740 37874 -28734
rect 37630 -28774 37642 -28740
rect 37862 -28774 37874 -28740
rect 37500 -28822 37546 -28821
rect 37366 -29118 37412 -29059
rect 37478 -28833 37546 -28822
rect 37478 -28909 37506 -28833
rect 37540 -28909 37546 -28833
rect 37478 -28921 37546 -28909
rect 37478 -29152 37522 -28921
rect 37630 -28968 37874 -28774
rect 37958 -28833 38004 -28642
rect 37958 -28909 37964 -28833
rect 37998 -28909 38004 -28833
rect 37958 -28921 38004 -28909
rect 37630 -29002 37642 -28968
rect 37862 -29002 37874 -28968
rect 37630 -29008 37874 -29002
rect 37168 -29212 37548 -29152
rect 37766 -29200 37806 -29008
rect 37168 -29463 37208 -29212
rect 37504 -29270 37548 -29212
rect 37398 -29276 37548 -29270
rect 37398 -29334 37404 -29276
rect 37542 -29334 37548 -29276
rect 37750 -29210 37970 -29200
rect 37750 -29290 37760 -29210
rect 37960 -29290 37970 -29210
rect 37750 -29300 37970 -29290
rect 37398 -29340 37548 -29334
rect 37386 -29420 37438 -29408
rect 37157 -29469 37221 -29463
rect 37157 -29503 37169 -29469
rect 37209 -29503 37221 -29469
rect 37157 -29509 37221 -29503
rect 37064 -29553 37133 -29541
rect 37064 -29729 37093 -29553
rect 37127 -29729 37133 -29553
rect 37064 -29741 37133 -29729
rect 37064 -29742 37108 -29741
rect 37168 -29773 37208 -29509
rect 37268 -29541 37312 -29538
rect 37245 -29553 37312 -29541
rect 37245 -29729 37251 -29553
rect 37285 -29729 37312 -29553
rect 37245 -29741 37312 -29729
rect 37157 -29779 37221 -29773
rect 37157 -29813 37169 -29779
rect 37209 -29813 37221 -29779
rect 37157 -29819 37221 -29813
rect 37168 -29820 37208 -29819
rect 37268 -29900 37312 -29741
rect 37386 -29862 37398 -29420
rect 37432 -29862 37438 -29420
rect 37504 -29540 37548 -29340
rect 37608 -29463 37648 -29446
rect 37766 -29463 37806 -29300
rect 37848 -29378 37994 -29376
rect 37848 -29430 37854 -29378
rect 37988 -29430 37994 -29378
rect 37848 -29432 37994 -29430
rect 37596 -29464 37660 -29463
rect 37754 -29464 37818 -29463
rect 37596 -29469 37818 -29464
rect 37596 -29503 37608 -29469
rect 37648 -29503 37766 -29469
rect 37806 -29503 37818 -29469
rect 37596 -29508 37818 -29503
rect 37596 -29509 37660 -29508
rect 37754 -29509 37818 -29508
rect 37472 -29546 37572 -29540
rect 37472 -29736 37478 -29546
rect 37566 -29736 37572 -29546
rect 37472 -29742 37572 -29736
rect 37608 -29773 37648 -29509
rect 37684 -29553 37730 -29541
rect 37684 -29729 37690 -29553
rect 37724 -29729 37730 -29553
rect 37684 -29741 37730 -29729
rect 37596 -29779 37660 -29773
rect 37596 -29813 37608 -29779
rect 37648 -29813 37660 -29779
rect 37596 -29819 37660 -29813
rect 37386 -29900 37438 -29862
rect 37688 -29900 37726 -29741
rect 37766 -29773 37806 -29509
rect 37848 -29541 37882 -29432
rect 37924 -29463 37964 -29462
rect 37912 -29469 37976 -29463
rect 37912 -29503 37924 -29469
rect 37964 -29503 37976 -29469
rect 37912 -29509 37976 -29503
rect 37842 -29553 37888 -29541
rect 37842 -29729 37848 -29553
rect 37882 -29729 37888 -29553
rect 37842 -29741 37888 -29729
rect 37924 -29773 37964 -29509
rect 38000 -29542 38046 -29541
rect 38000 -29553 38058 -29542
rect 38000 -29729 38006 -29553
rect 38040 -29729 38058 -29553
rect 38000 -29741 38058 -29729
rect 37754 -29774 37818 -29773
rect 37912 -29774 37976 -29773
rect 37754 -29779 37976 -29774
rect 37754 -29813 37766 -29779
rect 37806 -29813 37924 -29779
rect 37964 -29813 37976 -29779
rect 37754 -29814 37976 -29813
rect 37754 -29819 37818 -29814
rect 37912 -29819 37976 -29814
rect 38012 -29900 38058 -29741
rect 29790 -29904 33756 -29900
rect 33830 -29904 35956 -29900
rect 36030 -29904 38156 -29900
rect 29790 -29917 38192 -29904
rect 27610 -29930 27690 -29920
rect 28767 -29929 28814 -29917
rect 27370 -29985 27450 -29975
rect 27370 -30012 27380 -29985
rect 27260 -30058 27380 -30012
rect 27370 -30075 27380 -30058
rect 27440 -30012 27450 -29985
rect 28767 -29983 28774 -29929
rect 28808 -29983 28814 -29929
rect 28767 -29990 28814 -29983
rect 29070 -29930 29150 -29920
rect 29070 -29990 29080 -29930
rect 28767 -29995 29080 -29990
rect 27440 -30018 28736 -30012
rect 27440 -30052 27948 -30018
rect 28724 -30052 28736 -30018
rect 27440 -30058 28736 -30052
rect 27440 -30075 27450 -30058
rect 28770 -30075 29080 -29995
rect 27370 -30085 27450 -30075
rect 28767 -30080 29080 -30075
rect 28767 -30087 28814 -30080
rect 27610 -30145 27690 -30135
rect 27610 -30170 27620 -30145
rect 27260 -30216 27620 -30170
rect 27610 -30235 27620 -30216
rect 27680 -30170 27690 -30145
rect 28767 -30141 28774 -30087
rect 28808 -30141 28814 -30087
rect 29070 -30130 29080 -30080
rect 29140 -30130 29150 -29930
rect 29070 -30140 29150 -30130
rect 29790 -29951 31713 -29917
rect 32105 -29951 32192 -29917
rect 32506 -29951 32593 -29917
rect 32985 -29951 33103 -29917
rect 33669 -29951 33913 -29917
rect 34305 -29951 34392 -29917
rect 34706 -29951 34793 -29917
rect 35185 -29951 35303 -29917
rect 35869 -29951 36113 -29917
rect 36505 -29951 36592 -29917
rect 36906 -29951 36993 -29917
rect 37385 -29920 37503 -29917
rect 38069 -29951 38192 -29917
rect 29790 -30073 37250 -29951
rect 37690 -30073 38192 -29951
rect 29790 -30107 31753 -30073
rect 32319 -30107 32437 -30073
rect 32829 -30107 32916 -30073
rect 33230 -30107 33317 -30073
rect 33709 -30107 33953 -30073
rect 34519 -30107 34637 -30073
rect 35029 -30107 35116 -30073
rect 35430 -30107 35517 -30073
rect 35909 -30107 36153 -30073
rect 36719 -30107 36837 -30073
rect 37229 -30107 37250 -30073
rect 37690 -30107 37717 -30073
rect 38109 -30107 38192 -30073
rect 29790 -30110 37250 -30107
rect 37690 -30110 38192 -30107
rect 29790 -30120 38192 -30110
rect 28767 -30153 28814 -30141
rect 27680 -30176 28736 -30170
rect 27680 -30210 27948 -30176
rect 28724 -30210 28736 -30176
rect 27680 -30216 28736 -30210
rect 27680 -30235 27690 -30216
rect 28770 -30233 28810 -30153
rect 27610 -30245 27690 -30235
rect 28767 -30245 28814 -30233
rect 27370 -30300 27450 -30290
rect 27370 -30328 27380 -30300
rect 27260 -30374 27380 -30328
rect 27370 -30390 27380 -30374
rect 27440 -30328 27450 -30300
rect 28767 -30299 28774 -30245
rect 28808 -30299 28814 -30245
rect 28767 -30311 28814 -30299
rect 27440 -30334 28736 -30328
rect 27440 -30368 27948 -30334
rect 28724 -30368 28736 -30334
rect 27440 -30374 28736 -30368
rect 27440 -30390 27450 -30374
rect 27370 -30400 27450 -30390
rect 27910 -30468 28815 -30462
rect 27910 -30502 27931 -30468
rect 28803 -30480 28815 -30468
rect 29790 -30480 29990 -30120
rect 31608 -30124 38192 -30120
rect 28803 -30502 29990 -30480
rect 31764 -30283 31810 -30124
rect 31846 -30210 31910 -30205
rect 32004 -30210 32068 -30205
rect 31846 -30211 32068 -30210
rect 31846 -30245 31858 -30211
rect 31898 -30245 32016 -30211
rect 32056 -30245 32068 -30211
rect 31846 -30250 32068 -30245
rect 31846 -30251 31910 -30250
rect 32004 -30251 32068 -30250
rect 31764 -30295 31822 -30283
rect 31764 -30471 31782 -30295
rect 31816 -30471 31822 -30295
rect 31764 -30482 31822 -30471
rect 31776 -30483 31822 -30482
rect 27910 -30508 29990 -30502
rect 27930 -30602 29990 -30508
rect 31858 -30515 31898 -30251
rect 31934 -30295 31980 -30283
rect 31934 -30471 31940 -30295
rect 31974 -30471 31980 -30295
rect 31934 -30483 31980 -30471
rect 31846 -30521 31910 -30515
rect 31846 -30555 31858 -30521
rect 31898 -30555 31910 -30521
rect 31846 -30561 31910 -30555
rect 31858 -30562 31898 -30561
rect 31940 -30592 31974 -30483
rect 32016 -30515 32056 -30251
rect 32096 -30283 32134 -30124
rect 32384 -30162 32436 -30124
rect 32162 -30211 32226 -30205
rect 32162 -30245 32174 -30211
rect 32214 -30245 32226 -30211
rect 32162 -30251 32226 -30245
rect 32092 -30295 32138 -30283
rect 32092 -30471 32098 -30295
rect 32132 -30471 32138 -30295
rect 32092 -30483 32138 -30471
rect 32174 -30515 32214 -30251
rect 32250 -30288 32350 -30282
rect 32250 -30478 32256 -30288
rect 32344 -30478 32350 -30288
rect 32250 -30484 32350 -30478
rect 32004 -30516 32068 -30515
rect 32162 -30516 32226 -30515
rect 32004 -30521 32226 -30516
rect 32004 -30555 32016 -30521
rect 32056 -30555 32174 -30521
rect 32214 -30555 32226 -30521
rect 32004 -30560 32226 -30555
rect 32004 -30561 32068 -30560
rect 32162 -30561 32226 -30560
rect 27910 -30608 29990 -30602
rect 27910 -30642 27931 -30608
rect 28803 -30610 29990 -30608
rect 28803 -30642 28815 -30610
rect 27910 -30648 28815 -30642
rect 27370 -30710 27450 -30700
rect 27370 -30736 27380 -30710
rect 27260 -30782 27380 -30736
rect 27370 -30800 27380 -30782
rect 27440 -30736 27450 -30710
rect 27440 -30742 28736 -30736
rect 27440 -30776 27948 -30742
rect 28724 -30776 28736 -30742
rect 27440 -30782 28736 -30776
rect 27440 -30800 27450 -30782
rect 27370 -30810 27450 -30800
rect 28767 -30811 28814 -30799
rect 27490 -30870 27570 -30860
rect 27490 -30894 27500 -30870
rect 27260 -30940 27500 -30894
rect 27490 -30960 27500 -30940
rect 27560 -30894 27570 -30870
rect 28767 -30865 28774 -30811
rect 28808 -30865 28814 -30811
rect 28767 -30877 28814 -30865
rect 27560 -30900 28736 -30894
rect 27560 -30934 27948 -30900
rect 28724 -30934 28736 -30900
rect 27560 -30940 28736 -30934
rect 27560 -30960 27570 -30940
rect 28770 -30957 28810 -30877
rect 27490 -30970 27570 -30960
rect 28767 -30960 28814 -30957
rect 29060 -30960 29300 -30950
rect 28767 -30969 29070 -30960
rect 27370 -31025 27450 -31015
rect 27370 -31052 27380 -31025
rect 27260 -31098 27380 -31052
rect 27370 -31115 27380 -31098
rect 27440 -31052 27450 -31025
rect 28767 -31023 28774 -30969
rect 28808 -31023 29070 -30969
rect 28767 -31030 29070 -31023
rect 29290 -31030 29300 -30960
rect 28767 -31035 28814 -31030
rect 27440 -31058 28736 -31052
rect 27440 -31092 27948 -31058
rect 28724 -31092 28736 -31058
rect 27440 -31098 28736 -31092
rect 27440 -31115 27450 -31098
rect 28770 -31115 28810 -31035
rect 29060 -31040 29300 -31030
rect 27370 -31125 27450 -31115
rect 28767 -31127 28814 -31115
rect 27490 -31185 27570 -31175
rect 27490 -31210 27500 -31185
rect 27260 -31256 27500 -31210
rect 27490 -31275 27500 -31256
rect 27560 -31210 27570 -31185
rect 28767 -31181 28774 -31127
rect 28808 -31181 28814 -31127
rect 28767 -31193 28814 -31181
rect 27560 -31216 28736 -31210
rect 27560 -31250 27948 -31216
rect 28724 -31250 28736 -31216
rect 27560 -31256 28736 -31250
rect 27560 -31275 27570 -31256
rect 28770 -31273 28810 -31193
rect 27490 -31285 27570 -31275
rect 28767 -31285 28814 -31273
rect 27370 -31340 27450 -31330
rect 27370 -31368 27380 -31340
rect 27260 -31414 27380 -31368
rect 27370 -31430 27380 -31414
rect 27440 -31368 27450 -31340
rect 28767 -31339 28774 -31285
rect 28808 -31339 28814 -31285
rect 28767 -31351 28814 -31339
rect 27440 -31374 28736 -31368
rect 27440 -31408 27948 -31374
rect 28724 -31408 28736 -31374
rect 27440 -31414 28736 -31408
rect 27440 -31430 27450 -31414
rect 27370 -31440 27450 -31430
rect 27910 -31508 28815 -31502
rect 27910 -31542 27931 -31508
rect 28803 -31520 28815 -31508
rect 29790 -31520 29990 -30610
rect 31828 -30594 31974 -30592
rect 31828 -30646 31834 -30594
rect 31968 -30646 31974 -30594
rect 31828 -30648 31974 -30646
rect 32016 -30720 32056 -30561
rect 32174 -30578 32214 -30561
rect 32274 -30684 32318 -30484
rect 32384 -30604 32390 -30162
rect 32424 -30604 32436 -30162
rect 32510 -30283 32554 -30124
rect 32614 -30205 32654 -30204
rect 32601 -30211 32665 -30205
rect 32601 -30245 32613 -30211
rect 32653 -30245 32665 -30211
rect 32601 -30251 32665 -30245
rect 32510 -30295 32577 -30283
rect 32510 -30471 32537 -30295
rect 32571 -30471 32577 -30295
rect 32510 -30483 32577 -30471
rect 32510 -30486 32554 -30483
rect 32614 -30515 32654 -30251
rect 32714 -30283 32758 -30282
rect 32689 -30295 32758 -30283
rect 32689 -30471 32695 -30295
rect 32729 -30471 32758 -30295
rect 32689 -30483 32758 -30471
rect 32601 -30521 32665 -30515
rect 32601 -30555 32613 -30521
rect 32653 -30555 32665 -30521
rect 32601 -30561 32665 -30555
rect 32384 -30616 32436 -30604
rect 32274 -30690 32424 -30684
rect 31840 -30730 32060 -30720
rect 31840 -30810 31850 -30730
rect 32050 -30810 32060 -30730
rect 31840 -30820 32060 -30810
rect 32274 -30748 32280 -30690
rect 32418 -30748 32424 -30690
rect 32274 -30754 32424 -30748
rect 32274 -30812 32318 -30754
rect 32614 -30812 32654 -30561
rect 32016 -31016 32056 -30820
rect 32274 -30872 32654 -30812
rect 31948 -31022 32192 -31016
rect 31948 -31056 31960 -31022
rect 32180 -31056 32192 -31022
rect 31818 -31115 31864 -31103
rect 31818 -31191 31824 -31115
rect 31858 -31191 31864 -31115
rect 31818 -31382 31864 -31191
rect 31948 -31250 32192 -31056
rect 32300 -31103 32344 -30872
rect 32276 -31115 32344 -31103
rect 32276 -31191 32282 -31115
rect 32316 -31191 32344 -31115
rect 32276 -31202 32344 -31191
rect 32410 -30965 32456 -30906
rect 32276 -31203 32322 -31202
rect 31948 -31284 31960 -31250
rect 32180 -31284 32192 -31250
rect 31948 -31290 32192 -31284
rect 32410 -31341 32416 -30965
rect 32450 -31341 32456 -30965
rect 32614 -31016 32654 -30872
rect 32714 -30812 32758 -30483
rect 32950 -30283 32994 -30124
rect 33262 -30162 33320 -30124
rect 33054 -30205 33094 -30204
rect 33027 -30211 33119 -30205
rect 33027 -30245 33039 -30211
rect 33107 -30245 33119 -30211
rect 33027 -30251 33119 -30245
rect 32950 -30295 33017 -30283
rect 32950 -30471 32977 -30295
rect 33011 -30471 33017 -30295
rect 32950 -30483 33017 -30471
rect 32950 -30486 32994 -30483
rect 33054 -30515 33094 -30251
rect 33152 -30283 33222 -30282
rect 33129 -30288 33222 -30283
rect 33129 -30295 33158 -30288
rect 33129 -30471 33135 -30295
rect 33129 -30474 33158 -30471
rect 33216 -30474 33222 -30288
rect 33129 -30480 33222 -30474
rect 33129 -30482 33196 -30480
rect 33129 -30483 33175 -30482
rect 33027 -30521 33119 -30515
rect 33027 -30555 33039 -30521
rect 33107 -30555 33119 -30521
rect 33027 -30561 33119 -30555
rect 33054 -30684 33094 -30561
rect 33262 -30604 33269 -30162
rect 33303 -30604 33320 -30162
rect 33494 -30205 33534 -30204
rect 33467 -30211 33559 -30205
rect 33467 -30245 33479 -30211
rect 33547 -30245 33559 -30211
rect 33467 -30251 33559 -30245
rect 33411 -30284 33457 -30283
rect 33364 -30290 33457 -30284
rect 33364 -30476 33370 -30290
rect 33428 -30295 33457 -30290
rect 33451 -30471 33457 -30295
rect 33428 -30476 33457 -30471
rect 33364 -30482 33457 -30476
rect 33411 -30483 33457 -30482
rect 33494 -30515 33534 -30251
rect 33592 -30283 33636 -30124
rect 33569 -30295 33636 -30283
rect 33569 -30471 33575 -30295
rect 33609 -30471 33636 -30295
rect 33569 -30483 33636 -30471
rect 33964 -30283 34010 -30124
rect 34046 -30210 34110 -30205
rect 34204 -30210 34268 -30205
rect 34046 -30211 34268 -30210
rect 34046 -30245 34058 -30211
rect 34098 -30245 34216 -30211
rect 34256 -30245 34268 -30211
rect 34046 -30250 34268 -30245
rect 34046 -30251 34110 -30250
rect 34204 -30251 34268 -30250
rect 33964 -30295 34022 -30283
rect 33964 -30471 33982 -30295
rect 34016 -30471 34022 -30295
rect 33964 -30482 34022 -30471
rect 33976 -30483 34022 -30482
rect 33592 -30486 33636 -30483
rect 34058 -30515 34098 -30251
rect 34134 -30295 34180 -30283
rect 34134 -30471 34140 -30295
rect 34174 -30471 34180 -30295
rect 34134 -30483 34180 -30471
rect 33467 -30521 33559 -30515
rect 33467 -30555 33479 -30521
rect 33547 -30555 33559 -30521
rect 33467 -30561 33559 -30555
rect 34046 -30521 34110 -30515
rect 34046 -30555 34058 -30521
rect 34098 -30555 34110 -30521
rect 34046 -30561 34110 -30555
rect 33262 -30616 33320 -30604
rect 32944 -30690 33094 -30684
rect 32944 -30748 32950 -30690
rect 33088 -30748 33094 -30690
rect 32944 -30754 33094 -30748
rect 33494 -30812 33534 -30561
rect 34058 -30562 34098 -30561
rect 34140 -30592 34174 -30483
rect 34216 -30515 34256 -30251
rect 34296 -30283 34334 -30124
rect 34584 -30162 34636 -30124
rect 34362 -30211 34426 -30205
rect 34362 -30245 34374 -30211
rect 34414 -30245 34426 -30211
rect 34362 -30251 34426 -30245
rect 34292 -30295 34338 -30283
rect 34292 -30471 34298 -30295
rect 34332 -30471 34338 -30295
rect 34292 -30483 34338 -30471
rect 34374 -30515 34414 -30251
rect 34450 -30288 34550 -30282
rect 34450 -30478 34456 -30288
rect 34544 -30478 34550 -30288
rect 34450 -30484 34550 -30478
rect 34204 -30516 34268 -30515
rect 34362 -30516 34426 -30515
rect 34204 -30521 34426 -30516
rect 34204 -30555 34216 -30521
rect 34256 -30555 34374 -30521
rect 34414 -30555 34426 -30521
rect 34204 -30560 34426 -30555
rect 34204 -30561 34268 -30560
rect 34362 -30561 34426 -30560
rect 34028 -30594 34174 -30592
rect 34028 -30646 34034 -30594
rect 34168 -30646 34174 -30594
rect 34028 -30648 34174 -30646
rect 34216 -30720 34256 -30561
rect 34374 -30578 34414 -30561
rect 34474 -30684 34518 -30484
rect 34584 -30604 34590 -30162
rect 34624 -30604 34636 -30162
rect 34710 -30283 34754 -30124
rect 34814 -30205 34854 -30204
rect 34801 -30211 34865 -30205
rect 34801 -30245 34813 -30211
rect 34853 -30245 34865 -30211
rect 34801 -30251 34865 -30245
rect 34710 -30295 34777 -30283
rect 34710 -30471 34737 -30295
rect 34771 -30471 34777 -30295
rect 34710 -30483 34777 -30471
rect 34710 -30486 34754 -30483
rect 34814 -30515 34854 -30251
rect 34914 -30283 34958 -30282
rect 34889 -30295 34958 -30283
rect 34889 -30471 34895 -30295
rect 34929 -30471 34958 -30295
rect 34889 -30483 34958 -30471
rect 34801 -30521 34865 -30515
rect 34801 -30555 34813 -30521
rect 34853 -30555 34865 -30521
rect 34801 -30561 34865 -30555
rect 34584 -30616 34636 -30604
rect 34474 -30690 34624 -30684
rect 32714 -30872 33534 -30812
rect 34050 -30730 34270 -30720
rect 34050 -30810 34060 -30730
rect 34260 -30810 34270 -30730
rect 34050 -30820 34270 -30810
rect 34474 -30748 34480 -30690
rect 34618 -30748 34624 -30690
rect 34474 -30754 34624 -30748
rect 34474 -30812 34518 -30754
rect 34814 -30812 34854 -30561
rect 32602 -31022 32666 -31016
rect 32602 -31056 32614 -31022
rect 32654 -31056 32666 -31022
rect 32602 -31062 32666 -31056
rect 32532 -31104 32578 -31103
rect 32410 -31382 32456 -31341
rect 28803 -31542 29990 -31520
rect 27910 -31548 29990 -31542
rect 27940 -31650 29990 -31548
rect 27024 -31668 27070 -31656
rect 26347 -31901 26909 -31895
rect 29790 -31940 29990 -31650
rect 31712 -31388 32456 -31382
rect 31712 -31422 31793 -31388
rect 32347 -31416 32456 -31388
rect 32512 -31115 32578 -31104
rect 32347 -31422 32428 -31416
rect 31712 -31664 32428 -31422
rect 32512 -31491 32538 -31115
rect 32572 -31491 32578 -31115
rect 32512 -31503 32578 -31491
rect 32512 -31664 32556 -31503
rect 32614 -31544 32654 -31062
rect 32714 -31103 32758 -30872
rect 33054 -31016 33094 -31004
rect 33494 -31016 33534 -31004
rect 34216 -31016 34256 -30820
rect 34474 -30872 34854 -30812
rect 33042 -31022 33318 -31016
rect 33042 -31056 33054 -31022
rect 33094 -31056 33318 -31022
rect 33042 -31062 33318 -31056
rect 33482 -31022 33546 -31016
rect 33482 -31056 33494 -31022
rect 33534 -31056 33546 -31022
rect 33482 -31062 33546 -31056
rect 34148 -31022 34392 -31016
rect 34148 -31056 34160 -31022
rect 34380 -31056 34392 -31022
rect 32690 -31115 32758 -31103
rect 32972 -31104 33018 -31103
rect 32690 -31491 32696 -31115
rect 32730 -31491 32758 -31115
rect 32690 -31502 32758 -31491
rect 32950 -31115 33018 -31104
rect 32950 -31491 32978 -31115
rect 33012 -31491 33018 -31115
rect 32690 -31503 32736 -31502
rect 32950 -31503 33018 -31491
rect 32602 -31550 32666 -31544
rect 32602 -31584 32614 -31550
rect 32654 -31584 32666 -31550
rect 32602 -31590 32666 -31584
rect 32950 -31664 32994 -31503
rect 33054 -31544 33094 -31062
rect 33130 -31104 33176 -31103
rect 33270 -31104 33318 -31062
rect 33412 -31104 33458 -31103
rect 33130 -31110 33222 -31104
rect 33130 -31115 33158 -31110
rect 33130 -31491 33136 -31115
rect 33216 -31454 33222 -31110
rect 33270 -31110 33458 -31104
rect 33270 -31150 33370 -31110
rect 33428 -31115 33458 -31110
rect 33130 -31496 33158 -31491
rect 33216 -31496 33318 -31454
rect 33130 -31500 33318 -31496
rect 33130 -31502 33222 -31500
rect 33130 -31503 33176 -31502
rect 33270 -31544 33318 -31500
rect 33364 -31496 33370 -31150
rect 33452 -31491 33458 -31115
rect 33428 -31496 33458 -31491
rect 33364 -31502 33458 -31496
rect 33412 -31503 33458 -31502
rect 33494 -31544 33534 -31062
rect 33570 -31104 33616 -31103
rect 33570 -31115 33638 -31104
rect 33570 -31491 33576 -31115
rect 33610 -31491 33638 -31115
rect 34018 -31115 34064 -31103
rect 34018 -31191 34024 -31115
rect 34058 -31191 34064 -31115
rect 34018 -31382 34064 -31191
rect 34148 -31250 34392 -31056
rect 34500 -31103 34544 -30872
rect 34476 -31115 34544 -31103
rect 34476 -31191 34482 -31115
rect 34516 -31191 34544 -31115
rect 34476 -31202 34544 -31191
rect 34610 -30965 34656 -30906
rect 34476 -31203 34522 -31202
rect 34148 -31284 34160 -31250
rect 34380 -31284 34392 -31250
rect 34148 -31290 34392 -31284
rect 34610 -31341 34616 -30965
rect 34650 -31341 34656 -30965
rect 34814 -31016 34854 -30872
rect 34914 -30812 34958 -30483
rect 35150 -30283 35194 -30124
rect 35462 -30162 35520 -30124
rect 35254 -30205 35294 -30204
rect 35227 -30211 35319 -30205
rect 35227 -30245 35239 -30211
rect 35307 -30245 35319 -30211
rect 35227 -30251 35319 -30245
rect 35150 -30295 35217 -30283
rect 35150 -30471 35177 -30295
rect 35211 -30471 35217 -30295
rect 35150 -30483 35217 -30471
rect 35150 -30486 35194 -30483
rect 35254 -30515 35294 -30251
rect 35352 -30283 35422 -30282
rect 35329 -30288 35422 -30283
rect 35329 -30295 35358 -30288
rect 35329 -30471 35335 -30295
rect 35329 -30474 35358 -30471
rect 35416 -30474 35422 -30288
rect 35329 -30480 35422 -30474
rect 35329 -30482 35396 -30480
rect 35329 -30483 35375 -30482
rect 35227 -30521 35319 -30515
rect 35227 -30555 35239 -30521
rect 35307 -30555 35319 -30521
rect 35227 -30561 35319 -30555
rect 35254 -30684 35294 -30561
rect 35462 -30604 35469 -30162
rect 35503 -30604 35520 -30162
rect 35694 -30205 35734 -30204
rect 35667 -30211 35759 -30205
rect 35667 -30245 35679 -30211
rect 35747 -30245 35759 -30211
rect 35667 -30251 35759 -30245
rect 35611 -30284 35657 -30283
rect 35564 -30290 35657 -30284
rect 35564 -30476 35570 -30290
rect 35628 -30295 35657 -30290
rect 35651 -30471 35657 -30295
rect 35628 -30476 35657 -30471
rect 35564 -30482 35657 -30476
rect 35611 -30483 35657 -30482
rect 35694 -30515 35734 -30251
rect 35792 -30283 35836 -30124
rect 35769 -30295 35836 -30283
rect 35769 -30471 35775 -30295
rect 35809 -30471 35836 -30295
rect 35769 -30483 35836 -30471
rect 36164 -30283 36210 -30124
rect 36246 -30210 36310 -30205
rect 36404 -30210 36468 -30205
rect 36246 -30211 36468 -30210
rect 36246 -30245 36258 -30211
rect 36298 -30245 36416 -30211
rect 36456 -30245 36468 -30211
rect 36246 -30250 36468 -30245
rect 36246 -30251 36310 -30250
rect 36404 -30251 36468 -30250
rect 36164 -30295 36222 -30283
rect 36164 -30471 36182 -30295
rect 36216 -30471 36222 -30295
rect 36164 -30482 36222 -30471
rect 36176 -30483 36222 -30482
rect 35792 -30486 35836 -30483
rect 36258 -30515 36298 -30251
rect 36334 -30295 36380 -30283
rect 36334 -30471 36340 -30295
rect 36374 -30471 36380 -30295
rect 36334 -30483 36380 -30471
rect 35667 -30521 35759 -30515
rect 35667 -30555 35679 -30521
rect 35747 -30555 35759 -30521
rect 35667 -30561 35759 -30555
rect 36246 -30521 36310 -30515
rect 36246 -30555 36258 -30521
rect 36298 -30555 36310 -30521
rect 36246 -30561 36310 -30555
rect 35462 -30616 35520 -30604
rect 35144 -30690 35294 -30684
rect 35144 -30748 35150 -30690
rect 35288 -30748 35294 -30690
rect 35144 -30754 35294 -30748
rect 35694 -30812 35734 -30561
rect 36258 -30562 36298 -30561
rect 36340 -30592 36374 -30483
rect 36416 -30515 36456 -30251
rect 36496 -30283 36534 -30124
rect 36784 -30162 36836 -30124
rect 36562 -30211 36626 -30205
rect 36562 -30245 36574 -30211
rect 36614 -30245 36626 -30211
rect 36562 -30251 36626 -30245
rect 36492 -30295 36538 -30283
rect 36492 -30471 36498 -30295
rect 36532 -30471 36538 -30295
rect 36492 -30483 36538 -30471
rect 36574 -30515 36614 -30251
rect 36650 -30288 36750 -30282
rect 36650 -30478 36656 -30288
rect 36744 -30478 36750 -30288
rect 36650 -30484 36750 -30478
rect 36404 -30516 36468 -30515
rect 36562 -30516 36626 -30515
rect 36404 -30521 36626 -30516
rect 36404 -30555 36416 -30521
rect 36456 -30555 36574 -30521
rect 36614 -30555 36626 -30521
rect 36404 -30560 36626 -30555
rect 36404 -30561 36468 -30560
rect 36562 -30561 36626 -30560
rect 36228 -30594 36374 -30592
rect 36228 -30646 36234 -30594
rect 36368 -30646 36374 -30594
rect 36228 -30648 36374 -30646
rect 36416 -30730 36456 -30561
rect 36574 -30578 36614 -30561
rect 36674 -30684 36718 -30484
rect 36784 -30604 36790 -30162
rect 36824 -30604 36836 -30162
rect 36910 -30283 36954 -30124
rect 37014 -30205 37054 -30204
rect 37001 -30211 37065 -30205
rect 37001 -30245 37013 -30211
rect 37053 -30245 37065 -30211
rect 37001 -30251 37065 -30245
rect 36910 -30295 36977 -30283
rect 36910 -30471 36937 -30295
rect 36971 -30471 36977 -30295
rect 36910 -30483 36977 -30471
rect 36910 -30486 36954 -30483
rect 37014 -30515 37054 -30251
rect 37114 -30283 37158 -30282
rect 37089 -30295 37158 -30283
rect 37089 -30471 37095 -30295
rect 37129 -30471 37158 -30295
rect 37089 -30483 37158 -30471
rect 37001 -30521 37065 -30515
rect 37001 -30555 37013 -30521
rect 37053 -30555 37065 -30521
rect 37001 -30561 37065 -30555
rect 36784 -30616 36836 -30604
rect 36674 -30690 36824 -30684
rect 34914 -30872 35734 -30812
rect 36250 -30740 36470 -30730
rect 36250 -30820 36260 -30740
rect 36460 -30820 36470 -30740
rect 36250 -30830 36470 -30820
rect 36674 -30748 36680 -30690
rect 36818 -30748 36824 -30690
rect 36674 -30754 36824 -30748
rect 36674 -30812 36718 -30754
rect 37014 -30812 37054 -30561
rect 34802 -31022 34866 -31016
rect 34802 -31056 34814 -31022
rect 34854 -31056 34866 -31022
rect 34802 -31062 34866 -31056
rect 34732 -31104 34778 -31103
rect 34610 -31382 34656 -31341
rect 33570 -31503 33638 -31491
rect 33042 -31550 33106 -31544
rect 33042 -31584 33054 -31550
rect 33094 -31584 33106 -31550
rect 33042 -31590 33106 -31584
rect 33270 -31550 33546 -31544
rect 33270 -31584 33494 -31550
rect 33534 -31584 33546 -31550
rect 33270 -31590 33546 -31584
rect 33594 -31664 33638 -31503
rect 33912 -31388 34656 -31382
rect 33912 -31422 33993 -31388
rect 34547 -31416 34656 -31388
rect 34712 -31115 34778 -31104
rect 34547 -31422 34628 -31416
rect 33912 -31664 34628 -31422
rect 34712 -31491 34738 -31115
rect 34772 -31491 34778 -31115
rect 34712 -31503 34778 -31491
rect 34712 -31664 34756 -31503
rect 34814 -31544 34854 -31062
rect 34914 -31103 34958 -30872
rect 35254 -31016 35294 -31004
rect 35694 -31016 35734 -31004
rect 36416 -31016 36456 -30830
rect 36674 -30872 37054 -30812
rect 35242 -31022 35518 -31016
rect 35242 -31056 35254 -31022
rect 35294 -31056 35518 -31022
rect 35242 -31062 35518 -31056
rect 35682 -31022 35746 -31016
rect 35682 -31056 35694 -31022
rect 35734 -31056 35746 -31022
rect 35682 -31062 35746 -31056
rect 36348 -31022 36592 -31016
rect 36348 -31056 36360 -31022
rect 36580 -31056 36592 -31022
rect 34890 -31115 34958 -31103
rect 35172 -31104 35218 -31103
rect 34890 -31491 34896 -31115
rect 34930 -31491 34958 -31115
rect 34890 -31502 34958 -31491
rect 35150 -31115 35218 -31104
rect 35150 -31491 35178 -31115
rect 35212 -31491 35218 -31115
rect 34890 -31503 34936 -31502
rect 35150 -31503 35218 -31491
rect 34802 -31550 34866 -31544
rect 34802 -31584 34814 -31550
rect 34854 -31584 34866 -31550
rect 34802 -31590 34866 -31584
rect 35150 -31664 35194 -31503
rect 35254 -31544 35294 -31062
rect 35330 -31104 35376 -31103
rect 35470 -31104 35518 -31062
rect 35612 -31104 35658 -31103
rect 35330 -31110 35422 -31104
rect 35330 -31115 35358 -31110
rect 35330 -31491 35336 -31115
rect 35416 -31454 35422 -31110
rect 35470 -31110 35658 -31104
rect 35470 -31150 35570 -31110
rect 35628 -31115 35658 -31110
rect 35330 -31496 35358 -31491
rect 35416 -31496 35518 -31454
rect 35330 -31500 35518 -31496
rect 35330 -31502 35422 -31500
rect 35330 -31503 35376 -31502
rect 35470 -31544 35518 -31500
rect 35564 -31496 35570 -31150
rect 35652 -31491 35658 -31115
rect 35628 -31496 35658 -31491
rect 35564 -31502 35658 -31496
rect 35612 -31503 35658 -31502
rect 35694 -31544 35734 -31062
rect 35770 -31104 35816 -31103
rect 35770 -31115 35838 -31104
rect 35770 -31491 35776 -31115
rect 35810 -31491 35838 -31115
rect 36218 -31115 36264 -31103
rect 36218 -31191 36224 -31115
rect 36258 -31191 36264 -31115
rect 36218 -31382 36264 -31191
rect 36348 -31250 36592 -31056
rect 36700 -31103 36744 -30872
rect 36676 -31115 36744 -31103
rect 36676 -31191 36682 -31115
rect 36716 -31191 36744 -31115
rect 36676 -31202 36744 -31191
rect 36810 -30965 36856 -30906
rect 36676 -31203 36722 -31202
rect 36348 -31284 36360 -31250
rect 36580 -31284 36592 -31250
rect 36348 -31290 36592 -31284
rect 36810 -31341 36816 -30965
rect 36850 -31341 36856 -30965
rect 37014 -31016 37054 -30872
rect 37114 -30812 37158 -30483
rect 37350 -30283 37394 -30124
rect 37662 -30162 37720 -30124
rect 37454 -30205 37494 -30204
rect 37427 -30211 37519 -30205
rect 37427 -30245 37439 -30211
rect 37507 -30245 37519 -30211
rect 37427 -30251 37519 -30245
rect 37350 -30295 37417 -30283
rect 37350 -30471 37377 -30295
rect 37411 -30471 37417 -30295
rect 37350 -30483 37417 -30471
rect 37350 -30486 37394 -30483
rect 37454 -30515 37494 -30251
rect 37552 -30283 37622 -30282
rect 37529 -30288 37622 -30283
rect 37529 -30295 37558 -30288
rect 37529 -30471 37535 -30295
rect 37529 -30474 37558 -30471
rect 37616 -30474 37622 -30288
rect 37529 -30480 37622 -30474
rect 37529 -30482 37596 -30480
rect 37529 -30483 37575 -30482
rect 37427 -30521 37519 -30515
rect 37427 -30555 37439 -30521
rect 37507 -30555 37519 -30521
rect 37427 -30561 37519 -30555
rect 37454 -30684 37494 -30561
rect 37662 -30604 37669 -30162
rect 37703 -30604 37720 -30162
rect 37894 -30205 37934 -30204
rect 37867 -30211 37959 -30205
rect 37867 -30245 37879 -30211
rect 37947 -30245 37959 -30211
rect 37867 -30251 37959 -30245
rect 37811 -30284 37857 -30283
rect 37764 -30290 37857 -30284
rect 37764 -30476 37770 -30290
rect 37828 -30295 37857 -30290
rect 37851 -30471 37857 -30295
rect 37828 -30476 37857 -30471
rect 37764 -30482 37857 -30476
rect 37811 -30483 37857 -30482
rect 37894 -30515 37934 -30251
rect 37992 -30283 38036 -30124
rect 37969 -30295 38036 -30283
rect 37969 -30471 37975 -30295
rect 38009 -30471 38036 -30295
rect 37969 -30483 38036 -30471
rect 37992 -30486 38036 -30483
rect 37867 -30521 37959 -30515
rect 37867 -30555 37879 -30521
rect 37947 -30555 37959 -30521
rect 37867 -30561 37959 -30555
rect 37662 -30616 37720 -30604
rect 37344 -30690 37494 -30684
rect 37344 -30748 37350 -30690
rect 37488 -30748 37494 -30690
rect 37344 -30754 37494 -30748
rect 37894 -30812 37934 -30561
rect 37114 -30872 37934 -30812
rect 37002 -31022 37066 -31016
rect 37002 -31056 37014 -31022
rect 37054 -31056 37066 -31022
rect 37002 -31062 37066 -31056
rect 36932 -31104 36978 -31103
rect 36810 -31382 36856 -31341
rect 35770 -31503 35838 -31491
rect 35242 -31550 35306 -31544
rect 35242 -31584 35254 -31550
rect 35294 -31584 35306 -31550
rect 35242 -31590 35306 -31584
rect 35470 -31550 35746 -31544
rect 35470 -31584 35694 -31550
rect 35734 -31584 35746 -31550
rect 35470 -31590 35746 -31584
rect 35794 -31664 35838 -31503
rect 36112 -31388 36856 -31382
rect 36112 -31422 36193 -31388
rect 36747 -31416 36856 -31388
rect 36912 -31115 36978 -31104
rect 36747 -31422 36828 -31416
rect 36112 -31664 36828 -31422
rect 36912 -31491 36938 -31115
rect 36972 -31491 36978 -31115
rect 36912 -31503 36978 -31491
rect 36912 -31664 36956 -31503
rect 37014 -31544 37054 -31062
rect 37114 -31103 37158 -30872
rect 37454 -31016 37494 -31004
rect 37894 -31016 37934 -31004
rect 37442 -31022 37718 -31016
rect 37442 -31056 37454 -31022
rect 37494 -31056 37718 -31022
rect 37442 -31062 37718 -31056
rect 37882 -31022 37946 -31016
rect 37882 -31056 37894 -31022
rect 37934 -31056 37946 -31022
rect 37882 -31062 37946 -31056
rect 37090 -31115 37158 -31103
rect 37372 -31104 37418 -31103
rect 37090 -31491 37096 -31115
rect 37130 -31491 37158 -31115
rect 37090 -31502 37158 -31491
rect 37350 -31115 37418 -31104
rect 37350 -31491 37378 -31115
rect 37412 -31491 37418 -31115
rect 37090 -31503 37136 -31502
rect 37350 -31503 37418 -31491
rect 37002 -31550 37066 -31544
rect 37002 -31584 37014 -31550
rect 37054 -31584 37066 -31550
rect 37002 -31590 37066 -31584
rect 37350 -31664 37394 -31503
rect 37454 -31544 37494 -31062
rect 37530 -31104 37576 -31103
rect 37670 -31104 37718 -31062
rect 37812 -31104 37858 -31103
rect 37530 -31110 37622 -31104
rect 37530 -31115 37558 -31110
rect 37530 -31491 37536 -31115
rect 37616 -31454 37622 -31110
rect 37670 -31110 37858 -31104
rect 37670 -31150 37770 -31110
rect 37828 -31115 37858 -31110
rect 37530 -31496 37558 -31491
rect 37616 -31496 37718 -31454
rect 37530 -31500 37718 -31496
rect 37530 -31502 37622 -31500
rect 37530 -31503 37576 -31502
rect 37670 -31544 37718 -31500
rect 37764 -31496 37770 -31150
rect 37852 -31491 37858 -31115
rect 37828 -31496 37858 -31491
rect 37764 -31502 37858 -31496
rect 37812 -31503 37858 -31502
rect 37894 -31544 37934 -31062
rect 37970 -31104 38016 -31103
rect 37970 -31115 38038 -31104
rect 37970 -31491 37976 -31115
rect 38010 -31491 38038 -31115
rect 37970 -31503 38038 -31491
rect 37442 -31550 37506 -31544
rect 37442 -31584 37454 -31550
rect 37494 -31584 37506 -31550
rect 37442 -31590 37506 -31584
rect 37670 -31550 37946 -31544
rect 37670 -31584 37894 -31550
rect 37934 -31584 37946 -31550
rect 37670 -31590 37946 -31584
rect 37994 -31664 38038 -31503
rect 31712 -31688 33792 -31664
rect 31712 -31690 32438 -31688
rect 31660 -31722 32438 -31690
rect 32830 -31722 32878 -31688
rect 33270 -31722 33318 -31688
rect 33710 -31690 33792 -31688
rect 33912 -31688 35992 -31664
rect 33912 -31690 34638 -31688
rect 33710 -31722 34638 -31690
rect 35030 -31722 35078 -31688
rect 35470 -31722 35518 -31688
rect 35910 -31690 35992 -31688
rect 36112 -31688 38192 -31664
rect 36112 -31690 36838 -31688
rect 35910 -31722 36838 -31690
rect 37230 -31722 37278 -31688
rect 37670 -31722 37718 -31688
rect 38110 -31722 38192 -31688
rect 31660 -31730 38192 -31722
rect 31660 -31950 32540 -31730
rect 33690 -31764 38192 -31730
rect 33690 -31950 38190 -31764
rect 31660 -31990 38190 -31950
rect 22458 -32030 26802 -32024
rect 22458 -32064 22470 -32030
rect 26790 -32064 26802 -32030
rect 22458 -32070 26802 -32064
<< via1 >>
rect 2510 11180 2690 11240
rect 3170 11180 3350 11240
rect 3830 11180 4010 11240
rect 4710 11180 4890 11240
rect 5370 11180 5550 11240
rect 6030 11180 6210 11240
rect 6910 11040 7090 11100
rect 7570 11040 7750 11100
rect 8230 11040 8410 11100
rect 9110 11040 9290 11100
rect 9770 11040 9950 11100
rect 10430 11040 10610 11100
rect 11310 11040 11490 11100
rect 11970 11040 12150 11100
rect 12630 11040 12810 11100
rect 13510 11040 13690 11100
rect 14170 11040 14350 11100
rect 14830 11040 15010 11100
rect 15710 11180 15890 11240
rect 16370 11180 16550 11240
rect 17030 11180 17210 11240
rect 17910 11180 18090 11240
rect 18570 11180 18750 11240
rect 19230 11180 19410 11240
rect -70 10870 -10 10930
rect 2130 10870 2190 10930
rect 2020 10650 2080 10710
rect 4330 10870 4390 10930
rect 4220 10760 4280 10820
rect 4220 10650 4280 10710
rect 6530 10870 6590 10930
rect 6420 10760 6480 10820
rect 6640 10650 6700 10710
rect 8730 10870 8790 10930
rect 8840 10760 8900 10820
rect 8840 10650 8900 10710
rect 10930 10870 10990 10930
rect 11040 10760 11100 10820
rect 11040 10650 11100 10710
rect 13130 10870 13190 10930
rect 13240 10760 13300 10820
rect 13240 10650 13300 10710
rect 15330 10870 15390 10930
rect 15440 10760 15500 10820
rect 15220 10650 15280 10710
rect 17530 10870 17590 10930
rect 17420 10760 17480 10820
rect 17420 10650 17480 10710
rect 19730 10870 19790 10930
rect 21930 10870 21990 10930
rect 19620 10740 19680 10800
rect 2510 10582 4010 10610
rect 2510 10550 4010 10582
rect 4710 10582 6210 10610
rect 4710 10550 6210 10582
rect 6910 10582 8410 10610
rect 6910 10550 8410 10582
rect 9110 10582 10610 10610
rect 9110 10550 10610 10582
rect 11310 10582 12810 10610
rect 11310 10550 12810 10582
rect 13510 10582 15010 10610
rect 13510 10550 15010 10582
rect 15710 10582 17210 10610
rect 15710 10550 17210 10582
rect 17910 10582 19410 10610
rect 17910 10550 19410 10582
rect 2510 10240 2690 10300
rect 3170 10240 3350 10300
rect 3830 10240 4010 10300
rect 4710 10240 4890 10300
rect 5370 10240 5550 10300
rect 6030 10240 6210 10300
rect 6910 10380 7090 10440
rect 7570 10380 7750 10440
rect 8230 10380 8410 10440
rect 9110 10380 9290 10440
rect 9770 10380 9950 10440
rect 10430 10380 10610 10440
rect 11310 10380 11490 10440
rect 11970 10380 12150 10440
rect 12630 10380 12810 10440
rect 13510 10380 13690 10440
rect 14170 10380 14350 10440
rect 14830 10380 15010 10440
rect 15710 10240 15890 10300
rect 16370 10240 16550 10300
rect 17030 10240 17210 10300
rect 17910 10240 18090 10300
rect 18570 10240 18750 10300
rect 19230 10240 19410 10300
rect -70 10070 -10 10130
rect 2130 10070 2190 10130
rect 2240 9850 2300 9910
rect 4330 10070 4390 10130
rect 4440 9960 4500 10020
rect 4440 9850 4500 9910
rect 6530 10070 6590 10130
rect 6640 9960 6700 10020
rect 6420 9850 6480 9910
rect 8730 10070 8790 10130
rect 8620 9960 8680 10020
rect 8620 9850 8680 9910
rect 10930 10070 10990 10130
rect 10820 9960 10880 10020
rect 10820 9850 10880 9910
rect 13130 10070 13190 10130
rect 13020 9960 13080 10020
rect 13020 9850 13080 9910
rect 15330 10070 15390 10130
rect 15220 9960 15280 10020
rect 15440 9850 15500 9910
rect 17530 10070 17590 10130
rect 17640 9960 17700 10020
rect 17640 9850 17700 9910
rect 19730 10070 19790 10130
rect 21930 10070 21990 10130
rect 19840 9940 19900 10000
rect 2510 9782 4010 9810
rect 2510 9750 4010 9782
rect 4710 9782 6210 9810
rect 4710 9750 6210 9782
rect 6910 9782 8410 9810
rect 6910 9750 8410 9782
rect 9110 9782 10610 9810
rect 9110 9750 10610 9782
rect 11310 9782 12810 9810
rect 11310 9750 12810 9782
rect 13510 9782 15010 9810
rect 13510 9750 15010 9782
rect 15710 9782 17210 9810
rect 15710 9750 17210 9782
rect 17910 9782 19410 9810
rect 17910 9750 19410 9782
rect 2510 9580 2690 9640
rect 3170 9580 3350 9640
rect 3830 9580 4010 9640
rect 4710 9580 4890 9640
rect 5370 9580 5550 9640
rect 6030 9580 6210 9640
rect 6910 9440 7090 9500
rect 7570 9440 7750 9500
rect 8230 9440 8410 9500
rect 9110 9440 9290 9500
rect 9770 9440 9950 9500
rect 10430 9440 10610 9500
rect 11310 9440 11490 9500
rect 11970 9440 12150 9500
rect 12630 9440 12810 9500
rect 13510 9440 13690 9500
rect 14170 9440 14350 9500
rect 14830 9440 15010 9500
rect 15710 9580 15890 9640
rect 16370 9580 16550 9640
rect 17030 9580 17210 9640
rect 17910 9580 18090 9640
rect 18570 9580 18750 9640
rect 19230 9580 19410 9640
rect -70 9270 -10 9330
rect 2130 9270 2190 9330
rect 1420 9060 1480 9210
rect 4330 9270 4390 9330
rect 4220 9050 4280 9110
rect 6530 9270 6590 9330
rect 6420 9160 6480 9220
rect 6640 9050 6700 9110
rect 8730 9270 8790 9330
rect 8840 9160 8900 9220
rect 8840 9050 8900 9110
rect 10930 9270 10990 9330
rect 11040 9160 11100 9220
rect 11040 9050 11100 9110
rect 13130 9270 13190 9330
rect 13240 9160 13300 9220
rect 13240 9050 13300 9110
rect 15330 9270 15390 9330
rect 15440 9160 15500 9220
rect 15220 9050 15280 9110
rect 17530 9270 17590 9330
rect 17420 9160 17480 9220
rect 19730 9270 19790 9330
rect 20240 9150 20300 9300
rect 21930 9270 21990 9330
rect 430 8910 610 8990
rect 4710 8982 6210 9010
rect 4710 8950 6210 8982
rect 6910 8982 8410 9010
rect 6910 8950 8410 8982
rect 9110 8982 10610 9010
rect 9110 8950 10610 8982
rect 11310 8982 12810 9010
rect 11310 8950 12810 8982
rect 13510 8982 15010 9010
rect 13510 8950 15010 8982
rect 15710 8982 17210 9010
rect 15710 8950 17210 8982
rect 21310 8910 21490 8990
rect 2510 8640 2690 8700
rect 3170 8640 3350 8700
rect 3830 8640 4010 8700
rect 4710 8640 4890 8700
rect 5370 8640 5550 8700
rect 6030 8640 6210 8700
rect 6910 8780 7090 8840
rect 7570 8780 7750 8840
rect 8230 8780 8410 8840
rect 9110 8780 9290 8840
rect 9770 8780 9950 8840
rect 10430 8780 10610 8840
rect 11310 8780 11490 8840
rect 11970 8780 12150 8840
rect 12630 8780 12810 8840
rect 13510 8780 13690 8840
rect 14170 8780 14350 8840
rect 14830 8780 15010 8840
rect 15710 8640 15890 8700
rect 16370 8640 16550 8700
rect 17030 8640 17210 8700
rect 17910 8640 18090 8700
rect 18570 8640 18750 8700
rect 19230 8640 19410 8700
rect -70 8470 -10 8530
rect 2130 8470 2190 8530
rect 1620 8260 1680 8410
rect 4330 8470 4390 8530
rect 4440 8250 4500 8310
rect 6530 8470 6590 8530
rect 6640 8360 6700 8420
rect 6420 8250 6480 8310
rect 8730 8470 8790 8530
rect 8620 8360 8680 8420
rect 8620 8250 8680 8310
rect 10930 8470 10990 8530
rect 10820 8360 10880 8420
rect 10820 8250 10880 8310
rect 13130 8470 13190 8530
rect 13020 8360 13080 8420
rect 13020 8250 13080 8310
rect 15330 8470 15390 8530
rect 15220 8360 15280 8420
rect 15440 8250 15500 8310
rect 17530 8470 17590 8530
rect 17640 8360 17700 8420
rect 19730 8470 19790 8530
rect 20440 8350 20500 8500
rect 21930 8470 21990 8530
rect 430 8110 610 8190
rect 4710 8182 6210 8210
rect 4710 8150 6210 8182
rect 6910 8182 8410 8210
rect 6910 8150 8410 8182
rect 9110 8182 10610 8210
rect 9110 8150 10610 8182
rect 11310 8182 12810 8210
rect 11310 8150 12810 8182
rect 13510 8182 15010 8210
rect 13510 8150 15010 8182
rect 15710 8182 17210 8210
rect 15710 8150 17210 8182
rect 21310 8110 21490 8190
rect 2510 7840 2690 7900
rect 3170 7840 3350 7900
rect 3830 7840 4010 7900
rect 4710 7840 4890 7900
rect 5370 7840 5550 7900
rect 6030 7840 6210 7900
rect 6910 7980 7090 8040
rect 7570 7980 7750 8040
rect 8230 7980 8410 8040
rect 9110 7980 9290 8040
rect 9770 7980 9950 8040
rect 10430 7980 10610 8040
rect 11310 7980 11490 8040
rect 11970 7980 12150 8040
rect 12630 7980 12810 8040
rect 13510 7980 13690 8040
rect 14170 7980 14350 8040
rect 14830 7980 15010 8040
rect 15710 7840 15890 7900
rect 16370 7840 16550 7900
rect 17030 7840 17210 7900
rect 17910 7840 18090 7900
rect 18570 7840 18750 7900
rect 19230 7840 19410 7900
rect -70 7670 -10 7730
rect 2130 7670 2190 7730
rect 1620 7460 1680 7610
rect 4330 7670 4390 7730
rect 4440 7450 4500 7510
rect 6530 7670 6590 7730
rect 6640 7560 6700 7620
rect 6420 7450 6480 7510
rect 8730 7670 8790 7730
rect 8620 7560 8680 7620
rect 8620 7450 8680 7510
rect 10930 7670 10990 7730
rect 10820 7560 10880 7620
rect 10820 7450 10880 7510
rect 13130 7670 13190 7730
rect 13020 7560 13080 7620
rect 13020 7450 13080 7510
rect 15330 7670 15390 7730
rect 15220 7560 15280 7620
rect 15440 7450 15500 7510
rect 17530 7670 17590 7730
rect 17640 7560 17700 7620
rect 19730 7670 19790 7730
rect 20440 7550 20500 7700
rect 21930 7670 21990 7730
rect 430 7310 610 7390
rect 4710 7382 6210 7410
rect 4710 7350 6210 7382
rect 6910 7382 8410 7410
rect 6910 7350 8410 7382
rect 9110 7382 10610 7410
rect 9110 7350 10610 7382
rect 11310 7382 12810 7410
rect 11310 7350 12810 7382
rect 13510 7382 15010 7410
rect 13510 7350 15010 7382
rect 15710 7382 17210 7410
rect 15710 7350 17210 7382
rect 21310 7310 21490 7390
rect 2510 7180 2690 7240
rect 3170 7180 3350 7240
rect 3830 7180 4010 7240
rect 4710 7180 4890 7240
rect 5370 7180 5550 7240
rect 6030 7180 6210 7240
rect 6910 7040 7090 7100
rect 7570 7040 7750 7100
rect 8230 7040 8410 7100
rect 9110 7040 9290 7100
rect 9770 7040 9950 7100
rect 10430 7040 10610 7100
rect 11310 7040 11490 7100
rect 11970 7040 12150 7100
rect 12630 7040 12810 7100
rect 13510 7040 13690 7100
rect 14170 7040 14350 7100
rect 14830 7040 15010 7100
rect 15710 7180 15890 7240
rect 16370 7180 16550 7240
rect 17030 7180 17210 7240
rect 17910 7180 18090 7240
rect 18570 7180 18750 7240
rect 19230 7180 19410 7240
rect -70 6870 -10 6930
rect 2130 6870 2190 6930
rect 1420 6660 1480 6810
rect 4330 6870 4390 6930
rect 4220 6650 4280 6710
rect 6530 6870 6590 6930
rect 6420 6760 6480 6820
rect 6640 6650 6700 6710
rect 8730 6870 8790 6930
rect 8840 6760 8900 6820
rect 8840 6650 8900 6710
rect 10930 6870 10990 6930
rect 11040 6760 11100 6820
rect 11040 6650 11100 6710
rect 13130 6870 13190 6930
rect 13240 6760 13300 6820
rect 13240 6650 13300 6710
rect 15330 6870 15390 6930
rect 15440 6760 15500 6820
rect 15220 6650 15280 6710
rect 17530 6870 17590 6930
rect 17420 6760 17480 6820
rect 19730 6870 19790 6930
rect 20240 6750 20300 6900
rect 21930 6870 21990 6930
rect 430 6510 610 6590
rect 4710 6582 6210 6610
rect 4710 6550 6210 6582
rect 6910 6582 8410 6610
rect 6910 6550 8410 6582
rect 9110 6582 10610 6610
rect 9110 6550 10610 6582
rect 11310 6582 12810 6610
rect 11310 6550 12810 6582
rect 13510 6582 15010 6610
rect 13510 6550 15010 6582
rect 15710 6582 17210 6610
rect 15710 6550 17210 6582
rect 21310 6510 21490 6590
rect 2510 6240 2690 6300
rect 3170 6240 3350 6300
rect 3830 6240 4010 6300
rect 4710 6240 4890 6300
rect 5370 6240 5550 6300
rect 6030 6240 6210 6300
rect 6910 6380 7090 6440
rect 7570 6380 7750 6440
rect 8230 6380 8410 6440
rect 9110 6380 9290 6440
rect 9770 6380 9950 6440
rect 10430 6380 10610 6440
rect 11310 6380 11490 6440
rect 11970 6380 12150 6440
rect 12630 6380 12810 6440
rect 13510 6380 13690 6440
rect 14170 6380 14350 6440
rect 14830 6380 15010 6440
rect 15710 6240 15890 6300
rect 16370 6240 16550 6300
rect 17030 6240 17210 6300
rect 17910 6240 18090 6300
rect 18570 6240 18750 6300
rect 19230 6240 19410 6300
rect -70 6070 -10 6130
rect 2130 6070 2190 6130
rect 2240 5850 2300 5910
rect 4330 6070 4390 6130
rect 4440 5960 4500 6020
rect 4440 5850 4500 5910
rect 6530 6070 6590 6130
rect 6640 5960 6700 6020
rect 6420 5850 6480 5910
rect 8730 6070 8790 6130
rect 8620 5960 8680 6020
rect 8620 5850 8680 5910
rect 10930 6070 10990 6130
rect 10820 5960 10880 6020
rect 10820 5850 10880 5910
rect 13130 6070 13190 6130
rect 13020 5960 13080 6020
rect 13020 5850 13080 5910
rect 15330 6070 15390 6130
rect 15220 5960 15280 6020
rect 15440 5850 15500 5910
rect 17530 6070 17590 6130
rect 17640 5960 17700 6020
rect 17640 5850 17700 5910
rect 19730 6070 19790 6130
rect 21930 6070 21990 6130
rect 19840 5940 19900 6000
rect 2510 5782 4010 5810
rect 2510 5750 4010 5782
rect 4710 5782 6210 5810
rect 4710 5750 6210 5782
rect 6910 5782 8410 5810
rect 6910 5750 8410 5782
rect 9110 5782 10610 5810
rect 9110 5750 10610 5782
rect 11310 5782 12810 5810
rect 11310 5750 12810 5782
rect 13510 5782 15010 5810
rect 13510 5750 15010 5782
rect 15710 5782 17210 5810
rect 15710 5750 17210 5782
rect 17910 5782 19410 5810
rect 17910 5750 19410 5782
rect 2510 5580 2690 5640
rect 3170 5580 3350 5640
rect 3830 5580 4010 5640
rect 4710 5580 4890 5640
rect 5370 5580 5550 5640
rect 6030 5580 6210 5640
rect 6910 5440 7090 5500
rect 7570 5440 7750 5500
rect 8230 5440 8410 5500
rect 9110 5440 9290 5500
rect 9770 5440 9950 5500
rect 10430 5440 10610 5500
rect 11310 5440 11490 5500
rect 11970 5440 12150 5500
rect 12630 5440 12810 5500
rect 13510 5440 13690 5500
rect 14170 5440 14350 5500
rect 14830 5440 15010 5500
rect 15710 5580 15890 5640
rect 16370 5580 16550 5640
rect 17030 5580 17210 5640
rect 17910 5580 18090 5640
rect 18570 5580 18750 5640
rect 19230 5580 19410 5640
rect -70 5270 -10 5330
rect 2130 5270 2190 5330
rect 2020 5050 2080 5110
rect 4330 5270 4390 5330
rect 4220 5160 4280 5220
rect 4220 5050 4280 5110
rect 6530 5270 6590 5330
rect 6420 5160 6480 5220
rect 6640 5050 6700 5110
rect 8730 5270 8790 5330
rect 8840 5160 8900 5220
rect 8840 5050 8900 5110
rect 10930 5270 10990 5330
rect 11040 5160 11100 5220
rect 11040 5050 11100 5110
rect 13130 5270 13190 5330
rect 13240 5160 13300 5220
rect 13240 5050 13300 5110
rect 15330 5270 15390 5330
rect 15440 5160 15500 5220
rect 15220 5050 15280 5110
rect 17530 5270 17590 5330
rect 17420 5160 17480 5220
rect 17420 5050 17480 5110
rect 19730 5270 19790 5330
rect 21930 5270 21990 5330
rect 19620 5140 19680 5200
rect 2510 4982 4010 5010
rect 2510 4950 4010 4982
rect 4710 4982 6210 5010
rect 4710 4950 6210 4982
rect 6910 4982 8410 5010
rect 6910 4950 8410 4982
rect 9110 4982 10610 5010
rect 9110 4950 10610 4982
rect 11310 4982 12810 5010
rect 11310 4950 12810 4982
rect 13510 4982 15010 5010
rect 13510 4950 15010 4982
rect 15710 4982 17210 5010
rect 15710 4950 17210 4982
rect 17910 4982 19410 5010
rect 17910 4950 19410 4982
rect 25720 11410 26240 11780
rect 7800 4540 7940 4680
rect 23050 4600 23580 4970
rect 27260 11400 27320 11490
rect 30576 11715 30664 11722
rect 30576 11539 30610 11715
rect 30610 11539 30664 11715
rect 30576 11532 30664 11539
rect 27740 11240 27800 11330
rect 30154 11364 30288 11416
rect 28780 11231 28840 11260
rect 27260 11080 27320 11170
rect 28780 11177 28807 11231
rect 28807 11177 28840 11231
rect 28780 11073 28840 11177
rect 27740 10925 27800 11015
rect 28780 11040 28807 11073
rect 28807 11040 28840 11073
rect 30190 11190 30390 11270
rect 30600 11262 30738 11320
rect 27260 10765 27320 10855
rect 31478 11715 31536 11722
rect 31478 11539 31489 11715
rect 31489 11539 31536 11715
rect 31478 11536 31536 11539
rect 31690 11715 31748 11720
rect 31690 11539 31737 11715
rect 31737 11539 31748 11715
rect 31690 11534 31748 11539
rect 31270 11262 31408 11320
rect 32776 11715 32864 11722
rect 32776 11539 32810 11715
rect 32810 11539 32864 11715
rect 32776 11532 32864 11539
rect 32354 11364 32488 11416
rect 32390 11190 32590 11270
rect 32800 11262 32938 11320
rect 27740 10360 27800 10450
rect 27380 10200 27440 10290
rect 31478 10895 31536 10900
rect 31478 10519 31490 10895
rect 31490 10519 31536 10895
rect 31690 10895 31748 10900
rect 31478 10514 31536 10519
rect 31690 10519 31738 10895
rect 31738 10519 31748 10895
rect 31690 10514 31748 10519
rect 33678 11715 33736 11722
rect 33678 11539 33689 11715
rect 33689 11539 33736 11715
rect 33678 11536 33736 11539
rect 33890 11715 33948 11720
rect 33890 11539 33937 11715
rect 33937 11539 33948 11715
rect 33890 11534 33948 11539
rect 33470 11262 33608 11320
rect 34976 11715 35064 11722
rect 34976 11539 35010 11715
rect 35010 11539 35064 11715
rect 34976 11532 35064 11539
rect 34554 11364 34688 11416
rect 34570 11190 34770 11270
rect 35000 11262 35138 11320
rect 33678 10895 33736 10900
rect 33678 10519 33690 10895
rect 33690 10519 33736 10895
rect 33890 10895 33948 10900
rect 33678 10514 33736 10519
rect 33890 10519 33938 10895
rect 33938 10519 33948 10895
rect 33890 10514 33948 10519
rect 35878 11715 35936 11722
rect 35878 11539 35889 11715
rect 35889 11539 35936 11715
rect 35878 11536 35936 11539
rect 36090 11715 36148 11720
rect 36090 11539 36137 11715
rect 36137 11539 36148 11715
rect 36090 11534 36148 11539
rect 36480 11510 36810 11980
rect 35670 11262 35808 11320
rect 35878 10895 35936 10900
rect 35878 10519 35890 10895
rect 35890 10519 35936 10895
rect 36090 10895 36148 10900
rect 35878 10514 35936 10519
rect 36090 10519 36138 10895
rect 36138 10519 36148 10895
rect 36090 10514 36148 10519
rect 27740 10040 27800 10130
rect 27380 9885 27440 9975
rect 29140 9970 29200 10190
rect 27740 9725 27800 9815
rect 27260 9315 27320 9405
rect 27500 9160 27560 9250
rect 27260 9000 27320 9090
rect 27500 8845 27560 8935
rect 28880 8940 28940 9160
rect 31460 9220 31482 9410
rect 31482 9243 31582 9410
rect 31582 9243 31616 9410
rect 31616 9243 31670 9410
rect 31482 9220 31670 9243
rect 27260 8685 27320 8775
rect 31450 8780 31680 8990
rect 32070 8990 32200 9120
rect 27260 8280 27320 8370
rect 27620 8120 27680 8210
rect 27260 7960 27320 8050
rect 27620 7800 27680 7890
rect 29010 7890 29070 8110
rect 27260 7650 27320 7740
rect 30570 8210 30590 8580
rect 30590 8210 30624 8580
rect 30624 8210 30640 8580
rect 30890 8112 31280 8120
rect 30890 8038 31280 8112
rect 30890 8030 31280 8038
rect 30570 7570 30590 7940
rect 30590 7570 30624 7940
rect 30624 7570 30640 7940
rect 33670 8071 33750 8830
rect 33750 8071 33770 8830
rect 33670 8030 33770 8071
rect 34500 8880 35520 8940
rect 34510 8440 34590 8600
rect 34590 8440 34610 8600
rect 34930 8440 35010 8600
rect 35010 8440 35030 8600
rect 35350 8450 35430 8610
rect 35430 8450 35450 8610
rect 32300 7890 32460 7970
rect 34290 7930 34360 7990
rect 34290 7850 34610 7930
rect 34290 7790 34360 7850
rect 32260 7570 32320 7770
rect 27380 7240 27440 7330
rect 27620 7080 27680 7170
rect 27380 6925 27440 7015
rect 27620 6765 27680 6855
rect 28880 6860 28940 7080
rect 27380 6610 27440 6700
rect 30470 7064 30850 7150
rect 30470 7050 30545 7064
rect 30545 7050 30850 7064
rect 30120 6410 30420 6470
rect 27380 6200 27440 6290
rect 27500 6040 27560 6130
rect 27380 5885 27440 5975
rect 27500 5725 27560 5815
rect 29010 5820 29070 6040
rect 27380 5570 27440 5660
rect 27180 5110 27310 5240
rect 30060 5670 30240 5730
rect 8620 4250 8680 4310
rect 10820 4360 10880 4420
rect 11040 4250 11100 4310
rect 13240 4360 13300 4420
rect 30040 5070 30320 5170
rect 29770 4682 30546 4710
rect 30546 4682 30550 4710
rect 29770 4640 30550 4682
rect 33460 6966 33548 6990
rect 33548 6966 33588 6990
rect 33588 6966 33590 6990
rect 33460 6930 33590 6966
rect 33700 6966 33706 6990
rect 33706 6966 33746 6990
rect 33746 6966 33864 6990
rect 33864 6966 33904 6990
rect 33904 6966 33910 6990
rect 33700 6930 33910 6966
rect 34750 7960 34890 8180
rect 35170 7760 35310 7980
rect 34500 7150 34590 7310
rect 34590 7150 34600 7310
rect 34920 7150 35010 7310
rect 35010 7150 35020 7310
rect 35340 7150 35430 7310
rect 35430 7150 35440 7310
rect 34020 6966 34022 6990
rect 34022 6966 34062 6990
rect 34062 6966 34190 6990
rect 34020 6930 34190 6966
rect 34500 6830 35540 6920
rect 31080 6250 31380 6310
rect 36230 6080 36410 6260
rect 36530 6080 36710 6260
rect 31380 5680 31560 5740
rect 36300 5820 36376 5890
rect 36376 5820 36390 5890
rect 37680 5820 37706 5890
rect 37706 5820 37770 5890
rect 36300 5560 36376 5630
rect 36376 5560 36390 5630
rect 33330 5020 33630 5290
rect 36300 5300 36376 5370
rect 36376 5300 36390 5370
rect 37680 5560 37706 5630
rect 37706 5560 37770 5630
rect 37680 5300 37706 5370
rect 37706 5300 37770 5370
rect 36300 5040 36376 5110
rect 36376 5040 36390 5110
rect 32260 4650 32320 4880
rect 10890 3960 11030 4100
rect 30080 3860 30260 4040
rect 36300 4780 36376 4850
rect 36376 4780 36390 4850
rect 37680 5040 37706 5110
rect 37706 5040 37770 5110
rect 37680 4780 37706 4850
rect 37706 4780 37770 4850
rect 36300 4520 36376 4590
rect 36376 4520 36390 4590
rect 31680 3860 31860 4040
rect 32810 4030 32980 4070
rect 32810 4010 32835 4030
rect 32835 4010 32959 4030
rect 32959 4010 32980 4030
rect 16910 2640 17102 2780
rect 17102 2640 17130 2780
rect 17380 2640 17418 2780
rect 17418 2640 17452 2780
rect 17452 2640 17490 2780
rect 33130 4030 33300 4070
rect 33130 4010 33151 4030
rect 33151 4010 33275 4030
rect 33275 4010 33300 4030
rect 33440 4030 33610 4070
rect 33440 4010 33467 4030
rect 33467 4010 33591 4030
rect 33591 4010 33610 4030
rect 33760 4030 33930 4070
rect 33760 4010 33783 4030
rect 33783 4010 33907 4030
rect 33907 4010 33930 4030
rect 34870 4030 35190 4090
rect 34870 4010 34991 4030
rect 34991 4010 35025 4030
rect 35025 4010 35149 4030
rect 35149 4010 35183 4030
rect 35183 4010 35190 4030
rect 32850 3350 33870 3430
rect 36300 4260 36376 4330
rect 36376 4260 36390 4330
rect 37680 4520 37706 4590
rect 37706 4520 37770 4590
rect 37680 4260 37706 4330
rect 37706 4260 37770 4330
rect 36300 4000 36376 4070
rect 36376 4000 36390 4070
rect 35070 3350 35410 3430
rect 36380 3440 36520 3580
rect 37680 4000 37706 4070
rect 37706 4000 37770 4070
rect 18060 2870 18200 3010
rect 17740 2640 17768 2780
rect 17768 2640 17960 2780
rect 32466 3100 32668 3156
rect 32466 3068 32471 3100
rect 32471 3068 32505 3100
rect 32505 3068 32629 3100
rect 32629 3068 32663 3100
rect 32663 3068 32668 3100
rect 34066 3100 34268 3156
rect 34066 3068 34071 3100
rect 34071 3068 34105 3100
rect 34105 3068 34229 3100
rect 34229 3068 34263 3100
rect 34263 3068 34268 3100
rect 32450 2430 32690 2510
rect 34050 2430 34290 2510
rect 35666 3100 35868 3156
rect 35666 3068 35671 3100
rect 35671 3068 35705 3100
rect 35705 3068 35829 3100
rect 35829 3068 35863 3100
rect 35863 3068 35868 3100
rect 35650 2430 35890 2510
rect 480 2195 660 2220
rect 480 1995 660 2195
rect 32450 2095 32690 2130
rect 34050 2095 34290 2130
rect 32450 2070 32689 2095
rect 32689 2070 32690 2095
rect 34050 2070 34289 2095
rect 34289 2070 34290 2095
rect 35650 2095 35890 2130
rect 35650 2070 35889 2095
rect 35889 2070 35890 2095
rect 480 1303 497 1995
rect 497 1303 531 1995
rect 531 1303 605 1995
rect 605 1303 639 1995
rect 639 1303 660 1995
rect 480 870 660 1303
rect 2110 1310 2131 1990
rect 2131 1310 2205 1990
rect 2205 1310 2230 1990
rect 3710 1310 3731 1990
rect 3731 1310 3805 1990
rect 3805 1310 3830 1990
rect 5310 1310 5331 1990
rect 5331 1310 5405 1990
rect 5405 1310 5430 1990
rect 6910 1310 6931 1990
rect 6931 1310 7005 1990
rect 7005 1310 7030 1990
rect 8510 1310 8531 1990
rect 8531 1310 8605 1990
rect 8605 1310 8630 1990
rect 10110 1310 10131 1990
rect 10131 1310 10205 1990
rect 10205 1310 10230 1990
rect 11030 1330 11150 1950
rect 12610 1330 12730 1950
rect 13990 1330 14110 1950
rect 14910 1320 14931 1980
rect 14931 1320 15005 1980
rect 15005 1320 15030 1980
rect 16510 1310 16531 1990
rect 16531 1310 16605 1990
rect 16605 1310 16630 1990
rect 18110 1310 18131 1990
rect 18131 1310 18205 1990
rect 18205 1310 18230 1990
rect 19710 1310 19731 1990
rect 19731 1310 19805 1990
rect 19805 1310 19830 1990
rect 21310 1310 21331 1990
rect 21331 1310 21405 1990
rect 21405 1310 21430 1990
rect 22910 1310 22931 1990
rect 22931 1310 23005 1990
rect 23005 1310 23030 1990
rect 24510 1310 24531 1990
rect 24531 1310 24605 1990
rect 24605 1310 24630 1990
rect 26110 1310 26131 1990
rect 26131 1310 26205 1990
rect 26205 1310 26230 1990
rect 27710 1310 27731 1990
rect 27731 1310 27805 1990
rect 27805 1310 27830 1990
rect 29310 1310 29331 1990
rect 29331 1310 29405 1990
rect 29405 1310 29430 1990
rect 30910 1310 30931 1990
rect 30931 1310 31005 1990
rect 31005 1310 31030 1990
rect 32510 1310 32531 1990
rect 32531 1310 32605 1990
rect 32605 1310 32630 1990
rect 34110 1310 34131 1990
rect 34131 1310 34205 1990
rect 34205 1310 34230 1990
rect 35710 1310 35731 1990
rect 35731 1310 35805 1990
rect 35805 1310 35830 1990
rect 37310 1310 37331 1990
rect 37331 1310 37405 1990
rect 37405 1310 37430 1990
rect 1410 1030 1530 1150
rect 3010 1030 3130 1150
rect 4610 1030 4730 1150
rect 6210 1030 6330 1150
rect 7810 1030 7930 1150
rect 9410 1030 9530 1150
rect 11250 1203 11271 1230
rect 11271 1203 11647 1230
rect 11647 1203 11670 1230
rect 11250 1070 11670 1203
rect 15600 1030 15700 1150
rect 17200 1030 17300 1150
rect 18800 1030 18900 1150
rect 20400 1030 20500 1150
rect 22000 1030 22100 1150
rect 23600 1030 23700 1150
rect 26800 1030 26900 1150
rect 28400 1030 28500 1150
rect 480 736 497 870
rect 497 736 531 870
rect 531 736 605 870
rect 605 736 639 870
rect 639 736 660 870
rect 480 429 660 736
rect 12390 750 12510 870
rect 1190 560 1310 680
rect 2790 560 2910 680
rect 4390 560 4510 680
rect 5990 560 6110 680
rect 7590 560 7710 680
rect 9190 560 9310 680
rect 15820 560 15920 680
rect 17420 560 17520 680
rect 19020 560 19120 680
rect 20620 560 20720 680
rect 22220 560 22320 680
rect 23820 560 23920 680
rect 27020 560 27120 680
rect 28620 560 28720 680
rect 31820 560 31920 680
rect 36600 550 36720 670
rect 37850 530 37970 650
rect 480 395 660 429
rect 480 195 660 395
rect 480 -497 497 195
rect 497 -497 531 195
rect 531 -497 605 195
rect 605 -497 639 195
rect 639 -497 660 195
rect 480 -930 660 -497
rect 2110 -490 2131 190
rect 2131 -490 2205 190
rect 2205 -490 2230 190
rect 3710 -490 3731 190
rect 3731 -490 3805 190
rect 3805 -490 3830 190
rect 5310 -490 5331 190
rect 5331 -490 5405 190
rect 5405 -490 5430 190
rect 6910 -490 6931 190
rect 6931 -490 7005 190
rect 7005 -490 7030 190
rect 8510 -490 8531 190
rect 8531 -490 8605 190
rect 8605 -490 8630 190
rect 10110 -490 10131 190
rect 10131 -490 10205 190
rect 10205 -490 10230 190
rect 11710 -497 11731 190
rect 11731 -497 11805 190
rect 11805 -497 11830 190
rect 11710 -570 11830 -497
rect 13310 -490 13331 190
rect 13331 -490 13405 190
rect 13405 -490 13430 190
rect 11270 -597 11271 -570
rect 11271 -597 11647 -570
rect 11647 -597 11889 -570
rect 11889 -597 12265 -570
rect 12265 -597 12270 -570
rect 1410 -770 1530 -650
rect 3010 -770 3130 -650
rect 4610 -770 4730 -650
rect 6210 -770 6330 -650
rect 7810 -770 7930 -650
rect 9410 -770 9530 -650
rect 11270 -730 12270 -597
rect 14910 -497 14931 190
rect 14931 -497 15005 190
rect 15005 -497 15030 190
rect 14910 -570 15030 -497
rect 16510 -490 16531 190
rect 16531 -490 16605 190
rect 16605 -490 16630 190
rect 18110 -490 18131 190
rect 18131 -490 18205 190
rect 18205 -490 18230 190
rect 19710 -490 19731 190
rect 19731 -490 19805 190
rect 19805 -490 19830 190
rect 21310 -490 21331 190
rect 21331 -490 21405 190
rect 21405 -490 21430 190
rect 22910 -490 22931 190
rect 22931 -490 23005 190
rect 23005 -490 23030 190
rect 24510 -490 24531 190
rect 24531 -490 24605 190
rect 24605 -490 24630 190
rect 26110 -490 26131 190
rect 26131 -490 26205 190
rect 26205 -490 26230 190
rect 27710 -490 27731 190
rect 27731 -490 27805 190
rect 27805 -490 27830 190
rect 29310 -490 29331 190
rect 29331 -490 29405 190
rect 29405 -490 29430 190
rect 30910 -490 30931 190
rect 30931 -490 31005 190
rect 31005 -490 31030 190
rect 32510 -490 32531 190
rect 32531 -490 32605 190
rect 32605 -490 32630 190
rect 34110 -490 34131 190
rect 34131 -490 34205 190
rect 34205 -490 34230 190
rect 35710 -490 35731 190
rect 35731 -490 35805 190
rect 35805 -490 35830 190
rect 12390 -810 12510 -650
rect 14470 -597 14471 -570
rect 14471 -597 14847 -570
rect 14847 -597 15089 -570
rect 15089 -597 15465 -570
rect 15465 -597 15470 -570
rect 14470 -730 15470 -597
rect 15600 -770 15700 -650
rect 17200 -770 17300 -650
rect 18800 -770 18900 -650
rect 20400 -770 20500 -650
rect 22000 -770 22100 -650
rect 23600 -770 23700 -650
rect 26800 -770 26900 -650
rect 28400 -770 28500 -650
rect 480 -1064 497 -930
rect 497 -1064 531 -930
rect 531 -1064 605 -930
rect 605 -1064 639 -930
rect 639 -1064 660 -930
rect 480 -1371 660 -1064
rect 12390 -1050 12510 -980
rect 12630 -1070 12750 -930
rect 13970 -1070 14090 -930
rect 1190 -1240 1310 -1120
rect 2790 -1240 2910 -1120
rect 4390 -1240 4510 -1120
rect 5990 -1240 6110 -1120
rect 7590 -1240 7710 -1120
rect 9190 -1240 9310 -1120
rect 12880 -1143 13240 -1110
rect 12880 -1260 13240 -1143
rect 15820 -1240 15920 -1120
rect 17420 -1240 17520 -1120
rect 19020 -1240 19120 -1120
rect 20620 -1240 20720 -1120
rect 22220 -1240 22320 -1120
rect 23820 -1240 23920 -1120
rect 27020 -1240 27120 -1120
rect 28620 -1240 28720 -1120
rect 31600 -1240 31700 -1120
rect 480 -1405 660 -1371
rect 480 -1605 660 -1405
rect 480 -2297 497 -1605
rect 497 -2297 531 -1605
rect 531 -2297 605 -1605
rect 605 -2297 639 -1605
rect 639 -2297 660 -1605
rect 480 -2730 660 -2297
rect 33360 -1590 33480 -1470
rect 2110 -2290 2131 -1610
rect 2131 -2290 2205 -1610
rect 2205 -2290 2230 -1610
rect 3710 -2290 3731 -1610
rect 3731 -2290 3805 -1610
rect 3805 -2290 3830 -1610
rect 5310 -2290 5331 -1610
rect 5331 -2290 5405 -1610
rect 5405 -2290 5430 -1610
rect 6910 -2290 6931 -1610
rect 6931 -2290 7005 -1610
rect 7005 -2290 7030 -1610
rect 8510 -2290 8531 -1610
rect 8531 -2290 8605 -1610
rect 8605 -2290 8630 -1610
rect 10110 -2290 10131 -1610
rect 10131 -2290 10205 -1610
rect 10205 -2290 10230 -1610
rect 11710 -2290 11731 -1610
rect 11731 -2290 11805 -1610
rect 11805 -2290 11830 -1610
rect 13310 -2290 13331 -1610
rect 13331 -2290 13405 -1610
rect 13405 -2290 13430 -1610
rect 14910 -2290 14931 -1610
rect 14931 -2290 15005 -1610
rect 15005 -2290 15030 -1610
rect 16510 -2290 16531 -1610
rect 16531 -2290 16605 -1610
rect 16605 -2290 16630 -1610
rect 18110 -2290 18131 -1610
rect 18131 -2290 18205 -1610
rect 18205 -2290 18230 -1610
rect 19710 -2290 19731 -1610
rect 19731 -2290 19805 -1610
rect 19805 -2290 19830 -1610
rect 21310 -2290 21331 -1610
rect 21331 -2290 21405 -1610
rect 21405 -2290 21430 -1610
rect 22910 -2290 22931 -1610
rect 22931 -2290 23005 -1610
rect 23005 -2290 23030 -1610
rect 24510 -2290 24531 -1610
rect 24531 -2290 24605 -1610
rect 24605 -2290 24630 -1610
rect 26110 -2290 26131 -1610
rect 26131 -2290 26205 -1610
rect 26205 -2290 26230 -1610
rect 27710 -2290 27731 -1610
rect 27731 -2290 27805 -1610
rect 27805 -2290 27830 -1610
rect 29310 -2290 29331 -1610
rect 29331 -2290 29405 -1610
rect 29405 -2290 29430 -1610
rect 30910 -2290 30931 -1610
rect 30931 -2290 31005 -1610
rect 31005 -2290 31030 -1610
rect 32510 -2290 32531 -1610
rect 32531 -2290 32605 -1610
rect 32605 -2290 32630 -1610
rect 35020 -1590 35140 -1470
rect 34110 -2290 34131 -1610
rect 34131 -2290 34205 -1610
rect 34205 -2290 34230 -1610
rect 35690 -1605 35750 -1600
rect 35690 -2297 35697 -1605
rect 35697 -2297 35731 -1605
rect 35731 -2297 35750 -1605
rect 35690 -2310 35750 -2297
rect 1410 -2570 1530 -2450
rect 3010 -2570 3130 -2450
rect 4610 -2570 4730 -2450
rect 6210 -2570 6330 -2450
rect 7810 -2570 7930 -2450
rect 9410 -2570 9530 -2450
rect 15600 -2570 15700 -2450
rect 17200 -2570 17300 -2450
rect 18800 -2570 18900 -2450
rect 20400 -2570 20500 -2450
rect 22000 -2570 22100 -2450
rect 23600 -2570 23700 -2450
rect 25200 -2570 25300 -2450
rect 26800 -2570 26900 -2450
rect 28400 -2570 28500 -2450
rect 30000 -2570 30100 -2450
rect 33180 -2570 33300 -2450
rect 480 -2864 497 -2730
rect 497 -2864 531 -2730
rect 531 -2864 605 -2730
rect 605 -2864 639 -2730
rect 639 -2864 660 -2730
rect 480 -3171 660 -2864
rect 12390 -2850 12510 -2730
rect 1190 -3040 1310 -2920
rect 2790 -3040 2910 -2920
rect 4390 -3040 4510 -2920
rect 5990 -3040 6110 -2920
rect 7590 -3040 7710 -2920
rect 9190 -3040 9310 -2920
rect 11010 -3040 11130 -2920
rect 14210 -3040 14330 -2920
rect 14430 -2943 14471 -2920
rect 14471 -2943 14550 -2920
rect 14430 -3040 14550 -2943
rect 15820 -3040 15920 -2920
rect 17420 -3040 17520 -2920
rect 19020 -3040 19120 -2920
rect 20620 -3040 20720 -2920
rect 22220 -3040 22320 -2920
rect 23820 -3040 23920 -2920
rect 25420 -3040 25520 -2920
rect 27020 -3040 27120 -2920
rect 28620 -3040 28720 -2920
rect 30220 -3040 30320 -2920
rect 36400 -3030 36500 -2910
rect 480 -3205 660 -3171
rect 480 -3405 660 -3205
rect 480 -4097 497 -3405
rect 497 -4097 531 -3405
rect 531 -4097 605 -3405
rect 605 -4097 639 -3405
rect 639 -4097 660 -3405
rect 480 -4530 660 -4097
rect 12610 -3390 12730 -3290
rect 2110 -4090 2131 -3410
rect 2131 -4090 2205 -3410
rect 2205 -4090 2230 -3410
rect 3710 -4090 3731 -3410
rect 3731 -4090 3805 -3410
rect 3805 -4090 3830 -3410
rect 5310 -4090 5331 -3410
rect 5331 -4090 5405 -3410
rect 5405 -4090 5430 -3410
rect 6910 -4090 6931 -3410
rect 6931 -4090 7005 -3410
rect 7005 -4090 7030 -3410
rect 8510 -4090 8531 -3410
rect 8531 -4090 8605 -3410
rect 8605 -4090 8630 -3410
rect 10110 -4090 10131 -3410
rect 10131 -4090 10205 -3410
rect 10205 -4090 10230 -3410
rect 11710 -4090 11731 -3410
rect 11731 -4090 11805 -3410
rect 11805 -4090 11830 -3410
rect 13310 -4090 13331 -3410
rect 13331 -4090 13405 -3410
rect 13405 -4090 13430 -3410
rect 14210 -3410 14330 -3290
rect 14910 -4090 14931 -3410
rect 14931 -4090 15005 -3410
rect 15005 -4090 15030 -3410
rect 16510 -4090 16531 -3410
rect 16531 -4090 16605 -3410
rect 16605 -4090 16630 -3410
rect 18110 -4090 18131 -3410
rect 18131 -4090 18205 -3410
rect 18205 -4090 18230 -3410
rect 19710 -4090 19731 -3410
rect 19731 -4090 19805 -3410
rect 19805 -4090 19830 -3410
rect 21310 -4090 21331 -3410
rect 21331 -4090 21405 -3410
rect 21405 -4090 21430 -3410
rect 22910 -4090 22931 -3410
rect 22931 -4090 23005 -3410
rect 23005 -4090 23030 -3410
rect 24510 -4090 24531 -3410
rect 24531 -4090 24605 -3410
rect 24605 -4090 24630 -3410
rect 26110 -4090 26131 -3410
rect 26131 -4090 26205 -3410
rect 26205 -4090 26230 -3410
rect 27710 -4090 27731 -3410
rect 27731 -4090 27805 -3410
rect 27805 -4090 27830 -3410
rect 29310 -4090 29331 -3410
rect 29331 -4090 29405 -3410
rect 29405 -4090 29430 -3410
rect 30910 -4090 30931 -3410
rect 30931 -4090 31005 -3410
rect 31005 -4090 31030 -3410
rect 32510 -4090 32531 -3410
rect 32531 -4090 32605 -3410
rect 32605 -4090 32630 -3410
rect 33400 -3400 33530 -3280
rect 34110 -4090 34131 -3410
rect 34131 -4090 34205 -3410
rect 34205 -4090 34230 -3410
rect 35710 -4090 35731 -3410
rect 35731 -4090 35805 -3410
rect 35805 -4090 35830 -3410
rect 1410 -4370 1530 -4250
rect 3010 -4370 3130 -4250
rect 4610 -4370 4730 -4250
rect 6210 -4370 6330 -4250
rect 7810 -4370 7930 -4250
rect 9410 -4370 9530 -4250
rect 15600 -4370 15700 -4250
rect 17200 -4370 17300 -4250
rect 18800 -4370 18900 -4250
rect 20400 -4370 20500 -4250
rect 22000 -4370 22100 -4250
rect 23600 -4370 23700 -4250
rect 25200 -4370 25300 -4250
rect 26800 -4370 26900 -4250
rect 28400 -4370 28500 -4250
rect 30000 -4370 30100 -4250
rect 33180 -4370 33300 -4250
rect 480 -4664 497 -4530
rect 497 -4664 531 -4530
rect 531 -4664 605 -4530
rect 605 -4664 639 -4530
rect 639 -4664 660 -4530
rect 480 -4780 660 -4664
rect 12390 -4650 12510 -4530
rect 1190 -4840 1310 -4720
rect 2790 -4840 2910 -4720
rect 4390 -4840 4510 -4720
rect 5990 -4840 6110 -4720
rect 7590 -4840 7710 -4720
rect 9190 -4840 9310 -4720
rect 11710 -4930 11830 -4810
rect 12610 -4850 12730 -4730
rect 13630 -4910 13750 -4790
rect 14210 -4850 14330 -4730
rect 15230 -4910 15350 -4790
rect 15820 -4840 15920 -4720
rect 17420 -4840 17520 -4720
rect 19020 -4840 19120 -4720
rect 20620 -4840 20720 -4720
rect 22220 -4840 22320 -4720
rect 23820 -4840 23920 -4720
rect 25420 -4840 25520 -4720
rect 27020 -4840 27120 -4720
rect 28620 -4840 28720 -4720
rect 30220 -4840 30320 -4720
rect 36400 -4830 36500 -4710
rect 11710 -5950 11830 -5830
rect 13310 -5950 13430 -5830
rect 11710 -6170 11830 -6050
rect 13630 -6170 13750 -6050
rect 14230 -6170 14350 -6050
rect 15230 -6170 15350 -6050
rect 12630 -6390 12750 -6270
rect 16510 -6390 16630 -6270
rect 12410 -6610 12530 -6490
rect 14910 -6610 15030 -6490
rect 12950 -6990 13110 -6830
rect 7810 -7990 7930 -7870
rect 14910 -8000 15040 -7880
rect 490 -8257 670 -8090
rect 1210 -8190 1330 -8070
rect 2810 -8190 2930 -8070
rect 4410 -8190 4530 -8070
rect 6010 -8190 6130 -8070
rect 7610 -8190 7730 -8070
rect 9210 -8190 9330 -8070
rect 490 -8375 504 -8257
rect 504 -8375 538 -8257
rect 538 -8375 612 -8257
rect 612 -8375 646 -8257
rect 646 -8375 670 -8257
rect 490 -8796 670 -8375
rect 11710 -8230 11840 -8110
rect 15830 -8190 15950 -8070
rect 17430 -8190 17550 -8070
rect 19030 -8190 19150 -8070
rect 20630 -8190 20750 -8070
rect 22230 -8190 22350 -8070
rect 23830 -8190 23950 -8070
rect 25430 -8190 25550 -8070
rect 27030 -8190 27150 -8070
rect 28630 -8190 28750 -8070
rect 30230 -8190 30350 -8070
rect 31830 -8190 31950 -8070
rect 34810 -8190 34930 -8070
rect 10810 -8380 10930 -8260
rect 16510 -8375 16538 -8260
rect 16538 -8375 16612 -8260
rect 16612 -8375 16640 -8260
rect 16510 -8380 16640 -8375
rect 1430 -8630 1550 -8510
rect 3030 -8630 3150 -8510
rect 4630 -8630 4750 -8510
rect 6230 -8630 6350 -8510
rect 7830 -8630 7950 -8510
rect 9430 -8630 9550 -8510
rect 490 -9488 504 -8796
rect 504 -9488 538 -8796
rect 538 -9488 612 -8796
rect 612 -9488 646 -8796
rect 646 -9488 670 -8796
rect 490 -9688 670 -9488
rect 2130 -9470 2138 -8810
rect 2138 -9470 2212 -8810
rect 2212 -9470 2230 -8810
rect 3730 -9470 3738 -8810
rect 3738 -9470 3812 -8810
rect 3812 -9470 3830 -8810
rect 5330 -9470 5338 -8810
rect 5338 -9470 5412 -8810
rect 5412 -9470 5430 -8810
rect 6930 -9470 6938 -8810
rect 6938 -9470 7012 -8810
rect 7012 -9470 7030 -8810
rect 8530 -9470 8538 -8810
rect 8538 -9470 8612 -8810
rect 8612 -9470 8630 -8810
rect 10130 -9470 10138 -8810
rect 10138 -9470 10212 -8810
rect 10212 -9470 10230 -8810
rect 11720 -9470 11738 -8810
rect 11738 -9470 11812 -8810
rect 11812 -9470 11830 -8810
rect 15610 -8640 15730 -8520
rect 17210 -8640 17330 -8520
rect 18810 -8640 18930 -8520
rect 20410 -8640 20530 -8520
rect 22010 -8640 22130 -8520
rect 23610 -8640 23730 -8520
rect 25210 -8640 25330 -8520
rect 26810 -8640 26930 -8520
rect 28410 -8640 28530 -8520
rect 30010 -8640 30130 -8520
rect 13320 -9470 13338 -8810
rect 13338 -9470 13412 -8810
rect 13412 -9470 13430 -8810
rect 16520 -9480 16538 -8800
rect 16538 -9480 16612 -8800
rect 16612 -9480 16630 -8800
rect 18120 -9480 18138 -8800
rect 18138 -9480 18212 -8800
rect 18212 -9480 18230 -8800
rect 19720 -9480 19738 -8800
rect 19738 -9480 19812 -8800
rect 19812 -9480 19830 -8800
rect 21320 -9480 21338 -8800
rect 21338 -9480 21412 -8800
rect 21412 -9480 21430 -8800
rect 22920 -9480 22938 -8800
rect 22938 -9480 23012 -8800
rect 23012 -9480 23030 -8800
rect 24520 -9480 24538 -8800
rect 24538 -9480 24612 -8800
rect 24612 -9480 24630 -8800
rect 26120 -9480 26138 -8800
rect 26138 -9480 26212 -8800
rect 26212 -9480 26230 -8800
rect 27720 -9480 27738 -8800
rect 27738 -9480 27812 -8800
rect 27812 -9480 27830 -8800
rect 29320 -9480 29338 -8800
rect 29338 -9480 29412 -8800
rect 29412 -9480 29430 -8800
rect 30920 -9480 30938 -8800
rect 30938 -9480 31012 -8800
rect 31012 -9480 31030 -8800
rect 32520 -9360 32538 -8800
rect 32538 -9360 32612 -8800
rect 32612 -9360 32630 -8800
rect 34120 -9360 34138 -8800
rect 34138 -9360 34212 -8800
rect 34212 -9360 34230 -8800
rect 35720 -9360 35738 -8800
rect 35738 -9360 35812 -8800
rect 35812 -9360 35830 -8800
rect 490 -9722 670 -9688
rect 33410 -9630 33530 -9510
rect 490 -10057 670 -9722
rect 1210 -9990 1330 -9870
rect 2810 -9990 2930 -9870
rect 4410 -9990 4530 -9870
rect 6010 -9990 6130 -9870
rect 7610 -9990 7730 -9870
rect 9210 -9990 9330 -9870
rect 15830 -9990 15950 -9870
rect 17430 -9990 17550 -9870
rect 19030 -9990 19150 -9870
rect 20630 -9990 20750 -9870
rect 22230 -9990 22350 -9870
rect 23830 -9990 23950 -9870
rect 25430 -9990 25550 -9870
rect 27030 -9990 27150 -9870
rect 28630 -9990 28750 -9870
rect 30230 -9990 30350 -9870
rect 31830 -9990 31950 -9870
rect 34810 -9990 34930 -9870
rect 490 -10175 504 -10057
rect 504 -10175 538 -10057
rect 538 -10175 612 -10057
rect 612 -10175 646 -10057
rect 646 -10175 670 -10057
rect 490 -10596 670 -10175
rect 10810 -10180 10930 -10060
rect 1430 -10430 1550 -10310
rect 3030 -10430 3150 -10310
rect 4630 -10430 4750 -10310
rect 6230 -10430 6350 -10310
rect 7830 -10430 7950 -10310
rect 9430 -10430 9550 -10310
rect 11030 -10530 11150 -10410
rect 15610 -10440 15730 -10320
rect 17210 -10440 17330 -10320
rect 18810 -10440 18930 -10320
rect 20410 -10440 20530 -10320
rect 22010 -10440 22130 -10320
rect 23610 -10440 23730 -10320
rect 25210 -10440 25330 -10320
rect 26810 -10440 26930 -10320
rect 28410 -10440 28530 -10320
rect 30010 -10440 30130 -10320
rect 31610 -10440 31730 -10320
rect 490 -11288 504 -10596
rect 504 -11288 538 -10596
rect 538 -11288 612 -10596
rect 612 -11288 646 -10596
rect 646 -11288 670 -10596
rect 490 -11488 670 -11288
rect 2130 -11270 2138 -10610
rect 2138 -11270 2212 -10610
rect 2212 -11270 2230 -10610
rect 3730 -11270 3738 -10610
rect 3738 -11270 3812 -10610
rect 3812 -11270 3830 -10610
rect 5330 -11270 5338 -10610
rect 5338 -11270 5412 -10610
rect 5412 -11270 5430 -10610
rect 6930 -11270 6938 -10610
rect 6938 -11270 7012 -10610
rect 7012 -11270 7030 -10610
rect 8530 -11270 8538 -10610
rect 8538 -11270 8612 -10610
rect 8612 -11270 8630 -10610
rect 10130 -11270 10138 -10610
rect 10138 -11270 10212 -10610
rect 10212 -11270 10230 -10610
rect 11720 -11270 11738 -10610
rect 11738 -11270 11812 -10610
rect 11812 -11270 11830 -10610
rect 13320 -11270 13338 -10610
rect 13338 -11270 13412 -10610
rect 13412 -11270 13430 -10610
rect 16520 -11280 16538 -10600
rect 16538 -11280 16612 -10600
rect 16612 -11280 16630 -10600
rect 18120 -11280 18138 -10600
rect 18138 -11280 18212 -10600
rect 18212 -11280 18230 -10600
rect 19720 -11280 19738 -10600
rect 19738 -11280 19812 -10600
rect 19812 -11280 19830 -10600
rect 21320 -11280 21338 -10600
rect 21338 -11280 21412 -10600
rect 21412 -11280 21430 -10600
rect 22920 -11280 22938 -10600
rect 22938 -11280 23012 -10600
rect 23012 -11280 23030 -10600
rect 24520 -11280 24538 -10600
rect 24538 -11280 24612 -10600
rect 24612 -11280 24630 -10600
rect 26120 -11280 26138 -10600
rect 26138 -11280 26212 -10600
rect 26212 -11280 26230 -10600
rect 27720 -11280 27738 -10600
rect 27738 -11280 27812 -10600
rect 27812 -11280 27830 -10600
rect 29320 -11280 29338 -10600
rect 29338 -11280 29412 -10600
rect 29412 -11280 29430 -10600
rect 30920 -11280 30938 -10600
rect 30938 -11280 31012 -10600
rect 31012 -11280 31030 -10600
rect 32520 -11110 32538 -10600
rect 32538 -11110 32612 -10600
rect 32612 -11110 32630 -10600
rect 34120 -11110 34138 -10600
rect 34138 -11110 34212 -10600
rect 34212 -11110 34230 -10600
rect 35720 -11110 35738 -10600
rect 35738 -11110 35812 -10600
rect 35812 -11110 35830 -10600
rect 35010 -11430 35130 -11310
rect 490 -11522 670 -11488
rect 490 -11857 670 -11522
rect 1210 -11790 1330 -11670
rect 2810 -11790 2930 -11670
rect 4410 -11790 4530 -11670
rect 6010 -11790 6130 -11670
rect 7610 -11790 7730 -11670
rect 9210 -11790 9330 -11670
rect 13310 -11790 13430 -11670
rect 14230 -11790 14350 -11670
rect 15830 -11790 15950 -11670
rect 17430 -11790 17550 -11670
rect 19030 -11790 19150 -11670
rect 20630 -11790 20750 -11670
rect 22230 -11790 22350 -11670
rect 23830 -11790 23950 -11670
rect 25430 -11790 25550 -11670
rect 27030 -11790 27150 -11670
rect 28630 -11790 28750 -11670
rect 30230 -11790 30350 -11670
rect 31830 -11790 31950 -11670
rect 34810 -11790 34930 -11670
rect 490 -11975 504 -11857
rect 504 -11975 538 -11857
rect 538 -11975 612 -11857
rect 612 -11975 646 -11857
rect 646 -11975 670 -11857
rect 490 -12396 670 -11975
rect 10810 -11980 10930 -11860
rect 1430 -12230 1550 -12110
rect 3030 -12230 3150 -12110
rect 4630 -12230 4750 -12110
rect 6230 -12230 6350 -12110
rect 7830 -12230 7950 -12110
rect 9430 -12230 9550 -12110
rect 14910 -12230 15040 -12100
rect 15610 -12240 15730 -12120
rect 17210 -12240 17330 -12120
rect 18810 -12240 18930 -12120
rect 20410 -12240 20530 -12120
rect 22010 -12240 22130 -12120
rect 23610 -12240 23730 -12120
rect 25210 -12240 25330 -12120
rect 26810 -12240 26930 -12120
rect 28410 -12240 28530 -12120
rect 30010 -12240 30130 -12120
rect 31610 -12240 31730 -12120
rect 490 -13088 504 -12396
rect 504 -13088 538 -12396
rect 538 -13088 612 -12396
rect 612 -13088 646 -12396
rect 646 -13088 670 -12396
rect 490 -13288 670 -13088
rect 2130 -13070 2138 -12410
rect 2138 -13070 2212 -12410
rect 2212 -13070 2230 -12410
rect 3730 -13070 3738 -12410
rect 3738 -13070 3812 -12410
rect 3812 -13070 3830 -12410
rect 5330 -13070 5338 -12410
rect 5338 -13070 5412 -12410
rect 5412 -13070 5430 -12410
rect 6930 -13070 6938 -12410
rect 6938 -13070 7012 -12410
rect 7012 -13070 7030 -12410
rect 8530 -13070 8538 -12410
rect 8538 -13070 8612 -12410
rect 8612 -13070 8630 -12410
rect 10130 -13070 10138 -12410
rect 10138 -13070 10212 -12410
rect 10212 -13070 10230 -12410
rect 11720 -13070 11738 -12410
rect 11738 -13070 11812 -12410
rect 11812 -13070 11830 -12410
rect 13320 -13070 13338 -12410
rect 13338 -13070 13412 -12410
rect 13412 -13070 13430 -12410
rect 14920 -13070 14938 -12410
rect 14938 -13070 15012 -12410
rect 15012 -13070 15030 -12410
rect 16520 -13080 16538 -12400
rect 16538 -13080 16612 -12400
rect 16612 -13080 16630 -12400
rect 18120 -13080 18138 -12400
rect 18138 -13080 18212 -12400
rect 18212 -13080 18230 -12400
rect 19720 -13080 19738 -12400
rect 19738 -13080 19812 -12400
rect 19812 -13080 19830 -12400
rect 21320 -13080 21338 -12400
rect 21338 -13080 21412 -12400
rect 21412 -13080 21430 -12400
rect 22920 -13080 22938 -12400
rect 22938 -13080 23012 -12400
rect 23012 -13080 23030 -12400
rect 24520 -13080 24538 -12400
rect 24538 -13080 24612 -12400
rect 24612 -13080 24630 -12400
rect 26120 -13080 26138 -12400
rect 26138 -13080 26212 -12400
rect 26212 -13080 26230 -12400
rect 27720 -13080 27738 -12400
rect 27738 -13080 27812 -12400
rect 27812 -13080 27830 -12400
rect 29320 -13080 29338 -12400
rect 29338 -13080 29412 -12400
rect 29412 -13080 29430 -12400
rect 30920 -13080 30938 -12400
rect 30938 -13080 31012 -12400
rect 31012 -13080 31030 -12400
rect 32520 -12910 32538 -12400
rect 32538 -12910 32612 -12400
rect 32612 -12910 32630 -12400
rect 34120 -12910 34138 -12400
rect 34138 -12910 34212 -12400
rect 34212 -12910 34230 -12400
rect 35720 -12910 35738 -12400
rect 35738 -12910 35812 -12400
rect 35812 -12910 35830 -12400
rect 11270 -13154 11650 -13150
rect 11270 -13188 11645 -13154
rect 11645 -13188 11650 -13154
rect 11270 -13210 11650 -13188
rect 490 -13322 670 -13288
rect 35010 -13230 35130 -13110
rect 490 -13657 670 -13322
rect 1210 -13590 1330 -13470
rect 2810 -13590 2930 -13470
rect 4410 -13590 4530 -13470
rect 6010 -13590 6130 -13470
rect 7610 -13590 7730 -13470
rect 9210 -13590 9330 -13470
rect 14010 -13600 14130 -13480
rect 15830 -13590 15950 -13470
rect 17430 -13590 17550 -13470
rect 19030 -13590 19150 -13470
rect 20630 -13590 20750 -13470
rect 22230 -13590 22350 -13470
rect 23830 -13590 23950 -13470
rect 25430 -13590 25550 -13470
rect 27030 -13590 27150 -13470
rect 28630 -13590 28750 -13470
rect 30230 -13590 30350 -13470
rect 31830 -13590 31950 -13470
rect 34810 -13590 34930 -13470
rect 490 -13775 504 -13657
rect 504 -13775 538 -13657
rect 538 -13775 612 -13657
rect 612 -13775 646 -13657
rect 646 -13775 670 -13657
rect 490 -14196 670 -13775
rect 10810 -13780 10930 -13660
rect 1430 -14030 1550 -13910
rect 3030 -14030 3150 -13910
rect 4630 -14030 4750 -13910
rect 6230 -14030 6350 -13910
rect 7830 -14030 7950 -13910
rect 9430 -14030 9550 -13910
rect 11270 -14096 11650 -14060
rect 11270 -14120 11645 -14096
rect 11645 -14120 11650 -14096
rect 15610 -14040 15730 -13920
rect 17210 -14040 17330 -13920
rect 18810 -14040 18930 -13920
rect 20410 -14040 20530 -13920
rect 22010 -14040 22130 -13920
rect 23610 -14040 23730 -13920
rect 25210 -14040 25330 -13920
rect 26810 -14040 26930 -13920
rect 28410 -14040 28530 -13920
rect 30010 -14040 30130 -13920
rect 31610 -14040 31730 -13920
rect 490 -14888 504 -14196
rect 504 -14888 538 -14196
rect 538 -14888 612 -14196
rect 612 -14888 646 -14196
rect 646 -14888 670 -14196
rect 490 -15088 670 -14888
rect 2130 -14870 2138 -14210
rect 2138 -14870 2212 -14210
rect 2212 -14870 2230 -14210
rect 3730 -14870 3738 -14210
rect 3738 -14870 3812 -14210
rect 3812 -14870 3830 -14210
rect 5330 -14870 5338 -14210
rect 5338 -14870 5412 -14210
rect 5412 -14870 5430 -14210
rect 6930 -14870 6938 -14210
rect 6938 -14870 7012 -14210
rect 7012 -14870 7030 -14210
rect 8530 -14870 8538 -14210
rect 8538 -14870 8612 -14210
rect 8612 -14870 8630 -14210
rect 10130 -14870 10138 -14210
rect 10138 -14870 10212 -14210
rect 10212 -14870 10230 -14210
rect 11720 -14870 11738 -14210
rect 11738 -14870 11812 -14210
rect 11812 -14870 11830 -14210
rect 13320 -14870 13338 -14210
rect 13338 -14870 13412 -14210
rect 13412 -14870 13430 -14210
rect 14920 -14870 14938 -14210
rect 14938 -14870 15012 -14210
rect 15012 -14870 15030 -14210
rect 16520 -14880 16538 -14200
rect 16538 -14880 16612 -14200
rect 16612 -14880 16630 -14200
rect 18120 -14880 18138 -14200
rect 18138 -14880 18212 -14200
rect 18212 -14880 18230 -14200
rect 19720 -14880 19738 -14200
rect 19738 -14880 19812 -14200
rect 19812 -14880 19830 -14200
rect 21320 -14880 21338 -14200
rect 21338 -14880 21412 -14200
rect 21412 -14880 21430 -14200
rect 22920 -14880 22938 -14200
rect 22938 -14880 23012 -14200
rect 23012 -14880 23030 -14200
rect 24520 -14880 24538 -14200
rect 24538 -14880 24612 -14200
rect 24612 -14880 24630 -14200
rect 26120 -14880 26138 -14200
rect 26138 -14880 26212 -14200
rect 26212 -14880 26230 -14200
rect 27720 -14880 27738 -14200
rect 27738 -14880 27812 -14200
rect 27812 -14880 27830 -14200
rect 29320 -14880 29338 -14200
rect 29338 -14880 29412 -14200
rect 29412 -14880 29430 -14200
rect 30920 -14880 30938 -14200
rect 30938 -14880 31012 -14200
rect 31012 -14880 31030 -14200
rect 32520 -14710 32538 -14200
rect 32538 -14710 32612 -14200
rect 32612 -14710 32630 -14200
rect 34120 -14710 34138 -14200
rect 34138 -14710 34212 -14200
rect 34212 -14710 34230 -14200
rect 35720 -14710 35738 -14200
rect 35738 -14710 35812 -14200
rect 35812 -14710 35830 -14200
rect 35010 -15030 35130 -14910
rect 490 -15122 670 -15088
rect 490 -15457 670 -15122
rect 1210 -15390 1330 -15270
rect 2810 -15390 2930 -15270
rect 4410 -15390 4530 -15270
rect 6010 -15390 6130 -15270
rect 7610 -15390 7730 -15270
rect 9210 -15390 9330 -15270
rect 13330 -15390 13430 -15290
rect 14020 -15410 14120 -15310
rect 14930 -15390 15030 -15290
rect 15830 -15390 15950 -15270
rect 17430 -15390 17550 -15270
rect 19030 -15390 19150 -15270
rect 20630 -15390 20750 -15270
rect 22230 -15390 22350 -15270
rect 23830 -15390 23950 -15270
rect 27030 -15390 27150 -15270
rect 28630 -15390 28750 -15270
rect 31850 -15400 31970 -15280
rect 490 -15575 504 -15457
rect 504 -15575 538 -15457
rect 538 -15575 612 -15457
rect 612 -15575 646 -15457
rect 646 -15575 670 -15457
rect 490 -15996 670 -15575
rect 10810 -15580 10930 -15460
rect 1430 -15830 1550 -15710
rect 3030 -15830 3150 -15710
rect 4630 -15830 4750 -15710
rect 6230 -15830 6350 -15710
rect 7830 -15830 7950 -15710
rect 9430 -15830 9550 -15710
rect 15610 -15840 15730 -15720
rect 17210 -15840 17330 -15720
rect 18810 -15840 18930 -15720
rect 20410 -15840 20530 -15720
rect 22010 -15840 22130 -15720
rect 23610 -15840 23730 -15720
rect 26810 -15840 26930 -15720
rect 28410 -15840 28530 -15720
rect 31590 -15840 31710 -15720
rect 490 -16688 504 -15996
rect 504 -16688 538 -15996
rect 538 -16688 612 -15996
rect 612 -16688 646 -15996
rect 646 -16688 670 -15996
rect 490 -16888 670 -16688
rect 2130 -16670 2138 -16010
rect 2138 -16670 2212 -16010
rect 2212 -16670 2230 -16010
rect 3730 -16670 3738 -16010
rect 3738 -16670 3812 -16010
rect 3812 -16670 3830 -16010
rect 5330 -16670 5338 -16010
rect 5338 -16670 5412 -16010
rect 5412 -16670 5430 -16010
rect 6930 -16670 6938 -16010
rect 6938 -16670 7012 -16010
rect 7012 -16670 7030 -16010
rect 8530 -16670 8538 -16010
rect 8538 -16670 8612 -16010
rect 8612 -16670 8630 -16010
rect 10130 -16670 10138 -16010
rect 10138 -16670 10212 -16010
rect 10212 -16670 10230 -16010
rect 13320 -16670 13338 -16010
rect 13338 -16670 13412 -16010
rect 13412 -16670 13430 -16010
rect 14920 -16670 14938 -16010
rect 14938 -16670 15012 -16010
rect 15012 -16670 15030 -16010
rect 16520 -16680 16538 -16000
rect 16538 -16680 16612 -16000
rect 16612 -16680 16630 -16000
rect 18120 -16680 18138 -16000
rect 18138 -16680 18212 -16000
rect 18212 -16680 18230 -16000
rect 19720 -16680 19738 -16000
rect 19738 -16680 19812 -16000
rect 19812 -16680 19830 -16000
rect 21320 -16680 21338 -16000
rect 21338 -16680 21412 -16000
rect 21412 -16680 21430 -16000
rect 22920 -16680 22938 -16000
rect 22938 -16680 23012 -16000
rect 23012 -16680 23030 -16000
rect 24520 -16680 24538 -16000
rect 24538 -16680 24612 -16000
rect 24612 -16680 24630 -16000
rect 26120 -16680 26138 -16000
rect 26138 -16680 26212 -16000
rect 26212 -16680 26230 -16000
rect 27720 -16680 27738 -16000
rect 27738 -16680 27812 -16000
rect 27812 -16680 27830 -16000
rect 29320 -16680 29338 -16000
rect 29338 -16680 29412 -16000
rect 29412 -16680 29430 -16000
rect 30920 -16680 30938 -16000
rect 30938 -16680 31012 -16000
rect 31012 -16680 31030 -16000
rect 32520 -16680 32538 -16000
rect 32538 -16680 32612 -16000
rect 32612 -16680 32630 -16000
rect 34120 -16680 34138 -16000
rect 34138 -16680 34212 -16000
rect 34212 -16680 34230 -16000
rect 35720 -16680 35738 -16000
rect 35738 -16680 35812 -16000
rect 35812 -16680 35830 -16000
rect 490 -16922 670 -16888
rect 490 -17257 670 -16922
rect 1210 -17190 1330 -17070
rect 2810 -17190 2930 -17070
rect 4410 -17190 4530 -17070
rect 6010 -17190 6130 -17070
rect 7610 -17190 7730 -17070
rect 9210 -17190 9330 -17070
rect 12630 -17200 12750 -17080
rect 15830 -17190 15950 -17070
rect 17430 -17190 17550 -17070
rect 19030 -17190 19150 -17070
rect 20630 -17190 20750 -17070
rect 22230 -17190 22350 -17070
rect 23830 -17190 23950 -17070
rect 27030 -17190 27150 -17070
rect 28630 -17190 28750 -17070
rect 31850 -17200 31970 -17080
rect 490 -17375 504 -17257
rect 504 -17375 538 -17257
rect 538 -17375 612 -17257
rect 612 -17375 646 -17257
rect 646 -17375 670 -17257
rect 490 -17796 670 -17375
rect 10810 -17380 10930 -17260
rect 1430 -17630 1550 -17510
rect 3030 -17630 3150 -17510
rect 4630 -17630 4750 -17510
rect 6230 -17630 6350 -17510
rect 7830 -17630 7950 -17510
rect 9430 -17630 9550 -17510
rect 15610 -17640 15730 -17520
rect 17210 -17640 17330 -17520
rect 18810 -17640 18930 -17520
rect 20410 -17640 20530 -17520
rect 22010 -17640 22130 -17520
rect 23610 -17640 23730 -17520
rect 26810 -17640 26930 -17520
rect 28410 -17640 28530 -17520
rect 31590 -17640 31710 -17520
rect 490 -18488 504 -17796
rect 504 -18488 538 -17796
rect 538 -18488 612 -17796
rect 612 -18488 646 -17796
rect 646 -18488 670 -17796
rect 490 -18688 670 -18488
rect 2130 -18470 2138 -17810
rect 2138 -18470 2212 -17810
rect 2212 -18470 2230 -17810
rect 3730 -18470 3738 -17810
rect 3738 -18470 3812 -17810
rect 3812 -18470 3830 -17810
rect 5330 -18470 5338 -17810
rect 5338 -18470 5412 -17810
rect 5412 -18470 5430 -17810
rect 6930 -18470 6938 -17810
rect 6938 -18470 7012 -17810
rect 7012 -18470 7030 -17810
rect 8530 -18470 8538 -17810
rect 8538 -18470 8612 -17810
rect 8612 -18470 8630 -17810
rect 10130 -18470 10138 -17810
rect 10138 -18470 10212 -17810
rect 10212 -18470 10230 -17810
rect 13320 -18470 13338 -17810
rect 13338 -18470 13412 -17810
rect 13412 -18470 13430 -17810
rect 14920 -18470 14938 -17810
rect 14938 -18470 15012 -17810
rect 15012 -18470 15030 -17810
rect 16520 -18480 16538 -17800
rect 16538 -18480 16612 -17800
rect 16612 -18480 16630 -17800
rect 18120 -18480 18138 -17800
rect 18138 -18480 18212 -17800
rect 18212 -18480 18230 -17800
rect 19720 -18480 19738 -17800
rect 19738 -18480 19812 -17800
rect 19812 -18480 19830 -17800
rect 21320 -18480 21338 -17800
rect 21338 -18480 21412 -17800
rect 21412 -18480 21430 -17800
rect 22920 -18480 22938 -17800
rect 22938 -18480 23012 -17800
rect 23012 -18480 23030 -17800
rect 24520 -18480 24538 -17800
rect 24538 -18480 24612 -17800
rect 24612 -18480 24630 -17800
rect 26120 -18480 26138 -17800
rect 26138 -18480 26212 -17800
rect 26212 -18480 26230 -17800
rect 27720 -18480 27738 -17800
rect 27738 -18480 27812 -17800
rect 27812 -18480 27830 -17800
rect 29320 -18480 29338 -17800
rect 29338 -18480 29412 -17800
rect 29412 -18480 29430 -17800
rect 30920 -18480 30938 -17800
rect 30938 -18480 31012 -17800
rect 31012 -18480 31030 -17800
rect 32520 -18480 32538 -17800
rect 32538 -18480 32612 -17800
rect 32612 -18480 32630 -17800
rect 34120 -18480 34138 -17800
rect 34138 -18480 34212 -17800
rect 34212 -18480 34230 -17800
rect 35720 -18480 35738 -17800
rect 35738 -18480 35812 -17800
rect 35812 -18480 35830 -17800
rect 490 -18722 670 -18688
rect 490 -19057 670 -18722
rect 1210 -18990 1330 -18870
rect 2810 -18990 2930 -18870
rect 4410 -18990 4530 -18870
rect 6010 -18990 6130 -18870
rect 7610 -18990 7730 -18870
rect 9210 -18990 9330 -18870
rect 12410 -19000 12530 -18880
rect 15830 -18990 15950 -18870
rect 17430 -18990 17550 -18870
rect 19030 -18990 19150 -18870
rect 20630 -18990 20750 -18870
rect 22230 -18990 22350 -18870
rect 23830 -18990 23950 -18870
rect 27030 -18990 27150 -18870
rect 28630 -18990 28750 -18870
rect 31590 -19000 31710 -18880
rect 490 -19175 504 -19057
rect 504 -19175 538 -19057
rect 538 -19175 612 -19057
rect 612 -19175 646 -19057
rect 646 -19175 670 -19057
rect 490 -19596 670 -19175
rect 10810 -19180 10930 -19060
rect 1430 -19430 1550 -19310
rect 3030 -19430 3150 -19310
rect 4630 -19430 4750 -19310
rect 6230 -19430 6350 -19310
rect 7830 -19430 7950 -19310
rect 9430 -19430 9550 -19310
rect 15610 -19440 15730 -19320
rect 17210 -19440 17330 -19320
rect 18810 -19440 18930 -19320
rect 20410 -19440 20530 -19320
rect 22010 -19440 22130 -19320
rect 23610 -19440 23730 -19320
rect 26810 -19440 26930 -19320
rect 28410 -19440 28530 -19320
rect 31750 -19520 31810 -19240
rect 490 -20288 504 -19596
rect 504 -20288 538 -19596
rect 538 -20288 612 -19596
rect 612 -20288 646 -19596
rect 646 -20288 670 -19596
rect 490 -20488 670 -20288
rect 2130 -20270 2138 -19610
rect 2138 -20270 2212 -19610
rect 2212 -20270 2230 -19610
rect 3730 -20270 3738 -19610
rect 3738 -20270 3812 -19610
rect 3812 -20270 3830 -19610
rect 5330 -20270 5338 -19610
rect 5338 -20270 5412 -19610
rect 5412 -20270 5430 -19610
rect 6930 -20270 6938 -19610
rect 6938 -20270 7012 -19610
rect 7012 -20270 7030 -19610
rect 8530 -20270 8538 -19610
rect 8538 -20270 8612 -19610
rect 8612 -20270 8630 -19610
rect 10130 -20270 10138 -19610
rect 10138 -20270 10212 -19610
rect 10212 -20270 10230 -19610
rect 13320 -20270 13338 -19610
rect 13338 -20270 13412 -19610
rect 13412 -20270 13430 -19610
rect 14920 -20270 14938 -19610
rect 14938 -20270 15012 -19610
rect 15012 -20270 15030 -19610
rect 16520 -20280 16538 -19600
rect 16538 -20280 16612 -19600
rect 16612 -20280 16630 -19600
rect 18120 -20280 18138 -19600
rect 18138 -20280 18212 -19600
rect 18212 -20280 18230 -19600
rect 19720 -20280 19738 -19600
rect 19738 -20280 19812 -19600
rect 19812 -20280 19830 -19600
rect 21320 -20280 21338 -19600
rect 21338 -20280 21412 -19600
rect 21412 -20280 21430 -19600
rect 22920 -20280 22938 -19600
rect 22938 -20280 23012 -19600
rect 23012 -20280 23030 -19600
rect 24520 -20280 24538 -19600
rect 24538 -20280 24612 -19600
rect 24612 -20280 24630 -19600
rect 26120 -20280 26138 -19600
rect 26138 -20280 26212 -19600
rect 26212 -20280 26230 -19600
rect 27720 -20280 27738 -19600
rect 27738 -20280 27812 -19600
rect 27812 -20280 27830 -19600
rect 29320 -20280 29338 -19600
rect 29338 -20280 29412 -19600
rect 29412 -20280 29430 -19600
rect 30920 -20280 30938 -19600
rect 30938 -20280 31012 -19600
rect 31012 -20280 31030 -19600
rect 32520 -20280 32538 -19600
rect 32538 -20280 32612 -19600
rect 32612 -20280 32630 -19600
rect 34120 -20280 34138 -19600
rect 34138 -20280 34212 -19600
rect 34212 -20280 34230 -19600
rect 35720 -20280 35738 -19600
rect 35738 -20280 35812 -19600
rect 35812 -20280 35830 -19600
rect 33190 -20460 33310 -20340
rect 490 -20522 670 -20488
rect 490 -20857 670 -20522
rect 1210 -20790 1330 -20670
rect 2810 -20790 2930 -20670
rect 4410 -20790 4530 -20670
rect 6010 -20790 6130 -20670
rect 7610 -20790 7730 -20670
rect 9210 -20790 9330 -20670
rect 12410 -20800 12530 -20680
rect 15830 -20790 15950 -20670
rect 17430 -20790 17550 -20670
rect 19030 -20790 19150 -20670
rect 20630 -20790 20750 -20670
rect 22230 -20790 22350 -20670
rect 23830 -20790 23950 -20670
rect 27030 -20790 27150 -20670
rect 28630 -20790 28750 -20670
rect 31590 -20800 31710 -20680
rect 490 -20975 504 -20857
rect 504 -20975 538 -20857
rect 538 -20975 612 -20857
rect 612 -20975 646 -20857
rect 646 -20975 670 -20857
rect 490 -21396 670 -20975
rect 10810 -20980 10930 -20860
rect 1430 -21230 1550 -21110
rect 3030 -21230 3150 -21110
rect 4630 -21230 4750 -21110
rect 6230 -21230 6350 -21110
rect 7830 -21230 7950 -21110
rect 9430 -21230 9550 -21110
rect 15610 -21240 15730 -21120
rect 17210 -21240 17330 -21120
rect 18810 -21240 18930 -21120
rect 20410 -21240 20530 -21120
rect 22010 -21240 22130 -21120
rect 23610 -21240 23730 -21120
rect 26810 -21240 26930 -21120
rect 28410 -21240 28530 -21120
rect 31750 -21320 31810 -21040
rect 490 -22088 504 -21396
rect 504 -22088 538 -21396
rect 538 -22088 612 -21396
rect 612 -22088 646 -21396
rect 646 -22088 670 -21396
rect 490 -22288 670 -22088
rect 2130 -22070 2138 -21410
rect 2138 -22070 2212 -21410
rect 2212 -22070 2230 -21410
rect 3730 -22070 3738 -21410
rect 3738 -22070 3812 -21410
rect 3812 -22070 3830 -21410
rect 5330 -22070 5338 -21410
rect 5338 -22070 5412 -21410
rect 5412 -22070 5430 -21410
rect 6930 -22070 6938 -21410
rect 6938 -22070 7012 -21410
rect 7012 -22070 7030 -21410
rect 8530 -22070 8538 -21410
rect 8538 -22070 8612 -21410
rect 8612 -22070 8630 -21410
rect 10130 -22070 10138 -21410
rect 10138 -22070 10212 -21410
rect 10212 -22070 10230 -21410
rect 11710 -22080 11738 -21400
rect 11738 -22080 11812 -21400
rect 11812 -22080 11840 -21400
rect 16520 -22080 16538 -21400
rect 16538 -22080 16612 -21400
rect 16612 -22080 16630 -21400
rect 18120 -22080 18138 -21400
rect 18138 -22080 18212 -21400
rect 18212 -22080 18230 -21400
rect 19720 -22080 19738 -21400
rect 19738 -22080 19812 -21400
rect 19812 -22080 19830 -21400
rect 21320 -22080 21338 -21400
rect 21338 -22080 21412 -21400
rect 21412 -22080 21430 -21400
rect 22920 -22080 22938 -21400
rect 22938 -22080 23012 -21400
rect 23012 -22080 23030 -21400
rect 24520 -22080 24538 -21400
rect 24538 -22080 24612 -21400
rect 24612 -22080 24630 -21400
rect 26120 -22080 26138 -21400
rect 26138 -22080 26212 -21400
rect 26212 -22080 26230 -21400
rect 27720 -22080 27738 -21400
rect 27738 -22080 27812 -21400
rect 27812 -22080 27830 -21400
rect 29320 -22080 29338 -21400
rect 29338 -22080 29412 -21400
rect 29412 -22080 29430 -21400
rect 30920 -22080 30938 -21400
rect 30938 -22080 31012 -21400
rect 31012 -22080 31030 -21400
rect 32520 -22080 32538 -21400
rect 32538 -22080 32612 -21400
rect 32612 -22080 32630 -21400
rect 34120 -22080 34138 -21400
rect 34138 -22080 34212 -21400
rect 34212 -22080 34230 -21400
rect 35720 -22080 35738 -21400
rect 35738 -22080 35812 -21400
rect 35812 -22080 35830 -21400
rect 33210 -22240 33290 -22140
rect 34020 -22188 34045 -22170
rect 34045 -22188 34305 -22170
rect 34305 -22188 34360 -22170
rect 34020 -22240 34360 -22188
rect 490 -22322 670 -22288
rect 490 -22380 670 -22322
rect 28150 -22870 28352 -22730
rect 28352 -22870 28370 -22730
rect 28630 -22870 28668 -22740
rect 28668 -22870 28702 -22740
rect 28702 -22870 28740 -22740
rect 29000 -22870 29018 -22730
rect 29018 -22870 29220 -22730
rect 32630 -22490 33300 -22430
rect 34040 -22490 34310 -22430
rect 32700 -23104 32711 -23070
rect 32711 -23104 32745 -23070
rect 32745 -23104 32869 -23070
rect 32869 -23104 32903 -23070
rect 32903 -23104 32910 -23070
rect 32700 -23150 32910 -23104
rect 33020 -23104 33027 -23070
rect 33027 -23104 33061 -23070
rect 33061 -23104 33185 -23070
rect 33185 -23104 33219 -23070
rect 33219 -23104 33230 -23070
rect 33020 -23150 33230 -23104
rect 34070 -23124 34081 -23100
rect 34081 -23124 34115 -23100
rect 34115 -23124 34239 -23100
rect 34239 -23124 34273 -23100
rect 34273 -23124 34300 -23100
rect 34070 -23160 34300 -23124
rect 29750 -23590 29880 -23520
rect 33410 -23620 33910 -23560
rect 35000 -23620 37020 -23560
rect 33170 -24246 33249 -24220
rect 33249 -24246 33280 -24220
rect 33170 -24280 33280 -24246
rect 33410 -24246 33441 -24220
rect 33441 -24246 33565 -24220
rect 33565 -24246 33599 -24220
rect 33599 -24246 33600 -24220
rect 33410 -24280 33600 -24246
rect 33730 -24246 33757 -24220
rect 33757 -24246 33881 -24220
rect 33881 -24246 33915 -24220
rect 33915 -24246 33920 -24220
rect 33730 -24280 33920 -24246
rect 34040 -24246 34073 -24220
rect 34073 -24246 34140 -24220
rect 34040 -24280 34140 -24246
rect 34620 -24244 34621 -24220
rect 34621 -24244 34655 -24220
rect 34655 -24244 34770 -24220
rect 34620 -24280 34770 -24244
rect 34990 -24244 35095 -24220
rect 35095 -24244 35129 -24220
rect 35129 -24244 35130 -24220
rect 34990 -24280 35130 -24244
rect 35260 -24244 35287 -24220
rect 35287 -24244 35411 -24220
rect 35411 -24244 35445 -24220
rect 35445 -24244 35450 -24220
rect 35260 -24280 35450 -24244
rect 35570 -24244 35603 -24220
rect 35603 -24244 35727 -24220
rect 35727 -24244 35760 -24220
rect 35570 -24280 35760 -24244
rect 35890 -24244 35919 -24220
rect 35919 -24244 36043 -24220
rect 36043 -24244 36077 -24220
rect 36077 -24244 36080 -24220
rect 35890 -24280 36080 -24244
rect 36200 -24244 36201 -24220
rect 36201 -24244 36235 -24220
rect 36235 -24244 36359 -24220
rect 36359 -24244 36390 -24220
rect 36200 -24280 36390 -24244
rect 36520 -24244 36551 -24220
rect 36551 -24244 36675 -24220
rect 36675 -24244 36709 -24220
rect 36709 -24244 36710 -24220
rect 36520 -24280 36710 -24244
rect 36830 -24244 36833 -24220
rect 36833 -24244 36867 -24220
rect 36867 -24244 36991 -24220
rect 36991 -24244 37020 -24220
rect 36830 -24280 37020 -24244
rect 2510 -25106 4010 -25070
rect 2510 -25130 4010 -25106
rect 4710 -25106 6210 -25070
rect 4710 -25130 6210 -25106
rect 6910 -25106 8410 -25070
rect 6910 -25130 8410 -25106
rect 9110 -25106 10610 -25070
rect 9110 -25130 10610 -25106
rect 11310 -25106 12810 -25070
rect 11310 -25130 12810 -25106
rect 13510 -25106 15010 -25070
rect 13510 -25130 15010 -25106
rect 15710 -25106 17210 -25070
rect 15710 -25130 17210 -25106
rect 17910 -25106 19410 -25070
rect 17910 -25130 19410 -25106
rect 2240 -25320 2300 -25260
rect 4440 -25230 4500 -25170
rect 4440 -25340 4500 -25280
rect 6640 -25230 6700 -25170
rect 6420 -25340 6480 -25280
rect 8620 -25230 8680 -25170
rect 8620 -25340 8680 -25280
rect 10820 -25230 10880 -25170
rect 10820 -25340 10880 -25280
rect 13020 -25230 13080 -25170
rect 13020 -25340 13080 -25280
rect 15220 -25230 15280 -25170
rect 15440 -25340 15500 -25280
rect 17640 -25230 17700 -25170
rect 17640 -25340 17700 -25280
rect 19840 -25230 19900 -25170
rect 2510 -25760 2690 -25700
rect 3170 -25760 3350 -25700
rect 3830 -25760 4010 -25700
rect 4710 -25760 4890 -25700
rect 5370 -25760 5550 -25700
rect 6030 -25760 6210 -25700
rect 6910 -25620 7090 -25560
rect 7570 -25620 7750 -25560
rect 8230 -25620 8410 -25560
rect 9110 -25620 9290 -25560
rect 9770 -25620 9950 -25560
rect 10430 -25620 10610 -25560
rect 11310 -25620 11490 -25560
rect 11970 -25620 12150 -25560
rect 12630 -25620 12810 -25560
rect 13510 -25620 13690 -25560
rect 14170 -25620 14350 -25560
rect 14830 -25620 15010 -25560
rect 15710 -25760 15890 -25700
rect 16370 -25760 16550 -25700
rect 17030 -25760 17210 -25700
rect 17910 -25760 18090 -25700
rect 18570 -25760 18750 -25700
rect 19230 -25760 19410 -25700
rect 2510 -25906 4010 -25870
rect 2510 -25930 4010 -25906
rect 4710 -25906 6210 -25870
rect 4710 -25930 6210 -25906
rect 6910 -25906 8410 -25870
rect 6910 -25930 8410 -25906
rect 9110 -25906 10610 -25870
rect 9110 -25930 10610 -25906
rect 11310 -25906 12810 -25870
rect 11310 -25930 12810 -25906
rect 13510 -25906 15010 -25870
rect 13510 -25930 15010 -25906
rect 15710 -25906 17210 -25870
rect 15710 -25930 17210 -25906
rect 17910 -25906 19410 -25870
rect 17910 -25930 19410 -25906
rect 2020 -26120 2080 -26060
rect 4220 -26030 4280 -25970
rect 4220 -26140 4280 -26080
rect 6420 -26030 6480 -25970
rect 6640 -26140 6700 -26080
rect 8840 -26030 8900 -25970
rect 8840 -26140 8900 -26080
rect 11040 -26030 11100 -25970
rect 11040 -26140 11100 -26080
rect 13240 -26030 13300 -25970
rect 13240 -26140 13300 -26080
rect 15440 -26030 15500 -25970
rect 15220 -26140 15280 -26080
rect 17420 -26030 17480 -25970
rect 17420 -26140 17480 -26080
rect 19620 -26030 19680 -25970
rect 2510 -26420 2690 -26360
rect 3170 -26420 3350 -26360
rect 3830 -26420 4010 -26360
rect 4710 -26420 4890 -26360
rect 5370 -26420 5550 -26360
rect 6030 -26420 6210 -26360
rect 6910 -26560 7090 -26500
rect 7570 -26560 7750 -26500
rect 8230 -26560 8410 -26500
rect 9110 -26560 9290 -26500
rect 9770 -26560 9950 -26500
rect 10430 -26560 10610 -26500
rect 11310 -26560 11490 -26500
rect 11970 -26560 12150 -26500
rect 12630 -26560 12810 -26500
rect 13510 -26560 13690 -26500
rect 14170 -26560 14350 -26500
rect 14830 -26560 15010 -26500
rect 15710 -26420 15890 -26360
rect 16370 -26420 16550 -26360
rect 17030 -26420 17210 -26360
rect 17910 -26420 18090 -26360
rect 18570 -26420 18750 -26360
rect 19230 -26420 19410 -26360
rect 430 -26710 610 -26630
rect 4710 -26706 6210 -26670
rect 4710 -26730 6210 -26706
rect 6910 -26706 8410 -26670
rect 6910 -26730 8410 -26706
rect 9110 -26706 10610 -26670
rect 9110 -26730 10610 -26706
rect 11310 -26706 12810 -26670
rect 11310 -26730 12810 -26706
rect 13510 -26706 15010 -26670
rect 13510 -26730 15010 -26706
rect 15710 -26706 17210 -26670
rect 15710 -26730 17210 -26706
rect 21310 -26710 21490 -26630
rect 1420 -27020 1480 -26870
rect 4440 -26940 4500 -26880
rect 6640 -26830 6700 -26770
rect 6420 -26940 6480 -26880
rect 8620 -26830 8680 -26770
rect 8620 -26940 8680 -26880
rect 10820 -26830 10880 -26770
rect 10820 -26940 10880 -26880
rect 13020 -26830 13080 -26770
rect 13020 -26940 13080 -26880
rect 15220 -26830 15280 -26770
rect 15440 -26940 15500 -26880
rect 17640 -26830 17700 -26770
rect 20240 -26930 20300 -26780
rect 2510 -27360 2690 -27300
rect 3170 -27360 3350 -27300
rect 3830 -27360 4010 -27300
rect 4710 -27360 4890 -27300
rect 5370 -27360 5550 -27300
rect 6030 -27360 6210 -27300
rect 6910 -27220 7090 -27160
rect 7570 -27220 7750 -27160
rect 8230 -27220 8410 -27160
rect 9110 -27220 9290 -27160
rect 9770 -27220 9950 -27160
rect 10430 -27220 10610 -27160
rect 11310 -27220 11490 -27160
rect 11970 -27220 12150 -27160
rect 12630 -27220 12810 -27160
rect 13510 -27220 13690 -27160
rect 14170 -27220 14350 -27160
rect 14830 -27220 15010 -27160
rect 15710 -27360 15890 -27300
rect 16370 -27360 16550 -27300
rect 17030 -27360 17210 -27300
rect 17910 -27360 18090 -27300
rect 18570 -27360 18750 -27300
rect 19230 -27360 19410 -27300
rect 430 -27510 610 -27430
rect 4710 -27506 6210 -27470
rect 4710 -27530 6210 -27506
rect 6910 -27506 8410 -27470
rect 6910 -27530 8410 -27506
rect 9110 -27506 10610 -27470
rect 9110 -27530 10610 -27506
rect 11310 -27506 12810 -27470
rect 11310 -27530 12810 -27506
rect 13510 -27506 15010 -27470
rect 13510 -27530 15010 -27506
rect 15710 -27506 17210 -27470
rect 15710 -27530 17210 -27506
rect 21310 -27510 21490 -27430
rect 1620 -27820 1680 -27670
rect 4220 -27740 4280 -27680
rect 6420 -27630 6480 -27570
rect 6640 -27740 6700 -27680
rect 8840 -27630 8900 -27570
rect 8840 -27740 8900 -27680
rect 11040 -27630 11100 -27570
rect 11040 -27740 11100 -27680
rect 13240 -27630 13300 -27570
rect 13240 -27740 13300 -27680
rect 15440 -27630 15500 -27570
rect 15220 -27740 15280 -27680
rect 17420 -27630 17480 -27570
rect 20440 -27730 20500 -27580
rect 2510 -28020 2690 -27960
rect 3170 -28020 3350 -27960
rect 3830 -28020 4010 -27960
rect 4710 -28020 4890 -27960
rect 5370 -28020 5550 -27960
rect 6030 -28020 6210 -27960
rect 6910 -28160 7090 -28100
rect 7570 -28160 7750 -28100
rect 8230 -28160 8410 -28100
rect 9110 -28160 9290 -28100
rect 9770 -28160 9950 -28100
rect 10430 -28160 10610 -28100
rect 11310 -28160 11490 -28100
rect 11970 -28160 12150 -28100
rect 12630 -28160 12810 -28100
rect 13510 -28160 13690 -28100
rect 14170 -28160 14350 -28100
rect 14830 -28160 15010 -28100
rect 15710 -28020 15890 -27960
rect 16370 -28020 16550 -27960
rect 17030 -28020 17210 -27960
rect 17910 -28020 18090 -27960
rect 18570 -28020 18750 -27960
rect 19230 -28020 19410 -27960
rect 430 -28310 610 -28230
rect 4710 -28306 6210 -28270
rect 4710 -28330 6210 -28306
rect 6910 -28306 8410 -28270
rect 6910 -28330 8410 -28306
rect 9110 -28306 10610 -28270
rect 9110 -28330 10610 -28306
rect 11310 -28306 12810 -28270
rect 11310 -28330 12810 -28306
rect 13510 -28306 15010 -28270
rect 13510 -28330 15010 -28306
rect 15710 -28306 17210 -28270
rect 15710 -28330 17210 -28306
rect 21310 -28310 21490 -28230
rect 1620 -28620 1680 -28470
rect 4220 -28540 4280 -28480
rect 6420 -28430 6480 -28370
rect 6640 -28540 6700 -28480
rect 8840 -28430 8900 -28370
rect 8840 -28540 8900 -28480
rect 11040 -28430 11100 -28370
rect 11040 -28540 11100 -28480
rect 13240 -28430 13300 -28370
rect 13240 -28540 13300 -28480
rect 15440 -28430 15500 -28370
rect 15220 -28540 15280 -28480
rect 17420 -28430 17480 -28370
rect 20440 -28530 20500 -28380
rect 2510 -28820 2690 -28760
rect 3170 -28820 3350 -28760
rect 3830 -28820 4010 -28760
rect 4710 -28820 4890 -28760
rect 5370 -28820 5550 -28760
rect 6030 -28820 6210 -28760
rect 6910 -28960 7090 -28900
rect 7570 -28960 7750 -28900
rect 8230 -28960 8410 -28900
rect 9110 -28960 9290 -28900
rect 9770 -28960 9950 -28900
rect 10430 -28960 10610 -28900
rect 11310 -28960 11490 -28900
rect 11970 -28960 12150 -28900
rect 12630 -28960 12810 -28900
rect 13510 -28960 13690 -28900
rect 14170 -28960 14350 -28900
rect 14830 -28960 15010 -28900
rect 15710 -28820 15890 -28760
rect 16370 -28820 16550 -28760
rect 17030 -28820 17210 -28760
rect 17910 -28820 18090 -28760
rect 18570 -28820 18750 -28760
rect 19230 -28820 19410 -28760
rect 430 -29110 610 -29030
rect 4710 -29106 6210 -29070
rect 4710 -29130 6210 -29106
rect 6910 -29106 8410 -29070
rect 6910 -29130 8410 -29106
rect 9110 -29106 10610 -29070
rect 9110 -29130 10610 -29106
rect 11310 -29106 12810 -29070
rect 11310 -29130 12810 -29106
rect 13510 -29106 15010 -29070
rect 13510 -29130 15010 -29106
rect 15710 -29106 17210 -29070
rect 15710 -29130 17210 -29106
rect 21310 -29110 21490 -29030
rect 1420 -29420 1480 -29270
rect 4440 -29340 4500 -29280
rect 6640 -29230 6700 -29170
rect 6420 -29340 6480 -29280
rect 8620 -29230 8680 -29170
rect 8620 -29340 8680 -29280
rect 10820 -29230 10880 -29170
rect 10820 -29340 10880 -29280
rect 13020 -29230 13080 -29170
rect 13020 -29340 13080 -29280
rect 15220 -29230 15280 -29170
rect 15440 -29340 15500 -29280
rect 17640 -29230 17700 -29170
rect 20240 -29330 20300 -29180
rect 2510 -29760 2690 -29700
rect 3170 -29760 3350 -29700
rect 3830 -29760 4010 -29700
rect 4710 -29760 4890 -29700
rect 5370 -29760 5550 -29700
rect 6030 -29760 6210 -29700
rect 6910 -29620 7090 -29560
rect 7570 -29620 7750 -29560
rect 8230 -29620 8410 -29560
rect 9110 -29620 9290 -29560
rect 9770 -29620 9950 -29560
rect 10430 -29620 10610 -29560
rect 11310 -29620 11490 -29560
rect 11970 -29620 12150 -29560
rect 12630 -29620 12810 -29560
rect 13510 -29620 13690 -29560
rect 14170 -29620 14350 -29560
rect 14830 -29620 15010 -29560
rect 15710 -29760 15890 -29700
rect 16370 -29760 16550 -29700
rect 17030 -29760 17210 -29700
rect 17910 -29760 18090 -29700
rect 18570 -29760 18750 -29700
rect 19230 -29760 19410 -29700
rect 2510 -29906 4010 -29870
rect 2510 -29930 4010 -29906
rect 4710 -29906 6210 -29870
rect 4710 -29930 6210 -29906
rect 6910 -29906 8410 -29870
rect 6910 -29930 8410 -29906
rect 9110 -29906 10610 -29870
rect 9110 -29930 10610 -29906
rect 11310 -29906 12810 -29870
rect 11310 -29930 12810 -29906
rect 13510 -29906 15010 -29870
rect 13510 -29930 15010 -29906
rect 15710 -29906 17210 -29870
rect 15710 -29930 17210 -29906
rect 17910 -29906 19410 -29870
rect 17910 -29930 19410 -29906
rect 2020 -30120 2080 -30060
rect 4220 -30030 4280 -29970
rect 4220 -30140 4280 -30080
rect 6420 -30030 6480 -29970
rect 6640 -30140 6700 -30080
rect 8840 -30030 8900 -29970
rect 8840 -30140 8900 -30080
rect 11040 -30030 11100 -29970
rect 11040 -30140 11100 -30080
rect 13240 -30030 13300 -29970
rect 13240 -30140 13300 -30080
rect 15440 -30030 15500 -29970
rect 15220 -30140 15280 -30080
rect 17420 -30030 17480 -29970
rect 17420 -30140 17480 -30080
rect 19620 -30030 19680 -29970
rect 2510 -30420 2690 -30360
rect 3170 -30420 3350 -30360
rect 3830 -30420 4010 -30360
rect 4710 -30420 4890 -30360
rect 5370 -30420 5550 -30360
rect 6030 -30420 6210 -30360
rect 6910 -30560 7090 -30500
rect 7570 -30560 7750 -30500
rect 8230 -30560 8410 -30500
rect 9110 -30560 9290 -30500
rect 9770 -30560 9950 -30500
rect 10430 -30560 10610 -30500
rect 11310 -30560 11490 -30500
rect 11970 -30560 12150 -30500
rect 12630 -30560 12810 -30500
rect 13510 -30560 13690 -30500
rect 14170 -30560 14350 -30500
rect 14830 -30560 15010 -30500
rect 15710 -30420 15890 -30360
rect 16370 -30420 16550 -30360
rect 17030 -30420 17210 -30360
rect 17910 -30420 18090 -30360
rect 18570 -30420 18750 -30360
rect 19230 -30420 19410 -30360
rect 2510 -30706 4010 -30670
rect 2510 -30730 4010 -30706
rect 4710 -30706 6210 -30670
rect 4710 -30730 6210 -30706
rect 6910 -30706 8410 -30670
rect 6910 -30730 8410 -30706
rect 9110 -30706 10610 -30670
rect 9110 -30730 10610 -30706
rect 11310 -30706 12810 -30670
rect 11310 -30730 12810 -30706
rect 13510 -30706 15010 -30670
rect 13510 -30730 15010 -30706
rect 15710 -30706 17210 -30670
rect 15710 -30730 17210 -30706
rect 17910 -30706 19410 -30670
rect 17910 -30730 19410 -30706
rect 2240 -30920 2300 -30860
rect 4440 -30830 4500 -30770
rect 4440 -30940 4500 -30880
rect 6640 -30830 6700 -30770
rect 6420 -30940 6480 -30880
rect 8620 -30830 8680 -30770
rect 8620 -30940 8680 -30880
rect 10820 -30830 10880 -30770
rect 10820 -30940 10880 -30880
rect 13020 -30830 13080 -30770
rect 13020 -30940 13080 -30880
rect 15220 -30830 15280 -30770
rect 15440 -30940 15500 -30880
rect 17640 -30830 17700 -30770
rect 17640 -30940 17700 -30880
rect 19840 -30830 19900 -30770
rect 2510 -31360 2690 -31300
rect 3170 -31360 3350 -31300
rect 3830 -31360 4010 -31300
rect 4710 -31360 4890 -31300
rect 5370 -31360 5550 -31300
rect 6030 -31360 6210 -31300
rect 6910 -31220 7090 -31160
rect 7570 -31220 7750 -31160
rect 8230 -31220 8410 -31160
rect 9110 -31220 9290 -31160
rect 9770 -31220 9950 -31160
rect 10430 -31220 10610 -31160
rect 11310 -31220 11490 -31160
rect 11970 -31220 12150 -31160
rect 12630 -31220 12810 -31160
rect 13510 -31220 13690 -31160
rect 14170 -31220 14350 -31160
rect 14830 -31220 15010 -31160
rect 15710 -31360 15890 -31300
rect 16370 -31360 16550 -31300
rect 17030 -31360 17210 -31300
rect 17910 -31360 18090 -31300
rect 18570 -31360 18750 -31300
rect 19230 -31360 19410 -31300
rect 23040 -25070 23560 -24690
rect 25700 -31880 26220 -31510
rect 34810 -24610 34930 -24490
rect 27260 -25600 27320 -25510
rect 27740 -25760 27800 -25670
rect 27260 -25920 27320 -25830
rect 27740 -26075 27800 -25985
rect 29380 -25970 29440 -25770
rect 27260 -26235 27320 -26145
rect 27740 -26640 27800 -26550
rect 27380 -26800 27440 -26710
rect 27740 -26960 27800 -26870
rect 27380 -27115 27440 -27025
rect 29530 -27010 29590 -26810
rect 27740 -27275 27800 -27185
rect 34810 -25010 34896 -24940
rect 34896 -25010 34900 -24940
rect 37190 -25010 37198 -24940
rect 37198 -25010 37280 -24940
rect 34810 -25270 34896 -25200
rect 34896 -25270 34900 -25200
rect 34810 -25530 34896 -25460
rect 34896 -25530 34900 -25460
rect 37190 -25270 37198 -25200
rect 37198 -25270 37280 -25200
rect 37190 -25530 37198 -25460
rect 37198 -25530 37280 -25460
rect 34810 -25790 34896 -25720
rect 34896 -25790 34900 -25720
rect 34810 -26050 34896 -25980
rect 34896 -26050 34900 -25980
rect 37190 -25790 37198 -25720
rect 37198 -25790 37280 -25720
rect 37190 -26050 37198 -25980
rect 37198 -26050 37280 -25980
rect 34810 -26310 34896 -26240
rect 34896 -26310 34900 -26240
rect 34810 -26570 34896 -26500
rect 34896 -26570 34900 -26500
rect 37190 -26310 37198 -26240
rect 37198 -26310 37280 -26240
rect 37190 -26570 37198 -26500
rect 37198 -26570 37280 -26500
rect 34810 -26830 34896 -26760
rect 34896 -26830 34900 -26760
rect 37190 -26830 37198 -26760
rect 37198 -26830 37280 -26760
rect 36030 -27140 36410 -27010
rect 36530 -27140 36910 -27010
rect 27260 -27685 27320 -27595
rect 27500 -27840 27560 -27750
rect 27260 -28000 27320 -27910
rect 27500 -28155 27560 -28065
rect 29080 -28050 29140 -27850
rect 27260 -28315 27320 -28225
rect 31820 -28290 33160 -28050
rect 27260 -28720 27320 -28630
rect 27620 -28880 27680 -28790
rect 27260 -29040 27320 -28950
rect 27620 -29200 27680 -29110
rect 29230 -29090 29290 -28890
rect 27260 -29350 27320 -29260
rect 31994 -28533 32052 -28528
rect 31994 -28909 32004 -28533
rect 32004 -28909 32052 -28533
rect 32206 -28533 32264 -28528
rect 31994 -28914 32052 -28909
rect 32206 -28909 32252 -28533
rect 32252 -28909 32264 -28533
rect 32206 -28914 32264 -28909
rect 32334 -29334 32472 -29276
rect 27380 -29760 27440 -29670
rect 27620 -29920 27680 -29830
rect 31994 -29553 32052 -29548
rect 31994 -29729 32005 -29553
rect 32005 -29729 32052 -29553
rect 31994 -29734 32052 -29729
rect 32206 -29553 32264 -29550
rect 32206 -29729 32253 -29553
rect 32253 -29729 32264 -29553
rect 32206 -29736 32264 -29729
rect 34194 -28533 34252 -28528
rect 34194 -28909 34204 -28533
rect 34204 -28909 34252 -28533
rect 34406 -28533 34464 -28528
rect 34194 -28914 34252 -28909
rect 34406 -28909 34452 -28533
rect 34452 -28909 34464 -28533
rect 34406 -28914 34464 -28909
rect 33004 -29334 33142 -29276
rect 33360 -29290 33560 -29210
rect 33454 -29430 33588 -29378
rect 33078 -29553 33166 -29546
rect 33078 -29729 33132 -29553
rect 33132 -29729 33166 -29553
rect 33078 -29736 33166 -29729
rect 34534 -29334 34672 -29276
rect 34194 -29553 34252 -29548
rect 34194 -29729 34205 -29553
rect 34205 -29729 34252 -29553
rect 34194 -29734 34252 -29729
rect 34406 -29553 34464 -29550
rect 34406 -29729 34453 -29553
rect 34453 -29729 34464 -29553
rect 34406 -29736 34464 -29729
rect 36394 -28533 36452 -28528
rect 36394 -28909 36404 -28533
rect 36404 -28909 36452 -28533
rect 36606 -28533 36664 -28528
rect 36394 -28914 36452 -28909
rect 36606 -28909 36652 -28533
rect 36652 -28909 36664 -28533
rect 36606 -28914 36664 -28909
rect 35204 -29334 35342 -29276
rect 35560 -29290 35760 -29210
rect 35654 -29430 35788 -29378
rect 35278 -29553 35366 -29546
rect 35278 -29729 35332 -29553
rect 35332 -29729 35366 -29553
rect 35278 -29736 35366 -29729
rect 36734 -29334 36872 -29276
rect 36394 -29553 36452 -29548
rect 36394 -29729 36405 -29553
rect 36405 -29729 36452 -29553
rect 36394 -29734 36452 -29729
rect 36606 -29553 36664 -29550
rect 36606 -29729 36653 -29553
rect 36653 -29729 36664 -29553
rect 36606 -29736 36664 -29729
rect 37404 -29334 37542 -29276
rect 37760 -29290 37960 -29210
rect 37854 -29430 37988 -29378
rect 37478 -29553 37566 -29546
rect 37478 -29729 37532 -29553
rect 37532 -29729 37566 -29553
rect 37478 -29736 37566 -29729
rect 27380 -30075 27440 -29985
rect 27620 -30235 27680 -30145
rect 29080 -30130 29140 -29930
rect 37250 -29951 37385 -29920
rect 37385 -29951 37503 -29920
rect 37503 -29951 37690 -29920
rect 37250 -30073 37690 -29951
rect 37250 -30107 37316 -30073
rect 37316 -30107 37630 -30073
rect 37630 -30107 37690 -30073
rect 37250 -30110 37690 -30107
rect 27380 -30390 27440 -30300
rect 32256 -30295 32344 -30288
rect 32256 -30471 32290 -30295
rect 32290 -30471 32344 -30295
rect 32256 -30478 32344 -30471
rect 27380 -30800 27440 -30710
rect 27500 -30960 27560 -30870
rect 27380 -31115 27440 -31025
rect 29070 -31030 29290 -30960
rect 27500 -31275 27560 -31185
rect 27380 -31430 27440 -31340
rect 31834 -30646 31968 -30594
rect 31850 -30810 32050 -30730
rect 32280 -30748 32418 -30690
rect 33158 -30295 33216 -30288
rect 33158 -30471 33169 -30295
rect 33169 -30471 33216 -30295
rect 33158 -30474 33216 -30471
rect 33370 -30295 33428 -30290
rect 33370 -30471 33417 -30295
rect 33417 -30471 33428 -30295
rect 33370 -30476 33428 -30471
rect 32950 -30748 33088 -30690
rect 34456 -30295 34544 -30288
rect 34456 -30471 34490 -30295
rect 34490 -30471 34544 -30295
rect 34456 -30478 34544 -30471
rect 34034 -30646 34168 -30594
rect 34060 -30810 34260 -30730
rect 34480 -30748 34618 -30690
rect 33158 -31115 33216 -31110
rect 33158 -31491 33170 -31115
rect 33170 -31491 33216 -31115
rect 33370 -31115 33428 -31110
rect 33158 -31496 33216 -31491
rect 33370 -31491 33418 -31115
rect 33418 -31491 33428 -31115
rect 33370 -31496 33428 -31491
rect 35358 -30295 35416 -30288
rect 35358 -30471 35369 -30295
rect 35369 -30471 35416 -30295
rect 35358 -30474 35416 -30471
rect 35570 -30295 35628 -30290
rect 35570 -30471 35617 -30295
rect 35617 -30471 35628 -30295
rect 35570 -30476 35628 -30471
rect 35150 -30748 35288 -30690
rect 36656 -30295 36744 -30288
rect 36656 -30471 36690 -30295
rect 36690 -30471 36744 -30295
rect 36656 -30478 36744 -30471
rect 36234 -30646 36368 -30594
rect 36260 -30820 36460 -30740
rect 36680 -30748 36818 -30690
rect 35358 -31115 35416 -31110
rect 35358 -31491 35370 -31115
rect 35370 -31491 35416 -31115
rect 35570 -31115 35628 -31110
rect 35358 -31496 35416 -31491
rect 35570 -31491 35618 -31115
rect 35618 -31491 35628 -31115
rect 35570 -31496 35628 -31491
rect 37558 -30295 37616 -30288
rect 37558 -30471 37569 -30295
rect 37569 -30471 37616 -30295
rect 37558 -30474 37616 -30471
rect 37770 -30295 37828 -30290
rect 37770 -30471 37817 -30295
rect 37817 -30471 37828 -30295
rect 37770 -30476 37828 -30471
rect 37350 -30748 37488 -30690
rect 37558 -31115 37616 -31110
rect 37558 -31491 37570 -31115
rect 37570 -31491 37616 -31115
rect 37770 -31115 37828 -31110
rect 37558 -31496 37616 -31491
rect 37770 -31491 37818 -31115
rect 37818 -31491 37828 -31115
rect 37770 -31496 37828 -31491
rect 32540 -31950 33690 -31730
<< metal2 >>
rect -360 11990 -160 12000
rect -360 11610 -350 11990
rect -170 11610 -160 11990
rect 2020 11720 2080 12020
rect 2200 12010 2340 12020
rect 2200 11890 2210 12010
rect 2330 11890 2340 12010
rect 2200 11880 2340 11890
rect 1980 11710 2120 11720
rect -360 -31450 -160 11610
rect 80 11690 280 11700
rect 80 11310 90 11690
rect 270 11310 280 11690
rect 1980 11590 1990 11710
rect 2110 11590 2120 11710
rect 1980 11580 2120 11590
rect -70 10930 -10 10940
rect -70 10860 -10 10870
rect -70 10130 -10 10140
rect -70 10060 -10 10070
rect -70 9330 -10 9340
rect -70 9260 -10 9270
rect -70 8530 -10 8540
rect -70 8460 -10 8470
rect -70 7730 -10 7740
rect -70 7660 -10 7670
rect -70 6930 -10 6940
rect -70 6860 -10 6870
rect -70 6130 -10 6140
rect -70 6060 -10 6070
rect -70 5330 -10 5340
rect -70 5260 -10 5270
rect -360 -31830 -350 -31450
rect -170 -31830 -160 -31450
rect -360 -32120 -160 -31830
rect 80 -31730 280 11310
rect 2020 10830 2080 11580
rect 2130 10930 2190 10940
rect 2130 10860 2190 10870
rect 2240 10830 2300 11880
rect 4220 11720 4280 12020
rect 4400 12010 4540 12020
rect 4400 11890 4410 12010
rect 4530 11890 4540 12010
rect 4400 11880 4540 11890
rect 4180 11710 4320 11720
rect 4180 11590 4190 11710
rect 4310 11590 4320 11710
rect 4180 11580 4320 11590
rect 2500 11240 2700 11250
rect 2500 11180 2510 11240
rect 2690 11180 2700 11240
rect 2500 11170 2700 11180
rect 3160 11240 3360 11250
rect 3160 11180 3170 11240
rect 3350 11180 3360 11240
rect 3160 11170 3360 11180
rect 3820 11240 4020 11250
rect 3820 11180 3830 11240
rect 4010 11180 4020 11240
rect 3820 11170 4020 11180
rect 2500 11030 2700 11110
rect 3160 11030 3360 11110
rect 3820 11030 4020 11110
rect 4220 10830 4280 11580
rect 4330 10930 4390 10940
rect 4330 10860 4390 10870
rect 4440 10830 4500 11880
rect 6420 11720 6480 12020
rect 6600 12010 6740 12020
rect 6600 11890 6610 12010
rect 6730 11890 6740 12010
rect 6600 11880 6740 11890
rect 6380 11710 6520 11720
rect 6380 11590 6390 11710
rect 6510 11590 6520 11710
rect 6380 11580 6520 11590
rect 4700 11240 4900 11250
rect 4700 11180 4710 11240
rect 4890 11180 4900 11240
rect 4700 11170 4900 11180
rect 5360 11240 5560 11250
rect 5360 11180 5370 11240
rect 5550 11180 5560 11240
rect 5360 11170 5560 11180
rect 6020 11240 6220 11250
rect 6020 11180 6030 11240
rect 6210 11180 6220 11240
rect 6020 11170 6220 11180
rect 4700 11030 4900 11110
rect 5360 11030 5560 11110
rect 6020 11030 6220 11110
rect 6420 10830 6480 11580
rect 6530 10930 6590 10940
rect 6530 10860 6590 10870
rect 6640 10830 6700 11880
rect 8620 11720 8680 12020
rect 8800 12010 8940 12020
rect 8800 11890 8810 12010
rect 8930 11890 8940 12010
rect 8800 11880 8940 11890
rect 8580 11710 8720 11720
rect 8580 11590 8590 11710
rect 8710 11590 8720 11710
rect 8580 11580 8720 11590
rect 6900 11170 7100 11250
rect 7560 11170 7760 11250
rect 8220 11170 8420 11250
rect 6900 11100 7100 11110
rect 6900 11040 6910 11100
rect 7090 11040 7100 11100
rect 6900 11030 7100 11040
rect 7560 11100 7760 11110
rect 7560 11040 7570 11100
rect 7750 11040 7760 11100
rect 7560 11030 7760 11040
rect 8220 11100 8420 11110
rect 8220 11040 8230 11100
rect 8410 11040 8420 11100
rect 8220 11030 8420 11040
rect 8620 10830 8680 11580
rect 8730 10930 8790 10940
rect 8730 10860 8790 10870
rect 8840 10830 8900 11880
rect 10820 11720 10880 12020
rect 11000 12010 11140 12020
rect 11000 11890 11010 12010
rect 11130 11890 11140 12010
rect 11000 11880 11140 11890
rect 10780 11710 10920 11720
rect 10780 11590 10790 11710
rect 10910 11590 10920 11710
rect 10780 11580 10920 11590
rect 9100 11170 9300 11250
rect 9760 11170 9960 11250
rect 10420 11170 10620 11250
rect 9100 11100 9300 11110
rect 9100 11040 9110 11100
rect 9290 11040 9300 11100
rect 9100 11030 9300 11040
rect 9760 11100 9960 11110
rect 9760 11040 9770 11100
rect 9950 11040 9960 11100
rect 9760 11030 9960 11040
rect 10420 11100 10620 11110
rect 10420 11040 10430 11100
rect 10610 11040 10620 11100
rect 10420 11030 10620 11040
rect 10820 10830 10880 11580
rect 10930 10930 10990 10940
rect 10930 10860 10990 10870
rect 11040 10830 11100 11880
rect 13020 11720 13080 12020
rect 13200 12010 13340 12020
rect 13200 11890 13210 12010
rect 13330 11890 13340 12010
rect 13200 11880 13340 11890
rect 12980 11710 13120 11720
rect 12980 11590 12990 11710
rect 13110 11590 13120 11710
rect 12980 11580 13120 11590
rect 11300 11170 11500 11250
rect 11960 11170 12160 11250
rect 12620 11170 12820 11250
rect 11300 11100 11500 11110
rect 11300 11040 11310 11100
rect 11490 11040 11500 11100
rect 11300 11030 11500 11040
rect 11960 11100 12160 11110
rect 11960 11040 11970 11100
rect 12150 11040 12160 11100
rect 11960 11030 12160 11040
rect 12620 11100 12820 11110
rect 12620 11040 12630 11100
rect 12810 11040 12820 11100
rect 12620 11030 12820 11040
rect 13020 10830 13080 11580
rect 13130 10930 13190 10940
rect 13130 10860 13190 10870
rect 13240 10830 13300 11880
rect 15220 11720 15280 12020
rect 15400 12010 15540 12020
rect 15400 11890 15410 12010
rect 15530 11890 15540 12010
rect 15400 11880 15540 11890
rect 15180 11710 15320 11720
rect 15180 11590 15190 11710
rect 15310 11590 15320 11710
rect 15180 11580 15320 11590
rect 13500 11170 13700 11250
rect 14160 11170 14360 11250
rect 14820 11170 15020 11250
rect 13500 11100 13700 11110
rect 13500 11040 13510 11100
rect 13690 11040 13700 11100
rect 13500 11030 13700 11040
rect 14160 11100 14360 11110
rect 14160 11040 14170 11100
rect 14350 11040 14360 11100
rect 14160 11030 14360 11040
rect 14820 11100 15020 11110
rect 14820 11040 14830 11100
rect 15010 11040 15020 11100
rect 14820 11030 15020 11040
rect 15220 10830 15280 11580
rect 15330 10930 15390 10940
rect 15330 10860 15390 10870
rect 15440 10830 15500 11880
rect 17420 11720 17480 12020
rect 17600 12010 17740 12020
rect 17600 11890 17610 12010
rect 17730 11890 17740 12010
rect 17600 11880 17740 11890
rect 17380 11710 17520 11720
rect 17380 11590 17390 11710
rect 17510 11590 17520 11710
rect 17380 11580 17520 11590
rect 15700 11240 15900 11250
rect 15700 11180 15710 11240
rect 15890 11180 15900 11240
rect 15700 11170 15900 11180
rect 16360 11240 16560 11250
rect 16360 11180 16370 11240
rect 16550 11180 16560 11240
rect 16360 11170 16560 11180
rect 17020 11240 17220 11250
rect 17020 11180 17030 11240
rect 17210 11180 17220 11240
rect 17020 11170 17220 11180
rect 15700 11030 15900 11110
rect 16360 11030 16560 11110
rect 17020 11030 17220 11110
rect 17420 10830 17480 11580
rect 17530 10930 17590 10940
rect 17530 10860 17590 10870
rect 17640 10830 17700 11880
rect 19620 11720 19680 12020
rect 19800 12010 19940 12020
rect 19800 11890 19810 12010
rect 19930 11890 19940 12010
rect 19800 11880 19940 11890
rect 36470 11980 36820 11990
rect 19580 11710 19720 11720
rect 19580 11590 19590 11710
rect 19710 11590 19720 11710
rect 19580 11580 19720 11590
rect 17900 11240 18100 11250
rect 17900 11180 17910 11240
rect 18090 11180 18100 11240
rect 17900 11170 18100 11180
rect 18560 11240 18760 11250
rect 18560 11180 18570 11240
rect 18750 11180 18760 11240
rect 18560 11170 18760 11180
rect 19220 11240 19420 11250
rect 19220 11180 19230 11240
rect 19410 11180 19420 11240
rect 19220 11170 19420 11180
rect 17900 11030 18100 11110
rect 18560 11030 18760 11110
rect 19220 11030 19420 11110
rect 2010 10710 2090 10830
rect 2010 10650 2020 10710
rect 2080 10650 2090 10710
rect 2010 10640 2090 10650
rect 2230 10640 2310 10830
rect 4210 10820 4290 10830
rect 4210 10760 4220 10820
rect 4280 10760 4290 10820
rect 4210 10710 4290 10760
rect 4210 10650 4220 10710
rect 4280 10650 4290 10710
rect 4210 10640 4290 10650
rect 4430 10640 4510 10830
rect 6410 10820 6490 10830
rect 6410 10760 6420 10820
rect 6480 10760 6490 10820
rect 6410 10640 6490 10760
rect 6630 10710 6710 10830
rect 6630 10650 6640 10710
rect 6700 10650 6710 10710
rect 6630 10640 6710 10650
rect 8610 10640 8690 10830
rect 8830 10820 8910 10830
rect 8830 10760 8840 10820
rect 8900 10760 8910 10820
rect 8830 10710 8910 10760
rect 8830 10650 8840 10710
rect 8900 10650 8910 10710
rect 8830 10640 8910 10650
rect 10810 10640 10890 10830
rect 11030 10820 11110 10830
rect 11030 10760 11040 10820
rect 11100 10760 11110 10820
rect 11030 10710 11110 10760
rect 11030 10650 11040 10710
rect 11100 10650 11110 10710
rect 11030 10640 11110 10650
rect 13010 10640 13090 10830
rect 13230 10820 13310 10830
rect 13230 10760 13240 10820
rect 13300 10760 13310 10820
rect 13230 10710 13310 10760
rect 13230 10650 13240 10710
rect 13300 10650 13310 10710
rect 13230 10640 13310 10650
rect 15210 10710 15290 10830
rect 15210 10650 15220 10710
rect 15280 10650 15290 10710
rect 15210 10640 15290 10650
rect 15430 10820 15510 10830
rect 15430 10760 15440 10820
rect 15500 10760 15510 10820
rect 15430 10640 15510 10760
rect 17410 10820 17490 10830
rect 17410 10760 17420 10820
rect 17480 10760 17490 10820
rect 17410 10710 17490 10760
rect 17410 10650 17420 10710
rect 17480 10650 17490 10710
rect 17410 10640 17490 10650
rect 17630 10640 17710 10830
rect 19620 10810 19680 11580
rect 19730 10930 19790 10940
rect 19730 10860 19790 10870
rect 19840 10810 19900 11880
rect 25710 11780 26250 11790
rect 25710 11410 25720 11780
rect 26240 11690 26250 11780
rect 30570 11722 30670 11728
rect 26240 11500 27320 11690
rect 30570 11532 30576 11722
rect 30664 11532 30670 11722
rect 26240 11490 27330 11500
rect 26240 11410 26250 11490
rect 25710 11400 26250 11410
rect 21930 10930 21990 10940
rect 21930 10860 21990 10870
rect 19610 10800 19690 10810
rect 19610 10740 19620 10800
rect 19680 10740 19690 10800
rect 19610 10640 19690 10740
rect 19830 10640 19910 10810
rect 2020 10030 2080 10640
rect 2130 10130 2190 10140
rect 2130 10060 2190 10070
rect 2240 10030 2300 10640
rect 2500 10610 4020 10620
rect 2500 10550 2510 10610
rect 4010 10550 4020 10610
rect 2500 10540 4020 10550
rect 2500 10370 2700 10450
rect 3160 10370 3360 10450
rect 3820 10370 4020 10450
rect 2500 10300 2700 10310
rect 2500 10240 2510 10300
rect 2690 10240 2700 10300
rect 2500 10230 2700 10240
rect 3160 10300 3360 10310
rect 3160 10240 3170 10300
rect 3350 10240 3360 10300
rect 3160 10230 3360 10240
rect 3820 10300 4020 10310
rect 3820 10240 3830 10300
rect 4010 10240 4020 10300
rect 3820 10230 4020 10240
rect 4220 10030 4280 10640
rect 4330 10130 4390 10140
rect 4330 10060 4390 10070
rect 4440 10030 4500 10640
rect 4700 10610 6220 10620
rect 4700 10550 4710 10610
rect 6210 10550 6220 10610
rect 4700 10540 6220 10550
rect 4700 10370 4900 10450
rect 5360 10370 5560 10450
rect 6020 10370 6220 10450
rect 4700 10300 4900 10310
rect 4700 10240 4710 10300
rect 4890 10240 4900 10300
rect 4700 10230 4900 10240
rect 5360 10300 5560 10310
rect 5360 10240 5370 10300
rect 5550 10240 5560 10300
rect 5360 10230 5560 10240
rect 6020 10300 6220 10310
rect 6020 10240 6030 10300
rect 6210 10240 6220 10300
rect 6020 10230 6220 10240
rect 6420 10030 6480 10640
rect 6530 10130 6590 10140
rect 6530 10060 6590 10070
rect 6640 10030 6700 10640
rect 6900 10610 8420 10620
rect 6900 10550 6910 10610
rect 8410 10550 8420 10610
rect 6900 10540 8420 10550
rect 6900 10440 7100 10450
rect 6900 10380 6910 10440
rect 7090 10380 7100 10440
rect 6900 10370 7100 10380
rect 7560 10440 7760 10450
rect 7560 10380 7570 10440
rect 7750 10380 7760 10440
rect 7560 10370 7760 10380
rect 8220 10440 8420 10450
rect 8220 10380 8230 10440
rect 8410 10380 8420 10440
rect 8220 10370 8420 10380
rect 6900 10230 7100 10310
rect 7560 10230 7760 10310
rect 8220 10230 8420 10310
rect 8620 10030 8680 10640
rect 8730 10130 8790 10140
rect 8730 10060 8790 10070
rect 8840 10030 8900 10640
rect 9100 10610 10620 10620
rect 9100 10550 9110 10610
rect 10610 10550 10620 10610
rect 9100 10540 10620 10550
rect 9100 10440 9300 10450
rect 9100 10380 9110 10440
rect 9290 10380 9300 10440
rect 9100 10370 9300 10380
rect 9760 10440 9960 10450
rect 9760 10380 9770 10440
rect 9950 10380 9960 10440
rect 9760 10370 9960 10380
rect 10420 10440 10620 10450
rect 10420 10380 10430 10440
rect 10610 10380 10620 10440
rect 10420 10370 10620 10380
rect 9100 10230 9300 10310
rect 9760 10230 9960 10310
rect 10420 10230 10620 10310
rect 10820 10030 10880 10640
rect 10930 10130 10990 10140
rect 10930 10060 10990 10070
rect 11040 10030 11100 10640
rect 11300 10610 12820 10620
rect 11300 10550 11310 10610
rect 12810 10550 12820 10610
rect 11300 10540 12820 10550
rect 11300 10440 11500 10450
rect 11300 10380 11310 10440
rect 11490 10380 11500 10440
rect 11300 10370 11500 10380
rect 11960 10440 12160 10450
rect 11960 10380 11970 10440
rect 12150 10380 12160 10440
rect 11960 10370 12160 10380
rect 12620 10440 12820 10450
rect 12620 10380 12630 10440
rect 12810 10380 12820 10440
rect 12620 10370 12820 10380
rect 11300 10230 11500 10310
rect 11960 10230 12160 10310
rect 12620 10230 12820 10310
rect 13020 10030 13080 10640
rect 13130 10130 13190 10140
rect 13130 10060 13190 10070
rect 13240 10030 13300 10640
rect 13500 10610 15020 10620
rect 13500 10550 13510 10610
rect 15010 10550 15020 10610
rect 13500 10540 15020 10550
rect 13500 10440 13700 10450
rect 13500 10380 13510 10440
rect 13690 10380 13700 10440
rect 13500 10370 13700 10380
rect 14160 10440 14360 10450
rect 14160 10380 14170 10440
rect 14350 10380 14360 10440
rect 14160 10370 14360 10380
rect 14820 10440 15020 10450
rect 14820 10380 14830 10440
rect 15010 10380 15020 10440
rect 14820 10370 15020 10380
rect 13500 10230 13700 10310
rect 14160 10230 14360 10310
rect 14820 10230 15020 10310
rect 15220 10030 15280 10640
rect 15330 10130 15390 10140
rect 15330 10060 15390 10070
rect 15440 10030 15500 10640
rect 15700 10610 17220 10620
rect 15700 10550 15710 10610
rect 17210 10550 17220 10610
rect 15700 10540 17220 10550
rect 15700 10370 15900 10450
rect 16360 10370 16560 10450
rect 17020 10370 17220 10450
rect 15700 10300 15900 10310
rect 15700 10240 15710 10300
rect 15890 10240 15900 10300
rect 15700 10230 15900 10240
rect 16360 10300 16560 10310
rect 16360 10240 16370 10300
rect 16550 10240 16560 10300
rect 16360 10230 16560 10240
rect 17020 10300 17220 10310
rect 17020 10240 17030 10300
rect 17210 10240 17220 10300
rect 17020 10230 17220 10240
rect 17420 10030 17480 10640
rect 17530 10130 17590 10140
rect 17530 10060 17590 10070
rect 17640 10030 17700 10640
rect 17900 10610 19420 10620
rect 17900 10550 17910 10610
rect 19410 10550 19420 10610
rect 17900 10540 19420 10550
rect 17900 10370 18100 10450
rect 18560 10370 18760 10450
rect 19220 10370 19420 10450
rect 17900 10300 18100 10310
rect 17900 10240 17910 10300
rect 18090 10240 18100 10300
rect 17900 10230 18100 10240
rect 18560 10300 18760 10310
rect 18560 10240 18570 10300
rect 18750 10240 18760 10300
rect 18560 10230 18760 10240
rect 19220 10300 19420 10310
rect 19220 10240 19230 10300
rect 19410 10240 19420 10300
rect 19220 10230 19420 10240
rect 2010 9840 2090 10030
rect 2230 9910 2310 10030
rect 2230 9850 2240 9910
rect 2300 9850 2310 9910
rect 2230 9840 2310 9850
rect 4210 9840 4290 10030
rect 4430 10020 4510 10030
rect 4430 9960 4440 10020
rect 4500 9960 4510 10020
rect 4430 9910 4510 9960
rect 4430 9850 4440 9910
rect 4500 9850 4510 9910
rect 4430 9840 4510 9850
rect 6410 9910 6490 10030
rect 6410 9850 6420 9910
rect 6480 9850 6490 9910
rect 6410 9840 6490 9850
rect 6630 10020 6710 10030
rect 6630 9960 6640 10020
rect 6700 9960 6710 10020
rect 6630 9840 6710 9960
rect 8610 10020 8690 10030
rect 8610 9960 8620 10020
rect 8680 9960 8690 10020
rect 8610 9910 8690 9960
rect 8610 9850 8620 9910
rect 8680 9850 8690 9910
rect 8610 9840 8690 9850
rect 8830 9840 8910 10030
rect 10810 10020 10890 10030
rect 10810 9960 10820 10020
rect 10880 9960 10890 10020
rect 10810 9910 10890 9960
rect 10810 9850 10820 9910
rect 10880 9850 10890 9910
rect 10810 9840 10890 9850
rect 11030 9840 11110 10030
rect 13010 10020 13090 10030
rect 13010 9960 13020 10020
rect 13080 9960 13090 10020
rect 13010 9910 13090 9960
rect 13010 9850 13020 9910
rect 13080 9850 13090 9910
rect 13010 9840 13090 9850
rect 13230 9840 13310 10030
rect 15210 10020 15290 10030
rect 15210 9960 15220 10020
rect 15280 9960 15290 10020
rect 15210 9840 15290 9960
rect 15430 9910 15510 10030
rect 15430 9850 15440 9910
rect 15500 9850 15510 9910
rect 15430 9840 15510 9850
rect 17410 9840 17490 10030
rect 17630 10020 17710 10030
rect 17630 9960 17640 10020
rect 17700 9960 17710 10020
rect 19620 10010 19680 10640
rect 19730 10130 19790 10140
rect 19730 10060 19790 10070
rect 19840 10010 19900 10640
rect 21930 10130 21990 10140
rect 21930 10060 21990 10070
rect 17630 9910 17710 9960
rect 17630 9850 17640 9910
rect 17700 9850 17710 9910
rect 17630 9840 17710 9850
rect 19610 9840 19690 10010
rect 19830 10000 19910 10010
rect 19830 9940 19840 10000
rect 19900 9940 19910 10000
rect 19830 9840 19910 9940
rect 2020 9230 2080 9840
rect 2130 9330 2190 9340
rect 2130 9260 2190 9270
rect 2240 9230 2300 9840
rect 2500 9810 4020 9820
rect 2500 9750 2510 9810
rect 4010 9750 4020 9810
rect 2500 9740 4020 9750
rect 2500 9640 2700 9650
rect 2500 9580 2510 9640
rect 2690 9580 2700 9640
rect 2500 9570 2700 9580
rect 3160 9640 3360 9650
rect 3160 9580 3170 9640
rect 3350 9580 3360 9640
rect 3160 9570 3360 9580
rect 3820 9640 4020 9650
rect 3820 9580 3830 9640
rect 4010 9580 4020 9640
rect 3820 9570 4020 9580
rect 2500 9430 2700 9510
rect 3160 9430 3360 9510
rect 3820 9430 4020 9510
rect 4220 9230 4280 9840
rect 4330 9330 4390 9340
rect 4330 9260 4390 9270
rect 4440 9230 4500 9840
rect 4700 9810 6220 9820
rect 4700 9750 4710 9810
rect 6210 9750 6220 9810
rect 4700 9740 6220 9750
rect 4700 9640 4900 9650
rect 4700 9580 4710 9640
rect 4890 9580 4900 9640
rect 4700 9570 4900 9580
rect 5360 9640 5560 9650
rect 5360 9580 5370 9640
rect 5550 9580 5560 9640
rect 5360 9570 5560 9580
rect 6020 9640 6220 9650
rect 6020 9580 6030 9640
rect 6210 9580 6220 9640
rect 6020 9570 6220 9580
rect 4700 9430 4900 9510
rect 5360 9430 5560 9510
rect 6020 9430 6220 9510
rect 6420 9230 6480 9840
rect 6530 9330 6590 9340
rect 6530 9260 6590 9270
rect 6640 9230 6700 9840
rect 6900 9810 8420 9820
rect 6900 9750 6910 9810
rect 8410 9750 8420 9810
rect 6900 9740 8420 9750
rect 6900 9570 7100 9650
rect 7560 9570 7760 9650
rect 8220 9570 8420 9650
rect 6900 9500 7100 9510
rect 6900 9440 6910 9500
rect 7090 9440 7100 9500
rect 6900 9430 7100 9440
rect 7560 9500 7760 9510
rect 7560 9440 7570 9500
rect 7750 9440 7760 9500
rect 7560 9430 7760 9440
rect 8220 9500 8420 9510
rect 8220 9440 8230 9500
rect 8410 9440 8420 9500
rect 8220 9430 8420 9440
rect 8620 9230 8680 9840
rect 8730 9330 8790 9340
rect 8730 9260 8790 9270
rect 8840 9230 8900 9840
rect 9100 9810 10620 9820
rect 9100 9750 9110 9810
rect 10610 9750 10620 9810
rect 9100 9740 10620 9750
rect 9100 9570 9300 9650
rect 9760 9570 9960 9650
rect 10420 9570 10620 9650
rect 9100 9500 9300 9510
rect 9100 9440 9110 9500
rect 9290 9440 9300 9500
rect 9100 9430 9300 9440
rect 9760 9500 9960 9510
rect 9760 9440 9770 9500
rect 9950 9440 9960 9500
rect 9760 9430 9960 9440
rect 10420 9500 10620 9510
rect 10420 9440 10430 9500
rect 10610 9440 10620 9500
rect 10420 9430 10620 9440
rect 10820 9230 10880 9840
rect 10930 9330 10990 9340
rect 10930 9260 10990 9270
rect 11040 9230 11100 9840
rect 11300 9810 12820 9820
rect 11300 9750 11310 9810
rect 12810 9750 12820 9810
rect 11300 9740 12820 9750
rect 11300 9570 11500 9650
rect 11960 9570 12160 9650
rect 12620 9570 12820 9650
rect 11300 9500 11500 9510
rect 11300 9440 11310 9500
rect 11490 9440 11500 9500
rect 11300 9430 11500 9440
rect 11960 9500 12160 9510
rect 11960 9440 11970 9500
rect 12150 9440 12160 9500
rect 11960 9430 12160 9440
rect 12620 9500 12820 9510
rect 12620 9440 12630 9500
rect 12810 9440 12820 9500
rect 12620 9430 12820 9440
rect 13020 9230 13080 9840
rect 13130 9330 13190 9340
rect 13130 9260 13190 9270
rect 13240 9230 13300 9840
rect 13500 9810 15020 9820
rect 13500 9750 13510 9810
rect 15010 9750 15020 9810
rect 13500 9740 15020 9750
rect 13500 9570 13700 9650
rect 14160 9570 14360 9650
rect 14820 9570 15020 9650
rect 13500 9500 13700 9510
rect 13500 9440 13510 9500
rect 13690 9440 13700 9500
rect 13500 9430 13700 9440
rect 14160 9500 14360 9510
rect 14160 9440 14170 9500
rect 14350 9440 14360 9500
rect 14160 9430 14360 9440
rect 14820 9500 15020 9510
rect 14820 9440 14830 9500
rect 15010 9440 15020 9500
rect 14820 9430 15020 9440
rect 15220 9230 15280 9840
rect 15330 9330 15390 9340
rect 15330 9260 15390 9270
rect 15440 9230 15500 9840
rect 15700 9810 17220 9820
rect 15700 9750 15710 9810
rect 17210 9750 17220 9810
rect 15700 9740 17220 9750
rect 15700 9640 15900 9650
rect 15700 9580 15710 9640
rect 15890 9580 15900 9640
rect 15700 9570 15900 9580
rect 16360 9640 16560 9650
rect 16360 9580 16370 9640
rect 16550 9580 16560 9640
rect 16360 9570 16560 9580
rect 17020 9640 17220 9650
rect 17020 9580 17030 9640
rect 17210 9580 17220 9640
rect 17020 9570 17220 9580
rect 15700 9430 15900 9510
rect 16360 9430 16560 9510
rect 17020 9430 17220 9510
rect 17420 9230 17480 9840
rect 17530 9330 17590 9340
rect 17530 9260 17590 9270
rect 17640 9230 17700 9840
rect 17900 9810 19420 9820
rect 17900 9750 17910 9810
rect 19410 9750 19420 9810
rect 17900 9740 19420 9750
rect 17900 9640 18100 9650
rect 17900 9580 17910 9640
rect 18090 9580 18100 9640
rect 17900 9570 18100 9580
rect 18560 9640 18760 9650
rect 18560 9580 18570 9640
rect 18750 9580 18760 9640
rect 18560 9570 18760 9580
rect 19220 9640 19420 9650
rect 19220 9580 19230 9640
rect 19410 9580 19420 9640
rect 19220 9570 19420 9580
rect 17900 9430 18100 9510
rect 18560 9430 18760 9510
rect 19220 9430 19420 9510
rect 1410 9210 1490 9220
rect 1410 9060 1420 9210
rect 1480 9060 1490 9210
rect 1410 9050 1490 9060
rect 420 8990 620 9000
rect 420 8910 430 8990
rect 610 8910 620 8990
rect 420 8900 620 8910
rect 420 8190 620 8200
rect 420 8110 430 8190
rect 610 8110 620 8190
rect 420 8100 620 8110
rect 420 7390 620 7400
rect 420 7310 430 7390
rect 610 7310 620 7390
rect 420 7300 620 7310
rect 1420 6820 1480 9050
rect 1620 8420 1680 9220
rect 2010 9040 2090 9230
rect 2230 9040 2310 9230
rect 4210 9110 4290 9230
rect 4210 9050 4220 9110
rect 4280 9050 4290 9110
rect 4210 9040 4290 9050
rect 4430 9040 4510 9230
rect 6410 9220 6490 9230
rect 6410 9160 6420 9220
rect 6480 9160 6490 9220
rect 6410 9040 6490 9160
rect 6630 9110 6710 9230
rect 6630 9050 6640 9110
rect 6700 9050 6710 9110
rect 6630 9040 6710 9050
rect 8610 9040 8690 9230
rect 8830 9220 8910 9230
rect 8830 9160 8840 9220
rect 8900 9160 8910 9220
rect 8830 9110 8910 9160
rect 8830 9050 8840 9110
rect 8900 9050 8910 9110
rect 8830 9040 8910 9050
rect 10810 9040 10890 9230
rect 11030 9220 11110 9230
rect 11030 9160 11040 9220
rect 11100 9160 11110 9220
rect 11030 9110 11110 9160
rect 11030 9050 11040 9110
rect 11100 9050 11110 9110
rect 11030 9040 11110 9050
rect 13010 9040 13090 9230
rect 13230 9220 13310 9230
rect 13230 9160 13240 9220
rect 13300 9160 13310 9220
rect 13230 9110 13310 9160
rect 13230 9050 13240 9110
rect 13300 9050 13310 9110
rect 13230 9040 13310 9050
rect 15210 9110 15290 9230
rect 15210 9050 15220 9110
rect 15280 9050 15290 9110
rect 15210 9040 15290 9050
rect 15430 9220 15510 9230
rect 15430 9160 15440 9220
rect 15500 9160 15510 9220
rect 15430 9040 15510 9160
rect 17410 9220 17490 9230
rect 17410 9160 17420 9220
rect 17480 9160 17490 9220
rect 17410 9040 17490 9160
rect 17630 9040 17710 9230
rect 19620 9210 19680 9840
rect 19730 9330 19790 9340
rect 19730 9260 19790 9270
rect 19840 9210 19900 9840
rect 21930 9330 21990 9340
rect 20230 9300 20310 9310
rect 19610 9040 19690 9210
rect 19830 9040 19910 9210
rect 20230 9150 20240 9300
rect 20300 9150 20310 9300
rect 20230 9140 20310 9150
rect 2020 8430 2080 9040
rect 2130 8530 2190 8540
rect 2130 8460 2190 8470
rect 2240 8430 2300 9040
rect 2500 8770 2700 8850
rect 3160 8770 3360 8850
rect 3820 8770 4020 8850
rect 2500 8700 2700 8710
rect 2500 8640 2510 8700
rect 2690 8640 2700 8700
rect 2500 8630 2700 8640
rect 3160 8700 3360 8710
rect 3160 8640 3170 8700
rect 3350 8640 3360 8700
rect 3160 8630 3360 8640
rect 3820 8700 4020 8710
rect 3820 8640 3830 8700
rect 4010 8640 4020 8700
rect 3820 8630 4020 8640
rect 4220 8430 4280 9040
rect 4330 8530 4390 8540
rect 4330 8460 4390 8470
rect 4440 8430 4500 9040
rect 4700 9010 6220 9020
rect 4700 8950 4710 9010
rect 6210 8950 6220 9010
rect 4700 8940 6220 8950
rect 4700 8770 4900 8850
rect 5360 8770 5560 8850
rect 6020 8770 6220 8850
rect 4700 8700 4900 8710
rect 4700 8640 4710 8700
rect 4890 8640 4900 8700
rect 4700 8630 4900 8640
rect 5360 8700 5560 8710
rect 5360 8640 5370 8700
rect 5550 8640 5560 8700
rect 5360 8630 5560 8640
rect 6020 8700 6220 8710
rect 6020 8640 6030 8700
rect 6210 8640 6220 8700
rect 6020 8630 6220 8640
rect 6420 8430 6480 9040
rect 6530 8530 6590 8540
rect 6530 8460 6590 8470
rect 6640 8430 6700 9040
rect 6900 9010 8420 9020
rect 6900 8950 6910 9010
rect 8410 8950 8420 9010
rect 6900 8940 8420 8950
rect 6900 8840 7100 8850
rect 6900 8780 6910 8840
rect 7090 8780 7100 8840
rect 6900 8770 7100 8780
rect 7560 8840 7760 8850
rect 7560 8780 7570 8840
rect 7750 8780 7760 8840
rect 7560 8770 7760 8780
rect 8220 8840 8420 8850
rect 8220 8780 8230 8840
rect 8410 8780 8420 8840
rect 8220 8770 8420 8780
rect 6900 8630 7100 8710
rect 7560 8630 7760 8710
rect 8220 8630 8420 8710
rect 8620 8430 8680 9040
rect 8730 8530 8790 8540
rect 8730 8460 8790 8470
rect 8840 8430 8900 9040
rect 9100 9010 10620 9020
rect 9100 8950 9110 9010
rect 10610 8950 10620 9010
rect 9100 8940 10620 8950
rect 9100 8840 9300 8850
rect 9100 8780 9110 8840
rect 9290 8780 9300 8840
rect 9100 8770 9300 8780
rect 9760 8840 9960 8850
rect 9760 8780 9770 8840
rect 9950 8780 9960 8840
rect 9760 8770 9960 8780
rect 10420 8840 10620 8850
rect 10420 8780 10430 8840
rect 10610 8780 10620 8840
rect 10420 8770 10620 8780
rect 9100 8630 9300 8710
rect 9760 8630 9960 8710
rect 10420 8630 10620 8710
rect 10820 8430 10880 9040
rect 10930 8530 10990 8540
rect 10930 8460 10990 8470
rect 11040 8430 11100 9040
rect 11300 9010 12820 9020
rect 11300 8950 11310 9010
rect 12810 8950 12820 9010
rect 11300 8940 12820 8950
rect 11300 8840 11500 8850
rect 11300 8780 11310 8840
rect 11490 8780 11500 8840
rect 11300 8770 11500 8780
rect 11960 8840 12160 8850
rect 11960 8780 11970 8840
rect 12150 8780 12160 8840
rect 11960 8770 12160 8780
rect 12620 8840 12820 8850
rect 12620 8780 12630 8840
rect 12810 8780 12820 8840
rect 12620 8770 12820 8780
rect 11300 8630 11500 8710
rect 11960 8630 12160 8710
rect 12620 8630 12820 8710
rect 13020 8430 13080 9040
rect 13130 8530 13190 8540
rect 13130 8460 13190 8470
rect 13240 8430 13300 9040
rect 13500 9010 15020 9020
rect 13500 8950 13510 9010
rect 15010 8950 15020 9010
rect 13500 8940 15020 8950
rect 13500 8840 13700 8850
rect 13500 8780 13510 8840
rect 13690 8780 13700 8840
rect 13500 8770 13700 8780
rect 14160 8840 14360 8850
rect 14160 8780 14170 8840
rect 14350 8780 14360 8840
rect 14160 8770 14360 8780
rect 14820 8840 15020 8850
rect 14820 8780 14830 8840
rect 15010 8780 15020 8840
rect 14820 8770 15020 8780
rect 13500 8630 13700 8710
rect 14160 8630 14360 8710
rect 14820 8630 15020 8710
rect 15220 8430 15280 9040
rect 15330 8530 15390 8540
rect 15330 8460 15390 8470
rect 15440 8430 15500 9040
rect 15700 9010 17220 9020
rect 15700 8950 15710 9010
rect 17210 8950 17220 9010
rect 15700 8940 17220 8950
rect 15700 8770 15900 8850
rect 16360 8770 16560 8850
rect 17020 8770 17220 8850
rect 15700 8700 15900 8710
rect 15700 8640 15710 8700
rect 15890 8640 15900 8700
rect 15700 8630 15900 8640
rect 16360 8700 16560 8710
rect 16360 8640 16370 8700
rect 16550 8640 16560 8700
rect 16360 8630 16560 8640
rect 17020 8700 17220 8710
rect 17020 8640 17030 8700
rect 17210 8640 17220 8700
rect 17020 8630 17220 8640
rect 17420 8430 17480 9040
rect 17530 8530 17590 8540
rect 17530 8460 17590 8470
rect 17640 8430 17700 9040
rect 17900 8770 18100 8850
rect 18560 8770 18760 8850
rect 19220 8770 19420 8850
rect 17900 8700 18100 8710
rect 17900 8640 17910 8700
rect 18090 8640 18100 8700
rect 17900 8630 18100 8640
rect 18560 8700 18760 8710
rect 18560 8640 18570 8700
rect 18750 8640 18760 8700
rect 18560 8630 18760 8640
rect 19220 8700 19420 8710
rect 19220 8640 19230 8700
rect 19410 8640 19420 8700
rect 19220 8630 19420 8640
rect 1610 8410 1690 8420
rect 1610 8260 1620 8410
rect 1680 8260 1690 8410
rect 1610 8250 1690 8260
rect 1620 7620 1680 8250
rect 2010 8240 2090 8430
rect 2230 8240 2310 8430
rect 4210 8240 4290 8430
rect 4430 8310 4510 8430
rect 4430 8250 4440 8310
rect 4500 8250 4510 8310
rect 4430 8240 4510 8250
rect 6410 8310 6490 8430
rect 6410 8250 6420 8310
rect 6480 8250 6490 8310
rect 6410 8240 6490 8250
rect 6630 8420 6710 8430
rect 6630 8360 6640 8420
rect 6700 8360 6710 8420
rect 6630 8240 6710 8360
rect 8610 8420 8690 8430
rect 8610 8360 8620 8420
rect 8680 8360 8690 8420
rect 8610 8310 8690 8360
rect 8610 8250 8620 8310
rect 8680 8250 8690 8310
rect 8610 8240 8690 8250
rect 8830 8240 8910 8430
rect 10810 8420 10890 8430
rect 10810 8360 10820 8420
rect 10880 8360 10890 8420
rect 10810 8310 10890 8360
rect 10810 8250 10820 8310
rect 10880 8250 10890 8310
rect 10810 8240 10890 8250
rect 11030 8240 11110 8430
rect 13010 8420 13090 8430
rect 13010 8360 13020 8420
rect 13080 8360 13090 8420
rect 13010 8310 13090 8360
rect 13010 8250 13020 8310
rect 13080 8250 13090 8310
rect 13010 8240 13090 8250
rect 13230 8240 13310 8430
rect 15210 8420 15290 8430
rect 15210 8360 15220 8420
rect 15280 8360 15290 8420
rect 15210 8240 15290 8360
rect 15430 8310 15510 8430
rect 15430 8250 15440 8310
rect 15500 8250 15510 8310
rect 15430 8240 15510 8250
rect 17410 8240 17490 8430
rect 17630 8420 17710 8430
rect 17630 8360 17640 8420
rect 17700 8360 17710 8420
rect 19620 8410 19680 9040
rect 19730 8530 19790 8540
rect 19730 8460 19790 8470
rect 19840 8410 19900 9040
rect 17630 8240 17710 8360
rect 19610 8240 19690 8410
rect 19830 8240 19910 8410
rect 2020 7630 2080 8240
rect 2130 7730 2190 7740
rect 2130 7660 2190 7670
rect 2240 7630 2300 8240
rect 2500 7970 2700 8050
rect 3160 7970 3360 8050
rect 3820 7970 4020 8050
rect 2500 7900 2700 7910
rect 2500 7840 2510 7900
rect 2690 7840 2700 7900
rect 2500 7830 2700 7840
rect 3160 7900 3360 7910
rect 3160 7840 3170 7900
rect 3350 7840 3360 7900
rect 3160 7830 3360 7840
rect 3820 7900 4020 7910
rect 3820 7840 3830 7900
rect 4010 7840 4020 7900
rect 3820 7830 4020 7840
rect 4220 7630 4280 8240
rect 4330 7730 4390 7740
rect 4330 7660 4390 7670
rect 4440 7630 4500 8240
rect 4700 8210 6220 8220
rect 4700 8150 4710 8210
rect 6210 8150 6220 8210
rect 4700 8140 6220 8150
rect 4700 7970 4900 8050
rect 5360 7970 5560 8050
rect 6020 7970 6220 8050
rect 4700 7900 4900 7910
rect 4700 7840 4710 7900
rect 4890 7840 4900 7900
rect 4700 7830 4900 7840
rect 5360 7900 5560 7910
rect 5360 7840 5370 7900
rect 5550 7840 5560 7900
rect 5360 7830 5560 7840
rect 6020 7900 6220 7910
rect 6020 7840 6030 7900
rect 6210 7840 6220 7900
rect 6020 7830 6220 7840
rect 6420 7630 6480 8240
rect 6530 7730 6590 7740
rect 6530 7660 6590 7670
rect 6640 7630 6700 8240
rect 6900 8210 8420 8220
rect 6900 8150 6910 8210
rect 8410 8150 8420 8210
rect 6900 8140 8420 8150
rect 6900 8040 7100 8050
rect 6900 7980 6910 8040
rect 7090 7980 7100 8040
rect 6900 7970 7100 7980
rect 7560 8040 7760 8050
rect 7560 7980 7570 8040
rect 7750 7980 7760 8040
rect 7560 7970 7760 7980
rect 8220 8040 8420 8050
rect 8220 7980 8230 8040
rect 8410 7980 8420 8040
rect 8220 7970 8420 7980
rect 6900 7830 7100 7910
rect 7560 7830 7760 7910
rect 8220 7830 8420 7910
rect 8620 7630 8680 8240
rect 8730 7730 8790 7740
rect 8730 7660 8790 7670
rect 8840 7630 8900 8240
rect 9100 8210 10620 8220
rect 9100 8150 9110 8210
rect 10610 8150 10620 8210
rect 9100 8140 10620 8150
rect 9100 8040 9300 8050
rect 9100 7980 9110 8040
rect 9290 7980 9300 8040
rect 9100 7970 9300 7980
rect 9760 8040 9960 8050
rect 9760 7980 9770 8040
rect 9950 7980 9960 8040
rect 9760 7970 9960 7980
rect 10420 8040 10620 8050
rect 10420 7980 10430 8040
rect 10610 7980 10620 8040
rect 10420 7970 10620 7980
rect 9100 7830 9300 7910
rect 9760 7830 9960 7910
rect 10420 7830 10620 7910
rect 10820 7630 10880 8240
rect 10930 7730 10990 7740
rect 10930 7660 10990 7670
rect 11040 7630 11100 8240
rect 11300 8210 12820 8220
rect 11300 8150 11310 8210
rect 12810 8150 12820 8210
rect 11300 8140 12820 8150
rect 11300 8040 11500 8050
rect 11300 7980 11310 8040
rect 11490 7980 11500 8040
rect 11300 7970 11500 7980
rect 11960 8040 12160 8050
rect 11960 7980 11970 8040
rect 12150 7980 12160 8040
rect 11960 7970 12160 7980
rect 12620 8040 12820 8050
rect 12620 7980 12630 8040
rect 12810 7980 12820 8040
rect 12620 7970 12820 7980
rect 11300 7830 11500 7910
rect 11960 7830 12160 7910
rect 12620 7830 12820 7910
rect 13020 7630 13080 8240
rect 13130 7730 13190 7740
rect 13130 7660 13190 7670
rect 13240 7630 13300 8240
rect 13500 8210 15020 8220
rect 13500 8150 13510 8210
rect 15010 8150 15020 8210
rect 13500 8140 15020 8150
rect 13500 8040 13700 8050
rect 13500 7980 13510 8040
rect 13690 7980 13700 8040
rect 13500 7970 13700 7980
rect 14160 8040 14360 8050
rect 14160 7980 14170 8040
rect 14350 7980 14360 8040
rect 14160 7970 14360 7980
rect 14820 8040 15020 8050
rect 14820 7980 14830 8040
rect 15010 7980 15020 8040
rect 14820 7970 15020 7980
rect 13500 7830 13700 7910
rect 14160 7830 14360 7910
rect 14820 7830 15020 7910
rect 15220 7630 15280 8240
rect 15330 7730 15390 7740
rect 15330 7660 15390 7670
rect 15440 7630 15500 8240
rect 15700 8210 17220 8220
rect 15700 8150 15710 8210
rect 17210 8150 17220 8210
rect 15700 8140 17220 8150
rect 15700 7970 15900 8050
rect 16360 7970 16560 8050
rect 17020 7970 17220 8050
rect 15700 7900 15900 7910
rect 15700 7840 15710 7900
rect 15890 7840 15900 7900
rect 15700 7830 15900 7840
rect 16360 7900 16560 7910
rect 16360 7840 16370 7900
rect 16550 7840 16560 7900
rect 16360 7830 16560 7840
rect 17020 7900 17220 7910
rect 17020 7840 17030 7900
rect 17210 7840 17220 7900
rect 17020 7830 17220 7840
rect 17420 7630 17480 8240
rect 17530 7730 17590 7740
rect 17530 7660 17590 7670
rect 17640 7630 17700 8240
rect 17900 7970 18100 8050
rect 18560 7970 18760 8050
rect 19220 7970 19420 8050
rect 17900 7900 18100 7910
rect 17900 7840 17910 7900
rect 18090 7840 18100 7900
rect 17900 7830 18100 7840
rect 18560 7900 18760 7910
rect 18560 7840 18570 7900
rect 18750 7840 18760 7900
rect 18560 7830 18760 7840
rect 19220 7900 19420 7910
rect 19220 7840 19230 7900
rect 19410 7840 19420 7900
rect 19220 7830 19420 7840
rect 1610 7610 1690 7620
rect 1610 7460 1620 7610
rect 1680 7460 1690 7610
rect 1610 7450 1690 7460
rect 1410 6810 1490 6820
rect 1410 6660 1420 6810
rect 1480 6660 1490 6810
rect 1410 6650 1490 6660
rect 420 6590 620 6600
rect 420 6510 430 6590
rect 610 6510 620 6590
rect 420 6500 620 6510
rect 1420 4540 1480 6650
rect 1280 4530 1480 4540
rect 1280 4350 1290 4530
rect 1470 4350 1480 4530
rect 1280 4340 1480 4350
rect 1620 4140 1680 7450
rect 2010 7440 2090 7630
rect 2230 7440 2310 7630
rect 4210 7440 4290 7630
rect 4430 7510 4510 7630
rect 4430 7450 4440 7510
rect 4500 7450 4510 7510
rect 4430 7440 4510 7450
rect 6410 7510 6490 7630
rect 6410 7450 6420 7510
rect 6480 7450 6490 7510
rect 6410 7440 6490 7450
rect 6630 7620 6710 7630
rect 6630 7560 6640 7620
rect 6700 7560 6710 7620
rect 6630 7440 6710 7560
rect 8610 7620 8690 7630
rect 8610 7560 8620 7620
rect 8680 7560 8690 7620
rect 8610 7510 8690 7560
rect 8610 7450 8620 7510
rect 8680 7450 8690 7510
rect 8610 7440 8690 7450
rect 8830 7440 8910 7630
rect 10810 7620 10890 7630
rect 10810 7560 10820 7620
rect 10880 7560 10890 7620
rect 10810 7510 10890 7560
rect 10810 7450 10820 7510
rect 10880 7450 10890 7510
rect 10810 7440 10890 7450
rect 11030 7440 11110 7630
rect 13010 7620 13090 7630
rect 13010 7560 13020 7620
rect 13080 7560 13090 7620
rect 13010 7510 13090 7560
rect 13010 7450 13020 7510
rect 13080 7450 13090 7510
rect 13010 7440 13090 7450
rect 13230 7440 13310 7630
rect 15210 7620 15290 7630
rect 15210 7560 15220 7620
rect 15280 7560 15290 7620
rect 15210 7440 15290 7560
rect 15430 7510 15510 7630
rect 15430 7450 15440 7510
rect 15500 7450 15510 7510
rect 15430 7440 15510 7450
rect 17410 7440 17490 7630
rect 17630 7620 17710 7630
rect 17630 7560 17640 7620
rect 17700 7560 17710 7620
rect 19620 7610 19680 8240
rect 19730 7730 19790 7740
rect 19730 7660 19790 7670
rect 19840 7610 19900 8240
rect 17630 7440 17710 7560
rect 19610 7440 19690 7610
rect 19830 7440 19910 7610
rect 2020 6830 2080 7440
rect 2130 6930 2190 6940
rect 2130 6860 2190 6870
rect 2240 6830 2300 7440
rect 2500 7240 2700 7250
rect 2500 7180 2510 7240
rect 2690 7180 2700 7240
rect 2500 7170 2700 7180
rect 3160 7240 3360 7250
rect 3160 7180 3170 7240
rect 3350 7180 3360 7240
rect 3160 7170 3360 7180
rect 3820 7240 4020 7250
rect 3820 7180 3830 7240
rect 4010 7180 4020 7240
rect 3820 7170 4020 7180
rect 2500 7030 2700 7110
rect 3160 7030 3360 7110
rect 3820 7030 4020 7110
rect 4220 6830 4280 7440
rect 4330 6930 4390 6940
rect 4330 6860 4390 6870
rect 4440 6830 4500 7440
rect 4700 7410 6220 7420
rect 4700 7350 4710 7410
rect 6210 7350 6220 7410
rect 4700 7340 6220 7350
rect 4700 7240 4900 7250
rect 4700 7180 4710 7240
rect 4890 7180 4900 7240
rect 4700 7170 4900 7180
rect 5360 7240 5560 7250
rect 5360 7180 5370 7240
rect 5550 7180 5560 7240
rect 5360 7170 5560 7180
rect 6020 7240 6220 7250
rect 6020 7180 6030 7240
rect 6210 7180 6220 7240
rect 6020 7170 6220 7180
rect 4700 7030 4900 7110
rect 5360 7030 5560 7110
rect 6020 7030 6220 7110
rect 6420 6830 6480 7440
rect 6530 6930 6590 6940
rect 6530 6860 6590 6870
rect 6640 6830 6700 7440
rect 6900 7410 8420 7420
rect 6900 7350 6910 7410
rect 8410 7350 8420 7410
rect 6900 7340 8420 7350
rect 6900 7170 7100 7250
rect 7560 7170 7760 7250
rect 8220 7170 8420 7250
rect 6900 7100 7100 7110
rect 6900 7040 6910 7100
rect 7090 7040 7100 7100
rect 6900 7030 7100 7040
rect 7560 7100 7760 7110
rect 7560 7040 7570 7100
rect 7750 7040 7760 7100
rect 7560 7030 7760 7040
rect 8220 7100 8420 7110
rect 8220 7040 8230 7100
rect 8410 7040 8420 7100
rect 8220 7030 8420 7040
rect 8620 6830 8680 7440
rect 8730 6930 8790 6940
rect 8730 6860 8790 6870
rect 8840 6830 8900 7440
rect 9100 7410 10620 7420
rect 9100 7350 9110 7410
rect 10610 7350 10620 7410
rect 9100 7340 10620 7350
rect 9100 7170 9300 7250
rect 9760 7170 9960 7250
rect 10420 7170 10620 7250
rect 9100 7100 9300 7110
rect 9100 7040 9110 7100
rect 9290 7040 9300 7100
rect 9100 7030 9300 7040
rect 9760 7100 9960 7110
rect 9760 7040 9770 7100
rect 9950 7040 9960 7100
rect 9760 7030 9960 7040
rect 10420 7100 10620 7110
rect 10420 7040 10430 7100
rect 10610 7040 10620 7100
rect 10420 7030 10620 7040
rect 10820 6830 10880 7440
rect 10930 6930 10990 6940
rect 10930 6860 10990 6870
rect 11040 6830 11100 7440
rect 11300 7410 12820 7420
rect 11300 7350 11310 7410
rect 12810 7350 12820 7410
rect 11300 7340 12820 7350
rect 11300 7170 11500 7250
rect 11960 7170 12160 7250
rect 12620 7170 12820 7250
rect 11300 7100 11500 7110
rect 11300 7040 11310 7100
rect 11490 7040 11500 7100
rect 11300 7030 11500 7040
rect 11960 7100 12160 7110
rect 11960 7040 11970 7100
rect 12150 7040 12160 7100
rect 11960 7030 12160 7040
rect 12620 7100 12820 7110
rect 12620 7040 12630 7100
rect 12810 7040 12820 7100
rect 12620 7030 12820 7040
rect 13020 6830 13080 7440
rect 13130 6930 13190 6940
rect 13130 6860 13190 6870
rect 13240 6830 13300 7440
rect 13500 7410 15020 7420
rect 13500 7350 13510 7410
rect 15010 7350 15020 7410
rect 13500 7340 15020 7350
rect 13500 7170 13700 7250
rect 14160 7170 14360 7250
rect 14820 7170 15020 7250
rect 13500 7100 13700 7110
rect 13500 7040 13510 7100
rect 13690 7040 13700 7100
rect 13500 7030 13700 7040
rect 14160 7100 14360 7110
rect 14160 7040 14170 7100
rect 14350 7040 14360 7100
rect 14160 7030 14360 7040
rect 14820 7100 15020 7110
rect 14820 7040 14830 7100
rect 15010 7040 15020 7100
rect 14820 7030 15020 7040
rect 15220 6830 15280 7440
rect 15330 6930 15390 6940
rect 15330 6860 15390 6870
rect 15440 6830 15500 7440
rect 15700 7410 17220 7420
rect 15700 7350 15710 7410
rect 17210 7350 17220 7410
rect 15700 7340 17220 7350
rect 15700 7240 15900 7250
rect 15700 7180 15710 7240
rect 15890 7180 15900 7240
rect 15700 7170 15900 7180
rect 16360 7240 16560 7250
rect 16360 7180 16370 7240
rect 16550 7180 16560 7240
rect 16360 7170 16560 7180
rect 17020 7240 17220 7250
rect 17020 7180 17030 7240
rect 17210 7180 17220 7240
rect 17020 7170 17220 7180
rect 15700 7030 15900 7110
rect 16360 7030 16560 7110
rect 17020 7030 17220 7110
rect 17420 6830 17480 7440
rect 17530 6930 17590 6940
rect 17530 6860 17590 6870
rect 17640 6830 17700 7440
rect 17900 7240 18100 7250
rect 17900 7180 17910 7240
rect 18090 7180 18100 7240
rect 17900 7170 18100 7180
rect 18560 7240 18760 7250
rect 18560 7180 18570 7240
rect 18750 7180 18760 7240
rect 18560 7170 18760 7180
rect 19220 7240 19420 7250
rect 19220 7180 19230 7240
rect 19410 7180 19420 7240
rect 19220 7170 19420 7180
rect 17900 7030 18100 7110
rect 18560 7030 18760 7110
rect 19220 7030 19420 7110
rect 2010 6640 2090 6830
rect 2230 6640 2310 6830
rect 4210 6710 4290 6830
rect 4210 6650 4220 6710
rect 4280 6650 4290 6710
rect 4210 6640 4290 6650
rect 4430 6640 4510 6830
rect 6410 6820 6490 6830
rect 6410 6760 6420 6820
rect 6480 6760 6490 6820
rect 6410 6640 6490 6760
rect 6630 6710 6710 6830
rect 6630 6650 6640 6710
rect 6700 6650 6710 6710
rect 6630 6640 6710 6650
rect 8610 6640 8690 6830
rect 8830 6820 8910 6830
rect 8830 6760 8840 6820
rect 8900 6760 8910 6820
rect 8830 6710 8910 6760
rect 8830 6650 8840 6710
rect 8900 6650 8910 6710
rect 8830 6640 8910 6650
rect 10810 6640 10890 6830
rect 11030 6820 11110 6830
rect 11030 6760 11040 6820
rect 11100 6760 11110 6820
rect 11030 6710 11110 6760
rect 11030 6650 11040 6710
rect 11100 6650 11110 6710
rect 11030 6640 11110 6650
rect 13010 6640 13090 6830
rect 13230 6820 13310 6830
rect 13230 6760 13240 6820
rect 13300 6760 13310 6820
rect 13230 6710 13310 6760
rect 13230 6650 13240 6710
rect 13300 6650 13310 6710
rect 13230 6640 13310 6650
rect 15210 6710 15290 6830
rect 15210 6650 15220 6710
rect 15280 6650 15290 6710
rect 15210 6640 15290 6650
rect 15430 6820 15510 6830
rect 15430 6760 15440 6820
rect 15500 6760 15510 6820
rect 15430 6640 15510 6760
rect 17410 6820 17490 6830
rect 17410 6760 17420 6820
rect 17480 6760 17490 6820
rect 17410 6640 17490 6760
rect 17630 6640 17710 6830
rect 19620 6810 19680 7440
rect 19730 6930 19790 6940
rect 19730 6860 19790 6870
rect 19840 6810 19900 7440
rect 20240 6910 20300 9140
rect 20440 8510 20500 9310
rect 21930 9260 21990 9270
rect 21300 8990 21500 9000
rect 21300 8910 21310 8990
rect 21490 8910 21500 8990
rect 21300 8900 21500 8910
rect 21930 8530 21990 8540
rect 20430 8500 20510 8510
rect 20430 8350 20440 8500
rect 20500 8350 20510 8500
rect 21930 8460 21990 8470
rect 20430 8340 20510 8350
rect 20440 7710 20500 8340
rect 21300 8190 21500 8200
rect 21300 8110 21310 8190
rect 21490 8110 21500 8190
rect 21300 8100 21500 8110
rect 21930 7730 21990 7740
rect 20430 7700 20510 7710
rect 20430 7550 20440 7700
rect 20500 7550 20510 7700
rect 21930 7660 21990 7670
rect 20430 7540 20510 7550
rect 20230 6900 20310 6910
rect 19610 6640 19690 6810
rect 19830 6640 19910 6810
rect 20230 6750 20240 6900
rect 20300 6750 20310 6900
rect 20230 6740 20310 6750
rect 2020 6030 2080 6640
rect 2130 6130 2190 6140
rect 2130 6060 2190 6070
rect 2240 6030 2300 6640
rect 2500 6370 2700 6450
rect 3160 6370 3360 6450
rect 3820 6370 4020 6450
rect 2500 6300 2700 6310
rect 2500 6240 2510 6300
rect 2690 6240 2700 6300
rect 2500 6230 2700 6240
rect 3160 6300 3360 6310
rect 3160 6240 3170 6300
rect 3350 6240 3360 6300
rect 3160 6230 3360 6240
rect 3820 6300 4020 6310
rect 3820 6240 3830 6300
rect 4010 6240 4020 6300
rect 3820 6230 4020 6240
rect 4220 6030 4280 6640
rect 4330 6130 4390 6140
rect 4330 6060 4390 6070
rect 4440 6030 4500 6640
rect 4700 6610 6220 6620
rect 4700 6550 4710 6610
rect 6210 6550 6220 6610
rect 4700 6540 6220 6550
rect 4700 6370 4900 6450
rect 5360 6370 5560 6450
rect 6020 6370 6220 6450
rect 4700 6300 4900 6310
rect 4700 6240 4710 6300
rect 4890 6240 4900 6300
rect 4700 6230 4900 6240
rect 5360 6300 5560 6310
rect 5360 6240 5370 6300
rect 5550 6240 5560 6300
rect 5360 6230 5560 6240
rect 6020 6300 6220 6310
rect 6020 6240 6030 6300
rect 6210 6240 6220 6300
rect 6020 6230 6220 6240
rect 6420 6030 6480 6640
rect 6530 6130 6590 6140
rect 6530 6060 6590 6070
rect 6640 6030 6700 6640
rect 6900 6610 8420 6620
rect 6900 6550 6910 6610
rect 8410 6550 8420 6610
rect 6900 6540 8420 6550
rect 6900 6440 7100 6450
rect 6900 6380 6910 6440
rect 7090 6380 7100 6440
rect 6900 6370 7100 6380
rect 7560 6440 7760 6450
rect 7560 6380 7570 6440
rect 7750 6380 7760 6440
rect 7560 6370 7760 6380
rect 8220 6440 8420 6450
rect 8220 6380 8230 6440
rect 8410 6380 8420 6440
rect 8220 6370 8420 6380
rect 6900 6230 7100 6310
rect 7560 6230 7760 6310
rect 8220 6230 8420 6310
rect 8620 6030 8680 6640
rect 8730 6130 8790 6140
rect 8730 6060 8790 6070
rect 8840 6030 8900 6640
rect 9100 6610 10620 6620
rect 9100 6550 9110 6610
rect 10610 6550 10620 6610
rect 9100 6540 10620 6550
rect 9100 6440 9300 6450
rect 9100 6380 9110 6440
rect 9290 6380 9300 6440
rect 9100 6370 9300 6380
rect 9760 6440 9960 6450
rect 9760 6380 9770 6440
rect 9950 6380 9960 6440
rect 9760 6370 9960 6380
rect 10420 6440 10620 6450
rect 10420 6380 10430 6440
rect 10610 6380 10620 6440
rect 10420 6370 10620 6380
rect 9100 6230 9300 6310
rect 9760 6230 9960 6310
rect 10420 6230 10620 6310
rect 10820 6030 10880 6640
rect 10930 6130 10990 6140
rect 10930 6060 10990 6070
rect 11040 6030 11100 6640
rect 11300 6610 12820 6620
rect 11300 6550 11310 6610
rect 12810 6550 12820 6610
rect 11300 6540 12820 6550
rect 11300 6440 11500 6450
rect 11300 6380 11310 6440
rect 11490 6380 11500 6440
rect 11300 6370 11500 6380
rect 11960 6440 12160 6450
rect 11960 6380 11970 6440
rect 12150 6380 12160 6440
rect 11960 6370 12160 6380
rect 12620 6440 12820 6450
rect 12620 6380 12630 6440
rect 12810 6380 12820 6440
rect 12620 6370 12820 6380
rect 11300 6230 11500 6310
rect 11960 6230 12160 6310
rect 12620 6230 12820 6310
rect 13020 6030 13080 6640
rect 13130 6130 13190 6140
rect 13130 6060 13190 6070
rect 13240 6030 13300 6640
rect 13500 6610 15020 6620
rect 13500 6550 13510 6610
rect 15010 6550 15020 6610
rect 13500 6540 15020 6550
rect 13500 6440 13700 6450
rect 13500 6380 13510 6440
rect 13690 6380 13700 6440
rect 13500 6370 13700 6380
rect 14160 6440 14360 6450
rect 14160 6380 14170 6440
rect 14350 6380 14360 6440
rect 14160 6370 14360 6380
rect 14820 6440 15020 6450
rect 14820 6380 14830 6440
rect 15010 6380 15020 6440
rect 14820 6370 15020 6380
rect 13500 6230 13700 6310
rect 14160 6230 14360 6310
rect 14820 6230 15020 6310
rect 15220 6030 15280 6640
rect 15330 6130 15390 6140
rect 15330 6060 15390 6070
rect 15440 6030 15500 6640
rect 15700 6610 17220 6620
rect 15700 6550 15710 6610
rect 17210 6550 17220 6610
rect 15700 6540 17220 6550
rect 15700 6370 15900 6450
rect 16360 6370 16560 6450
rect 17020 6370 17220 6450
rect 15700 6300 15900 6310
rect 15700 6240 15710 6300
rect 15890 6240 15900 6300
rect 15700 6230 15900 6240
rect 16360 6300 16560 6310
rect 16360 6240 16370 6300
rect 16550 6240 16560 6300
rect 16360 6230 16560 6240
rect 17020 6300 17220 6310
rect 17020 6240 17030 6300
rect 17210 6240 17220 6300
rect 17020 6230 17220 6240
rect 17420 6030 17480 6640
rect 17530 6130 17590 6140
rect 17530 6060 17590 6070
rect 17640 6030 17700 6640
rect 17900 6370 18100 6450
rect 18560 6370 18760 6450
rect 19220 6370 19420 6450
rect 17900 6300 18100 6310
rect 17900 6240 17910 6300
rect 18090 6240 18100 6300
rect 17900 6230 18100 6240
rect 18560 6300 18760 6310
rect 18560 6240 18570 6300
rect 18750 6240 18760 6300
rect 18560 6230 18760 6240
rect 19220 6300 19420 6310
rect 19220 6240 19230 6300
rect 19410 6240 19420 6300
rect 19220 6230 19420 6240
rect 2010 5840 2090 6030
rect 2230 5910 2310 6030
rect 2230 5850 2240 5910
rect 2300 5850 2310 5910
rect 2230 5840 2310 5850
rect 4210 5840 4290 6030
rect 4430 6020 4510 6030
rect 4430 5960 4440 6020
rect 4500 5960 4510 6020
rect 4430 5910 4510 5960
rect 4430 5850 4440 5910
rect 4500 5850 4510 5910
rect 4430 5840 4510 5850
rect 6410 5910 6490 6030
rect 6410 5850 6420 5910
rect 6480 5850 6490 5910
rect 6410 5840 6490 5850
rect 6630 6020 6710 6030
rect 6630 5960 6640 6020
rect 6700 5960 6710 6020
rect 6630 5840 6710 5960
rect 8610 6020 8690 6030
rect 8610 5960 8620 6020
rect 8680 5960 8690 6020
rect 8610 5910 8690 5960
rect 8610 5850 8620 5910
rect 8680 5850 8690 5910
rect 8610 5840 8690 5850
rect 8830 5840 8910 6030
rect 10810 6020 10890 6030
rect 10810 5960 10820 6020
rect 10880 5960 10890 6020
rect 10810 5910 10890 5960
rect 10810 5850 10820 5910
rect 10880 5850 10890 5910
rect 10810 5840 10890 5850
rect 11030 5840 11110 6030
rect 13010 6020 13090 6030
rect 13010 5960 13020 6020
rect 13080 5960 13090 6020
rect 13010 5910 13090 5960
rect 13010 5850 13020 5910
rect 13080 5850 13090 5910
rect 13010 5840 13090 5850
rect 13230 5840 13310 6030
rect 15210 6020 15290 6030
rect 15210 5960 15220 6020
rect 15280 5960 15290 6020
rect 15210 5840 15290 5960
rect 15430 5910 15510 6030
rect 15430 5850 15440 5910
rect 15500 5850 15510 5910
rect 15430 5840 15510 5850
rect 17410 5840 17490 6030
rect 17630 6020 17710 6030
rect 17630 5960 17640 6020
rect 17700 5960 17710 6020
rect 19620 6010 19680 6640
rect 19730 6130 19790 6140
rect 19730 6060 19790 6070
rect 19840 6010 19900 6640
rect 17630 5910 17710 5960
rect 17630 5850 17640 5910
rect 17700 5850 17710 5910
rect 17630 5840 17710 5850
rect 19610 5840 19690 6010
rect 19830 6000 19910 6010
rect 19830 5940 19840 6000
rect 19900 5940 19910 6000
rect 19830 5840 19910 5940
rect 2020 5230 2080 5840
rect 2130 5330 2190 5340
rect 2130 5260 2190 5270
rect 2240 5230 2300 5840
rect 2500 5810 4020 5820
rect 2500 5750 2510 5810
rect 4010 5750 4020 5810
rect 2500 5740 4020 5750
rect 2500 5640 2700 5650
rect 2500 5580 2510 5640
rect 2690 5580 2700 5640
rect 2500 5570 2700 5580
rect 3160 5640 3360 5650
rect 3160 5580 3170 5640
rect 3350 5580 3360 5640
rect 3160 5570 3360 5580
rect 3820 5640 4020 5650
rect 3820 5580 3830 5640
rect 4010 5580 4020 5640
rect 3820 5570 4020 5580
rect 2500 5430 2700 5510
rect 3160 5430 3360 5510
rect 3820 5430 4020 5510
rect 4220 5230 4280 5840
rect 4330 5330 4390 5340
rect 4330 5260 4390 5270
rect 4440 5230 4500 5840
rect 4700 5810 6220 5820
rect 4700 5750 4710 5810
rect 6210 5750 6220 5810
rect 4700 5740 6220 5750
rect 4700 5640 4900 5650
rect 4700 5580 4710 5640
rect 4890 5580 4900 5640
rect 4700 5570 4900 5580
rect 5360 5640 5560 5650
rect 5360 5580 5370 5640
rect 5550 5580 5560 5640
rect 5360 5570 5560 5580
rect 6020 5640 6220 5650
rect 6020 5580 6030 5640
rect 6210 5580 6220 5640
rect 6020 5570 6220 5580
rect 4700 5430 4900 5510
rect 5360 5430 5560 5510
rect 6020 5430 6220 5510
rect 6420 5230 6480 5840
rect 6530 5330 6590 5340
rect 6530 5260 6590 5270
rect 6640 5230 6700 5840
rect 6900 5810 8420 5820
rect 6900 5750 6910 5810
rect 8410 5750 8420 5810
rect 6900 5740 8420 5750
rect 6900 5570 7100 5650
rect 7560 5570 7760 5650
rect 8220 5570 8420 5650
rect 6900 5500 7100 5510
rect 6900 5440 6910 5500
rect 7090 5440 7100 5500
rect 6900 5430 7100 5440
rect 7560 5500 7760 5510
rect 7560 5440 7570 5500
rect 7750 5440 7760 5500
rect 7560 5430 7760 5440
rect 8220 5500 8420 5510
rect 8220 5440 8230 5500
rect 8410 5440 8420 5500
rect 8220 5430 8420 5440
rect 8620 5230 8680 5840
rect 8730 5330 8790 5340
rect 8730 5260 8790 5270
rect 8840 5230 8900 5840
rect 9100 5810 10620 5820
rect 9100 5750 9110 5810
rect 10610 5750 10620 5810
rect 9100 5740 10620 5750
rect 9100 5570 9300 5650
rect 9760 5570 9960 5650
rect 10420 5570 10620 5650
rect 9100 5500 9300 5510
rect 9100 5440 9110 5500
rect 9290 5440 9300 5500
rect 9100 5430 9300 5440
rect 9760 5500 9960 5510
rect 9760 5440 9770 5500
rect 9950 5440 9960 5500
rect 9760 5430 9960 5440
rect 10420 5500 10620 5510
rect 10420 5440 10430 5500
rect 10610 5440 10620 5500
rect 10420 5430 10620 5440
rect 10820 5230 10880 5840
rect 10930 5330 10990 5340
rect 10930 5260 10990 5270
rect 11040 5230 11100 5840
rect 11300 5810 12820 5820
rect 11300 5750 11310 5810
rect 12810 5750 12820 5810
rect 11300 5740 12820 5750
rect 11300 5570 11500 5650
rect 11960 5570 12160 5650
rect 12620 5570 12820 5650
rect 11300 5500 11500 5510
rect 11300 5440 11310 5500
rect 11490 5440 11500 5500
rect 11300 5430 11500 5440
rect 11960 5500 12160 5510
rect 11960 5440 11970 5500
rect 12150 5440 12160 5500
rect 11960 5430 12160 5440
rect 12620 5500 12820 5510
rect 12620 5440 12630 5500
rect 12810 5440 12820 5500
rect 12620 5430 12820 5440
rect 13020 5230 13080 5840
rect 13130 5330 13190 5340
rect 13130 5260 13190 5270
rect 13240 5230 13300 5840
rect 13500 5810 15020 5820
rect 13500 5750 13510 5810
rect 15010 5750 15020 5810
rect 13500 5740 15020 5750
rect 13500 5570 13700 5650
rect 14160 5570 14360 5650
rect 14820 5570 15020 5650
rect 13500 5500 13700 5510
rect 13500 5440 13510 5500
rect 13690 5440 13700 5500
rect 13500 5430 13700 5440
rect 14160 5500 14360 5510
rect 14160 5440 14170 5500
rect 14350 5440 14360 5500
rect 14160 5430 14360 5440
rect 14820 5500 15020 5510
rect 14820 5440 14830 5500
rect 15010 5440 15020 5500
rect 14820 5430 15020 5440
rect 15220 5230 15280 5840
rect 15330 5330 15390 5340
rect 15330 5260 15390 5270
rect 15440 5230 15500 5840
rect 15700 5810 17220 5820
rect 15700 5750 15710 5810
rect 17210 5750 17220 5810
rect 15700 5740 17220 5750
rect 15700 5640 15900 5650
rect 15700 5580 15710 5640
rect 15890 5580 15900 5640
rect 15700 5570 15900 5580
rect 16360 5640 16560 5650
rect 16360 5580 16370 5640
rect 16550 5580 16560 5640
rect 16360 5570 16560 5580
rect 17020 5640 17220 5650
rect 17020 5580 17030 5640
rect 17210 5580 17220 5640
rect 17020 5570 17220 5580
rect 15700 5430 15900 5510
rect 16360 5430 16560 5510
rect 17020 5430 17220 5510
rect 17420 5230 17480 5840
rect 17530 5330 17590 5340
rect 17530 5260 17590 5270
rect 17640 5230 17700 5840
rect 17900 5810 19420 5820
rect 17900 5750 17910 5810
rect 19410 5750 19420 5810
rect 17900 5740 19420 5750
rect 17900 5640 18100 5650
rect 17900 5580 17910 5640
rect 18090 5580 18100 5640
rect 17900 5570 18100 5580
rect 18560 5640 18760 5650
rect 18560 5580 18570 5640
rect 18750 5580 18760 5640
rect 18560 5570 18760 5580
rect 19220 5640 19420 5650
rect 19220 5580 19230 5640
rect 19410 5580 19420 5640
rect 19220 5570 19420 5580
rect 17900 5430 18100 5510
rect 18560 5430 18760 5510
rect 19220 5430 19420 5510
rect 2010 5110 2090 5230
rect 2010 5050 2020 5110
rect 2080 5050 2090 5110
rect 2010 5040 2090 5050
rect 2230 5040 2310 5230
rect 4210 5220 4290 5230
rect 4210 5160 4220 5220
rect 4280 5160 4290 5220
rect 4210 5110 4290 5160
rect 4210 5050 4220 5110
rect 4280 5050 4290 5110
rect 4210 5040 4290 5050
rect 4430 5040 4510 5230
rect 6410 5220 6490 5230
rect 6410 5160 6420 5220
rect 6480 5160 6490 5220
rect 6410 5040 6490 5160
rect 6630 5110 6710 5230
rect 6630 5050 6640 5110
rect 6700 5050 6710 5110
rect 6630 5040 6710 5050
rect 8610 5040 8690 5230
rect 8830 5220 8910 5230
rect 8830 5160 8840 5220
rect 8900 5160 8910 5220
rect 8830 5110 8910 5160
rect 8830 5050 8840 5110
rect 8900 5050 8910 5110
rect 8830 5040 8910 5050
rect 10810 5040 10890 5230
rect 11030 5220 11110 5230
rect 11030 5160 11040 5220
rect 11100 5160 11110 5220
rect 11030 5110 11110 5160
rect 11030 5050 11040 5110
rect 11100 5050 11110 5110
rect 11030 5040 11110 5050
rect 13010 5040 13090 5230
rect 13230 5220 13310 5230
rect 13230 5160 13240 5220
rect 13300 5160 13310 5220
rect 13230 5110 13310 5160
rect 13230 5050 13240 5110
rect 13300 5050 13310 5110
rect 13230 5040 13310 5050
rect 15210 5110 15290 5230
rect 15210 5050 15220 5110
rect 15280 5050 15290 5110
rect 15210 5040 15290 5050
rect 15430 5220 15510 5230
rect 15430 5160 15440 5220
rect 15500 5160 15510 5220
rect 15430 5040 15510 5160
rect 17410 5220 17490 5230
rect 17410 5160 17420 5220
rect 17480 5160 17490 5220
rect 17410 5110 17490 5160
rect 17410 5050 17420 5110
rect 17480 5050 17490 5110
rect 17410 5040 17490 5050
rect 17630 5040 17710 5230
rect 19620 5210 19680 5840
rect 19730 5330 19790 5340
rect 19730 5260 19790 5270
rect 19840 5210 19900 5840
rect 19610 5200 19690 5210
rect 19610 5140 19620 5200
rect 19680 5140 19690 5200
rect 19610 5040 19690 5140
rect 19830 5040 19910 5210
rect 2020 4830 2080 5040
rect 2240 4830 2300 5040
rect 2500 5010 4020 5020
rect 2500 4950 2510 5010
rect 4010 4950 4020 5010
rect 2500 4940 4020 4950
rect 4220 4830 4280 5040
rect 4440 4830 4500 5040
rect 4700 5010 6220 5020
rect 4700 4950 4710 5010
rect 6210 4950 6220 5010
rect 4700 4940 6220 4950
rect 6420 4830 6480 5040
rect 6640 4830 6700 5040
rect 6900 5010 8420 5020
rect 6900 4950 6910 5010
rect 8410 4950 8420 5010
rect 6900 4940 8420 4950
rect 7790 4680 7950 4690
rect 7790 4540 7800 4680
rect 7940 4540 7950 4680
rect 7790 4530 7950 4540
rect 1620 4130 1820 4140
rect 1620 3950 1630 4130
rect 1810 3950 1820 4130
rect 1620 3940 1820 3950
rect 1160 3330 1340 3340
rect 1160 3150 1170 3330
rect 1330 3150 1340 3330
rect 1160 3140 1340 3150
rect 2760 3330 2940 3340
rect 2760 3150 2770 3330
rect 2930 3150 2940 3330
rect 2760 3140 2940 3150
rect 4360 3330 4540 3340
rect 4360 3150 4370 3330
rect 4530 3150 4540 3330
rect 4360 3140 4540 3150
rect 5960 3330 6140 3340
rect 5960 3150 5970 3330
rect 6130 3150 6140 3330
rect 5960 3140 6140 3150
rect 7560 3330 7740 3340
rect 7560 3150 7570 3330
rect 7730 3150 7740 3330
rect 7560 3140 7740 3150
rect 470 2220 670 2240
rect 470 -4780 480 2220
rect 660 -4780 670 2220
rect 1200 690 1300 3140
rect 2100 2250 2240 2260
rect 2100 2090 2110 2250
rect 2230 2090 2240 2250
rect 2100 1990 2240 2090
rect 2100 1310 2110 1990
rect 2230 1310 2240 1990
rect 1420 1160 1520 1180
rect 1400 1150 1540 1160
rect 1400 1030 1410 1150
rect 1530 1030 1540 1150
rect 1400 1020 1540 1030
rect 1180 680 1320 690
rect 1180 560 1190 680
rect 1310 560 1320 680
rect 1180 550 1320 560
rect 1200 -1110 1300 550
rect 1420 -640 1520 1020
rect 2100 450 2240 1310
rect 2800 690 2900 3140
rect 3700 2250 3840 2260
rect 3700 2090 3710 2250
rect 3830 2090 3840 2250
rect 3700 1990 3840 2090
rect 3700 1310 3710 1990
rect 3830 1310 3840 1990
rect 3020 1160 3120 1180
rect 3000 1150 3140 1160
rect 3000 1030 3010 1150
rect 3130 1030 3140 1150
rect 3000 1020 3140 1030
rect 2780 680 2920 690
rect 2780 560 2790 680
rect 2910 560 2920 680
rect 2780 550 2920 560
rect 2100 290 2110 450
rect 2230 290 2240 450
rect 2100 190 2240 290
rect 2100 -490 2110 190
rect 2230 -490 2240 190
rect 1400 -650 1540 -640
rect 1400 -770 1410 -650
rect 1530 -770 1540 -650
rect 1400 -780 1540 -770
rect 1180 -1120 1320 -1110
rect 1180 -1240 1190 -1120
rect 1310 -1240 1320 -1120
rect 1180 -1250 1320 -1240
rect 1200 -2910 1300 -1250
rect 1420 -2440 1520 -780
rect 2100 -1350 2240 -490
rect 2800 -1110 2900 550
rect 3020 -640 3120 1020
rect 3700 450 3840 1310
rect 4400 690 4500 3140
rect 5300 2250 5440 2260
rect 5300 2090 5310 2250
rect 5430 2090 5440 2250
rect 5300 1990 5440 2090
rect 5300 1310 5310 1990
rect 5430 1310 5440 1990
rect 4620 1160 4720 1180
rect 4600 1150 4740 1160
rect 4600 1030 4610 1150
rect 4730 1030 4740 1150
rect 4600 1020 4740 1030
rect 4380 680 4520 690
rect 4380 560 4390 680
rect 4510 560 4520 680
rect 4380 550 4520 560
rect 3700 290 3710 450
rect 3830 290 3840 450
rect 3700 190 3840 290
rect 3700 -490 3710 190
rect 3830 -490 3840 190
rect 3000 -650 3140 -640
rect 3000 -770 3010 -650
rect 3130 -770 3140 -650
rect 3000 -780 3140 -770
rect 2780 -1120 2920 -1110
rect 2780 -1240 2790 -1120
rect 2910 -1240 2920 -1120
rect 2780 -1250 2920 -1240
rect 2100 -1510 2110 -1350
rect 2230 -1510 2240 -1350
rect 2100 -1610 2240 -1510
rect 2100 -2290 2110 -1610
rect 2230 -2290 2240 -1610
rect 1400 -2450 1540 -2440
rect 1400 -2570 1410 -2450
rect 1530 -2570 1540 -2450
rect 1400 -2580 1540 -2570
rect 1180 -2920 1320 -2910
rect 1180 -3040 1190 -2920
rect 1310 -3040 1320 -2920
rect 1180 -3050 1320 -3040
rect 1200 -4710 1300 -3050
rect 1420 -4240 1520 -2580
rect 2100 -3150 2240 -2290
rect 2800 -2910 2900 -1250
rect 3020 -2440 3120 -780
rect 3700 -1350 3840 -490
rect 4400 -1110 4500 550
rect 4620 -640 4720 1020
rect 5300 450 5440 1310
rect 6000 690 6100 3140
rect 6900 2250 7040 2260
rect 6900 2090 6910 2250
rect 7030 2090 7040 2250
rect 6900 1990 7040 2090
rect 6900 1310 6910 1990
rect 7030 1310 7040 1990
rect 6220 1160 6320 1180
rect 6200 1150 6340 1160
rect 6200 1030 6210 1150
rect 6330 1030 6340 1150
rect 6200 1020 6340 1030
rect 5980 680 6120 690
rect 5980 560 5990 680
rect 6110 560 6120 680
rect 5980 550 6120 560
rect 5300 290 5310 450
rect 5430 290 5440 450
rect 5300 190 5440 290
rect 5300 -490 5310 190
rect 5430 -490 5440 190
rect 4600 -650 4740 -640
rect 4600 -770 4610 -650
rect 4730 -770 4740 -650
rect 4600 -780 4740 -770
rect 4380 -1120 4520 -1110
rect 4380 -1240 4390 -1120
rect 4510 -1240 4520 -1120
rect 4380 -1250 4520 -1240
rect 3700 -1510 3710 -1350
rect 3830 -1510 3840 -1350
rect 3700 -1610 3840 -1510
rect 3700 -2290 3710 -1610
rect 3830 -2290 3840 -1610
rect 3000 -2450 3140 -2440
rect 3000 -2570 3010 -2450
rect 3130 -2570 3140 -2450
rect 3000 -2580 3140 -2570
rect 2780 -2920 2920 -2910
rect 2780 -3040 2790 -2920
rect 2910 -3040 2920 -2920
rect 2780 -3050 2920 -3040
rect 2100 -3310 2110 -3150
rect 2230 -3310 2240 -3150
rect 2100 -3410 2240 -3310
rect 2100 -4090 2110 -3410
rect 2230 -4090 2240 -3410
rect 2100 -4100 2240 -4090
rect 1400 -4250 1540 -4240
rect 1400 -4370 1410 -4250
rect 1530 -4370 1540 -4250
rect 1400 -4380 1540 -4370
rect 1420 -4400 1520 -4380
rect 2800 -4710 2900 -3050
rect 3020 -4240 3120 -2580
rect 3700 -3150 3840 -2290
rect 4400 -2910 4500 -1250
rect 4620 -2440 4720 -780
rect 5300 -1350 5440 -490
rect 6000 -1110 6100 550
rect 6220 -640 6320 1020
rect 6900 450 7040 1310
rect 7600 690 7700 3140
rect 7820 2940 7920 4530
rect 8620 4430 8680 5040
rect 8840 4430 8900 5040
rect 9100 5010 10620 5020
rect 9100 4950 9110 5010
rect 10610 4950 10620 5010
rect 9100 4940 10620 4950
rect 10820 4430 10880 5040
rect 11040 4430 11100 5040
rect 11300 5010 12820 5020
rect 11300 4950 11310 5010
rect 12810 4950 12820 5010
rect 11300 4940 12820 4950
rect 13020 4430 13080 5040
rect 13240 4430 13300 5040
rect 13500 5010 15020 5020
rect 13500 4950 13510 5010
rect 15010 4950 15020 5010
rect 13500 4940 15020 4950
rect 15220 4830 15280 5040
rect 15440 4830 15500 5040
rect 15700 5010 17220 5020
rect 15700 4950 15710 5010
rect 17210 4950 17220 5010
rect 15700 4940 17220 4950
rect 17420 4830 17480 5040
rect 17640 4830 17700 5040
rect 17900 5010 19420 5020
rect 17900 4950 17910 5010
rect 19410 4950 19420 5010
rect 17900 4940 19420 4950
rect 19620 4830 19680 5040
rect 19840 4830 19900 5040
rect 20240 4540 20300 6740
rect 20100 4530 20300 4540
rect 8610 4310 8690 4430
rect 8610 4250 8620 4310
rect 8680 4250 8690 4310
rect 8610 4240 8690 4250
rect 8830 4240 8910 4430
rect 10810 4420 10890 4430
rect 10810 4360 10820 4420
rect 10880 4360 10890 4420
rect 10810 4240 10890 4360
rect 11030 4310 11110 4430
rect 11030 4250 11040 4310
rect 11100 4250 11110 4310
rect 11030 4240 11110 4250
rect 13010 4240 13090 4430
rect 13230 4420 13310 4430
rect 13230 4360 13240 4420
rect 13300 4360 13310 4420
rect 13230 4240 13310 4360
rect 20100 4350 20110 4530
rect 20290 4350 20300 4530
rect 20100 4340 20300 4350
rect 8620 4230 8680 4240
rect 8840 4230 8900 4240
rect 10820 4230 10880 4240
rect 11040 4230 11100 4240
rect 13020 4230 13080 4240
rect 13240 4230 13300 4240
rect 20440 4140 20500 7540
rect 21300 7390 21500 7400
rect 21300 7310 21310 7390
rect 21490 7310 21500 7390
rect 21300 7300 21500 7310
rect 21930 6930 21990 6940
rect 21930 6860 21990 6870
rect 21300 6590 21500 6600
rect 21300 6510 21310 6590
rect 21490 6510 21500 6590
rect 21300 6500 21500 6510
rect 21930 6130 21990 6140
rect 21930 6060 21990 6070
rect 21930 5330 21990 5340
rect 21930 5260 21990 5270
rect 23040 4970 23590 4980
rect 23040 4600 23050 4970
rect 23580 4600 23590 4970
rect 23040 4590 23590 4600
rect 20440 4130 20640 4140
rect 10880 4100 11040 4110
rect 10880 3960 10890 4100
rect 11030 3960 11040 4100
rect 10880 3950 11040 3960
rect 20440 3950 20450 4130
rect 20630 3950 20640 4130
rect 9160 3330 9340 3340
rect 9160 3150 9170 3330
rect 9330 3150 9340 3330
rect 9160 3140 9340 3150
rect 7800 2930 7940 2940
rect 7800 2810 7810 2930
rect 7930 2810 7940 2930
rect 7820 2540 7920 2810
rect 8500 2250 8640 2260
rect 8500 2090 8510 2250
rect 8630 2090 8640 2250
rect 8500 1990 8640 2090
rect 8500 1310 8510 1990
rect 8630 1310 8640 1990
rect 7820 1160 7920 1180
rect 7800 1150 7940 1160
rect 7800 1030 7810 1150
rect 7930 1030 7940 1150
rect 7800 1020 7940 1030
rect 7580 680 7720 690
rect 7580 560 7590 680
rect 7710 560 7720 680
rect 7580 550 7720 560
rect 6900 290 6910 450
rect 7030 290 7040 450
rect 6900 190 7040 290
rect 6900 -490 6910 190
rect 7030 -490 7040 190
rect 6200 -650 6340 -640
rect 6200 -770 6210 -650
rect 6330 -770 6340 -650
rect 6200 -780 6340 -770
rect 5980 -1120 6120 -1110
rect 5980 -1240 5990 -1120
rect 6110 -1240 6120 -1120
rect 5980 -1250 6120 -1240
rect 5300 -1510 5310 -1350
rect 5430 -1510 5440 -1350
rect 5300 -1610 5440 -1510
rect 5300 -2290 5310 -1610
rect 5430 -2290 5440 -1610
rect 4600 -2450 4740 -2440
rect 4600 -2570 4610 -2450
rect 4730 -2570 4740 -2450
rect 4600 -2580 4740 -2570
rect 4380 -2920 4520 -2910
rect 4380 -3040 4390 -2920
rect 4510 -3040 4520 -2920
rect 4380 -3050 4520 -3040
rect 3700 -3310 3710 -3150
rect 3830 -3310 3840 -3150
rect 3700 -3410 3840 -3310
rect 3700 -4090 3710 -3410
rect 3830 -4090 3840 -3410
rect 3700 -4100 3840 -4090
rect 3000 -4250 3140 -4240
rect 3000 -4370 3010 -4250
rect 3130 -4370 3140 -4250
rect 3000 -4380 3140 -4370
rect 3020 -4400 3120 -4380
rect 4400 -4710 4500 -3050
rect 4620 -4240 4720 -2580
rect 5300 -3150 5440 -2290
rect 6000 -2910 6100 -1250
rect 6220 -2440 6320 -780
rect 6900 -1350 7040 -490
rect 7600 -1110 7700 550
rect 7820 -640 7920 1020
rect 8500 450 8640 1310
rect 9200 690 9300 3140
rect 10910 3020 11010 3950
rect 20440 3940 20640 3950
rect 23210 3090 23410 4590
rect 26590 3360 26790 11490
rect 27250 11400 27260 11490
rect 27320 11400 27330 11490
rect 27250 11390 27330 11400
rect 27260 11180 27320 11390
rect 27250 11170 27330 11180
rect 27250 11080 27260 11170
rect 27320 11080 27330 11170
rect 27250 11070 27330 11080
rect 27260 10865 27320 11070
rect 27250 10855 27330 10865
rect 27250 10765 27260 10855
rect 27320 10765 27330 10855
rect 27250 10755 27330 10765
rect 27260 9415 27320 10755
rect 27380 10300 27440 11480
rect 27370 10290 27450 10300
rect 27370 10200 27380 10290
rect 27440 10200 27450 10290
rect 27370 10190 27450 10200
rect 27380 9985 27440 10190
rect 27370 9975 27450 9985
rect 27370 9885 27380 9975
rect 27440 9885 27450 9975
rect 27370 9875 27450 9885
rect 27250 9405 27330 9415
rect 27250 9315 27260 9405
rect 27320 9315 27330 9405
rect 27250 9305 27330 9315
rect 27260 9100 27320 9305
rect 27250 9090 27330 9100
rect 27250 9000 27260 9090
rect 27320 9000 27330 9090
rect 27250 8990 27330 9000
rect 27260 8785 27320 8990
rect 27250 8775 27330 8785
rect 27250 8685 27260 8775
rect 27320 8685 27330 8775
rect 27250 8675 27330 8685
rect 27260 8380 27320 8675
rect 27250 8370 27330 8380
rect 27250 8280 27260 8370
rect 27320 8280 27330 8370
rect 27250 8270 27330 8280
rect 27260 8060 27320 8270
rect 27250 8050 27330 8060
rect 27250 7960 27260 8050
rect 27320 7960 27330 8050
rect 27250 7950 27330 7960
rect 27260 7750 27320 7950
rect 27250 7740 27330 7750
rect 27250 7650 27260 7740
rect 27320 7650 27330 7740
rect 27250 7640 27330 7650
rect 27260 5250 27320 7640
rect 27380 7340 27440 9875
rect 27500 9260 27560 11480
rect 27490 9250 27570 9260
rect 27490 9160 27500 9250
rect 27560 9160 27570 9250
rect 27490 9150 27570 9160
rect 27500 8945 27560 9150
rect 27490 8935 27570 8945
rect 27490 8845 27500 8935
rect 27560 8845 27570 8935
rect 27490 8835 27570 8845
rect 27370 7330 27450 7340
rect 27370 7240 27380 7330
rect 27440 7240 27450 7330
rect 27370 7230 27450 7240
rect 27380 7025 27440 7230
rect 27370 7015 27450 7025
rect 27370 6925 27380 7015
rect 27440 6925 27450 7015
rect 27370 6915 27450 6925
rect 27380 6710 27440 6915
rect 27370 6700 27450 6710
rect 27370 6610 27380 6700
rect 27440 6610 27450 6700
rect 27370 6600 27450 6610
rect 27380 6300 27440 6600
rect 27370 6290 27450 6300
rect 27370 6200 27380 6290
rect 27440 6200 27450 6290
rect 27370 6190 27450 6200
rect 27380 5985 27440 6190
rect 27500 6140 27560 8835
rect 27620 8220 27680 11480
rect 27740 11340 27800 11480
rect 30570 11418 30670 11532
rect 30148 11416 30670 11418
rect 30148 11364 30154 11416
rect 30288 11364 30670 11416
rect 30148 11362 30670 11364
rect 27730 11330 27810 11340
rect 27730 11240 27740 11330
rect 27800 11240 27810 11330
rect 30570 11326 30670 11362
rect 31472 11722 31542 11728
rect 31472 11536 31478 11722
rect 31536 11536 31542 11722
rect 30570 11320 31414 11326
rect 30180 11270 30400 11280
rect 27730 11230 27810 11240
rect 28770 11260 28850 11270
rect 27740 11025 27800 11230
rect 28770 11040 28780 11260
rect 28840 11040 28850 11260
rect 29270 11190 29520 11200
rect 29270 11120 29280 11190
rect 29510 11120 29520 11190
rect 30180 11190 30190 11270
rect 30390 11190 30400 11270
rect 30570 11262 30600 11320
rect 30738 11262 31270 11320
rect 31408 11262 31414 11320
rect 30570 11256 31414 11262
rect 31472 11210 31542 11536
rect 30180 11180 30400 11190
rect 31280 11200 31542 11210
rect 29270 11110 29520 11120
rect 28770 11030 28850 11040
rect 28950 11040 29200 11050
rect 27730 11015 27810 11025
rect 27730 10925 27740 11015
rect 27800 10925 27810 11015
rect 28950 10970 28960 11040
rect 29190 10970 29200 11040
rect 28950 10960 29200 10970
rect 27730 10915 27810 10925
rect 27740 10460 27800 10915
rect 28860 10880 28940 10890
rect 28860 10710 28870 10880
rect 28930 10710 28940 10880
rect 28860 10700 28940 10710
rect 27730 10450 27810 10460
rect 27730 10360 27740 10450
rect 27800 10360 27810 10450
rect 27730 10350 27810 10360
rect 27740 10140 27800 10350
rect 27730 10130 27810 10140
rect 27730 10040 27740 10130
rect 27800 10040 27810 10130
rect 27730 10030 27810 10040
rect 27740 9825 27800 10030
rect 27730 9815 27810 9825
rect 27730 9725 27740 9815
rect 27800 9725 27810 9815
rect 27730 9715 27810 9725
rect 28880 9170 28940 10700
rect 29010 10740 29090 10750
rect 29010 10570 29020 10740
rect 29080 10570 29090 10740
rect 29010 10560 29090 10570
rect 28870 9160 28950 9170
rect 28870 8940 28880 9160
rect 28940 8940 28950 9160
rect 28870 8930 28950 8940
rect 27610 8210 27690 8220
rect 27610 8120 27620 8210
rect 27680 8120 27690 8210
rect 27610 8110 27690 8120
rect 27620 7900 27680 8110
rect 27610 7890 27690 7900
rect 27610 7800 27620 7890
rect 27680 7800 27690 7890
rect 27610 7790 27690 7800
rect 27620 7180 27680 7790
rect 27610 7170 27690 7180
rect 27610 7080 27620 7170
rect 27680 7080 27690 7170
rect 28880 7090 28940 8930
rect 29010 8120 29070 10560
rect 29140 10200 29200 10960
rect 29130 10190 29210 10200
rect 29130 9970 29140 10190
rect 29200 9970 29210 10190
rect 29130 9960 29210 9970
rect 29000 8110 29080 8120
rect 29000 7890 29010 8110
rect 29070 7890 29080 8110
rect 29000 7880 29080 7890
rect 27610 7070 27690 7080
rect 28870 7080 28950 7090
rect 27620 6865 27680 7070
rect 27610 6855 27690 6865
rect 27610 6765 27620 6855
rect 27680 6765 27690 6855
rect 28870 6860 28880 7080
rect 28940 6860 28950 7080
rect 28870 6850 28950 6860
rect 27610 6755 27690 6765
rect 27490 6130 27570 6140
rect 27490 6040 27500 6130
rect 27560 6040 27570 6130
rect 27490 6030 27570 6040
rect 27370 5975 27450 5985
rect 27370 5885 27380 5975
rect 27440 5885 27450 5975
rect 27370 5875 27450 5885
rect 27380 5670 27440 5875
rect 27500 5825 27560 6030
rect 27490 5815 27570 5825
rect 27490 5725 27500 5815
rect 27560 5725 27570 5815
rect 27490 5715 27570 5725
rect 27370 5660 27450 5670
rect 27370 5570 27380 5660
rect 27440 5570 27450 5660
rect 27370 5560 27450 5570
rect 27170 5240 27320 5250
rect 27170 5110 27180 5240
rect 27310 5110 27320 5240
rect 27170 5100 27320 5110
rect 27380 5000 27440 5560
rect 27240 4930 27440 5000
rect 27240 4750 27250 4930
rect 27430 4750 27440 4930
rect 27240 4740 27440 4750
rect 27500 4600 27560 5715
rect 27360 4530 27560 4600
rect 27360 4350 27370 4530
rect 27550 4350 27560 4530
rect 27360 4340 27560 4350
rect 27620 4200 27680 6755
rect 29010 6050 29070 7880
rect 29000 6040 29080 6050
rect 29000 5820 29010 6040
rect 29070 5820 29080 6040
rect 29000 5810 29080 5820
rect 29140 4530 29200 9960
rect 29130 4520 29210 4530
rect 29130 4290 29140 4520
rect 29200 4290 29210 4520
rect 29130 4280 29210 4290
rect 29270 4270 29330 11110
rect 30310 10190 30390 11180
rect 31280 11110 31290 11200
rect 31530 11110 31542 11200
rect 31280 11100 31542 11110
rect 31472 10900 31542 11100
rect 31472 10514 31478 10900
rect 31536 10514 31542 10900
rect 31472 10508 31542 10514
rect 31684 11720 31754 11726
rect 31684 11534 31690 11720
rect 31748 11534 31754 11720
rect 31684 10900 31754 11534
rect 32770 11722 32870 11728
rect 32770 11532 32776 11722
rect 32864 11532 32870 11722
rect 32770 11418 32870 11532
rect 32348 11416 32870 11418
rect 32348 11364 32354 11416
rect 32488 11364 32870 11416
rect 32348 11362 32870 11364
rect 32770 11326 32870 11362
rect 33672 11722 33742 11728
rect 33672 11536 33678 11722
rect 33736 11536 33742 11722
rect 32770 11320 33614 11326
rect 32380 11270 32600 11280
rect 32380 11190 32390 11270
rect 32590 11190 32600 11270
rect 32770 11262 32800 11320
rect 32938 11262 33470 11320
rect 33608 11262 33614 11320
rect 32770 11256 33614 11262
rect 32380 11180 32600 11190
rect 31684 10514 31690 10900
rect 31748 10514 31754 10900
rect 31684 10508 31754 10514
rect 30290 10180 30410 10190
rect 30290 10080 30300 10180
rect 30400 10080 30410 10180
rect 30290 10070 30410 10080
rect 32390 10010 32470 11180
rect 33672 11070 33742 11536
rect 33480 11060 33742 11070
rect 33480 10970 33490 11060
rect 33730 10970 33742 11060
rect 33480 10960 33742 10970
rect 33672 10900 33742 10960
rect 33672 10514 33678 10900
rect 33736 10514 33742 10900
rect 33672 10508 33742 10514
rect 33884 11720 33954 11726
rect 33884 11534 33890 11720
rect 33948 11534 33954 11720
rect 33884 10900 33954 11534
rect 34970 11722 35070 11728
rect 34970 11532 34976 11722
rect 35064 11532 35070 11722
rect 34970 11418 35070 11532
rect 34548 11416 35070 11418
rect 34548 11364 34554 11416
rect 34688 11364 35070 11416
rect 34548 11362 35070 11364
rect 34970 11326 35070 11362
rect 35872 11722 35942 11728
rect 35872 11536 35878 11722
rect 35936 11536 35942 11722
rect 34970 11320 35814 11326
rect 34560 11270 34780 11280
rect 34560 11190 34570 11270
rect 34770 11190 34780 11270
rect 34970 11262 35000 11320
rect 35138 11262 35670 11320
rect 35808 11262 35814 11320
rect 34970 11256 35814 11262
rect 34560 11180 34780 11190
rect 33884 10514 33890 10900
rect 33948 10514 33954 10900
rect 33884 10508 33954 10514
rect 32370 10000 32490 10010
rect 32370 9900 32380 10000
rect 32480 9900 32490 10000
rect 32370 9890 32490 9900
rect 34570 9830 34650 11180
rect 35872 10930 35942 11536
rect 36084 11720 36154 11726
rect 36084 11534 36090 11720
rect 36148 11534 36154 11720
rect 35690 10920 35950 10930
rect 35690 10830 35700 10920
rect 35940 10830 35950 10920
rect 35690 10820 35878 10830
rect 35872 10514 35878 10820
rect 35936 10820 35950 10830
rect 36084 10900 36154 11534
rect 36470 11510 36480 11980
rect 36810 11510 36820 11980
rect 36470 11500 36820 11510
rect 35936 10514 35942 10820
rect 36084 10750 36090 10900
rect 36080 10640 36090 10750
rect 36148 10750 36154 10900
rect 36148 10740 36340 10750
rect 36330 10650 36340 10740
rect 35872 10508 35942 10514
rect 36084 10514 36090 10640
rect 36148 10640 36340 10650
rect 36148 10514 36154 10640
rect 36084 10508 36154 10514
rect 34550 9820 34670 9830
rect 34550 9720 34560 9820
rect 34660 9720 34670 9820
rect 34550 9710 34670 9720
rect 31450 9410 31680 9420
rect 31450 9220 31460 9410
rect 31670 9220 31680 9410
rect 31450 9210 31680 9220
rect 32060 9120 32210 9130
rect 31440 8990 31690 9000
rect 31440 8780 31450 8990
rect 31680 8780 31690 8990
rect 32060 8990 32070 9120
rect 32200 8990 32210 9120
rect 32060 8980 32210 8990
rect 31440 8770 31690 8780
rect 30560 8580 30650 8590
rect 30560 8210 30570 8580
rect 30640 8210 30650 8580
rect 30560 7940 30650 8210
rect 32090 8130 32180 8980
rect 34490 8940 35530 8950
rect 34490 8880 34500 8940
rect 35520 8880 35530 8940
rect 34490 8870 35530 8880
rect 30880 8120 32180 8130
rect 30880 8030 30890 8120
rect 31280 8030 32180 8120
rect 30880 8020 32180 8030
rect 33660 8830 33780 8840
rect 33660 8030 33670 8830
rect 33770 8030 33780 8830
rect 34540 8610 34600 8870
rect 34960 8610 35020 8870
rect 35370 8620 35430 8870
rect 35340 8610 35460 8620
rect 34500 8600 34620 8610
rect 34500 8440 34510 8600
rect 34610 8440 34620 8600
rect 34500 8430 34620 8440
rect 34920 8600 35040 8610
rect 34920 8440 34930 8600
rect 35030 8440 35040 8600
rect 35340 8450 35350 8610
rect 35450 8450 35460 8610
rect 35340 8440 35460 8450
rect 34920 8430 35040 8440
rect 33660 8020 33780 8030
rect 34740 8180 34900 8190
rect 30560 7570 30570 7940
rect 30640 7570 30650 7940
rect 30560 7160 30650 7570
rect 30460 7150 30790 7160
rect 30460 7050 30470 7150
rect 30850 7090 30870 7150
rect 30850 7050 30860 7090
rect 30460 7040 30860 7050
rect 30110 6470 31510 6480
rect 30110 6410 30120 6470
rect 30420 6410 31510 6470
rect 30110 6400 31510 6410
rect 30110 6310 31390 6320
rect 30110 6250 31080 6310
rect 31380 6250 31390 6310
rect 30110 6240 31390 6250
rect 30110 5740 30190 6240
rect 31430 5750 31510 6400
rect 31370 5740 31570 5750
rect 30050 5730 30250 5740
rect 30050 5670 30060 5730
rect 30240 5670 30250 5730
rect 31370 5680 31380 5740
rect 31560 5680 31570 5740
rect 31370 5670 31570 5680
rect 30050 5660 30250 5670
rect 30030 5170 30330 5180
rect 30030 5070 30040 5170
rect 30320 5070 30330 5170
rect 30030 5060 30330 5070
rect 29760 4710 30560 4720
rect 29760 4640 29770 4710
rect 30550 4640 30560 4710
rect 29760 4630 30560 4640
rect 29270 4260 29520 4270
rect 27620 4130 27820 4200
rect 29270 4190 29280 4260
rect 29510 4190 29520 4260
rect 29270 4180 29520 4190
rect 27620 3950 27630 4130
rect 27810 3950 27820 4130
rect 27620 3940 27820 3950
rect 30070 4040 30270 4050
rect 30070 3860 30080 4040
rect 30260 3860 30270 4040
rect 30070 3850 30270 3860
rect 31670 4040 31870 4050
rect 31670 3860 31680 4040
rect 31860 3860 31870 4040
rect 31670 3850 31870 3860
rect 32090 3750 32180 8020
rect 32290 7970 32470 7980
rect 32290 7890 32300 7970
rect 32460 7890 32470 7970
rect 32290 7880 32470 7890
rect 32250 7770 32330 7780
rect 32250 7570 32260 7770
rect 32320 7570 32330 7770
rect 32250 7560 32330 7570
rect 32260 4890 32320 7560
rect 32410 4890 32470 7880
rect 33670 7940 33770 8020
rect 34280 7990 34370 8000
rect 34280 7940 34290 7990
rect 33670 7840 34290 7940
rect 34360 7940 34370 7990
rect 34740 7960 34750 8180
rect 34890 7960 34900 8180
rect 34740 7950 34900 7960
rect 35160 7980 35320 7990
rect 34360 7930 34620 7940
rect 34610 7850 34620 7930
rect 34280 7790 34290 7840
rect 34360 7840 34620 7850
rect 34360 7790 34370 7840
rect 34280 7780 34370 7790
rect 35160 7760 35170 7980
rect 35310 7760 35320 7980
rect 35160 7750 35320 7760
rect 34490 7310 34610 7320
rect 34490 7150 34500 7310
rect 34600 7150 34610 7310
rect 34490 7140 34610 7150
rect 34910 7310 35030 7320
rect 34910 7150 34920 7310
rect 35020 7150 35030 7310
rect 34910 7140 35030 7150
rect 35330 7310 35450 7320
rect 35330 7150 35340 7310
rect 35440 7150 35450 7310
rect 35330 7140 35450 7150
rect 33450 6990 33600 7000
rect 33450 6980 33460 6990
rect 32560 6940 33460 6980
rect 32560 5520 32620 6940
rect 33450 6930 33460 6940
rect 33590 6980 33600 6990
rect 33690 6990 33920 7000
rect 33690 6980 33700 6990
rect 33590 6940 33700 6980
rect 33590 6930 33600 6940
rect 33450 6920 33600 6930
rect 33690 6930 33700 6940
rect 33910 6980 33920 6990
rect 34010 6990 34200 7000
rect 34010 6980 34020 6990
rect 33910 6940 34020 6980
rect 33910 6930 33920 6940
rect 33690 6920 33920 6930
rect 34010 6930 34020 6940
rect 34190 6930 34200 6990
rect 34520 6930 34590 7140
rect 34940 6930 35010 7140
rect 35360 6930 35430 7140
rect 34010 6920 34200 6930
rect 34490 6920 35550 6930
rect 34490 6830 34500 6920
rect 35540 6830 35550 6920
rect 34490 6820 35550 6830
rect 36220 6260 36420 6270
rect 36220 6080 36230 6260
rect 36410 6080 36420 6260
rect 36220 6070 36420 6080
rect 36520 6260 36720 6270
rect 36520 6080 36530 6260
rect 36710 6080 36720 6260
rect 36520 6070 36720 6080
rect 36290 5890 36400 5900
rect 36290 5820 36300 5890
rect 36390 5820 36400 5890
rect 36290 5630 36400 5820
rect 36290 5560 36300 5630
rect 36390 5560 36400 5630
rect 32550 5510 32630 5520
rect 32550 5280 32560 5510
rect 32620 5280 32630 5510
rect 36290 5370 36400 5560
rect 32550 5270 32630 5280
rect 33320 5290 33640 5300
rect 33320 5020 33330 5290
rect 33630 5020 33640 5290
rect 33320 5010 33640 5020
rect 36290 5040 36300 5370
rect 36390 5040 36400 5370
rect 32250 4880 32330 4890
rect 32250 4650 32260 4880
rect 32320 4650 32330 4880
rect 32250 4640 32330 4650
rect 32400 4880 32480 4890
rect 32400 4650 32410 4880
rect 32470 4650 32480 4880
rect 32400 4640 32480 4650
rect 36290 4850 36400 5040
rect 36290 4780 36300 4850
rect 36390 4780 36400 4850
rect 36290 4590 36400 4780
rect 36290 4520 36300 4590
rect 36390 4520 36400 4590
rect 32490 4480 32650 4490
rect 32490 4340 32500 4480
rect 32640 4340 32650 4480
rect 32490 4330 32650 4340
rect 34080 4480 34240 4490
rect 34080 4340 34090 4480
rect 34230 4340 34240 4480
rect 34080 4330 34240 4340
rect 36290 4330 36400 4520
rect 32070 3740 32220 3750
rect 31520 3730 31700 3740
rect 31520 3550 31530 3730
rect 31690 3550 31700 3730
rect 32070 3610 32080 3740
rect 32210 3610 32220 3740
rect 32070 3600 32220 3610
rect 31520 3540 31700 3550
rect 26590 3220 26620 3360
rect 26760 3220 26790 3360
rect 26590 3210 26790 3220
rect 14180 3030 14360 3040
rect 10880 3010 11040 3020
rect 10880 2870 10890 3010
rect 11030 2870 11040 3010
rect 10880 2860 11040 2870
rect 14180 2870 14190 3030
rect 14350 2870 14360 3030
rect 14180 2860 14360 2870
rect 18050 3010 18210 3020
rect 18050 2870 18060 3010
rect 18200 2870 18210 3010
rect 23210 2910 23220 3090
rect 23400 2910 23410 3090
rect 23210 2900 23410 2910
rect 18050 2860 18210 2870
rect 11690 2770 11850 2780
rect 11690 2620 11700 2770
rect 11840 2620 11850 2770
rect 11690 2610 11850 2620
rect 10990 2540 11150 2550
rect 10990 2400 11000 2540
rect 11140 2400 11150 2540
rect 10990 2390 11150 2400
rect 10100 2250 10240 2260
rect 10100 2090 10110 2250
rect 10230 2090 10240 2250
rect 10100 1990 10240 2090
rect 10100 1310 10110 1990
rect 10230 1310 10240 1990
rect 11020 1960 11120 2390
rect 11700 2250 11840 2610
rect 12590 2540 12750 2550
rect 12590 2400 12600 2540
rect 12740 2400 12750 2540
rect 12590 2390 12750 2400
rect 13970 2540 14130 2550
rect 13970 2400 13980 2540
rect 14120 2400 14130 2540
rect 13970 2390 14130 2400
rect 11700 2090 11710 2250
rect 11830 2090 11840 2250
rect 11020 1950 11160 1960
rect 11020 1330 11030 1950
rect 11150 1330 11160 1950
rect 11020 1320 11160 1330
rect 9420 1160 9520 1180
rect 9400 1150 9540 1160
rect 9400 1030 9410 1150
rect 9530 1030 9540 1150
rect 9400 1020 9540 1030
rect 9180 680 9320 690
rect 9180 560 9190 680
rect 9310 560 9320 680
rect 9180 550 9320 560
rect 8500 290 8510 450
rect 8630 290 8640 450
rect 8500 190 8640 290
rect 8500 -490 8510 190
rect 8630 -490 8640 190
rect 7800 -650 7940 -640
rect 7800 -770 7810 -650
rect 7930 -770 7940 -650
rect 7800 -780 7940 -770
rect 7580 -1120 7720 -1110
rect 7580 -1240 7590 -1120
rect 7710 -1240 7720 -1120
rect 7580 -1250 7720 -1240
rect 6900 -1510 6910 -1350
rect 7030 -1510 7040 -1350
rect 6900 -1610 7040 -1510
rect 6900 -2290 6910 -1610
rect 7030 -2290 7040 -1610
rect 6200 -2450 6340 -2440
rect 6200 -2570 6210 -2450
rect 6330 -2570 6340 -2450
rect 6200 -2580 6340 -2570
rect 5980 -2920 6120 -2910
rect 5980 -3040 5990 -2920
rect 6110 -3040 6120 -2920
rect 5980 -3050 6120 -3040
rect 5300 -3310 5310 -3150
rect 5430 -3310 5440 -3150
rect 5300 -3410 5440 -3310
rect 5300 -4090 5310 -3410
rect 5430 -4090 5440 -3410
rect 5300 -4100 5440 -4090
rect 4600 -4250 4740 -4240
rect 4600 -4370 4610 -4250
rect 4730 -4370 4740 -4250
rect 4600 -4380 4740 -4370
rect 4620 -4400 4720 -4380
rect 6000 -4710 6100 -3050
rect 6220 -4240 6320 -2580
rect 6900 -3150 7040 -2290
rect 7600 -2910 7700 -1250
rect 7820 -2440 7920 -780
rect 8500 -1350 8640 -490
rect 9200 -1110 9300 550
rect 9420 -640 9520 1020
rect 10100 450 10240 1310
rect 11700 1240 11840 2090
rect 12620 1960 12720 2390
rect 13300 2250 13440 2260
rect 13300 2090 13310 2250
rect 13430 2090 13440 2250
rect 12600 1950 12740 1960
rect 12600 1330 12610 1950
rect 12730 1330 12740 1950
rect 12600 1320 12740 1330
rect 11240 1230 11840 1240
rect 11240 1070 11250 1230
rect 11670 1070 11840 1230
rect 11240 1060 11840 1070
rect 10100 290 10110 450
rect 10230 290 10240 450
rect 10100 190 10240 290
rect 10100 -490 10110 190
rect 10230 -490 10240 190
rect 9400 -650 9540 -640
rect 9400 -770 9410 -650
rect 9530 -770 9540 -650
rect 9400 -780 9540 -770
rect 9180 -1120 9320 -1110
rect 9180 -1240 9190 -1120
rect 9310 -1240 9320 -1120
rect 9180 -1250 9320 -1240
rect 8500 -1510 8510 -1350
rect 8630 -1510 8640 -1350
rect 8500 -1610 8640 -1510
rect 8500 -2290 8510 -1610
rect 8630 -2290 8640 -1610
rect 7800 -2450 7940 -2440
rect 7800 -2570 7810 -2450
rect 7930 -2570 7940 -2450
rect 7800 -2580 7940 -2570
rect 7580 -2920 7720 -2910
rect 7580 -3040 7590 -2920
rect 7710 -3040 7720 -2920
rect 7580 -3050 7720 -3040
rect 6900 -3310 6910 -3150
rect 7030 -3310 7040 -3150
rect 6900 -3410 7040 -3310
rect 6900 -4090 6910 -3410
rect 7030 -4090 7040 -3410
rect 6900 -4100 7040 -4090
rect 6200 -4250 6340 -4240
rect 6200 -4370 6210 -4250
rect 6330 -4370 6340 -4250
rect 6200 -4380 6340 -4370
rect 6220 -4400 6320 -4380
rect 7600 -4710 7700 -3050
rect 7820 -4240 7920 -2580
rect 8500 -3150 8640 -2290
rect 9200 -2910 9300 -1250
rect 9420 -2440 9520 -780
rect 10100 -1350 10240 -490
rect 11700 450 11840 1060
rect 12380 870 12520 880
rect 12380 750 12390 870
rect 12510 750 12520 870
rect 12380 740 12520 750
rect 11700 290 11710 450
rect 11830 290 11840 450
rect 11700 190 11840 290
rect 11700 -560 11710 190
rect 11260 -570 11710 -560
rect 11830 -560 11840 190
rect 11830 -570 12280 -560
rect 11260 -730 11270 -570
rect 12270 -730 12280 -570
rect 12400 -640 12500 740
rect 11260 -740 12280 -730
rect 12380 -650 12520 -640
rect 10100 -1510 10110 -1350
rect 10230 -1510 10240 -1350
rect 10100 -1610 10240 -1510
rect 10100 -2290 10110 -1610
rect 10230 -2290 10240 -1610
rect 9400 -2450 9540 -2440
rect 9400 -2570 9410 -2450
rect 9530 -2570 9540 -2450
rect 9400 -2580 9540 -2570
rect 9180 -2920 9320 -2910
rect 9180 -3040 9190 -2920
rect 9310 -3040 9320 -2920
rect 9180 -3050 9320 -3040
rect 8500 -3310 8510 -3150
rect 8630 -3310 8640 -3150
rect 8500 -3410 8640 -3310
rect 8500 -4090 8510 -3410
rect 8630 -4090 8640 -3410
rect 8500 -4100 8640 -4090
rect 7800 -4250 7940 -4240
rect 7800 -4370 7810 -4250
rect 7930 -4370 7940 -4250
rect 7800 -4380 7940 -4370
rect 7820 -4400 7920 -4380
rect 9200 -4710 9300 -3050
rect 9420 -4240 9520 -2580
rect 10100 -3150 10240 -2290
rect 11700 -1350 11840 -740
rect 12380 -810 12390 -650
rect 12510 -810 12520 -650
rect 12380 -980 12520 -810
rect 12380 -1050 12390 -980
rect 12510 -1050 12520 -980
rect 12380 -1060 12520 -1050
rect 12620 -710 12720 1320
rect 13300 450 13440 2090
rect 14000 1960 14100 2390
rect 13980 1950 14120 1960
rect 13980 1330 13990 1950
rect 14110 1330 14120 1950
rect 13980 1320 14120 1330
rect 13300 290 13310 450
rect 13430 290 13440 450
rect 13300 190 13440 290
rect 13300 -490 13310 190
rect 13430 -490 13440 190
rect 12620 -920 12721 -710
rect 12620 -930 12760 -920
rect 11700 -1510 11710 -1350
rect 11830 -1510 11840 -1350
rect 11700 -1610 11840 -1510
rect 11700 -2290 11710 -1610
rect 11830 -2290 11840 -1610
rect 11020 -2910 11120 -2900
rect 11000 -2920 11140 -2910
rect 11000 -3040 11010 -2920
rect 11130 -3040 11140 -2920
rect 11000 -3050 11140 -3040
rect 10100 -3310 10110 -3150
rect 10230 -3310 10240 -3150
rect 10100 -3410 10240 -3310
rect 10100 -4090 10110 -3410
rect 10230 -4090 10240 -3410
rect 10100 -4100 10240 -4090
rect 9400 -4250 9540 -4240
rect 9400 -4370 9410 -4250
rect 9530 -4370 9540 -4250
rect 9400 -4380 9540 -4370
rect 9420 -4400 9520 -4380
rect 470 -4800 670 -4780
rect 1180 -4720 1320 -4710
rect 1180 -4840 1190 -4720
rect 1310 -4840 1320 -4720
rect 1180 -4850 1320 -4840
rect 2780 -4720 2920 -4710
rect 2780 -4840 2790 -4720
rect 2910 -4840 2920 -4720
rect 2780 -4850 2920 -4840
rect 4380 -4720 4520 -4710
rect 4380 -4840 4390 -4720
rect 4510 -4840 4520 -4720
rect 4380 -4850 4520 -4840
rect 5980 -4720 6120 -4710
rect 5980 -4840 5990 -4720
rect 6110 -4840 6120 -4720
rect 5980 -4850 6120 -4840
rect 7580 -4720 7720 -4710
rect 7580 -4840 7590 -4720
rect 7710 -4840 7720 -4720
rect 7580 -4850 7720 -4840
rect 9180 -4720 9320 -4710
rect 9180 -4840 9190 -4720
rect 9310 -4840 9320 -4720
rect 9180 -4850 9320 -4840
rect 11020 -4750 11120 -3050
rect 11700 -3150 11840 -2290
rect 12400 -2720 12500 -1060
rect 12620 -1070 12630 -930
rect 12750 -1070 12760 -930
rect 12620 -1100 12760 -1070
rect 12870 -1110 13250 -1100
rect 12870 -1260 12880 -1110
rect 13240 -1260 13250 -1110
rect 12870 -1270 13250 -1260
rect 13300 -1350 13440 -490
rect 14000 -920 14100 1320
rect 13960 -930 14100 -920
rect 13960 -1070 13970 -930
rect 14090 -1070 14100 -930
rect 13960 -1100 14100 -1070
rect 13300 -1510 13310 -1350
rect 13430 -1510 13440 -1350
rect 13300 -1610 13440 -1510
rect 13300 -2290 13310 -1610
rect 13430 -2290 13440 -1610
rect 12380 -2730 12520 -2720
rect 12380 -2850 12390 -2730
rect 12510 -2850 12520 -2730
rect 12380 -2860 12520 -2850
rect 11700 -3310 11710 -3150
rect 11830 -3310 11840 -3150
rect 11700 -3410 11840 -3310
rect 11700 -4090 11710 -3410
rect 11830 -4090 11840 -3410
rect 11700 -4100 11840 -4090
rect 12400 -4520 12500 -2860
rect 13300 -3150 13440 -2290
rect 14220 -2910 14320 2860
rect 16900 2780 17140 2790
rect 16900 2640 16910 2780
rect 17130 2640 17140 2780
rect 16900 2630 17140 2640
rect 17370 2780 17500 2790
rect 17370 2640 17380 2780
rect 17490 2640 17500 2780
rect 17370 2630 17500 2640
rect 17730 2780 17970 2790
rect 17730 2640 17740 2780
rect 17960 2640 17970 2780
rect 17730 2630 17970 2640
rect 16500 2250 16640 2260
rect 16500 2090 16510 2250
rect 16630 2090 16640 2250
rect 14900 1980 15040 2010
rect 14900 1320 14910 1980
rect 15030 1320 15040 1980
rect 14900 1240 15040 1320
rect 16500 1990 16640 2090
rect 16500 1310 16510 1990
rect 16630 1310 16640 1990
rect 18100 2250 18240 2260
rect 18100 2090 18110 2250
rect 18230 2090 18240 2250
rect 18100 1990 18240 2090
rect 18100 1310 18110 1990
rect 18230 1310 18240 1990
rect 19700 2250 19840 2260
rect 19700 2090 19710 2250
rect 19830 2090 19840 2250
rect 19700 1990 19840 2090
rect 19700 1310 19710 1990
rect 19830 1310 19840 1990
rect 21300 2250 21440 2260
rect 21300 2090 21310 2250
rect 21430 2090 21440 2250
rect 21300 1990 21440 2090
rect 21300 1310 21310 1990
rect 21430 1310 21440 1990
rect 22900 2250 23040 2260
rect 22900 2090 22910 2250
rect 23030 2090 23040 2250
rect 22900 1990 23040 2090
rect 22900 1310 22910 1990
rect 23030 1310 23040 1990
rect 24500 2250 24640 2260
rect 24500 2090 24510 2250
rect 24630 2090 24640 2250
rect 24500 1990 24640 2090
rect 24500 1310 24510 1990
rect 24630 1310 24640 1990
rect 26100 2250 26240 2260
rect 26100 2090 26110 2250
rect 26230 2090 26240 2250
rect 26100 1990 26240 2090
rect 26100 1310 26110 1990
rect 26230 1310 26240 1990
rect 27700 2250 27840 2260
rect 27700 2070 27710 2250
rect 27830 2070 27840 2250
rect 27700 1990 27840 2070
rect 27700 1310 27710 1990
rect 27830 1310 27840 1990
rect 29300 2250 29440 2260
rect 29300 2070 29310 2250
rect 29430 2070 29440 2250
rect 29300 1990 29440 2070
rect 29300 1310 29310 1990
rect 29430 1310 29440 1990
rect 15600 1160 15700 1310
rect 15590 1150 15710 1160
rect 15590 1030 15600 1150
rect 15700 1030 15710 1150
rect 15590 1020 15710 1030
rect 14900 190 15040 460
rect 14900 -560 14910 190
rect 14460 -570 14910 -560
rect 15030 -560 15040 190
rect 15030 -570 15480 -560
rect 14460 -730 14470 -570
rect 15470 -730 15480 -570
rect 15600 -640 15700 1020
rect 15820 690 15920 1310
rect 15810 680 15930 690
rect 15810 560 15820 680
rect 15920 560 15930 680
rect 15810 550 15930 560
rect 14460 -740 15480 -730
rect 15590 -650 15710 -640
rect 14900 -1350 15040 -1340
rect 14900 -1510 14910 -1350
rect 15030 -1510 15040 -1350
rect 14900 -1610 15040 -1510
rect 15240 -1350 15380 -740
rect 15590 -770 15600 -650
rect 15700 -770 15710 -650
rect 15590 -780 15710 -770
rect 15240 -1510 15250 -1350
rect 15370 -1510 15380 -1350
rect 15240 -1520 15380 -1510
rect 14900 -2290 14910 -1610
rect 15030 -2290 15040 -1610
rect 14200 -2920 14340 -2910
rect 14200 -3040 14210 -2920
rect 14330 -3040 14340 -2920
rect 14200 -3050 14340 -3040
rect 14420 -2920 14560 -2910
rect 14420 -3040 14430 -2920
rect 14550 -3040 14560 -2920
rect 14420 -3050 14560 -3040
rect 14440 -3110 14540 -3050
rect 12600 -3290 12740 -3280
rect 12600 -3390 12610 -3290
rect 12730 -3390 12740 -3290
rect 12600 -3400 12740 -3390
rect 13300 -3310 13310 -3150
rect 13430 -3310 13440 -3150
rect 12380 -4530 12520 -4520
rect 12380 -4650 12390 -4530
rect 12510 -4650 12520 -4530
rect 12380 -4660 12520 -4650
rect 12620 -4720 12720 -3400
rect 13300 -3410 13440 -3310
rect 13300 -4090 13310 -3410
rect 13430 -4090 13440 -3410
rect 13300 -4100 13440 -4090
rect 14000 -3220 14540 -3110
rect 14900 -3150 15040 -2290
rect 15600 -2440 15700 -780
rect 15820 -1110 15920 550
rect 16500 450 16640 1310
rect 17200 1160 17300 1310
rect 17190 1150 17310 1160
rect 17190 1030 17200 1150
rect 17300 1030 17310 1150
rect 17190 1020 17310 1030
rect 16500 290 16510 450
rect 16630 290 16640 450
rect 16500 190 16640 290
rect 16500 -490 16510 190
rect 16630 -490 16640 190
rect 15810 -1120 15930 -1110
rect 15810 -1240 15820 -1120
rect 15920 -1240 15930 -1120
rect 15810 -1250 15930 -1240
rect 15590 -2450 15710 -2440
rect 15590 -2570 15600 -2450
rect 15700 -2570 15710 -2450
rect 15590 -2580 15710 -2570
rect 12600 -4730 12740 -4720
rect 11020 -4850 11140 -4750
rect 1200 -4860 1300 -4850
rect 2800 -4880 2900 -4850
rect 4400 -4880 4500 -4850
rect 6000 -4880 6100 -4850
rect 7600 -4880 7700 -4850
rect 9200 -4880 9300 -4850
rect 7800 -7870 7940 -7860
rect 7800 -7990 7810 -7870
rect 7930 -7990 7940 -7870
rect 7800 -8000 7940 -7990
rect 1220 -8060 1320 -8050
rect 1200 -8070 1340 -8060
rect 480 -8090 680 -8080
rect 480 -22380 490 -8090
rect 670 -22380 680 -8090
rect 1200 -8190 1210 -8070
rect 1330 -8190 1340 -8070
rect 1200 -8200 1340 -8190
rect 1220 -9860 1320 -8200
rect 1440 -8500 1540 -8050
rect 2820 -8060 2920 -8050
rect 2800 -8070 2940 -8060
rect 2800 -8190 2810 -8070
rect 2930 -8190 2940 -8070
rect 2800 -8200 2940 -8190
rect 1420 -8510 1560 -8500
rect 1420 -8630 1430 -8510
rect 1550 -8630 1560 -8510
rect 1420 -8640 1560 -8630
rect 1200 -9870 1340 -9860
rect 1200 -9990 1210 -9870
rect 1330 -9990 1340 -9870
rect 1200 -10000 1340 -9990
rect 1220 -11660 1320 -10000
rect 1440 -10300 1540 -8640
rect 2120 -8810 2240 -8780
rect 2120 -9470 2130 -8810
rect 2230 -9470 2240 -8810
rect 2120 -9590 2240 -9470
rect 2120 -9750 2130 -9590
rect 2230 -9750 2240 -9590
rect 1420 -10310 1560 -10300
rect 1420 -10430 1430 -10310
rect 1550 -10430 1560 -10310
rect 1420 -10440 1560 -10430
rect 1200 -11670 1340 -11660
rect 1200 -11790 1210 -11670
rect 1330 -11790 1340 -11670
rect 1200 -11800 1340 -11790
rect 1220 -13460 1320 -11800
rect 1440 -12100 1540 -10440
rect 2120 -10610 2240 -9750
rect 2820 -9860 2920 -8200
rect 3040 -8500 3140 -8050
rect 4420 -8060 4520 -8050
rect 4400 -8070 4540 -8060
rect 4400 -8190 4410 -8070
rect 4530 -8190 4540 -8070
rect 4400 -8200 4540 -8190
rect 3020 -8510 3160 -8500
rect 3020 -8630 3030 -8510
rect 3150 -8630 3160 -8510
rect 3020 -8640 3160 -8630
rect 2800 -9870 2940 -9860
rect 2800 -9990 2810 -9870
rect 2930 -9990 2940 -9870
rect 2800 -10000 2940 -9990
rect 2120 -11270 2130 -10610
rect 2230 -11270 2240 -10610
rect 2120 -11390 2240 -11270
rect 2120 -11550 2130 -11390
rect 2230 -11550 2240 -11390
rect 1420 -12110 1560 -12100
rect 1420 -12230 1430 -12110
rect 1550 -12230 1560 -12110
rect 1420 -12240 1560 -12230
rect 1200 -13470 1340 -13460
rect 1200 -13590 1210 -13470
rect 1330 -13590 1340 -13470
rect 1200 -13600 1340 -13590
rect 1220 -15260 1320 -13600
rect 1440 -13900 1540 -12240
rect 2120 -12410 2240 -11550
rect 2820 -11660 2920 -10000
rect 3040 -10300 3140 -8640
rect 3720 -8810 3840 -8780
rect 3720 -9470 3730 -8810
rect 3830 -9470 3840 -8810
rect 3720 -9590 3840 -9470
rect 3720 -9750 3730 -9590
rect 3830 -9750 3840 -9590
rect 3020 -10310 3160 -10300
rect 3020 -10430 3030 -10310
rect 3150 -10430 3160 -10310
rect 3020 -10440 3160 -10430
rect 2800 -11670 2940 -11660
rect 2800 -11790 2810 -11670
rect 2930 -11790 2940 -11670
rect 2800 -11800 2940 -11790
rect 2120 -13070 2130 -12410
rect 2230 -13070 2240 -12410
rect 2120 -13190 2240 -13070
rect 2120 -13350 2130 -13190
rect 2230 -13350 2240 -13190
rect 1420 -13910 1560 -13900
rect 1420 -14030 1430 -13910
rect 1550 -14030 1560 -13910
rect 1420 -14040 1560 -14030
rect 1200 -15270 1340 -15260
rect 1200 -15390 1210 -15270
rect 1330 -15390 1340 -15270
rect 1200 -15400 1340 -15390
rect 1220 -17060 1320 -15400
rect 1440 -15700 1540 -14040
rect 2120 -14210 2240 -13350
rect 2820 -13460 2920 -11800
rect 3040 -12100 3140 -10440
rect 3720 -10610 3840 -9750
rect 4420 -9860 4520 -8200
rect 4640 -8500 4740 -8050
rect 6020 -8060 6120 -8050
rect 6000 -8070 6140 -8060
rect 6000 -8190 6010 -8070
rect 6130 -8190 6140 -8070
rect 6000 -8200 6140 -8190
rect 4620 -8510 4760 -8500
rect 4620 -8630 4630 -8510
rect 4750 -8630 4760 -8510
rect 4620 -8640 4760 -8630
rect 4400 -9870 4540 -9860
rect 4400 -9990 4410 -9870
rect 4530 -9990 4540 -9870
rect 4400 -10000 4540 -9990
rect 3720 -11270 3730 -10610
rect 3830 -11270 3840 -10610
rect 3720 -11390 3840 -11270
rect 3720 -11550 3730 -11390
rect 3830 -11550 3840 -11390
rect 3020 -12110 3160 -12100
rect 3020 -12230 3030 -12110
rect 3150 -12230 3160 -12110
rect 3020 -12240 3160 -12230
rect 2800 -13470 2940 -13460
rect 2800 -13590 2810 -13470
rect 2930 -13590 2940 -13470
rect 2800 -13600 2940 -13590
rect 2120 -14870 2130 -14210
rect 2230 -14870 2240 -14210
rect 2120 -14990 2240 -14870
rect 2120 -15150 2130 -14990
rect 2230 -15150 2240 -14990
rect 1420 -15710 1560 -15700
rect 1420 -15830 1430 -15710
rect 1550 -15830 1560 -15710
rect 1420 -15840 1560 -15830
rect 1200 -17070 1340 -17060
rect 1200 -17190 1210 -17070
rect 1330 -17190 1340 -17070
rect 1200 -17200 1340 -17190
rect 1220 -18860 1320 -17200
rect 1440 -17500 1540 -15840
rect 2120 -16010 2240 -15150
rect 2820 -15260 2920 -13600
rect 3040 -13900 3140 -12240
rect 3720 -12410 3840 -11550
rect 4420 -11660 4520 -10000
rect 4640 -10300 4740 -8640
rect 5320 -8810 5440 -8780
rect 5320 -9470 5330 -8810
rect 5430 -9470 5440 -8810
rect 5320 -9590 5440 -9470
rect 5320 -9750 5330 -9590
rect 5430 -9750 5440 -9590
rect 4620 -10310 4760 -10300
rect 4620 -10430 4630 -10310
rect 4750 -10430 4760 -10310
rect 4620 -10440 4760 -10430
rect 4400 -11670 4540 -11660
rect 4400 -11790 4410 -11670
rect 4530 -11790 4540 -11670
rect 4400 -11800 4540 -11790
rect 3720 -13070 3730 -12410
rect 3830 -13070 3840 -12410
rect 3720 -13190 3840 -13070
rect 3720 -13350 3730 -13190
rect 3830 -13350 3840 -13190
rect 3020 -13910 3160 -13900
rect 3020 -14030 3030 -13910
rect 3150 -14030 3160 -13910
rect 3020 -14040 3160 -14030
rect 2800 -15270 2940 -15260
rect 2800 -15390 2810 -15270
rect 2930 -15390 2940 -15270
rect 2800 -15400 2940 -15390
rect 2120 -16670 2130 -16010
rect 2230 -16670 2240 -16010
rect 2120 -16790 2240 -16670
rect 2120 -16950 2130 -16790
rect 2230 -16950 2240 -16790
rect 1420 -17510 1560 -17500
rect 1420 -17630 1430 -17510
rect 1550 -17630 1560 -17510
rect 1420 -17640 1560 -17630
rect 1200 -18870 1340 -18860
rect 1200 -18990 1210 -18870
rect 1330 -18990 1340 -18870
rect 1200 -19000 1340 -18990
rect 1220 -20660 1320 -19000
rect 1440 -19300 1540 -17640
rect 2120 -17810 2240 -16950
rect 2820 -17060 2920 -15400
rect 3040 -15700 3140 -14040
rect 3720 -14210 3840 -13350
rect 4420 -13460 4520 -11800
rect 4640 -12100 4740 -10440
rect 5320 -10610 5440 -9750
rect 6020 -9860 6120 -8200
rect 6240 -8500 6340 -8050
rect 7620 -8060 7720 -8050
rect 9220 -8060 9320 -8050
rect 7600 -8070 7740 -8060
rect 7600 -8190 7610 -8070
rect 7730 -8190 7740 -8070
rect 7600 -8200 7740 -8190
rect 9200 -8070 9340 -8060
rect 9200 -8190 9210 -8070
rect 9330 -8190 9340 -8070
rect 9200 -8200 9340 -8190
rect 6220 -8510 6360 -8500
rect 6220 -8630 6230 -8510
rect 6350 -8630 6360 -8510
rect 6220 -8640 6360 -8630
rect 6000 -9870 6140 -9860
rect 6000 -9990 6010 -9870
rect 6130 -9990 6140 -9870
rect 6000 -10000 6140 -9990
rect 5320 -11270 5330 -10610
rect 5430 -11270 5440 -10610
rect 5320 -11390 5440 -11270
rect 5320 -11550 5330 -11390
rect 5430 -11550 5440 -11390
rect 4620 -12110 4760 -12100
rect 4620 -12230 4630 -12110
rect 4750 -12230 4760 -12110
rect 4620 -12240 4760 -12230
rect 4400 -13470 4540 -13460
rect 4400 -13590 4410 -13470
rect 4530 -13590 4540 -13470
rect 4400 -13600 4540 -13590
rect 3720 -14870 3730 -14210
rect 3830 -14870 3840 -14210
rect 3720 -14990 3840 -14870
rect 3720 -15150 3730 -14990
rect 3830 -15150 3840 -14990
rect 3020 -15710 3160 -15700
rect 3020 -15830 3030 -15710
rect 3150 -15830 3160 -15710
rect 3020 -15840 3160 -15830
rect 2800 -17070 2940 -17060
rect 2800 -17190 2810 -17070
rect 2930 -17190 2940 -17070
rect 2800 -17200 2940 -17190
rect 2120 -18470 2130 -17810
rect 2230 -18470 2240 -17810
rect 2120 -18590 2240 -18470
rect 2120 -18750 2130 -18590
rect 2230 -18750 2240 -18590
rect 1420 -19310 1560 -19300
rect 1420 -19430 1430 -19310
rect 1550 -19430 1560 -19310
rect 1420 -19440 1560 -19430
rect 1200 -20670 1340 -20660
rect 1200 -20790 1210 -20670
rect 1330 -20790 1340 -20670
rect 1200 -20800 1340 -20790
rect 480 -22400 680 -22380
rect 1220 -23260 1320 -20800
rect 1440 -21100 1540 -19440
rect 2120 -19610 2240 -18750
rect 2820 -18860 2920 -17200
rect 3040 -17500 3140 -15840
rect 3720 -16010 3840 -15150
rect 4420 -15260 4520 -13600
rect 4640 -13900 4740 -12240
rect 5320 -12410 5440 -11550
rect 6020 -11660 6120 -10000
rect 6240 -10300 6340 -8640
rect 6920 -8810 7040 -8780
rect 6920 -9470 6930 -8810
rect 7030 -9470 7040 -8810
rect 6920 -9590 7040 -9470
rect 6920 -9750 6930 -9590
rect 7030 -9750 7040 -9590
rect 6220 -10310 6360 -10300
rect 6220 -10430 6230 -10310
rect 6350 -10430 6360 -10310
rect 6220 -10440 6360 -10430
rect 6000 -11670 6140 -11660
rect 6000 -11790 6010 -11670
rect 6130 -11790 6140 -11670
rect 6000 -11800 6140 -11790
rect 5320 -13070 5330 -12410
rect 5430 -13070 5440 -12410
rect 5320 -13190 5440 -13070
rect 5320 -13350 5330 -13190
rect 5430 -13350 5440 -13190
rect 4620 -13910 4760 -13900
rect 4620 -14030 4630 -13910
rect 4750 -14030 4760 -13910
rect 4620 -14040 4760 -14030
rect 4400 -15270 4540 -15260
rect 4400 -15390 4410 -15270
rect 4530 -15390 4540 -15270
rect 4400 -15400 4540 -15390
rect 3720 -16670 3730 -16010
rect 3830 -16670 3840 -16010
rect 3720 -16790 3840 -16670
rect 3720 -16950 3730 -16790
rect 3830 -16950 3840 -16790
rect 3020 -17510 3160 -17500
rect 3020 -17630 3030 -17510
rect 3150 -17630 3160 -17510
rect 3020 -17640 3160 -17630
rect 2800 -18870 2940 -18860
rect 2800 -18990 2810 -18870
rect 2930 -18990 2940 -18870
rect 2800 -19000 2940 -18990
rect 2120 -20270 2130 -19610
rect 2230 -20270 2240 -19610
rect 2120 -20390 2240 -20270
rect 2120 -20550 2130 -20390
rect 2230 -20550 2240 -20390
rect 1420 -21110 1560 -21100
rect 1420 -21230 1430 -21110
rect 1550 -21230 1560 -21110
rect 1420 -21240 1560 -21230
rect 2120 -21410 2240 -20550
rect 2820 -20660 2920 -19000
rect 3040 -19300 3140 -17640
rect 3720 -17810 3840 -16950
rect 4420 -17060 4520 -15400
rect 4640 -15700 4740 -14040
rect 5320 -14210 5440 -13350
rect 6020 -13460 6120 -11800
rect 6240 -12100 6340 -10440
rect 6920 -10610 7040 -9750
rect 7620 -9860 7720 -8200
rect 7840 -8500 7940 -8220
rect 7820 -8510 7960 -8500
rect 7820 -8630 7830 -8510
rect 7950 -8630 7960 -8510
rect 7820 -8640 7960 -8630
rect 7600 -9870 7740 -9860
rect 7600 -9990 7610 -9870
rect 7730 -9990 7740 -9870
rect 7600 -10000 7740 -9990
rect 6920 -11270 6930 -10610
rect 7030 -11270 7040 -10610
rect 6920 -11390 7040 -11270
rect 6920 -11550 6930 -11390
rect 7030 -11550 7040 -11390
rect 6220 -12110 6360 -12100
rect 6220 -12230 6230 -12110
rect 6350 -12230 6360 -12110
rect 6220 -12240 6360 -12230
rect 6000 -13470 6140 -13460
rect 6000 -13590 6010 -13470
rect 6130 -13590 6140 -13470
rect 6000 -13600 6140 -13590
rect 5320 -14870 5330 -14210
rect 5430 -14870 5440 -14210
rect 5320 -14990 5440 -14870
rect 5320 -15150 5330 -14990
rect 5430 -15150 5440 -14990
rect 4620 -15710 4760 -15700
rect 4620 -15830 4630 -15710
rect 4750 -15830 4760 -15710
rect 4620 -15840 4760 -15830
rect 4400 -17070 4540 -17060
rect 4400 -17190 4410 -17070
rect 4530 -17190 4540 -17070
rect 4400 -17200 4540 -17190
rect 3720 -18470 3730 -17810
rect 3830 -18470 3840 -17810
rect 3720 -18590 3840 -18470
rect 3720 -18750 3730 -18590
rect 3830 -18750 3840 -18590
rect 3020 -19310 3160 -19300
rect 3020 -19430 3030 -19310
rect 3150 -19430 3160 -19310
rect 3020 -19440 3160 -19430
rect 2800 -20670 2940 -20660
rect 2800 -20790 2810 -20670
rect 2930 -20790 2940 -20670
rect 2800 -20800 2940 -20790
rect 2120 -22070 2130 -21410
rect 2230 -22070 2240 -21410
rect 2120 -22190 2240 -22070
rect 2120 -22350 2130 -22190
rect 2230 -22350 2240 -22190
rect 2120 -22360 2240 -22350
rect 2820 -23260 2920 -20800
rect 3040 -21100 3140 -19440
rect 3720 -19610 3840 -18750
rect 4420 -18860 4520 -17200
rect 4640 -17500 4740 -15840
rect 5320 -16010 5440 -15150
rect 6020 -15260 6120 -13600
rect 6240 -13900 6340 -12240
rect 6920 -12410 7040 -11550
rect 7620 -11660 7720 -10000
rect 7840 -10300 7940 -8640
rect 8520 -8810 8640 -8780
rect 8520 -9470 8530 -8810
rect 8630 -9470 8640 -8810
rect 8520 -9590 8640 -9470
rect 8520 -9750 8530 -9590
rect 8630 -9750 8640 -9590
rect 7820 -10310 7960 -10300
rect 7820 -10430 7830 -10310
rect 7950 -10430 7960 -10310
rect 7820 -10440 7960 -10430
rect 7600 -11670 7740 -11660
rect 7600 -11790 7610 -11670
rect 7730 -11790 7740 -11670
rect 7600 -11800 7740 -11790
rect 6920 -13070 6930 -12410
rect 7030 -13070 7040 -12410
rect 6920 -13190 7040 -13070
rect 6920 -13350 6930 -13190
rect 7030 -13350 7040 -13190
rect 6220 -13910 6360 -13900
rect 6220 -14030 6230 -13910
rect 6350 -14030 6360 -13910
rect 6220 -14040 6360 -14030
rect 6000 -15270 6140 -15260
rect 6000 -15390 6010 -15270
rect 6130 -15390 6140 -15270
rect 6000 -15400 6140 -15390
rect 5320 -16670 5330 -16010
rect 5430 -16670 5440 -16010
rect 5320 -16790 5440 -16670
rect 5320 -16950 5330 -16790
rect 5430 -16950 5440 -16790
rect 4620 -17510 4760 -17500
rect 4620 -17630 4630 -17510
rect 4750 -17630 4760 -17510
rect 4620 -17640 4760 -17630
rect 4400 -18870 4540 -18860
rect 4400 -18990 4410 -18870
rect 4530 -18990 4540 -18870
rect 4400 -19000 4540 -18990
rect 3720 -20270 3730 -19610
rect 3830 -20270 3840 -19610
rect 3720 -20390 3840 -20270
rect 3720 -20550 3730 -20390
rect 3830 -20550 3840 -20390
rect 3020 -21110 3160 -21100
rect 3020 -21230 3030 -21110
rect 3150 -21230 3160 -21110
rect 3020 -21240 3160 -21230
rect 3720 -21410 3840 -20550
rect 4420 -20660 4520 -19000
rect 4640 -19300 4740 -17640
rect 5320 -17810 5440 -16950
rect 6020 -17060 6120 -15400
rect 6240 -15700 6340 -14040
rect 6920 -14210 7040 -13350
rect 7620 -13460 7720 -11800
rect 7840 -12100 7940 -10440
rect 8520 -10610 8640 -9750
rect 9220 -9860 9320 -8200
rect 9440 -8500 9540 -8050
rect 10820 -8250 10920 -8030
rect 10800 -8260 10940 -8250
rect 10800 -8380 10810 -8260
rect 10930 -8380 10940 -8260
rect 10800 -8390 10940 -8380
rect 9420 -8510 9560 -8500
rect 9420 -8630 9430 -8510
rect 9550 -8630 9560 -8510
rect 9420 -8640 9560 -8630
rect 9200 -9870 9340 -9860
rect 9200 -9990 9210 -9870
rect 9330 -9990 9340 -9870
rect 9200 -10000 9340 -9990
rect 8520 -11270 8530 -10610
rect 8630 -11270 8640 -10610
rect 8520 -11390 8640 -11270
rect 8520 -11550 8530 -11390
rect 8630 -11550 8640 -11390
rect 7820 -12110 7960 -12100
rect 7820 -12230 7830 -12110
rect 7950 -12230 7960 -12110
rect 7820 -12240 7960 -12230
rect 7600 -13470 7740 -13460
rect 7600 -13590 7610 -13470
rect 7730 -13590 7740 -13470
rect 7600 -13600 7740 -13590
rect 6920 -14870 6930 -14210
rect 7030 -14870 7040 -14210
rect 6920 -14990 7040 -14870
rect 6920 -15150 6930 -14990
rect 7030 -15150 7040 -14990
rect 6220 -15710 6360 -15700
rect 6220 -15830 6230 -15710
rect 6350 -15830 6360 -15710
rect 6220 -15840 6360 -15830
rect 6000 -17070 6140 -17060
rect 6000 -17190 6010 -17070
rect 6130 -17190 6140 -17070
rect 6000 -17200 6140 -17190
rect 5320 -18470 5330 -17810
rect 5430 -18470 5440 -17810
rect 5320 -18590 5440 -18470
rect 5320 -18750 5330 -18590
rect 5430 -18750 5440 -18590
rect 4620 -19310 4760 -19300
rect 4620 -19430 4630 -19310
rect 4750 -19430 4760 -19310
rect 4620 -19440 4760 -19430
rect 4400 -20670 4540 -20660
rect 4400 -20790 4410 -20670
rect 4530 -20790 4540 -20670
rect 4400 -20800 4540 -20790
rect 3720 -22070 3730 -21410
rect 3830 -22070 3840 -21410
rect 3720 -22190 3840 -22070
rect 3720 -22350 3730 -22190
rect 3830 -22350 3840 -22190
rect 3720 -22360 3840 -22350
rect 4420 -23260 4520 -20800
rect 4640 -21100 4740 -19440
rect 5320 -19610 5440 -18750
rect 6020 -18860 6120 -17200
rect 6240 -17500 6340 -15840
rect 6920 -16010 7040 -15150
rect 7620 -15260 7720 -13600
rect 7840 -13900 7940 -12240
rect 8520 -12410 8640 -11550
rect 9220 -11660 9320 -10000
rect 9440 -10300 9540 -8640
rect 10120 -8810 10240 -8780
rect 10120 -9470 10130 -8810
rect 10230 -9470 10240 -8810
rect 10120 -9590 10240 -9470
rect 10120 -9750 10130 -9590
rect 10230 -9750 10240 -9590
rect 9420 -10310 9560 -10300
rect 9420 -10430 9430 -10310
rect 9550 -10430 9560 -10310
rect 9420 -10440 9560 -10430
rect 9200 -11670 9340 -11660
rect 9200 -11790 9210 -11670
rect 9330 -11790 9340 -11670
rect 9200 -11800 9340 -11790
rect 8520 -13070 8530 -12410
rect 8630 -13070 8640 -12410
rect 8520 -13190 8640 -13070
rect 8520 -13350 8530 -13190
rect 8630 -13350 8640 -13190
rect 7820 -13910 7960 -13900
rect 7820 -14030 7830 -13910
rect 7950 -14030 7960 -13910
rect 7820 -14040 7960 -14030
rect 7600 -15270 7740 -15260
rect 7600 -15390 7610 -15270
rect 7730 -15390 7740 -15270
rect 7600 -15400 7740 -15390
rect 6920 -16670 6930 -16010
rect 7030 -16670 7040 -16010
rect 6920 -16790 7040 -16670
rect 6920 -16950 6930 -16790
rect 7030 -16950 7040 -16790
rect 6220 -17510 6360 -17500
rect 6220 -17630 6230 -17510
rect 6350 -17630 6360 -17510
rect 6220 -17640 6360 -17630
rect 6000 -18870 6140 -18860
rect 6000 -18990 6010 -18870
rect 6130 -18990 6140 -18870
rect 6000 -19000 6140 -18990
rect 5320 -20270 5330 -19610
rect 5430 -20270 5440 -19610
rect 5320 -20390 5440 -20270
rect 5320 -20550 5330 -20390
rect 5430 -20550 5440 -20390
rect 4620 -21110 4760 -21100
rect 4620 -21230 4630 -21110
rect 4750 -21230 4760 -21110
rect 4620 -21240 4760 -21230
rect 5320 -21410 5440 -20550
rect 6020 -20660 6120 -19000
rect 6240 -19300 6340 -17640
rect 6920 -17810 7040 -16950
rect 7620 -17060 7720 -15400
rect 7840 -15700 7940 -14040
rect 8520 -14210 8640 -13350
rect 9220 -13460 9320 -11800
rect 9440 -12100 9540 -10440
rect 10120 -10610 10240 -9750
rect 10820 -10050 10920 -8390
rect 11040 -9580 11140 -4850
rect 11700 -4810 11840 -4800
rect 11700 -4930 11710 -4810
rect 11830 -4930 11840 -4810
rect 12600 -4850 12610 -4730
rect 12730 -4850 12740 -4730
rect 12600 -4860 12740 -4850
rect 13620 -4790 13760 -4780
rect 13620 -4910 13630 -4790
rect 13750 -4910 13760 -4790
rect 13620 -4920 13760 -4910
rect 11700 -4940 11840 -4930
rect 11720 -5820 11820 -4940
rect 11700 -5830 11840 -5820
rect 11700 -5950 11710 -5830
rect 11830 -5950 11840 -5830
rect 11700 -5960 11840 -5950
rect 13300 -5830 13440 -5820
rect 13300 -5950 13310 -5830
rect 13430 -5950 13440 -5830
rect 13300 -5960 13440 -5950
rect 11700 -6050 11840 -6040
rect 11700 -6170 11710 -6050
rect 11830 -6170 11840 -6050
rect 11700 -6180 11840 -6170
rect 11720 -8100 11820 -6180
rect 12620 -6270 12760 -6260
rect 12620 -6390 12630 -6270
rect 12750 -6390 12760 -6270
rect 12620 -6400 12760 -6390
rect 12400 -6490 12540 -6480
rect 12400 -6610 12410 -6490
rect 12530 -6610 12540 -6490
rect 12400 -6620 12540 -6610
rect 11700 -8110 11860 -8100
rect 11700 -8230 11710 -8110
rect 11840 -8140 11860 -8110
rect 11840 -8230 11850 -8140
rect 11700 -8240 11850 -8230
rect 11710 -8810 11840 -8240
rect 11710 -9470 11720 -8810
rect 11830 -9470 11840 -8810
rect 11710 -9480 11840 -9470
rect 11030 -9760 11150 -9580
rect 10800 -10060 10940 -10050
rect 10800 -10180 10810 -10060
rect 10930 -10180 10940 -10060
rect 10800 -10190 10940 -10180
rect 10120 -11270 10130 -10610
rect 10230 -11270 10240 -10610
rect 10120 -11390 10240 -11270
rect 10120 -11550 10130 -11390
rect 10230 -11550 10240 -11390
rect 9420 -12110 9560 -12100
rect 9420 -12230 9430 -12110
rect 9550 -12230 9560 -12110
rect 9420 -12240 9560 -12230
rect 9200 -13470 9340 -13460
rect 9200 -13590 9210 -13470
rect 9330 -13590 9340 -13470
rect 9200 -13600 9340 -13590
rect 8520 -14870 8530 -14210
rect 8630 -14870 8640 -14210
rect 8520 -14990 8640 -14870
rect 8520 -15150 8530 -14990
rect 8630 -15150 8640 -14990
rect 7820 -15710 7960 -15700
rect 7820 -15830 7830 -15710
rect 7950 -15830 7960 -15710
rect 7820 -15840 7960 -15830
rect 7600 -17070 7740 -17060
rect 7600 -17190 7610 -17070
rect 7730 -17190 7740 -17070
rect 7600 -17200 7740 -17190
rect 6920 -18470 6930 -17810
rect 7030 -18470 7040 -17810
rect 6920 -18590 7040 -18470
rect 6920 -18750 6930 -18590
rect 7030 -18750 7040 -18590
rect 6220 -19310 6360 -19300
rect 6220 -19430 6230 -19310
rect 6350 -19430 6360 -19310
rect 6220 -19440 6360 -19430
rect 6000 -20670 6140 -20660
rect 6000 -20790 6010 -20670
rect 6130 -20790 6140 -20670
rect 6000 -20800 6140 -20790
rect 5320 -22070 5330 -21410
rect 5430 -22070 5440 -21410
rect 5320 -22190 5440 -22070
rect 5320 -22350 5330 -22190
rect 5430 -22350 5440 -22190
rect 5320 -22360 5440 -22350
rect 6020 -23260 6120 -20800
rect 6240 -21100 6340 -19440
rect 6920 -19610 7040 -18750
rect 7620 -18860 7720 -17200
rect 7840 -17500 7940 -15840
rect 8520 -16010 8640 -15150
rect 9220 -15260 9320 -13600
rect 9440 -13900 9540 -12240
rect 10120 -12410 10240 -11550
rect 10820 -11850 10920 -10190
rect 11040 -10400 11140 -9760
rect 11020 -10410 11160 -10400
rect 11020 -10530 11030 -10410
rect 11150 -10530 11160 -10410
rect 11020 -10540 11160 -10530
rect 11040 -11380 11140 -10540
rect 11710 -10610 11840 -10600
rect 11710 -11270 11720 -10610
rect 11830 -11270 11840 -10610
rect 11030 -11560 11150 -11380
rect 10800 -11860 10940 -11850
rect 10800 -11980 10810 -11860
rect 10930 -11980 10940 -11860
rect 10800 -11990 10940 -11980
rect 10120 -13070 10130 -12410
rect 10230 -13070 10240 -12410
rect 10120 -13190 10240 -13070
rect 10120 -13350 10130 -13190
rect 10230 -13350 10240 -13190
rect 9420 -13910 9560 -13900
rect 9420 -14030 9430 -13910
rect 9550 -14030 9560 -13910
rect 9420 -14040 9560 -14030
rect 9200 -15270 9340 -15260
rect 9200 -15390 9210 -15270
rect 9330 -15390 9340 -15270
rect 9200 -15400 9340 -15390
rect 8520 -16670 8530 -16010
rect 8630 -16670 8640 -16010
rect 8520 -16790 8640 -16670
rect 8520 -16950 8530 -16790
rect 8630 -16950 8640 -16790
rect 7820 -17510 7960 -17500
rect 7820 -17630 7830 -17510
rect 7950 -17630 7960 -17510
rect 7820 -17640 7960 -17630
rect 7600 -18870 7740 -18860
rect 7600 -18990 7610 -18870
rect 7730 -18990 7740 -18870
rect 7600 -19000 7740 -18990
rect 6920 -20270 6930 -19610
rect 7030 -20270 7040 -19610
rect 6920 -20390 7040 -20270
rect 6920 -20550 6930 -20390
rect 7030 -20550 7040 -20390
rect 6220 -21110 6360 -21100
rect 6220 -21230 6230 -21110
rect 6350 -21230 6360 -21110
rect 6220 -21240 6360 -21230
rect 6920 -21410 7040 -20550
rect 7620 -20660 7720 -19000
rect 7840 -19300 7940 -17640
rect 8520 -17810 8640 -16950
rect 9220 -17060 9320 -15400
rect 9440 -15700 9540 -14040
rect 10120 -14210 10240 -13350
rect 10820 -13650 10920 -11990
rect 11040 -13180 11140 -11560
rect 11710 -12410 11840 -11270
rect 11710 -13070 11720 -12410
rect 11830 -13070 11840 -12410
rect 11030 -13360 11150 -13180
rect 11260 -13210 11270 -13150
rect 11650 -13210 11660 -13150
rect 10800 -13660 10940 -13650
rect 10800 -13780 10810 -13660
rect 10930 -13780 10940 -13660
rect 10800 -13790 10940 -13780
rect 10120 -14870 10130 -14210
rect 10230 -14870 10240 -14210
rect 10120 -14990 10240 -14870
rect 10120 -15150 10130 -14990
rect 10230 -15150 10240 -14990
rect 9420 -15710 9560 -15700
rect 9420 -15830 9430 -15710
rect 9550 -15830 9560 -15710
rect 9420 -15840 9560 -15830
rect 9200 -17070 9340 -17060
rect 9200 -17190 9210 -17070
rect 9330 -17190 9340 -17070
rect 9200 -17200 9340 -17190
rect 8520 -18470 8530 -17810
rect 8630 -18470 8640 -17810
rect 8520 -18590 8640 -18470
rect 8520 -18750 8530 -18590
rect 8630 -18750 8640 -18590
rect 7820 -19310 7960 -19300
rect 7820 -19430 7830 -19310
rect 7950 -19430 7960 -19310
rect 7820 -19440 7960 -19430
rect 7600 -20670 7740 -20660
rect 7600 -20790 7610 -20670
rect 7730 -20790 7740 -20670
rect 7600 -20800 7740 -20790
rect 6920 -22070 6930 -21410
rect 7030 -22070 7040 -21410
rect 6920 -22190 7040 -22070
rect 6920 -22350 6930 -22190
rect 7030 -22350 7040 -22190
rect 6920 -22360 7040 -22350
rect 7620 -23260 7720 -20800
rect 7840 -21100 7940 -19440
rect 8520 -19610 8640 -18750
rect 9220 -18860 9320 -17200
rect 9440 -17500 9540 -15840
rect 10120 -16010 10240 -15150
rect 10820 -15450 10920 -13790
rect 11040 -14980 11140 -13360
rect 11260 -14060 11660 -13210
rect 11260 -14120 11270 -14060
rect 11650 -14120 11660 -14060
rect 11260 -14130 11660 -14120
rect 11710 -14210 11840 -13070
rect 11710 -14870 11720 -14210
rect 11830 -14870 11840 -14210
rect 11710 -14880 11840 -14870
rect 11030 -15160 11150 -14980
rect 10800 -15460 10940 -15450
rect 10800 -15580 10810 -15460
rect 10930 -15580 10940 -15460
rect 10800 -15590 10940 -15580
rect 10120 -16670 10130 -16010
rect 10230 -16670 10240 -16010
rect 10120 -16790 10240 -16670
rect 10120 -16950 10130 -16790
rect 10230 -16950 10240 -16790
rect 9420 -17510 9560 -17500
rect 9420 -17630 9430 -17510
rect 9550 -17630 9560 -17510
rect 9420 -17640 9560 -17630
rect 9200 -18870 9340 -18860
rect 9200 -18990 9210 -18870
rect 9330 -18990 9340 -18870
rect 9200 -19000 9340 -18990
rect 8520 -20270 8530 -19610
rect 8630 -20270 8640 -19610
rect 8520 -20390 8640 -20270
rect 8520 -20550 8530 -20390
rect 8630 -20550 8640 -20390
rect 7820 -21110 7960 -21100
rect 7820 -21230 7830 -21110
rect 7950 -21230 7960 -21110
rect 7820 -21240 7960 -21230
rect 8520 -21410 8640 -20550
rect 9220 -20660 9320 -19000
rect 9440 -19300 9540 -17640
rect 10120 -17810 10240 -16950
rect 10820 -17250 10920 -15590
rect 11040 -16780 11140 -15160
rect 11030 -16960 11150 -16780
rect 10800 -17260 10940 -17250
rect 10800 -17380 10810 -17260
rect 10930 -17380 10940 -17260
rect 10800 -17390 10940 -17380
rect 10120 -18470 10130 -17810
rect 10230 -18470 10240 -17810
rect 10120 -18590 10240 -18470
rect 10120 -18750 10130 -18590
rect 10230 -18750 10240 -18590
rect 9420 -19310 9560 -19300
rect 9420 -19430 9430 -19310
rect 9550 -19430 9560 -19310
rect 9420 -19440 9560 -19430
rect 9200 -20670 9340 -20660
rect 9200 -20790 9210 -20670
rect 9330 -20790 9340 -20670
rect 9200 -20800 9340 -20790
rect 8520 -22070 8530 -21410
rect 8630 -22070 8640 -21410
rect 8520 -22190 8640 -22070
rect 8520 -22350 8530 -22190
rect 8630 -22350 8640 -22190
rect 8520 -22360 8640 -22350
rect 9220 -23260 9320 -20800
rect 9440 -21100 9540 -19440
rect 10120 -19610 10240 -18750
rect 10820 -19050 10920 -17390
rect 11040 -18580 11140 -16960
rect 11030 -18760 11150 -18580
rect 10800 -19060 10940 -19050
rect 10800 -19180 10810 -19060
rect 10930 -19180 10940 -19060
rect 10800 -19190 10940 -19180
rect 10120 -20270 10130 -19610
rect 10230 -20270 10240 -19610
rect 10120 -20390 10240 -20270
rect 10120 -20550 10130 -20390
rect 10230 -20550 10240 -20390
rect 9420 -21110 9560 -21100
rect 9420 -21230 9430 -21110
rect 9550 -21230 9560 -21110
rect 9420 -21240 9560 -21230
rect 10120 -21410 10240 -20550
rect 10820 -20850 10920 -19190
rect 11040 -20380 11140 -18760
rect 12420 -18870 12520 -6620
rect 12640 -17070 12740 -6400
rect 12940 -6830 13120 -6820
rect 12940 -6990 12950 -6830
rect 13110 -6990 13120 -6830
rect 12940 -7000 13120 -6990
rect 13310 -8240 13440 -5960
rect 13640 -6040 13740 -4920
rect 14000 -5070 14100 -3220
rect 14200 -3290 14340 -3280
rect 14200 -3410 14210 -3290
rect 14330 -3410 14340 -3290
rect 14200 -3420 14340 -3410
rect 14900 -3310 14910 -3150
rect 15030 -3310 15040 -3150
rect 14900 -3410 15040 -3310
rect 14220 -4720 14320 -3420
rect 14900 -4090 14910 -3410
rect 15030 -4090 15040 -3410
rect 14900 -4100 15040 -4090
rect 15600 -4240 15700 -2580
rect 15820 -2910 15920 -1250
rect 16500 -1350 16640 -490
rect 17200 -640 17300 1020
rect 17420 690 17520 1310
rect 17410 680 17530 690
rect 17410 560 17420 680
rect 17520 560 17530 680
rect 17410 550 17530 560
rect 17190 -650 17310 -640
rect 17190 -770 17200 -650
rect 17300 -770 17310 -650
rect 17190 -780 17310 -770
rect 16500 -1510 16510 -1350
rect 16630 -1510 16640 -1350
rect 16500 -1610 16640 -1510
rect 16500 -2290 16510 -1610
rect 16630 -2290 16640 -1610
rect 15810 -2920 15930 -2910
rect 15810 -3040 15820 -2920
rect 15920 -3040 15930 -2920
rect 15810 -3050 15930 -3040
rect 15590 -4250 15710 -4240
rect 15590 -4370 15600 -4250
rect 15700 -4370 15710 -4250
rect 15590 -4380 15710 -4370
rect 14200 -4730 14340 -4720
rect 14200 -4850 14210 -4730
rect 14330 -4850 14340 -4730
rect 14200 -4860 14340 -4850
rect 15220 -4790 15360 -4780
rect 15220 -4910 15230 -4790
rect 15350 -4910 15360 -4790
rect 15220 -4920 15360 -4910
rect 14000 -5200 14120 -5070
rect 13620 -6050 13760 -6040
rect 13620 -6170 13630 -6050
rect 13750 -6170 13760 -6050
rect 13620 -6180 13760 -6170
rect 13300 -8260 13450 -8240
rect 13300 -8380 13310 -8260
rect 13440 -8380 13450 -8260
rect 13300 -8390 13450 -8380
rect 13310 -8810 13440 -8390
rect 13310 -9470 13320 -8810
rect 13430 -9470 13440 -8810
rect 13310 -9480 13440 -9470
rect 13310 -10610 13440 -10600
rect 13310 -11270 13320 -10610
rect 13430 -11270 13440 -10610
rect 13310 -11280 13440 -11270
rect 13300 -11670 13440 -11660
rect 13300 -11790 13310 -11670
rect 13430 -11790 13440 -11670
rect 13300 -11800 13440 -11790
rect 13310 -12410 13440 -11800
rect 13310 -13070 13320 -12410
rect 13430 -13070 13440 -12410
rect 13310 -13160 13440 -13070
rect 13280 -13170 13470 -13160
rect 13280 -13330 13290 -13170
rect 13460 -13330 13470 -13170
rect 13280 -13340 13470 -13330
rect 13310 -14210 13440 -13340
rect 14020 -13470 14120 -5200
rect 15240 -6040 15340 -4920
rect 15600 -5160 15700 -4380
rect 15820 -4710 15920 -3050
rect 16500 -3150 16640 -2290
rect 17200 -2440 17300 -780
rect 17420 -1110 17520 550
rect 18100 450 18240 1310
rect 18800 1160 18900 1310
rect 18790 1150 18910 1160
rect 18790 1030 18800 1150
rect 18900 1030 18910 1150
rect 18790 1020 18910 1030
rect 18100 290 18110 450
rect 18230 290 18240 450
rect 18100 190 18240 290
rect 18100 -490 18110 190
rect 18230 -490 18240 190
rect 17410 -1120 17530 -1110
rect 17410 -1240 17420 -1120
rect 17520 -1240 17530 -1120
rect 17410 -1250 17530 -1240
rect 17190 -2450 17310 -2440
rect 17190 -2570 17200 -2450
rect 17300 -2570 17310 -2450
rect 17190 -2580 17310 -2570
rect 16500 -3310 16510 -3150
rect 16630 -3310 16640 -3150
rect 16500 -3410 16640 -3310
rect 16500 -4090 16510 -3410
rect 16630 -4090 16640 -3410
rect 15810 -4720 15930 -4710
rect 15810 -4840 15820 -4720
rect 15920 -4840 15930 -4720
rect 15810 -4850 15930 -4840
rect 15560 -5170 15740 -5160
rect 15560 -5350 15570 -5170
rect 15730 -5350 15740 -5170
rect 15560 -5360 15740 -5350
rect 15560 -5570 15740 -5560
rect 15560 -5750 15570 -5570
rect 15730 -5750 15740 -5570
rect 15560 -5760 15740 -5750
rect 14220 -6050 14360 -6040
rect 14220 -6170 14230 -6050
rect 14350 -6170 14360 -6050
rect 14220 -6180 14360 -6170
rect 15220 -6050 15360 -6040
rect 15220 -6170 15230 -6050
rect 15350 -6170 15360 -6050
rect 15220 -6180 15360 -6170
rect 14240 -11660 14340 -6180
rect 14900 -6490 15040 -6480
rect 14900 -6610 14910 -6490
rect 15030 -6610 15040 -6490
rect 14900 -6620 15040 -6610
rect 14900 -7880 15050 -7870
rect 14900 -8000 14910 -7880
rect 15040 -8000 15050 -7880
rect 14900 -8010 15050 -8000
rect 14220 -11670 14360 -11660
rect 14220 -11790 14230 -11670
rect 14350 -11790 14360 -11670
rect 14220 -11800 14360 -11790
rect 14000 -13480 14140 -13470
rect 14000 -13600 14010 -13480
rect 14130 -13600 14140 -13480
rect 14000 -13610 14140 -13600
rect 13310 -14870 13320 -14210
rect 13430 -14870 13440 -14210
rect 13310 -14960 13440 -14870
rect 13280 -14970 13470 -14960
rect 13280 -15130 13290 -14970
rect 13460 -15130 13470 -14970
rect 13280 -15140 13470 -15130
rect 13310 -15290 13440 -15280
rect 13310 -15390 13330 -15290
rect 13430 -15390 13440 -15290
rect 14020 -15300 14120 -13610
rect 13310 -16010 13440 -15390
rect 14010 -15310 14130 -15300
rect 14010 -15410 14020 -15310
rect 14120 -15410 14130 -15310
rect 14010 -15420 14130 -15410
rect 13310 -16670 13320 -16010
rect 13430 -16670 13440 -16010
rect 13310 -16680 13440 -16670
rect 13310 -16780 13430 -16680
rect 13290 -16790 13460 -16780
rect 13290 -16950 13300 -16790
rect 13450 -16950 13460 -16790
rect 13290 -16960 13460 -16950
rect 12620 -17080 12760 -17070
rect 12620 -17200 12630 -17080
rect 12750 -17200 12760 -17080
rect 12620 -17210 12760 -17200
rect 13310 -17800 13430 -16960
rect 13310 -17810 13440 -17800
rect 13310 -18470 13320 -17810
rect 13430 -18470 13440 -17810
rect 13310 -18580 13440 -18470
rect 13290 -18590 13460 -18580
rect 13290 -18750 13300 -18590
rect 13450 -18750 13460 -18590
rect 13290 -18760 13460 -18750
rect 12400 -18880 12540 -18870
rect 12400 -19000 12410 -18880
rect 12530 -19000 12540 -18880
rect 12400 -19010 12540 -19000
rect 14240 -19320 14340 -11800
rect 14910 -12090 15040 -8010
rect 15620 -8510 15720 -5760
rect 15820 -5960 15920 -4850
rect 15780 -5970 15960 -5960
rect 15780 -6150 15790 -5970
rect 15950 -6150 15960 -5970
rect 15780 -6160 15960 -6150
rect 15840 -8060 15940 -6160
rect 16500 -6270 16640 -4090
rect 17200 -4240 17300 -2580
rect 17420 -2910 17520 -1250
rect 18100 -1350 18240 -490
rect 18800 -640 18900 1020
rect 19020 690 19120 1310
rect 19010 680 19130 690
rect 19010 560 19020 680
rect 19120 560 19130 680
rect 19010 550 19130 560
rect 18790 -650 18910 -640
rect 18790 -770 18800 -650
rect 18900 -770 18910 -650
rect 18790 -780 18910 -770
rect 18100 -1510 18110 -1350
rect 18230 -1510 18240 -1350
rect 18100 -1610 18240 -1510
rect 18100 -2290 18110 -1610
rect 18230 -2290 18240 -1610
rect 17410 -2920 17530 -2910
rect 17410 -3040 17420 -2920
rect 17520 -3040 17530 -2920
rect 17410 -3050 17530 -3040
rect 17190 -4250 17310 -4240
rect 17190 -4370 17200 -4250
rect 17300 -4370 17310 -4250
rect 17190 -4380 17310 -4370
rect 16500 -6390 16510 -6270
rect 16630 -6390 16640 -6270
rect 16500 -6400 16640 -6390
rect 17200 -7160 17300 -4380
rect 17420 -4710 17520 -3050
rect 18100 -3150 18240 -2290
rect 18800 -2440 18900 -780
rect 19020 -1110 19120 550
rect 19700 450 19840 1310
rect 20400 1160 20500 1310
rect 20390 1150 20510 1160
rect 20390 1030 20400 1150
rect 20500 1030 20510 1150
rect 20390 1020 20510 1030
rect 19700 290 19710 450
rect 19830 290 19840 450
rect 19700 190 19840 290
rect 19700 -490 19710 190
rect 19830 -490 19840 190
rect 19010 -1120 19130 -1110
rect 19010 -1240 19020 -1120
rect 19120 -1240 19130 -1120
rect 19010 -1250 19130 -1240
rect 18790 -2450 18910 -2440
rect 18790 -2570 18800 -2450
rect 18900 -2570 18910 -2450
rect 18790 -2580 18910 -2570
rect 18100 -3310 18110 -3150
rect 18230 -3310 18240 -3150
rect 18100 -3410 18240 -3310
rect 18100 -4090 18110 -3410
rect 18230 -4090 18240 -3410
rect 18100 -4100 18240 -4090
rect 18800 -4240 18900 -2580
rect 19020 -2910 19120 -1250
rect 19700 -1350 19840 -490
rect 20400 -640 20500 1020
rect 20620 690 20720 1310
rect 20610 680 20730 690
rect 20610 560 20620 680
rect 20720 560 20730 680
rect 20610 550 20730 560
rect 20390 -650 20510 -640
rect 20390 -770 20400 -650
rect 20500 -770 20510 -650
rect 20390 -780 20510 -770
rect 19700 -1510 19710 -1350
rect 19830 -1510 19840 -1350
rect 19700 -1610 19840 -1510
rect 19700 -2290 19710 -1610
rect 19830 -2290 19840 -1610
rect 19010 -2920 19130 -2910
rect 19010 -3040 19020 -2920
rect 19120 -3040 19130 -2920
rect 19010 -3050 19130 -3040
rect 18790 -4250 18910 -4240
rect 18790 -4370 18800 -4250
rect 18900 -4370 18910 -4250
rect 18790 -4380 18910 -4370
rect 17410 -4720 17530 -4710
rect 17410 -4840 17420 -4720
rect 17520 -4840 17530 -4720
rect 17410 -4850 17530 -4840
rect 17420 -6760 17520 -4850
rect 18800 -5160 18900 -4380
rect 19020 -4710 19120 -3050
rect 19700 -3150 19840 -2290
rect 20400 -2440 20500 -780
rect 20620 -1110 20720 550
rect 21300 450 21440 1310
rect 22000 1160 22100 1310
rect 21990 1150 22110 1160
rect 21990 1030 22000 1150
rect 22100 1030 22110 1150
rect 21990 1020 22110 1030
rect 21300 290 21310 450
rect 21430 290 21440 450
rect 21300 190 21440 290
rect 21300 -490 21310 190
rect 21430 -490 21440 190
rect 20610 -1120 20730 -1110
rect 20610 -1240 20620 -1120
rect 20720 -1240 20730 -1120
rect 20610 -1250 20730 -1240
rect 20390 -2450 20510 -2440
rect 20390 -2570 20400 -2450
rect 20500 -2570 20510 -2450
rect 20390 -2580 20510 -2570
rect 19700 -3310 19710 -3150
rect 19830 -3310 19840 -3150
rect 19700 -3410 19840 -3310
rect 19700 -4090 19710 -3410
rect 19830 -4090 19840 -3410
rect 19700 -4100 19840 -4090
rect 20400 -4240 20500 -2580
rect 20620 -2910 20720 -1250
rect 21300 -1350 21440 -490
rect 22000 -640 22100 1020
rect 22220 690 22320 1310
rect 22210 680 22330 690
rect 22210 560 22220 680
rect 22320 560 22330 680
rect 22210 550 22330 560
rect 21990 -650 22110 -640
rect 21990 -770 22000 -650
rect 22100 -770 22110 -650
rect 21990 -780 22110 -770
rect 21300 -1510 21310 -1350
rect 21430 -1510 21440 -1350
rect 21300 -1610 21440 -1510
rect 21300 -2290 21310 -1610
rect 21430 -2290 21440 -1610
rect 20610 -2920 20730 -2910
rect 20610 -3040 20620 -2920
rect 20720 -3040 20730 -2920
rect 20610 -3050 20730 -3040
rect 20390 -4250 20510 -4240
rect 20390 -4370 20400 -4250
rect 20500 -4370 20510 -4250
rect 20390 -4380 20510 -4370
rect 19010 -4720 19130 -4710
rect 19010 -4840 19020 -4720
rect 19120 -4840 19130 -4720
rect 19010 -4850 19130 -4840
rect 18760 -5170 18940 -5160
rect 18760 -5350 18770 -5170
rect 18930 -5350 18940 -5170
rect 18760 -5360 18940 -5350
rect 18760 -5570 18940 -5560
rect 18760 -5750 18770 -5570
rect 18930 -5750 18940 -5570
rect 18760 -5760 18940 -5750
rect 17380 -6770 17560 -6760
rect 17380 -6950 17390 -6770
rect 17550 -6950 17560 -6770
rect 17380 -6960 17560 -6950
rect 17160 -7170 17340 -7160
rect 17160 -7350 17170 -7170
rect 17330 -7350 17340 -7170
rect 17160 -7360 17340 -7350
rect 17160 -7570 17340 -7560
rect 17160 -7750 17170 -7570
rect 17330 -7750 17340 -7570
rect 17160 -7760 17340 -7750
rect 15820 -8070 15960 -8060
rect 15820 -8190 15830 -8070
rect 15950 -8190 15960 -8070
rect 15820 -8200 15960 -8190
rect 15600 -8520 15740 -8510
rect 15600 -8640 15610 -8520
rect 15730 -8640 15740 -8520
rect 15600 -8650 15740 -8640
rect 15620 -10310 15720 -8650
rect 15840 -9860 15940 -8200
rect 16500 -8260 16650 -8250
rect 16500 -8380 16510 -8260
rect 16640 -8380 16650 -8260
rect 16500 -8390 16650 -8380
rect 17220 -8510 17320 -7760
rect 17440 -8060 17540 -6960
rect 17420 -8070 17560 -8060
rect 17420 -8190 17430 -8070
rect 17550 -8190 17560 -8070
rect 17420 -8200 17560 -8190
rect 17200 -8520 17340 -8510
rect 17200 -8640 17210 -8520
rect 17330 -8640 17340 -8520
rect 17200 -8650 17340 -8640
rect 16510 -8800 16640 -8790
rect 16510 -9480 16520 -8800
rect 16630 -9480 16640 -8800
rect 16510 -9560 16640 -9480
rect 16500 -9570 16650 -9560
rect 16500 -9730 16510 -9570
rect 16640 -9730 16650 -9570
rect 16500 -9740 16650 -9730
rect 15820 -9870 15960 -9860
rect 15820 -9990 15830 -9870
rect 15950 -9990 15960 -9870
rect 15820 -10000 15960 -9990
rect 15600 -10320 15740 -10310
rect 15600 -10440 15610 -10320
rect 15730 -10440 15740 -10320
rect 15600 -10450 15740 -10440
rect 14900 -12100 15050 -12090
rect 14900 -12230 14910 -12100
rect 15040 -12230 15050 -12100
rect 15620 -12110 15720 -10450
rect 15840 -11660 15940 -10000
rect 16510 -10600 16640 -9740
rect 17220 -10310 17320 -8650
rect 17440 -9860 17540 -8200
rect 18820 -8510 18920 -5760
rect 19020 -5960 19120 -4850
rect 18980 -5970 19160 -5960
rect 18980 -6150 18990 -5970
rect 19150 -6150 19160 -5970
rect 18980 -6160 19160 -6150
rect 19040 -8060 19140 -6160
rect 20400 -7160 20500 -4380
rect 20620 -4710 20720 -3050
rect 21300 -3150 21440 -2290
rect 22000 -2440 22100 -780
rect 22220 -1110 22320 550
rect 22900 450 23040 1310
rect 23600 1160 23700 1310
rect 23590 1150 23710 1160
rect 23590 1030 23600 1150
rect 23700 1030 23710 1150
rect 23590 1020 23710 1030
rect 22900 290 22910 450
rect 23030 290 23040 450
rect 22900 190 23040 290
rect 22900 -490 22910 190
rect 23030 -490 23040 190
rect 22210 -1120 22330 -1110
rect 22210 -1240 22220 -1120
rect 22320 -1240 22330 -1120
rect 22210 -1250 22330 -1240
rect 21990 -2450 22110 -2440
rect 21990 -2570 22000 -2450
rect 22100 -2570 22110 -2450
rect 21990 -2580 22110 -2570
rect 21300 -3310 21310 -3150
rect 21430 -3310 21440 -3150
rect 21300 -3410 21440 -3310
rect 21300 -4090 21310 -3410
rect 21430 -4090 21440 -3410
rect 21300 -4100 21440 -4090
rect 22000 -4240 22100 -2580
rect 22220 -2910 22320 -1250
rect 22900 -1350 23040 -490
rect 23600 -640 23700 1020
rect 23820 690 23920 1310
rect 23810 680 23930 690
rect 23810 560 23820 680
rect 23920 560 23930 680
rect 23810 550 23930 560
rect 23590 -650 23710 -640
rect 23590 -770 23600 -650
rect 23700 -770 23710 -650
rect 23590 -780 23710 -770
rect 22900 -1510 22910 -1350
rect 23030 -1510 23040 -1350
rect 22900 -1610 23040 -1510
rect 22900 -2290 22910 -1610
rect 23030 -2290 23040 -1610
rect 22210 -2920 22330 -2910
rect 22210 -3040 22220 -2920
rect 22320 -3040 22330 -2920
rect 22210 -3050 22330 -3040
rect 21990 -4250 22110 -4240
rect 21990 -4370 22000 -4250
rect 22100 -4370 22110 -4250
rect 21990 -4380 22110 -4370
rect 20610 -4720 20730 -4710
rect 20610 -4840 20620 -4720
rect 20720 -4840 20730 -4720
rect 20610 -4850 20730 -4840
rect 20620 -6760 20720 -4850
rect 22000 -5160 22100 -4380
rect 22220 -4710 22320 -3050
rect 22900 -3150 23040 -2290
rect 23600 -2440 23700 -780
rect 23820 -1110 23920 550
rect 24500 450 24640 1310
rect 24500 290 24510 450
rect 24630 290 24640 450
rect 24500 190 24640 290
rect 24500 -490 24510 190
rect 24630 -490 24640 190
rect 23810 -1120 23930 -1110
rect 23810 -1240 23820 -1120
rect 23920 -1240 23930 -1120
rect 23810 -1250 23930 -1240
rect 23590 -2450 23710 -2440
rect 23590 -2570 23600 -2450
rect 23700 -2570 23710 -2450
rect 23590 -2580 23710 -2570
rect 22900 -3310 22910 -3150
rect 23030 -3310 23040 -3150
rect 22900 -3410 23040 -3310
rect 22900 -4090 22910 -3410
rect 23030 -4090 23040 -3410
rect 22900 -4100 23040 -4090
rect 23600 -4240 23700 -2580
rect 23820 -2910 23920 -1250
rect 24500 -1350 24640 -490
rect 24500 -1510 24510 -1350
rect 24630 -1510 24640 -1350
rect 24500 -1610 24640 -1510
rect 24500 -2290 24510 -1610
rect 24630 -2290 24640 -1610
rect 23810 -2920 23930 -2910
rect 23810 -3040 23820 -2920
rect 23920 -3040 23930 -2920
rect 23810 -3050 23930 -3040
rect 23590 -4250 23710 -4240
rect 23590 -4370 23600 -4250
rect 23700 -4370 23710 -4250
rect 23590 -4380 23710 -4370
rect 22210 -4720 22330 -4710
rect 22210 -4840 22220 -4720
rect 22320 -4840 22330 -4720
rect 22210 -4850 22330 -4840
rect 21960 -5170 22140 -5160
rect 21960 -5350 21970 -5170
rect 22130 -5350 22140 -5170
rect 21960 -5360 22140 -5350
rect 21960 -5570 22140 -5560
rect 21960 -5750 21970 -5570
rect 22130 -5750 22140 -5570
rect 21960 -5760 22140 -5750
rect 20580 -6770 20760 -6760
rect 20580 -6950 20590 -6770
rect 20750 -6950 20760 -6770
rect 20580 -6960 20760 -6950
rect 20360 -7170 20540 -7160
rect 20360 -7350 20370 -7170
rect 20530 -7350 20540 -7170
rect 20360 -7360 20540 -7350
rect 20360 -7570 20540 -7560
rect 20360 -7750 20370 -7570
rect 20530 -7750 20540 -7570
rect 20360 -7760 20540 -7750
rect 19020 -8070 19160 -8060
rect 19020 -8190 19030 -8070
rect 19150 -8190 19160 -8070
rect 19020 -8200 19160 -8190
rect 18800 -8520 18940 -8510
rect 18800 -8640 18810 -8520
rect 18930 -8640 18940 -8520
rect 18800 -8650 18940 -8640
rect 18110 -8800 18240 -8790
rect 18110 -9480 18120 -8800
rect 18230 -9480 18240 -8800
rect 18110 -9560 18240 -9480
rect 18100 -9570 18250 -9560
rect 18100 -9730 18110 -9570
rect 18240 -9730 18250 -9570
rect 18100 -9740 18250 -9730
rect 17420 -9870 17560 -9860
rect 17420 -9990 17430 -9870
rect 17550 -9990 17560 -9870
rect 17420 -10000 17560 -9990
rect 17200 -10320 17340 -10310
rect 17200 -10440 17210 -10320
rect 17330 -10440 17340 -10320
rect 17200 -10450 17340 -10440
rect 16510 -11280 16520 -10600
rect 16630 -11280 16640 -10600
rect 16510 -11360 16640 -11280
rect 16500 -11370 16650 -11360
rect 16500 -11530 16510 -11370
rect 16640 -11530 16650 -11370
rect 16500 -11540 16650 -11530
rect 15820 -11670 15960 -11660
rect 15820 -11790 15830 -11670
rect 15950 -11790 15960 -11670
rect 15820 -11800 15960 -11790
rect 14900 -12240 15050 -12230
rect 15600 -12120 15740 -12110
rect 15600 -12240 15610 -12120
rect 15730 -12240 15740 -12120
rect 15600 -12250 15740 -12240
rect 14910 -12410 15040 -12400
rect 14910 -13070 14920 -12410
rect 15030 -13070 15040 -12410
rect 14910 -13160 15040 -13070
rect 14880 -13170 15070 -13160
rect 14880 -13330 14890 -13170
rect 15060 -13330 15070 -13170
rect 14880 -13340 15070 -13330
rect 14910 -14210 15040 -13340
rect 15620 -13910 15720 -12250
rect 15840 -13460 15940 -11800
rect 16510 -12400 16640 -11540
rect 17220 -12110 17320 -10450
rect 17440 -11660 17540 -10000
rect 18110 -10600 18240 -9740
rect 18820 -10310 18920 -8650
rect 19040 -9860 19140 -8200
rect 20420 -8510 20520 -7760
rect 20640 -8060 20740 -6960
rect 20620 -8070 20760 -8060
rect 20620 -8190 20630 -8070
rect 20750 -8190 20760 -8070
rect 20620 -8200 20760 -8190
rect 20400 -8520 20540 -8510
rect 20400 -8640 20410 -8520
rect 20530 -8640 20540 -8520
rect 20400 -8650 20540 -8640
rect 19710 -8800 19840 -8790
rect 19710 -9480 19720 -8800
rect 19830 -9480 19840 -8800
rect 19710 -9560 19840 -9480
rect 19700 -9570 19850 -9560
rect 19700 -9730 19710 -9570
rect 19840 -9730 19850 -9570
rect 19700 -9740 19850 -9730
rect 19020 -9870 19160 -9860
rect 19020 -9990 19030 -9870
rect 19150 -9990 19160 -9870
rect 19020 -10000 19160 -9990
rect 18800 -10320 18940 -10310
rect 18800 -10440 18810 -10320
rect 18930 -10440 18940 -10320
rect 18800 -10450 18940 -10440
rect 18110 -11280 18120 -10600
rect 18230 -11280 18240 -10600
rect 18110 -11360 18240 -11280
rect 18100 -11370 18250 -11360
rect 18100 -11530 18110 -11370
rect 18240 -11530 18250 -11370
rect 18100 -11540 18250 -11530
rect 17420 -11670 17560 -11660
rect 17420 -11790 17430 -11670
rect 17550 -11790 17560 -11670
rect 17420 -11800 17560 -11790
rect 17200 -12120 17340 -12110
rect 17200 -12240 17210 -12120
rect 17330 -12240 17340 -12120
rect 17200 -12250 17340 -12240
rect 16510 -13080 16520 -12400
rect 16630 -13080 16640 -12400
rect 16510 -13160 16640 -13080
rect 16500 -13170 16650 -13160
rect 16500 -13330 16510 -13170
rect 16640 -13330 16650 -13170
rect 16500 -13340 16650 -13330
rect 15820 -13470 15960 -13460
rect 15820 -13590 15830 -13470
rect 15950 -13590 15960 -13470
rect 15820 -13600 15960 -13590
rect 15600 -13920 15740 -13910
rect 15600 -14040 15610 -13920
rect 15730 -14040 15740 -13920
rect 15600 -14050 15740 -14040
rect 14910 -14870 14920 -14210
rect 15030 -14870 15040 -14210
rect 14910 -14960 15040 -14870
rect 14880 -14970 15070 -14960
rect 14880 -15130 14890 -14970
rect 15060 -15130 15070 -14970
rect 14880 -15140 15070 -15130
rect 14910 -15290 15040 -15280
rect 14910 -15390 14930 -15290
rect 15030 -15390 15040 -15290
rect 14910 -16010 15040 -15390
rect 15620 -15710 15720 -14050
rect 15840 -15260 15940 -13600
rect 16510 -14200 16640 -13340
rect 17220 -13910 17320 -12250
rect 17440 -13460 17540 -11800
rect 18110 -12400 18240 -11540
rect 18820 -12110 18920 -10450
rect 19040 -11660 19140 -10000
rect 19710 -10600 19840 -9740
rect 20420 -10310 20520 -8650
rect 20640 -9860 20740 -8200
rect 22020 -8510 22120 -5760
rect 22220 -5960 22320 -4850
rect 22180 -5970 22360 -5960
rect 22180 -6150 22190 -5970
rect 22350 -6150 22360 -5970
rect 22180 -6160 22360 -6150
rect 22240 -8060 22340 -6160
rect 23600 -7160 23700 -4380
rect 23820 -4710 23920 -3050
rect 24500 -3150 24640 -2290
rect 25200 -2440 25300 1310
rect 25190 -2450 25310 -2440
rect 25190 -2570 25200 -2450
rect 25300 -2570 25310 -2450
rect 25190 -2580 25310 -2570
rect 24500 -3310 24510 -3150
rect 24630 -3310 24640 -3150
rect 24500 -3410 24640 -3310
rect 24500 -4090 24510 -3410
rect 24630 -4090 24640 -3410
rect 24500 -4100 24640 -4090
rect 25200 -4240 25300 -2580
rect 25420 -2910 25520 1310
rect 26100 450 26240 1310
rect 26800 1160 26900 1310
rect 26790 1150 26910 1160
rect 26790 1030 26800 1150
rect 26900 1030 26910 1150
rect 26790 1020 26910 1030
rect 26100 290 26110 450
rect 26230 290 26240 450
rect 26100 190 26240 290
rect 26100 -490 26110 190
rect 26230 -490 26240 190
rect 26100 -1350 26240 -490
rect 26800 -640 26900 1020
rect 27020 690 27120 1310
rect 27010 680 27130 690
rect 27010 560 27020 680
rect 27120 560 27130 680
rect 27010 550 27130 560
rect 26790 -650 26910 -640
rect 26790 -770 26800 -650
rect 26900 -770 26910 -650
rect 26790 -780 26910 -770
rect 26100 -1510 26110 -1350
rect 26230 -1510 26240 -1350
rect 26100 -1610 26240 -1510
rect 26100 -2290 26110 -1610
rect 26230 -2290 26240 -1610
rect 25410 -2920 25530 -2910
rect 25410 -3040 25420 -2920
rect 25520 -3040 25530 -2920
rect 25410 -3050 25530 -3040
rect 25190 -4250 25310 -4240
rect 25190 -4370 25200 -4250
rect 25300 -4370 25310 -4250
rect 25190 -4380 25310 -4370
rect 23810 -4720 23930 -4710
rect 23810 -4840 23820 -4720
rect 23920 -4840 23930 -4720
rect 23810 -4850 23930 -4840
rect 23820 -6760 23920 -4850
rect 25200 -5160 25300 -4380
rect 25420 -4710 25520 -3050
rect 26100 -3150 26240 -2290
rect 26800 -2440 26900 -780
rect 27020 -1110 27120 550
rect 27700 450 27840 1310
rect 28400 1160 28500 1310
rect 28391 1150 28510 1160
rect 28391 1030 28400 1150
rect 28500 1030 28510 1150
rect 28391 1020 28510 1030
rect 27700 270 27710 450
rect 27830 270 27840 450
rect 27700 190 27840 270
rect 27700 -490 27710 190
rect 27830 -490 27840 190
rect 27010 -1120 27130 -1110
rect 27010 -1240 27020 -1120
rect 27120 -1240 27130 -1120
rect 27010 -1250 27130 -1240
rect 26791 -2450 26910 -2440
rect 26791 -2570 26800 -2450
rect 26900 -2570 26910 -2450
rect 26791 -2580 26910 -2570
rect 26100 -3310 26110 -3150
rect 26230 -3310 26240 -3150
rect 26100 -3410 26240 -3310
rect 26100 -4090 26110 -3410
rect 26230 -4090 26240 -3410
rect 26100 -4100 26240 -4090
rect 26800 -4240 26900 -2580
rect 27020 -2910 27120 -1250
rect 27700 -1350 27840 -490
rect 28400 -640 28500 1020
rect 28620 690 28720 1310
rect 28611 680 28730 690
rect 28611 560 28620 680
rect 28720 560 28730 680
rect 28611 550 28730 560
rect 28391 -650 28510 -640
rect 28391 -770 28400 -650
rect 28500 -770 28510 -650
rect 28391 -780 28510 -770
rect 27700 -1530 27710 -1350
rect 27830 -1530 27840 -1350
rect 27700 -1610 27840 -1530
rect 27700 -2290 27710 -1610
rect 27830 -2290 27840 -1610
rect 27011 -2920 27130 -2910
rect 27011 -3040 27020 -2920
rect 27120 -3040 27130 -2920
rect 27011 -3050 27130 -3040
rect 26791 -4250 26910 -4240
rect 26791 -4370 26800 -4250
rect 26900 -4370 26910 -4250
rect 26791 -4380 26910 -4370
rect 25410 -4720 25530 -4710
rect 25410 -4840 25420 -4720
rect 25520 -4840 25530 -4720
rect 25410 -4850 25530 -4840
rect 25160 -5170 25340 -5160
rect 25160 -5350 25170 -5170
rect 25330 -5350 25340 -5170
rect 25160 -5360 25340 -5350
rect 25160 -5570 25340 -5560
rect 25160 -5750 25170 -5570
rect 25330 -5750 25340 -5570
rect 25160 -5760 25340 -5750
rect 23780 -6770 23960 -6760
rect 23780 -6950 23790 -6770
rect 23950 -6950 23960 -6770
rect 23780 -6960 23960 -6950
rect 23560 -7170 23740 -7160
rect 23560 -7350 23570 -7170
rect 23730 -7350 23740 -7170
rect 23560 -7360 23740 -7350
rect 23560 -7570 23740 -7560
rect 23560 -7750 23570 -7570
rect 23730 -7750 23740 -7570
rect 23560 -7760 23740 -7750
rect 22220 -8070 22360 -8060
rect 22220 -8190 22230 -8070
rect 22350 -8190 22360 -8070
rect 22220 -8200 22360 -8190
rect 22000 -8520 22140 -8510
rect 22000 -8640 22010 -8520
rect 22130 -8640 22140 -8520
rect 22000 -8650 22140 -8640
rect 21310 -8800 21440 -8790
rect 21310 -9480 21320 -8800
rect 21430 -9480 21440 -8800
rect 21310 -9560 21440 -9480
rect 21300 -9570 21450 -9560
rect 21300 -9730 21310 -9570
rect 21440 -9730 21450 -9570
rect 21300 -9740 21450 -9730
rect 20620 -9870 20760 -9860
rect 20620 -9990 20630 -9870
rect 20750 -9990 20760 -9870
rect 20620 -10000 20760 -9990
rect 20400 -10320 20540 -10310
rect 20400 -10440 20410 -10320
rect 20530 -10440 20540 -10320
rect 20400 -10450 20540 -10440
rect 19710 -11280 19720 -10600
rect 19830 -11280 19840 -10600
rect 19710 -11360 19840 -11280
rect 19700 -11370 19850 -11360
rect 19700 -11530 19710 -11370
rect 19840 -11530 19850 -11370
rect 19700 -11540 19850 -11530
rect 19020 -11670 19160 -11660
rect 19020 -11790 19030 -11670
rect 19150 -11790 19160 -11670
rect 19020 -11800 19160 -11790
rect 18800 -12120 18940 -12110
rect 18800 -12240 18810 -12120
rect 18930 -12240 18940 -12120
rect 18800 -12250 18940 -12240
rect 18110 -13080 18120 -12400
rect 18230 -13080 18240 -12400
rect 18110 -13160 18240 -13080
rect 18100 -13170 18250 -13160
rect 18100 -13330 18110 -13170
rect 18240 -13330 18250 -13170
rect 18100 -13340 18250 -13330
rect 17420 -13470 17560 -13460
rect 17420 -13590 17430 -13470
rect 17550 -13590 17560 -13470
rect 17420 -13600 17560 -13590
rect 17200 -13920 17340 -13910
rect 17200 -14040 17210 -13920
rect 17330 -14040 17340 -13920
rect 17200 -14050 17340 -14040
rect 16510 -14880 16520 -14200
rect 16630 -14880 16640 -14200
rect 16510 -14960 16640 -14880
rect 16500 -14970 16650 -14960
rect 16500 -15130 16510 -14970
rect 16640 -15130 16650 -14970
rect 16500 -15140 16650 -15130
rect 15820 -15270 15960 -15260
rect 15820 -15390 15830 -15270
rect 15950 -15390 15960 -15270
rect 15820 -15400 15960 -15390
rect 15600 -15720 15740 -15710
rect 15600 -15840 15610 -15720
rect 15730 -15840 15740 -15720
rect 15600 -15850 15740 -15840
rect 14910 -16670 14920 -16010
rect 15030 -16670 15040 -16010
rect 14910 -16680 15040 -16670
rect 14910 -16780 15030 -16680
rect 14890 -16790 15060 -16780
rect 14890 -16950 14900 -16790
rect 15050 -16950 15060 -16790
rect 14890 -16960 15060 -16950
rect 14910 -17800 15030 -16960
rect 15620 -17510 15720 -15850
rect 15840 -17060 15940 -15400
rect 16510 -16000 16640 -15140
rect 17220 -15710 17320 -14050
rect 17440 -15260 17540 -13600
rect 18110 -14200 18240 -13340
rect 18820 -13910 18920 -12250
rect 19040 -13460 19140 -11800
rect 19710 -12400 19840 -11540
rect 20420 -12110 20520 -10450
rect 20640 -11660 20740 -10000
rect 21310 -10600 21440 -9740
rect 22020 -10310 22120 -8650
rect 22240 -9860 22340 -8200
rect 23620 -8510 23720 -7760
rect 23840 -8060 23940 -6960
rect 23820 -8070 23960 -8060
rect 23820 -8190 23830 -8070
rect 23950 -8190 23960 -8070
rect 23820 -8200 23960 -8190
rect 23600 -8520 23740 -8510
rect 23600 -8640 23610 -8520
rect 23730 -8640 23740 -8520
rect 23600 -8650 23740 -8640
rect 22910 -8800 23040 -8790
rect 22910 -9480 22920 -8800
rect 23030 -9480 23040 -8800
rect 22910 -9560 23040 -9480
rect 22900 -9570 23050 -9560
rect 22900 -9730 22910 -9570
rect 23040 -9730 23050 -9570
rect 22900 -9740 23050 -9730
rect 22220 -9870 22360 -9860
rect 22220 -9990 22230 -9870
rect 22350 -9990 22360 -9870
rect 22220 -10000 22360 -9990
rect 22000 -10320 22140 -10310
rect 22000 -10440 22010 -10320
rect 22130 -10440 22140 -10320
rect 22000 -10450 22140 -10440
rect 21310 -11280 21320 -10600
rect 21430 -11280 21440 -10600
rect 21310 -11360 21440 -11280
rect 21300 -11370 21450 -11360
rect 21300 -11530 21310 -11370
rect 21440 -11530 21450 -11370
rect 21300 -11540 21450 -11530
rect 20620 -11670 20760 -11660
rect 20620 -11790 20630 -11670
rect 20750 -11790 20760 -11670
rect 20620 -11800 20760 -11790
rect 20400 -12120 20540 -12110
rect 20400 -12240 20410 -12120
rect 20530 -12240 20540 -12120
rect 20400 -12250 20540 -12240
rect 19710 -13080 19720 -12400
rect 19830 -13080 19840 -12400
rect 19710 -13160 19840 -13080
rect 19700 -13170 19850 -13160
rect 19700 -13330 19710 -13170
rect 19840 -13330 19850 -13170
rect 19700 -13340 19850 -13330
rect 19020 -13470 19160 -13460
rect 19020 -13590 19030 -13470
rect 19150 -13590 19160 -13470
rect 19020 -13600 19160 -13590
rect 18800 -13920 18940 -13910
rect 18800 -14040 18810 -13920
rect 18930 -14040 18940 -13920
rect 18800 -14050 18940 -14040
rect 18110 -14880 18120 -14200
rect 18230 -14880 18240 -14200
rect 18110 -14960 18240 -14880
rect 18100 -14970 18250 -14960
rect 18100 -15130 18110 -14970
rect 18240 -15130 18250 -14970
rect 18100 -15140 18250 -15130
rect 17420 -15270 17560 -15260
rect 17420 -15390 17430 -15270
rect 17550 -15390 17560 -15270
rect 17420 -15400 17560 -15390
rect 17200 -15720 17340 -15710
rect 17200 -15840 17210 -15720
rect 17330 -15840 17340 -15720
rect 17200 -15850 17340 -15840
rect 16510 -16680 16520 -16000
rect 16630 -16680 16640 -16000
rect 16510 -16760 16640 -16680
rect 16500 -16770 16650 -16760
rect 16500 -16930 16510 -16770
rect 16640 -16930 16650 -16770
rect 16500 -16940 16650 -16930
rect 15820 -17070 15960 -17060
rect 15820 -17190 15830 -17070
rect 15950 -17190 15960 -17070
rect 15820 -17200 15960 -17190
rect 15600 -17520 15740 -17510
rect 15600 -17640 15610 -17520
rect 15730 -17640 15740 -17520
rect 15600 -17650 15740 -17640
rect 14910 -17810 15040 -17800
rect 14910 -18470 14920 -17810
rect 15030 -18470 15040 -17810
rect 14910 -18580 15040 -18470
rect 14890 -18590 15060 -18580
rect 14890 -18750 14900 -18590
rect 15050 -18750 15060 -18590
rect 14890 -18760 15060 -18750
rect 15620 -19310 15720 -17650
rect 15840 -18860 15940 -17200
rect 16510 -17800 16640 -16940
rect 17220 -17510 17320 -15850
rect 17440 -17060 17540 -15400
rect 18110 -16000 18240 -15140
rect 18820 -15710 18920 -14050
rect 19040 -15260 19140 -13600
rect 19710 -14200 19840 -13340
rect 20420 -13910 20520 -12250
rect 20640 -13460 20740 -11800
rect 21310 -12400 21440 -11540
rect 22020 -12110 22120 -10450
rect 22240 -11660 22340 -10000
rect 22910 -10600 23040 -9740
rect 23620 -10310 23720 -8650
rect 23840 -9860 23940 -8200
rect 25220 -8510 25320 -5760
rect 25420 -5960 25520 -4850
rect 25380 -5970 25560 -5960
rect 25380 -6150 25390 -5970
rect 25550 -6150 25560 -5970
rect 25380 -6160 25560 -6150
rect 25440 -8060 25540 -6160
rect 26800 -7160 26900 -4380
rect 27020 -4710 27120 -3050
rect 27700 -3150 27840 -2290
rect 28400 -2440 28500 -780
rect 28620 -1110 28720 550
rect 29300 450 29440 1310
rect 29300 270 29310 450
rect 29430 270 29440 450
rect 29300 190 29440 270
rect 29300 -490 29310 190
rect 29430 -490 29440 190
rect 28611 -1120 28730 -1110
rect 28611 -1240 28620 -1120
rect 28720 -1240 28730 -1120
rect 28611 -1250 28730 -1240
rect 28390 -2450 28510 -2440
rect 28390 -2570 28400 -2450
rect 28500 -2570 28510 -2450
rect 28390 -2580 28510 -2570
rect 27700 -3330 27710 -3150
rect 27830 -3330 27840 -3150
rect 27700 -3410 27840 -3330
rect 27700 -4090 27710 -3410
rect 27830 -4090 27840 -3410
rect 27011 -4720 27130 -4710
rect 27011 -4840 27020 -4720
rect 27120 -4840 27130 -4720
rect 27011 -4850 27130 -4840
rect 27020 -6760 27120 -4850
rect 27700 -5960 27840 -4090
rect 28400 -4240 28500 -2580
rect 28620 -2910 28720 -1250
rect 29300 -1350 29440 -490
rect 29300 -1530 29310 -1350
rect 29430 -1530 29440 -1350
rect 29300 -1610 29440 -1530
rect 29300 -2290 29310 -1610
rect 29430 -2290 29440 -1610
rect 28610 -2920 28730 -2910
rect 28610 -3040 28620 -2920
rect 28720 -3040 28730 -2920
rect 28610 -3050 28730 -3040
rect 28390 -4250 28510 -4240
rect 28390 -4370 28400 -4250
rect 28500 -4370 28510 -4250
rect 28390 -4380 28510 -4370
rect 28400 -5160 28500 -4380
rect 28620 -4710 28720 -3050
rect 29300 -3150 29440 -2290
rect 30900 2250 31040 2260
rect 30900 2070 30910 2250
rect 31030 2070 31040 2250
rect 30900 1990 31040 2070
rect 30900 1310 30910 1990
rect 31030 1310 31040 1990
rect 30900 450 31040 1310
rect 30900 270 30910 450
rect 31030 270 31040 450
rect 30900 190 31040 270
rect 30900 -490 30910 190
rect 31030 -490 31040 190
rect 30900 -1350 31040 -490
rect 31600 -1110 31700 3540
rect 32530 3162 32620 4330
rect 33120 4110 33300 4120
rect 33120 4080 33130 4110
rect 32800 4070 33130 4080
rect 33290 4080 33300 4110
rect 33290 4070 33940 4080
rect 32800 4010 32810 4070
rect 32980 4010 33130 4070
rect 33300 4010 33440 4070
rect 33610 4010 33760 4070
rect 33930 4010 33940 4070
rect 32800 4000 33940 4010
rect 32840 3430 33880 3440
rect 32840 3350 32850 3430
rect 33870 3350 33880 3430
rect 32840 3340 33880 3350
rect 32460 3156 32674 3162
rect 31820 3090 32000 3100
rect 31820 2910 31830 3090
rect 31990 2910 32000 3090
rect 32460 3068 32466 3156
rect 32668 3068 32674 3156
rect 32460 3062 32674 3068
rect 31820 2900 32000 2910
rect 31820 690 31920 2900
rect 33170 2550 33340 2560
rect 32440 2510 32700 2520
rect 32440 2430 32450 2510
rect 32690 2430 32700 2510
rect 32440 2130 32700 2430
rect 33170 2390 33180 2550
rect 33330 2390 33340 2550
rect 33170 2380 33340 2390
rect 32440 2070 32450 2130
rect 32690 2070 32700 2130
rect 32440 2060 32700 2070
rect 32500 1990 32640 2000
rect 32500 1310 32510 1990
rect 32630 1310 32640 1990
rect 32500 1150 32640 1310
rect 32500 1030 32510 1150
rect 32630 1030 32640 1150
rect 32500 1020 32640 1030
rect 31810 680 31930 690
rect 31810 560 31820 680
rect 31920 560 31930 680
rect 31810 550 31930 560
rect 33190 450 33320 2380
rect 33170 440 33340 450
rect 33170 280 33180 440
rect 33330 280 33340 440
rect 33170 270 33340 280
rect 32500 190 32640 200
rect 32500 -490 32510 190
rect 32630 -490 32640 190
rect 32500 -500 32640 -490
rect 31590 -1120 31710 -1110
rect 31590 -1240 31600 -1120
rect 31700 -1240 31710 -1120
rect 31590 -1250 31710 -1240
rect 30900 -1530 30910 -1350
rect 31030 -1530 31040 -1350
rect 33440 -1460 33560 3340
rect 34120 3162 34210 4330
rect 35690 4290 35850 4300
rect 35690 4150 35700 4290
rect 35840 4150 35850 4290
rect 35690 4140 35850 4150
rect 36290 4260 36300 4330
rect 36390 4260 36400 4330
rect 34860 4090 35200 4100
rect 34860 4010 34870 4090
rect 35190 4010 35200 4090
rect 34860 4000 35200 4010
rect 35040 3430 35420 3440
rect 35040 3350 35070 3430
rect 35410 3350 35420 3430
rect 35040 3340 35420 3350
rect 34060 3156 34274 3162
rect 34060 3068 34066 3156
rect 34268 3068 34274 3156
rect 34060 3062 34274 3068
rect 34770 2780 34940 2790
rect 34770 2620 34780 2780
rect 34930 2620 34940 2780
rect 34770 2610 34940 2620
rect 34040 2510 34300 2520
rect 34040 2430 34050 2510
rect 34290 2430 34300 2510
rect 34040 2130 34300 2430
rect 34040 2070 34050 2130
rect 34290 2070 34300 2130
rect 34040 2060 34300 2070
rect 34100 1990 34240 2000
rect 34100 1310 34110 1990
rect 34230 1310 34240 1990
rect 34100 1150 34240 1310
rect 34790 1160 34920 2610
rect 34100 1030 34110 1150
rect 34230 1030 34240 1150
rect 34100 1020 34240 1030
rect 34780 1150 34930 1160
rect 34780 1030 34790 1150
rect 34920 1030 34930 1150
rect 34780 1020 34930 1030
rect 34100 190 34240 200
rect 34100 -490 34110 190
rect 34230 -490 34240 190
rect 34100 -500 34240 -490
rect 30900 -1610 31040 -1530
rect 33350 -1470 33560 -1460
rect 33350 -1590 33360 -1470
rect 33480 -1590 33560 -1470
rect 33350 -1600 33560 -1590
rect 30900 -2290 30910 -1610
rect 31030 -2290 31040 -1610
rect 29990 -2450 30110 -2440
rect 29990 -2570 30000 -2450
rect 30100 -2570 30110 -2450
rect 29990 -2580 30110 -2570
rect 29300 -3330 29310 -3150
rect 29430 -3330 29440 -3150
rect 29300 -3410 29440 -3330
rect 29300 -4090 29310 -3410
rect 29430 -4090 29440 -3410
rect 28610 -4720 28730 -4710
rect 28610 -4840 28620 -4720
rect 28720 -4840 28730 -4720
rect 28610 -4850 28730 -4840
rect 28360 -5170 28540 -5160
rect 28360 -5350 28370 -5170
rect 28530 -5350 28540 -5170
rect 28360 -5360 28540 -5350
rect 28360 -5570 28540 -5560
rect 28360 -5750 28370 -5570
rect 28530 -5750 28540 -5570
rect 28360 -5760 28540 -5750
rect 27680 -5970 27860 -5960
rect 27680 -6150 27690 -5970
rect 27850 -6150 27860 -5970
rect 27680 -6160 27860 -6150
rect 26980 -6770 27160 -6760
rect 26980 -6950 26990 -6770
rect 27150 -6950 27160 -6770
rect 26980 -6960 27160 -6950
rect 26760 -7170 26940 -7160
rect 26760 -7350 26770 -7170
rect 26930 -7350 26940 -7170
rect 26760 -7360 26940 -7350
rect 26760 -7570 26940 -7560
rect 26760 -7750 26770 -7570
rect 26930 -7750 26940 -7570
rect 26760 -7760 26940 -7750
rect 25420 -8070 25560 -8060
rect 25420 -8190 25430 -8070
rect 25550 -8190 25560 -8070
rect 25420 -8200 25560 -8190
rect 25200 -8520 25340 -8510
rect 25200 -8640 25210 -8520
rect 25330 -8640 25340 -8520
rect 25200 -8650 25340 -8640
rect 24510 -8800 24640 -8790
rect 24510 -9480 24520 -8800
rect 24630 -9480 24640 -8800
rect 24510 -9560 24640 -9480
rect 24500 -9570 24650 -9560
rect 24500 -9730 24510 -9570
rect 24640 -9730 24650 -9570
rect 24500 -9740 24650 -9730
rect 23820 -9870 23960 -9860
rect 23820 -9990 23830 -9870
rect 23950 -9990 23960 -9870
rect 23820 -10000 23960 -9990
rect 23600 -10320 23740 -10310
rect 23600 -10440 23610 -10320
rect 23730 -10440 23740 -10320
rect 23600 -10450 23740 -10440
rect 22910 -11280 22920 -10600
rect 23030 -11280 23040 -10600
rect 22910 -11360 23040 -11280
rect 22900 -11370 23050 -11360
rect 22900 -11530 22910 -11370
rect 23040 -11530 23050 -11370
rect 22900 -11540 23050 -11530
rect 22220 -11670 22360 -11660
rect 22220 -11790 22230 -11670
rect 22350 -11790 22360 -11670
rect 22220 -11800 22360 -11790
rect 22000 -12120 22140 -12110
rect 22000 -12240 22010 -12120
rect 22130 -12240 22140 -12120
rect 22000 -12250 22140 -12240
rect 21310 -13080 21320 -12400
rect 21430 -13080 21440 -12400
rect 21310 -13160 21440 -13080
rect 21300 -13170 21450 -13160
rect 21300 -13330 21310 -13170
rect 21440 -13330 21450 -13170
rect 21300 -13340 21450 -13330
rect 20620 -13470 20760 -13460
rect 20620 -13590 20630 -13470
rect 20750 -13590 20760 -13470
rect 20620 -13600 20760 -13590
rect 20400 -13920 20540 -13910
rect 20400 -14040 20410 -13920
rect 20530 -14040 20540 -13920
rect 20400 -14050 20540 -14040
rect 19710 -14880 19720 -14200
rect 19830 -14880 19840 -14200
rect 19710 -14960 19840 -14880
rect 19700 -14970 19850 -14960
rect 19700 -15130 19710 -14970
rect 19840 -15130 19850 -14970
rect 19700 -15140 19850 -15130
rect 19020 -15270 19160 -15260
rect 19020 -15390 19030 -15270
rect 19150 -15390 19160 -15270
rect 19020 -15400 19160 -15390
rect 18800 -15720 18940 -15710
rect 18800 -15840 18810 -15720
rect 18930 -15840 18940 -15720
rect 18800 -15850 18940 -15840
rect 18110 -16680 18120 -16000
rect 18230 -16680 18240 -16000
rect 18110 -16760 18240 -16680
rect 18100 -16770 18250 -16760
rect 18100 -16930 18110 -16770
rect 18240 -16930 18250 -16770
rect 18100 -16940 18250 -16930
rect 17420 -17070 17560 -17060
rect 17420 -17190 17430 -17070
rect 17550 -17190 17560 -17070
rect 17420 -17200 17560 -17190
rect 17200 -17520 17340 -17510
rect 17200 -17640 17210 -17520
rect 17330 -17640 17340 -17520
rect 17200 -17650 17340 -17640
rect 16510 -18480 16520 -17800
rect 16630 -18480 16640 -17800
rect 16510 -18560 16640 -18480
rect 16500 -18570 16650 -18560
rect 16500 -18730 16510 -18570
rect 16640 -18730 16650 -18570
rect 16500 -18740 16650 -18730
rect 15820 -18870 15960 -18860
rect 15820 -18990 15830 -18870
rect 15950 -18990 15960 -18870
rect 15820 -19000 15960 -18990
rect 15600 -19320 15740 -19310
rect 13310 -19440 15040 -19320
rect 13310 -19610 13440 -19440
rect 13310 -20270 13320 -19610
rect 13430 -20270 13440 -19610
rect 13310 -20280 13440 -20270
rect 14910 -19610 15040 -19440
rect 15600 -19440 15610 -19320
rect 15730 -19440 15740 -19320
rect 15600 -19450 15740 -19440
rect 14910 -20270 14920 -19610
rect 15030 -20270 15040 -19610
rect 14910 -20280 15040 -20270
rect 11030 -20560 11150 -20380
rect 10800 -20860 10940 -20850
rect 10800 -20980 10810 -20860
rect 10930 -20980 10940 -20860
rect 10800 -20990 10940 -20980
rect 10120 -22070 10130 -21410
rect 10230 -22070 10240 -21410
rect 10120 -22190 10240 -22070
rect 10820 -22190 10920 -20990
rect 11040 -22180 11140 -20560
rect 12400 -20680 12540 -20670
rect 12400 -20800 12410 -20680
rect 12530 -20800 12540 -20680
rect 12400 -20810 12540 -20800
rect 11700 -21400 11850 -21390
rect 11700 -22080 11710 -21400
rect 11840 -22080 11850 -21400
rect 11700 -22090 11850 -22080
rect 10120 -22350 10130 -22190
rect 10230 -22350 10240 -22190
rect 10120 -22440 10240 -22350
rect 11030 -22360 11150 -22180
rect 10100 -22450 10260 -22440
rect 10100 -22590 10110 -22450
rect 10250 -22590 10260 -22450
rect 10100 -22600 10260 -22590
rect 11040 -22730 11150 -22360
rect 11720 -22730 11830 -22090
rect 11040 -22740 11160 -22730
rect 11040 -22850 11050 -22740
rect 11150 -22850 11160 -22740
rect 11040 -22860 11160 -22850
rect 11710 -22740 11830 -22730
rect 11710 -22850 11720 -22740
rect 11820 -22850 11830 -22740
rect 11710 -22860 11830 -22850
rect 12420 -22970 12520 -20810
rect 15620 -21110 15720 -19450
rect 15840 -20660 15940 -19000
rect 16510 -19600 16640 -18740
rect 17220 -19310 17320 -17650
rect 17440 -18860 17540 -17200
rect 18110 -17800 18240 -16940
rect 18820 -17510 18920 -15850
rect 19040 -17060 19140 -15400
rect 19710 -16000 19840 -15140
rect 20420 -15710 20520 -14050
rect 20640 -15260 20740 -13600
rect 21310 -14200 21440 -13340
rect 22020 -13910 22120 -12250
rect 22240 -13460 22340 -11800
rect 22910 -12400 23040 -11540
rect 23620 -12110 23720 -10450
rect 23840 -11660 23940 -10000
rect 24510 -10600 24640 -9740
rect 25220 -10310 25320 -8650
rect 25440 -9860 25540 -8200
rect 26820 -8510 26920 -7760
rect 27040 -8060 27140 -6960
rect 27020 -8070 27160 -8060
rect 27020 -8190 27030 -8070
rect 27150 -8190 27160 -8070
rect 27020 -8200 27160 -8190
rect 26800 -8520 26940 -8510
rect 26800 -8640 26810 -8520
rect 26930 -8640 26940 -8520
rect 26800 -8650 26940 -8640
rect 26110 -8800 26240 -8790
rect 26110 -9480 26120 -8800
rect 26230 -9480 26240 -8800
rect 26110 -9560 26240 -9480
rect 26100 -9570 26250 -9560
rect 26100 -9730 26110 -9570
rect 26240 -9730 26250 -9570
rect 26100 -9740 26250 -9730
rect 25420 -9870 25560 -9860
rect 25420 -9990 25430 -9870
rect 25550 -9990 25560 -9870
rect 25420 -10000 25560 -9990
rect 25200 -10320 25340 -10310
rect 25200 -10440 25210 -10320
rect 25330 -10440 25340 -10320
rect 25200 -10450 25340 -10440
rect 24510 -11280 24520 -10600
rect 24630 -11280 24640 -10600
rect 24510 -11360 24640 -11280
rect 24500 -11370 24650 -11360
rect 24500 -11530 24510 -11370
rect 24640 -11530 24650 -11370
rect 24500 -11540 24650 -11530
rect 23820 -11670 23960 -11660
rect 23820 -11790 23830 -11670
rect 23950 -11790 23960 -11670
rect 23820 -11800 23960 -11790
rect 23600 -12120 23740 -12110
rect 23600 -12240 23610 -12120
rect 23730 -12240 23740 -12120
rect 23600 -12250 23740 -12240
rect 22910 -13080 22920 -12400
rect 23030 -13080 23040 -12400
rect 22910 -13160 23040 -13080
rect 22900 -13170 23050 -13160
rect 22900 -13330 22910 -13170
rect 23040 -13330 23050 -13170
rect 22900 -13340 23050 -13330
rect 22220 -13470 22360 -13460
rect 22220 -13590 22230 -13470
rect 22350 -13590 22360 -13470
rect 22220 -13600 22360 -13590
rect 22000 -13920 22140 -13910
rect 22000 -14040 22010 -13920
rect 22130 -14040 22140 -13920
rect 22000 -14050 22140 -14040
rect 21310 -14880 21320 -14200
rect 21430 -14880 21440 -14200
rect 21310 -14960 21440 -14880
rect 21300 -14970 21450 -14960
rect 21300 -15130 21310 -14970
rect 21440 -15130 21450 -14970
rect 21300 -15140 21450 -15130
rect 20620 -15270 20760 -15260
rect 20620 -15390 20630 -15270
rect 20750 -15390 20760 -15270
rect 20620 -15400 20760 -15390
rect 20400 -15720 20540 -15710
rect 20400 -15840 20410 -15720
rect 20530 -15840 20540 -15720
rect 20400 -15850 20540 -15840
rect 19710 -16680 19720 -16000
rect 19830 -16680 19840 -16000
rect 19710 -16760 19840 -16680
rect 19700 -16770 19850 -16760
rect 19700 -16930 19710 -16770
rect 19840 -16930 19850 -16770
rect 19700 -16940 19850 -16930
rect 19020 -17070 19160 -17060
rect 19020 -17190 19030 -17070
rect 19150 -17190 19160 -17070
rect 19020 -17200 19160 -17190
rect 18800 -17520 18940 -17510
rect 18800 -17640 18810 -17520
rect 18930 -17640 18940 -17520
rect 18800 -17650 18940 -17640
rect 18110 -18480 18120 -17800
rect 18230 -18480 18240 -17800
rect 18110 -18560 18240 -18480
rect 18100 -18570 18250 -18560
rect 18100 -18730 18110 -18570
rect 18240 -18730 18250 -18570
rect 18100 -18740 18250 -18730
rect 17420 -18870 17560 -18860
rect 17420 -18990 17430 -18870
rect 17550 -18990 17560 -18870
rect 17420 -19000 17560 -18990
rect 17200 -19320 17340 -19310
rect 17200 -19440 17210 -19320
rect 17330 -19440 17340 -19320
rect 17200 -19450 17340 -19440
rect 16510 -20280 16520 -19600
rect 16630 -20280 16640 -19600
rect 16510 -20360 16640 -20280
rect 16500 -20370 16650 -20360
rect 16500 -20530 16510 -20370
rect 16640 -20530 16650 -20370
rect 16500 -20540 16650 -20530
rect 15820 -20670 15960 -20660
rect 15820 -20790 15830 -20670
rect 15950 -20790 15960 -20670
rect 15820 -20800 15960 -20790
rect 15600 -21120 15740 -21110
rect 15600 -21240 15610 -21120
rect 15730 -21240 15740 -21120
rect 15600 -21250 15740 -21240
rect 15620 -21370 15720 -21250
rect 15840 -21370 15940 -20800
rect 16510 -21400 16640 -20540
rect 17220 -21110 17320 -19450
rect 17440 -20660 17540 -19000
rect 18110 -19600 18240 -18740
rect 18820 -19310 18920 -17650
rect 19040 -18860 19140 -17200
rect 19710 -17800 19840 -16940
rect 20420 -17510 20520 -15850
rect 20640 -17060 20740 -15400
rect 21310 -16000 21440 -15140
rect 22020 -15710 22120 -14050
rect 22240 -15260 22340 -13600
rect 22910 -14200 23040 -13340
rect 23620 -13910 23720 -12250
rect 23840 -13460 23940 -11800
rect 24510 -12400 24640 -11540
rect 25220 -12110 25320 -10450
rect 25440 -11660 25540 -10000
rect 26110 -10600 26240 -9740
rect 26820 -10310 26920 -8650
rect 27040 -9860 27140 -8200
rect 28420 -8510 28520 -5760
rect 28620 -5960 28720 -4850
rect 29300 -5960 29440 -4090
rect 30000 -4240 30100 -2580
rect 30210 -2920 30330 -2910
rect 30210 -3040 30220 -2920
rect 30320 -3040 30330 -2920
rect 30210 -3050 30330 -3040
rect 29990 -4250 30110 -4240
rect 29990 -4370 30000 -4250
rect 30100 -4370 30110 -4250
rect 29990 -4380 30110 -4370
rect 28580 -5970 28760 -5960
rect 28580 -6150 28590 -5970
rect 28750 -6150 28760 -5970
rect 28580 -6160 28760 -6150
rect 29280 -5970 29460 -5960
rect 29280 -6150 29290 -5970
rect 29450 -6150 29460 -5970
rect 29280 -6160 29460 -6150
rect 28640 -8060 28740 -6160
rect 30000 -7160 30100 -4380
rect 30220 -4710 30320 -3050
rect 30900 -3150 31040 -2290
rect 30900 -3330 30910 -3150
rect 31030 -3330 31040 -3150
rect 30900 -3410 31040 -3330
rect 30900 -4090 30910 -3410
rect 31030 -4090 31040 -3410
rect 30210 -4720 30330 -4710
rect 30210 -4840 30220 -4720
rect 30320 -4840 30330 -4720
rect 30210 -4850 30330 -4840
rect 30220 -6760 30320 -4850
rect 30900 -5960 31040 -4090
rect 32500 -1610 32640 -1600
rect 32500 -2290 32510 -1610
rect 32630 -2290 32640 -1610
rect 32500 -2450 32640 -2290
rect 32500 -2570 32510 -2450
rect 32630 -2570 32640 -2450
rect 32500 -3410 32640 -2570
rect 32500 -4090 32510 -3410
rect 32630 -4090 32640 -3410
rect 32500 -4100 32640 -4090
rect 33170 -2450 33310 -2440
rect 33170 -2570 33180 -2450
rect 33300 -2570 33310 -2450
rect 33170 -4250 33310 -2570
rect 33440 -3270 33560 -1600
rect 33390 -3280 33560 -3270
rect 33390 -3400 33400 -3280
rect 33530 -3400 33560 -3280
rect 33390 -3410 33560 -3400
rect 33440 -3660 33560 -3410
rect 34100 -1610 34240 -1600
rect 34100 -2290 34110 -1610
rect 34230 -2290 34240 -1610
rect 34100 -2450 34240 -2290
rect 34790 -2440 34920 1020
rect 35040 -1460 35160 3340
rect 35720 3162 35810 4140
rect 36290 4070 36400 4260
rect 36290 4000 36300 4070
rect 36390 4000 36400 4070
rect 36290 3990 36400 4000
rect 37670 5890 37780 5900
rect 37670 5820 37680 5890
rect 37770 5820 37780 5890
rect 37670 5630 37780 5820
rect 37670 5560 37680 5630
rect 37770 5560 37780 5630
rect 37670 5370 37780 5560
rect 37670 5040 37680 5370
rect 37770 5040 37780 5370
rect 37670 4850 37780 5040
rect 37670 4780 37680 4850
rect 37770 4780 37780 4850
rect 37670 4590 37780 4780
rect 37670 4520 37680 4590
rect 37770 4520 37780 4590
rect 37670 4330 37780 4520
rect 37670 4260 37680 4330
rect 37770 4260 37780 4330
rect 37670 4070 37780 4260
rect 37670 4000 37680 4070
rect 37770 4000 37780 4070
rect 37670 3990 37780 4000
rect 37870 3710 38020 3720
rect 36370 3580 36530 3590
rect 36370 3440 36380 3580
rect 36520 3440 36530 3580
rect 37870 3580 37880 3710
rect 38010 3580 38020 3710
rect 37870 3570 38020 3580
rect 36370 3430 36530 3440
rect 35660 3156 35874 3162
rect 35660 3068 35666 3156
rect 35868 3068 35874 3156
rect 35660 3062 35874 3068
rect 35640 2510 35900 2520
rect 35640 2430 35650 2510
rect 35890 2430 35900 2510
rect 35640 2130 35900 2430
rect 35640 2070 35650 2130
rect 35890 2070 35900 2130
rect 35640 2060 35900 2070
rect 35700 1990 35840 2000
rect 35700 1310 35710 1990
rect 35830 1310 35840 1990
rect 35700 1150 35840 1310
rect 35700 1030 35710 1150
rect 35830 1030 35840 1150
rect 35700 1020 35840 1030
rect 35700 190 35840 200
rect 35700 -490 35710 190
rect 35830 -490 35840 190
rect 35700 -500 35840 -490
rect 35010 -1470 35160 -1460
rect 35010 -1590 35020 -1470
rect 35140 -1570 35160 -1470
rect 35140 -1590 35150 -1570
rect 35010 -1600 35150 -1590
rect 35680 -1600 35760 -1590
rect 35680 -2310 35690 -1600
rect 35750 -2310 35760 -1600
rect 35680 -2350 35760 -2310
rect 35700 -2360 35760 -2350
rect 34100 -2570 34110 -2450
rect 34230 -2570 34240 -2450
rect 34100 -3410 34240 -2570
rect 34780 -2450 34930 -2440
rect 34780 -2570 34790 -2450
rect 34920 -2570 34930 -2450
rect 34780 -2580 34930 -2570
rect 35700 -2450 35840 -2360
rect 35700 -2570 35710 -2450
rect 35830 -2570 35840 -2450
rect 34100 -4090 34110 -3410
rect 34230 -4090 34240 -3410
rect 34100 -4100 34240 -4090
rect 35700 -3410 35840 -2570
rect 36400 -2900 36500 3430
rect 36580 3360 36740 3370
rect 36580 3220 36590 3360
rect 36730 3220 36740 3360
rect 36580 3210 36740 3220
rect 36600 680 36720 3210
rect 37300 1990 37440 2000
rect 37300 1310 37310 1990
rect 37430 1310 37440 1990
rect 37300 1150 37440 1310
rect 37300 1030 37310 1150
rect 37430 1030 37440 1150
rect 37300 1020 37440 1030
rect 36590 670 36730 680
rect 36590 550 36600 670
rect 36720 550 36730 670
rect 37900 660 38020 3570
rect 36590 540 36730 550
rect 37840 650 38020 660
rect 37840 530 37850 650
rect 37970 530 38020 650
rect 37840 520 38020 530
rect 36390 -2910 36510 -2900
rect 36390 -3030 36400 -2910
rect 36500 -3030 36510 -2910
rect 36390 -3040 36510 -3030
rect 35700 -4090 35710 -3410
rect 35830 -4090 35840 -3410
rect 35700 -4100 35840 -4090
rect 33170 -4370 33180 -4250
rect 33300 -4370 33310 -4250
rect 33170 -4380 33310 -4370
rect 36400 -4700 36500 -3040
rect 36390 -4710 36510 -4700
rect 36390 -4830 36400 -4710
rect 36500 -4830 36510 -4710
rect 36390 -4840 36510 -4830
rect 30880 -5970 31060 -5960
rect 30880 -6150 30890 -5970
rect 31050 -6150 31060 -5970
rect 30880 -6160 31060 -6150
rect 30180 -6770 30360 -6760
rect 30180 -6950 30190 -6770
rect 30350 -6950 30360 -6770
rect 30180 -6960 30360 -6950
rect 29960 -7170 30140 -7160
rect 29960 -7350 29970 -7170
rect 30130 -7350 30140 -7170
rect 29960 -7360 30140 -7350
rect 29960 -7570 30140 -7560
rect 29960 -7750 29970 -7570
rect 30130 -7750 30140 -7570
rect 29960 -7760 30140 -7750
rect 28620 -8070 28760 -8060
rect 28620 -8190 28630 -8070
rect 28750 -8190 28760 -8070
rect 28620 -8200 28760 -8190
rect 28400 -8520 28540 -8510
rect 28400 -8640 28410 -8520
rect 28530 -8640 28540 -8520
rect 28400 -8650 28540 -8640
rect 27710 -8800 27840 -8790
rect 27710 -9480 27720 -8800
rect 27830 -9480 27840 -8800
rect 27710 -9560 27840 -9480
rect 27700 -9570 27850 -9560
rect 27700 -9730 27710 -9570
rect 27840 -9730 27850 -9570
rect 27700 -9740 27850 -9730
rect 27020 -9870 27160 -9860
rect 27020 -9990 27030 -9870
rect 27150 -9990 27160 -9870
rect 27020 -10000 27160 -9990
rect 26800 -10320 26940 -10310
rect 26800 -10440 26810 -10320
rect 26930 -10440 26940 -10320
rect 26800 -10450 26940 -10440
rect 26110 -11280 26120 -10600
rect 26230 -11280 26240 -10600
rect 26110 -11360 26240 -11280
rect 26100 -11370 26250 -11360
rect 26100 -11530 26110 -11370
rect 26240 -11530 26250 -11370
rect 26100 -11540 26250 -11530
rect 25420 -11670 25560 -11660
rect 25420 -11790 25430 -11670
rect 25550 -11790 25560 -11670
rect 25420 -11800 25560 -11790
rect 25200 -12120 25340 -12110
rect 25200 -12240 25210 -12120
rect 25330 -12240 25340 -12120
rect 25200 -12250 25340 -12240
rect 24510 -13080 24520 -12400
rect 24630 -13080 24640 -12400
rect 24510 -13160 24640 -13080
rect 24500 -13170 24650 -13160
rect 24500 -13330 24510 -13170
rect 24640 -13330 24650 -13170
rect 24500 -13340 24650 -13330
rect 23820 -13470 23960 -13460
rect 23820 -13590 23830 -13470
rect 23950 -13590 23960 -13470
rect 23820 -13600 23960 -13590
rect 23600 -13920 23740 -13910
rect 23600 -14040 23610 -13920
rect 23730 -14040 23740 -13920
rect 23600 -14050 23740 -14040
rect 22910 -14880 22920 -14200
rect 23030 -14880 23040 -14200
rect 22910 -14960 23040 -14880
rect 22900 -14970 23050 -14960
rect 22900 -15130 22910 -14970
rect 23040 -15130 23050 -14970
rect 22900 -15140 23050 -15130
rect 22220 -15270 22360 -15260
rect 22220 -15390 22230 -15270
rect 22350 -15390 22360 -15270
rect 22220 -15400 22360 -15390
rect 22000 -15720 22140 -15710
rect 22000 -15840 22010 -15720
rect 22130 -15840 22140 -15720
rect 22000 -15850 22140 -15840
rect 21310 -16680 21320 -16000
rect 21430 -16680 21440 -16000
rect 21310 -16760 21440 -16680
rect 21300 -16770 21450 -16760
rect 21300 -16930 21310 -16770
rect 21440 -16930 21450 -16770
rect 21300 -16940 21450 -16930
rect 20620 -17070 20760 -17060
rect 20620 -17190 20630 -17070
rect 20750 -17190 20760 -17070
rect 20620 -17200 20760 -17190
rect 20400 -17520 20540 -17510
rect 20400 -17640 20410 -17520
rect 20530 -17640 20540 -17520
rect 20400 -17650 20540 -17640
rect 19710 -18480 19720 -17800
rect 19830 -18480 19840 -17800
rect 19710 -18560 19840 -18480
rect 19700 -18570 19850 -18560
rect 19700 -18730 19710 -18570
rect 19840 -18730 19850 -18570
rect 19700 -18740 19850 -18730
rect 19020 -18870 19160 -18860
rect 19020 -18990 19030 -18870
rect 19150 -18990 19160 -18870
rect 19020 -19000 19160 -18990
rect 18800 -19320 18940 -19310
rect 18800 -19440 18810 -19320
rect 18930 -19440 18940 -19320
rect 18800 -19450 18940 -19440
rect 18110 -20280 18120 -19600
rect 18230 -20280 18240 -19600
rect 18110 -20360 18240 -20280
rect 18100 -20370 18250 -20360
rect 18100 -20530 18110 -20370
rect 18240 -20530 18250 -20370
rect 18100 -20540 18250 -20530
rect 17420 -20670 17560 -20660
rect 17420 -20790 17430 -20670
rect 17550 -20790 17560 -20670
rect 17420 -20800 17560 -20790
rect 17200 -21120 17340 -21110
rect 17200 -21240 17210 -21120
rect 17330 -21240 17340 -21120
rect 17200 -21250 17340 -21240
rect 17220 -21370 17320 -21250
rect 17440 -21370 17540 -20800
rect 16510 -22080 16520 -21400
rect 16630 -22080 16640 -21400
rect 16510 -22160 16640 -22080
rect 18110 -21400 18240 -20540
rect 18820 -21110 18920 -19450
rect 19040 -20660 19140 -19000
rect 19710 -19600 19840 -18740
rect 20420 -19310 20520 -17650
rect 20640 -18860 20740 -17200
rect 21310 -17800 21440 -16940
rect 22020 -17510 22120 -15850
rect 22240 -17060 22340 -15400
rect 22910 -16000 23040 -15140
rect 23620 -15710 23720 -14050
rect 23840 -15260 23940 -13600
rect 24510 -14200 24640 -13340
rect 25220 -13910 25320 -12250
rect 25440 -13460 25540 -11800
rect 26110 -12400 26240 -11540
rect 26820 -12110 26920 -10450
rect 27040 -11660 27140 -10000
rect 27710 -10600 27840 -9740
rect 28420 -10310 28520 -8650
rect 28640 -9860 28740 -8200
rect 30020 -8510 30120 -7760
rect 30240 -8060 30340 -6960
rect 30220 -8070 30360 -8060
rect 30220 -8190 30230 -8070
rect 30350 -8190 30360 -8070
rect 30220 -8200 30360 -8190
rect 30000 -8520 30140 -8510
rect 30000 -8640 30010 -8520
rect 30130 -8640 30140 -8520
rect 30000 -8650 30140 -8640
rect 29310 -8800 29440 -8790
rect 29310 -9480 29320 -8800
rect 29430 -9480 29440 -8800
rect 29310 -9560 29440 -9480
rect 29300 -9570 29450 -9560
rect 29300 -9730 29310 -9570
rect 29440 -9730 29450 -9570
rect 29300 -9740 29450 -9730
rect 28620 -9870 28760 -9860
rect 28620 -9990 28630 -9870
rect 28750 -9990 28760 -9870
rect 28620 -10000 28760 -9990
rect 28400 -10320 28540 -10310
rect 28400 -10440 28410 -10320
rect 28530 -10440 28540 -10320
rect 28400 -10450 28540 -10440
rect 27710 -11280 27720 -10600
rect 27830 -11280 27840 -10600
rect 27710 -11360 27840 -11280
rect 27700 -11370 27850 -11360
rect 27700 -11530 27710 -11370
rect 27840 -11530 27850 -11370
rect 27700 -11540 27850 -11530
rect 27020 -11670 27160 -11660
rect 27020 -11790 27030 -11670
rect 27150 -11790 27160 -11670
rect 27020 -11800 27160 -11790
rect 26800 -12120 26940 -12110
rect 26800 -12240 26810 -12120
rect 26930 -12240 26940 -12120
rect 26800 -12250 26940 -12240
rect 26110 -13080 26120 -12400
rect 26230 -13080 26240 -12400
rect 26110 -13160 26240 -13080
rect 26100 -13170 26250 -13160
rect 26100 -13330 26110 -13170
rect 26240 -13330 26250 -13170
rect 26100 -13340 26250 -13330
rect 25420 -13470 25560 -13460
rect 25420 -13590 25430 -13470
rect 25550 -13590 25560 -13470
rect 25420 -13600 25560 -13590
rect 25200 -13920 25340 -13910
rect 25200 -14040 25210 -13920
rect 25330 -14040 25340 -13920
rect 25200 -14050 25340 -14040
rect 24510 -14880 24520 -14200
rect 24630 -14880 24640 -14200
rect 24510 -14960 24640 -14880
rect 24500 -14970 24650 -14960
rect 24500 -15130 24510 -14970
rect 24640 -15130 24650 -14970
rect 24500 -15140 24650 -15130
rect 23820 -15270 23960 -15260
rect 23820 -15390 23830 -15270
rect 23950 -15390 23960 -15270
rect 23820 -15400 23960 -15390
rect 23600 -15720 23740 -15710
rect 23600 -15840 23610 -15720
rect 23730 -15840 23740 -15720
rect 23600 -15850 23740 -15840
rect 22910 -16680 22920 -16000
rect 23030 -16680 23040 -16000
rect 22910 -16760 23040 -16680
rect 22900 -16770 23050 -16760
rect 22900 -16930 22910 -16770
rect 23040 -16930 23050 -16770
rect 22900 -16940 23050 -16930
rect 22220 -17070 22360 -17060
rect 22220 -17190 22230 -17070
rect 22350 -17190 22360 -17070
rect 22220 -17200 22360 -17190
rect 22000 -17520 22140 -17510
rect 22000 -17640 22010 -17520
rect 22130 -17640 22140 -17520
rect 22000 -17650 22140 -17640
rect 21310 -18480 21320 -17800
rect 21430 -18480 21440 -17800
rect 21310 -18560 21440 -18480
rect 21300 -18570 21450 -18560
rect 21300 -18730 21310 -18570
rect 21440 -18730 21450 -18570
rect 21300 -18740 21450 -18730
rect 20620 -18870 20760 -18860
rect 20620 -18990 20630 -18870
rect 20750 -18990 20760 -18870
rect 20620 -19000 20760 -18990
rect 20400 -19320 20540 -19310
rect 20400 -19440 20410 -19320
rect 20530 -19440 20540 -19320
rect 20400 -19450 20540 -19440
rect 19710 -20280 19720 -19600
rect 19830 -20280 19840 -19600
rect 19710 -20360 19840 -20280
rect 19700 -20370 19850 -20360
rect 19700 -20530 19710 -20370
rect 19840 -20530 19850 -20370
rect 19700 -20540 19850 -20530
rect 19020 -20670 19160 -20660
rect 19020 -20790 19030 -20670
rect 19150 -20790 19160 -20670
rect 19020 -20800 19160 -20790
rect 18800 -21120 18940 -21110
rect 18800 -21240 18810 -21120
rect 18930 -21240 18940 -21120
rect 18800 -21250 18940 -21240
rect 18820 -21370 18920 -21250
rect 19040 -21370 19140 -20800
rect 18110 -22080 18120 -21400
rect 18230 -22080 18240 -21400
rect 18110 -22160 18240 -22080
rect 19710 -21400 19840 -20540
rect 20420 -21110 20520 -19450
rect 20640 -20660 20740 -19000
rect 21310 -19600 21440 -18740
rect 22020 -19310 22120 -17650
rect 22240 -18860 22340 -17200
rect 22910 -17800 23040 -16940
rect 23620 -17510 23720 -15850
rect 23840 -17060 23940 -15400
rect 24510 -16000 24640 -15140
rect 25220 -15220 25320 -14050
rect 25440 -15220 25540 -13600
rect 26110 -14200 26240 -13340
rect 26820 -13910 26920 -12250
rect 27040 -13460 27140 -11800
rect 27710 -12400 27840 -11540
rect 28420 -12110 28520 -10450
rect 28640 -11660 28740 -10000
rect 29310 -10600 29440 -9740
rect 30020 -10310 30120 -8650
rect 30240 -9860 30340 -8200
rect 30910 -8650 31040 -8030
rect 34820 -8060 34920 -8030
rect 31820 -8070 31960 -8060
rect 31820 -8190 31830 -8070
rect 31950 -8190 31960 -8070
rect 31820 -8200 31960 -8190
rect 34800 -8070 34940 -8060
rect 34800 -8190 34810 -8070
rect 34930 -8190 34940 -8070
rect 34800 -8200 34940 -8190
rect 30910 -8800 31040 -8790
rect 30910 -9480 30920 -8800
rect 31030 -9480 31040 -8800
rect 30910 -9560 31040 -9480
rect 30900 -9570 31050 -9560
rect 30900 -9730 30910 -9570
rect 31040 -9730 31050 -9570
rect 30900 -9740 31050 -9730
rect 30220 -9870 30360 -9860
rect 30220 -9990 30230 -9870
rect 30350 -9990 30360 -9870
rect 30220 -10000 30360 -9990
rect 30000 -10320 30140 -10310
rect 30000 -10440 30010 -10320
rect 30130 -10440 30140 -10320
rect 30000 -10450 30140 -10440
rect 29310 -11280 29320 -10600
rect 29430 -11280 29440 -10600
rect 29310 -11360 29440 -11280
rect 29300 -11370 29450 -11360
rect 29300 -11530 29310 -11370
rect 29440 -11530 29450 -11370
rect 29300 -11540 29450 -11530
rect 28620 -11670 28760 -11660
rect 28620 -11790 28630 -11670
rect 28750 -11790 28760 -11670
rect 28620 -11800 28760 -11790
rect 28400 -12120 28540 -12110
rect 28400 -12240 28410 -12120
rect 28530 -12240 28540 -12120
rect 28400 -12250 28540 -12240
rect 27710 -13080 27720 -12400
rect 27830 -13080 27840 -12400
rect 27710 -13160 27840 -13080
rect 27700 -13170 27850 -13160
rect 27700 -13330 27710 -13170
rect 27840 -13330 27850 -13170
rect 27700 -13340 27850 -13330
rect 27020 -13470 27160 -13460
rect 27020 -13590 27030 -13470
rect 27150 -13590 27160 -13470
rect 27020 -13600 27160 -13590
rect 26800 -13920 26940 -13910
rect 26800 -14040 26810 -13920
rect 26930 -14040 26940 -13920
rect 26800 -14050 26940 -14040
rect 26110 -14880 26120 -14200
rect 26230 -14880 26240 -14200
rect 26110 -14960 26240 -14880
rect 26100 -14970 26250 -14960
rect 26100 -15130 26110 -14970
rect 26240 -15130 26250 -14970
rect 26100 -15140 26250 -15130
rect 24510 -16680 24520 -16000
rect 24630 -16680 24640 -16000
rect 24510 -16760 24640 -16680
rect 26110 -16000 26240 -15140
rect 26820 -15710 26920 -14050
rect 27040 -15260 27140 -13600
rect 27710 -14200 27840 -13340
rect 28420 -13910 28520 -12250
rect 28640 -13460 28740 -11800
rect 29310 -12400 29440 -11540
rect 30020 -12110 30120 -10450
rect 30240 -11660 30340 -10000
rect 30910 -10600 31040 -9740
rect 31840 -9860 31940 -8200
rect 32510 -8800 32640 -8790
rect 32510 -9360 32520 -8800
rect 32630 -9360 32640 -8800
rect 32510 -9560 32640 -9360
rect 34110 -8800 34240 -8790
rect 34110 -9360 34120 -8800
rect 34230 -9360 34240 -8800
rect 33400 -9510 33540 -9500
rect 32500 -9570 32650 -9560
rect 32500 -9730 32510 -9570
rect 32640 -9730 32650 -9570
rect 33400 -9630 33410 -9510
rect 33530 -9630 33540 -9510
rect 34110 -9560 34240 -9360
rect 33400 -9640 33540 -9630
rect 32500 -9740 32650 -9730
rect 31820 -9870 31960 -9860
rect 31820 -9990 31830 -9870
rect 31950 -9990 31960 -9870
rect 31820 -10000 31960 -9990
rect 31600 -10320 31740 -10310
rect 31600 -10440 31610 -10320
rect 31730 -10440 31740 -10320
rect 31600 -10450 31740 -10440
rect 30910 -11280 30920 -10600
rect 31030 -11280 31040 -10600
rect 30910 -11360 31040 -11280
rect 30900 -11370 31050 -11360
rect 30900 -11530 30910 -11370
rect 31040 -11530 31050 -11370
rect 30900 -11540 31050 -11530
rect 30220 -11670 30360 -11660
rect 30220 -11790 30230 -11670
rect 30350 -11790 30360 -11670
rect 30220 -11800 30360 -11790
rect 30000 -12120 30140 -12110
rect 30000 -12240 30010 -12120
rect 30130 -12240 30140 -12120
rect 30000 -12250 30140 -12240
rect 29310 -13080 29320 -12400
rect 29430 -13080 29440 -12400
rect 29310 -13160 29440 -13080
rect 29300 -13170 29450 -13160
rect 29300 -13330 29310 -13170
rect 29440 -13330 29450 -13170
rect 29300 -13340 29450 -13330
rect 28620 -13470 28760 -13460
rect 28620 -13590 28630 -13470
rect 28750 -13590 28760 -13470
rect 28620 -13600 28760 -13590
rect 28400 -13920 28540 -13910
rect 28400 -14040 28410 -13920
rect 28530 -14040 28540 -13920
rect 28400 -14050 28540 -14040
rect 27710 -14880 27720 -14200
rect 27830 -14880 27840 -14200
rect 27710 -14960 27840 -14880
rect 27700 -14970 27850 -14960
rect 27700 -15130 27710 -14970
rect 27840 -15130 27850 -14970
rect 27700 -15140 27850 -15130
rect 27020 -15270 27160 -15260
rect 27020 -15390 27030 -15270
rect 27150 -15390 27160 -15270
rect 27020 -15400 27160 -15390
rect 26800 -15720 26940 -15710
rect 26800 -15840 26810 -15720
rect 26930 -15840 26940 -15720
rect 26800 -15850 26940 -15840
rect 26110 -16680 26120 -16000
rect 26230 -16680 26240 -16000
rect 26110 -16760 26240 -16680
rect 24500 -16770 24650 -16760
rect 24500 -16930 24510 -16770
rect 24640 -16930 24650 -16770
rect 24500 -16940 24650 -16930
rect 26100 -16770 26250 -16760
rect 26100 -16930 26110 -16770
rect 26240 -16930 26250 -16770
rect 26100 -16940 26250 -16930
rect 23820 -17070 23960 -17060
rect 23820 -17190 23830 -17070
rect 23950 -17190 23960 -17070
rect 23820 -17200 23960 -17190
rect 23600 -17520 23740 -17510
rect 23600 -17640 23610 -17520
rect 23730 -17640 23740 -17520
rect 23600 -17650 23740 -17640
rect 22910 -18480 22920 -17800
rect 23030 -18480 23040 -17800
rect 22910 -18560 23040 -18480
rect 22900 -18570 23050 -18560
rect 22900 -18730 22910 -18570
rect 23040 -18730 23050 -18570
rect 22900 -18740 23050 -18730
rect 22220 -18870 22360 -18860
rect 22220 -18990 22230 -18870
rect 22350 -18990 22360 -18870
rect 22220 -19000 22360 -18990
rect 22000 -19320 22140 -19310
rect 22000 -19440 22010 -19320
rect 22130 -19440 22140 -19320
rect 22000 -19450 22140 -19440
rect 21310 -20280 21320 -19600
rect 21430 -20280 21440 -19600
rect 21310 -20360 21440 -20280
rect 21300 -20370 21450 -20360
rect 21300 -20530 21310 -20370
rect 21440 -20530 21450 -20370
rect 21300 -20540 21450 -20530
rect 20620 -20670 20760 -20660
rect 20620 -20790 20630 -20670
rect 20750 -20790 20760 -20670
rect 20620 -20800 20760 -20790
rect 20400 -21120 20540 -21110
rect 20400 -21240 20410 -21120
rect 20530 -21240 20540 -21120
rect 20400 -21250 20540 -21240
rect 20420 -21370 20520 -21250
rect 20640 -21370 20740 -20800
rect 19710 -22080 19720 -21400
rect 19830 -22080 19840 -21400
rect 19710 -22160 19840 -22080
rect 21310 -21400 21440 -20540
rect 22020 -21110 22120 -19450
rect 22240 -20660 22340 -19000
rect 22910 -19600 23040 -18740
rect 23620 -19310 23720 -17650
rect 23840 -18860 23940 -17200
rect 24510 -17800 24640 -16940
rect 24510 -18480 24520 -17800
rect 24630 -18480 24640 -17800
rect 24510 -18560 24640 -18480
rect 26110 -17800 26240 -16940
rect 26820 -17510 26920 -15850
rect 27040 -17060 27140 -15400
rect 27710 -16000 27840 -15140
rect 28420 -15710 28520 -14050
rect 28640 -15260 28740 -13600
rect 29310 -14200 29440 -13340
rect 30020 -13910 30120 -12250
rect 30240 -13460 30340 -11800
rect 30910 -12400 31040 -11540
rect 31620 -12110 31720 -10450
rect 31840 -11660 31940 -10000
rect 32510 -10600 32640 -9740
rect 32510 -11110 32520 -10600
rect 32630 -11110 32640 -10600
rect 32510 -11360 32640 -11110
rect 32500 -11370 32650 -11360
rect 32500 -11530 32510 -11370
rect 32640 -11530 32650 -11370
rect 32500 -11540 32650 -11530
rect 31820 -11670 31960 -11660
rect 31820 -11790 31830 -11670
rect 31950 -11790 31960 -11670
rect 31820 -11800 31960 -11790
rect 31600 -12120 31740 -12110
rect 31600 -12240 31610 -12120
rect 31730 -12240 31740 -12120
rect 31600 -12250 31740 -12240
rect 30910 -13080 30920 -12400
rect 31030 -13080 31040 -12400
rect 30910 -13160 31040 -13080
rect 30900 -13170 31050 -13160
rect 30900 -13330 30910 -13170
rect 31040 -13330 31050 -13170
rect 30900 -13340 31050 -13330
rect 30220 -13470 30360 -13460
rect 30220 -13590 30230 -13470
rect 30350 -13590 30360 -13470
rect 30220 -13600 30360 -13590
rect 30000 -13920 30140 -13910
rect 30000 -14040 30010 -13920
rect 30130 -14040 30140 -13920
rect 30000 -14050 30140 -14040
rect 29310 -14880 29320 -14200
rect 29430 -14880 29440 -14200
rect 29310 -14960 29440 -14880
rect 29300 -14970 29450 -14960
rect 29300 -15130 29310 -14970
rect 29440 -15130 29450 -14970
rect 29300 -15140 29450 -15130
rect 28620 -15270 28760 -15260
rect 28620 -15390 28630 -15270
rect 28750 -15390 28760 -15270
rect 28620 -15400 28760 -15390
rect 28400 -15720 28540 -15710
rect 28400 -15840 28410 -15720
rect 28530 -15840 28540 -15720
rect 28400 -15850 28540 -15840
rect 27710 -16680 27720 -16000
rect 27830 -16680 27840 -16000
rect 27710 -16760 27840 -16680
rect 27700 -16770 27850 -16760
rect 27700 -16930 27710 -16770
rect 27840 -16930 27850 -16770
rect 27700 -16940 27850 -16930
rect 27020 -17070 27160 -17060
rect 27020 -17190 27030 -17070
rect 27150 -17190 27160 -17070
rect 27020 -17200 27160 -17190
rect 26800 -17520 26940 -17510
rect 26800 -17640 26810 -17520
rect 26930 -17640 26940 -17520
rect 26800 -17650 26940 -17640
rect 26110 -18480 26120 -17800
rect 26230 -18480 26240 -17800
rect 26110 -18560 26240 -18480
rect 24500 -18570 24650 -18560
rect 24500 -18730 24510 -18570
rect 24640 -18730 24650 -18570
rect 24500 -18740 24650 -18730
rect 26100 -18570 26250 -18560
rect 26100 -18730 26110 -18570
rect 26240 -18730 26250 -18570
rect 26100 -18740 26250 -18730
rect 23820 -18870 23960 -18860
rect 23820 -18990 23830 -18870
rect 23950 -18990 23960 -18870
rect 23820 -19000 23960 -18990
rect 23600 -19320 23740 -19310
rect 23600 -19440 23610 -19320
rect 23730 -19440 23740 -19320
rect 23600 -19450 23740 -19440
rect 22910 -20280 22920 -19600
rect 23030 -20280 23040 -19600
rect 22910 -20360 23040 -20280
rect 22900 -20370 23050 -20360
rect 22900 -20530 22910 -20370
rect 23040 -20530 23050 -20370
rect 22900 -20540 23050 -20530
rect 22220 -20670 22360 -20660
rect 22220 -20790 22230 -20670
rect 22350 -20790 22360 -20670
rect 22220 -20800 22360 -20790
rect 22000 -21120 22140 -21110
rect 22000 -21240 22010 -21120
rect 22130 -21240 22140 -21120
rect 22000 -21250 22140 -21240
rect 22020 -21370 22120 -21250
rect 22240 -21370 22340 -20800
rect 21310 -22080 21320 -21400
rect 21430 -22080 21440 -21400
rect 21310 -22160 21440 -22080
rect 22910 -21400 23040 -20540
rect 23620 -21110 23720 -19450
rect 23840 -20660 23940 -19000
rect 24510 -19600 24640 -18740
rect 24510 -20280 24520 -19600
rect 24630 -20280 24640 -19600
rect 24510 -20360 24640 -20280
rect 26110 -19600 26240 -18740
rect 26820 -19310 26920 -17650
rect 27040 -18860 27140 -17200
rect 27710 -17800 27840 -16940
rect 28420 -17510 28520 -15850
rect 28640 -17060 28740 -15400
rect 29310 -16000 29440 -15140
rect 29310 -16680 29320 -16000
rect 29430 -16680 29440 -16000
rect 29310 -16760 29440 -16680
rect 29300 -16770 29450 -16760
rect 29300 -16930 29310 -16770
rect 29440 -16930 29450 -16770
rect 29300 -16940 29450 -16930
rect 28620 -17070 28760 -17060
rect 28620 -17190 28630 -17070
rect 28750 -17190 28760 -17070
rect 28620 -17200 28760 -17190
rect 28400 -17520 28540 -17510
rect 28400 -17640 28410 -17520
rect 28530 -17640 28540 -17520
rect 28400 -17650 28540 -17640
rect 27710 -18480 27720 -17800
rect 27830 -18480 27840 -17800
rect 27710 -18560 27840 -18480
rect 27700 -18570 27850 -18560
rect 27700 -18730 27710 -18570
rect 27840 -18730 27850 -18570
rect 27700 -18740 27850 -18730
rect 27020 -18870 27160 -18860
rect 27020 -18990 27030 -18870
rect 27150 -18990 27160 -18870
rect 27020 -19000 27160 -18990
rect 26800 -19320 26940 -19310
rect 26800 -19440 26810 -19320
rect 26930 -19440 26940 -19320
rect 26800 -19450 26940 -19440
rect 26110 -20280 26120 -19600
rect 26230 -20280 26240 -19600
rect 26110 -20360 26240 -20280
rect 24500 -20370 24650 -20360
rect 24500 -20530 24510 -20370
rect 24640 -20530 24650 -20370
rect 24500 -20540 24650 -20530
rect 26100 -20370 26250 -20360
rect 26100 -20530 26110 -20370
rect 26240 -20530 26250 -20370
rect 26100 -20540 26250 -20530
rect 23820 -20670 23960 -20660
rect 23820 -20790 23830 -20670
rect 23950 -20790 23960 -20670
rect 23820 -20800 23960 -20790
rect 23600 -21120 23740 -21110
rect 23600 -21240 23610 -21120
rect 23730 -21240 23740 -21120
rect 23600 -21250 23740 -21240
rect 23620 -21370 23720 -21250
rect 23840 -21370 23940 -20800
rect 22910 -22080 22920 -21400
rect 23030 -22080 23040 -21400
rect 22910 -22160 23040 -22080
rect 24510 -21400 24640 -20540
rect 24510 -22080 24520 -21400
rect 24630 -22080 24640 -21400
rect 24510 -22160 24640 -22080
rect 26110 -21400 26240 -20540
rect 26820 -21110 26920 -19450
rect 27040 -20660 27140 -19000
rect 27710 -19600 27840 -18740
rect 28420 -19310 28520 -17650
rect 28640 -18860 28740 -17200
rect 29310 -17800 29440 -16940
rect 29310 -18480 29320 -17800
rect 29430 -18480 29440 -17800
rect 29310 -18560 29440 -18480
rect 29300 -18570 29450 -18560
rect 29300 -18730 29310 -18570
rect 29440 -18730 29450 -18570
rect 29300 -18740 29450 -18730
rect 28620 -18870 28760 -18860
rect 28620 -18990 28630 -18870
rect 28750 -18990 28760 -18870
rect 28620 -19000 28760 -18990
rect 28400 -19320 28540 -19310
rect 28400 -19440 28410 -19320
rect 28530 -19440 28540 -19320
rect 28400 -19450 28540 -19440
rect 27710 -20280 27720 -19600
rect 27830 -20280 27840 -19600
rect 27710 -20360 27840 -20280
rect 27700 -20370 27850 -20360
rect 27700 -20530 27710 -20370
rect 27840 -20530 27850 -20370
rect 27700 -20540 27850 -20530
rect 27020 -20670 27160 -20660
rect 27020 -20790 27030 -20670
rect 27150 -20790 27160 -20670
rect 27020 -20800 27160 -20790
rect 26800 -21120 26940 -21110
rect 26800 -21240 26810 -21120
rect 26930 -21240 26940 -21120
rect 26800 -21250 26940 -21240
rect 26820 -21370 26920 -21250
rect 27040 -21370 27140 -20800
rect 26110 -22080 26120 -21400
rect 26230 -22080 26240 -21400
rect 26110 -22160 26240 -22080
rect 27710 -21400 27840 -20540
rect 28420 -21110 28520 -19450
rect 28640 -20660 28740 -19000
rect 29310 -19600 29440 -18740
rect 29310 -20280 29320 -19600
rect 29430 -20280 29440 -19600
rect 29310 -20360 29440 -20280
rect 29300 -20370 29450 -20360
rect 29300 -20530 29310 -20370
rect 29440 -20530 29450 -20370
rect 29300 -20540 29450 -20530
rect 28620 -20670 28760 -20660
rect 28620 -20790 28630 -20670
rect 28750 -20790 28760 -20670
rect 28620 -20800 28760 -20790
rect 28400 -21120 28540 -21110
rect 28400 -21240 28410 -21120
rect 28530 -21240 28540 -21120
rect 28400 -21250 28540 -21240
rect 28420 -21370 28520 -21250
rect 28640 -21370 28740 -20800
rect 27710 -22080 27720 -21400
rect 27830 -22080 27840 -21400
rect 27710 -22160 27840 -22080
rect 29310 -21400 29440 -20540
rect 30020 -21370 30120 -14050
rect 30240 -21370 30340 -13600
rect 30910 -14200 31040 -13340
rect 31620 -13910 31720 -12250
rect 31840 -13460 31940 -11800
rect 32510 -12400 32640 -11540
rect 32510 -12910 32520 -12400
rect 32630 -12910 32640 -12400
rect 32510 -13160 32640 -12910
rect 32500 -13170 32650 -13160
rect 32500 -13330 32510 -13170
rect 32640 -13330 32650 -13170
rect 32500 -13340 32650 -13330
rect 31820 -13470 31960 -13460
rect 31820 -13590 31830 -13470
rect 31950 -13590 31960 -13470
rect 31820 -13600 31960 -13590
rect 31600 -13920 31740 -13910
rect 31600 -14040 31610 -13920
rect 31730 -14040 31740 -13920
rect 31600 -14050 31740 -14040
rect 30910 -14880 30920 -14200
rect 31030 -14880 31040 -14200
rect 30910 -14960 31040 -14880
rect 32510 -14200 32640 -13340
rect 32510 -14710 32520 -14200
rect 32630 -14710 32640 -14200
rect 32510 -14890 32640 -14710
rect 30900 -14970 31050 -14960
rect 30900 -15130 30910 -14970
rect 31040 -15130 31050 -14970
rect 30900 -15140 31050 -15130
rect 30910 -16000 31040 -15140
rect 31840 -15280 31980 -15270
rect 31840 -15400 31850 -15280
rect 31970 -15400 31980 -15280
rect 31840 -15410 31980 -15400
rect 31580 -15720 31720 -15710
rect 31580 -15840 31590 -15720
rect 31710 -15840 31720 -15720
rect 31580 -15850 31720 -15840
rect 30910 -16680 30920 -16000
rect 31030 -16680 31040 -16000
rect 30910 -16760 31040 -16680
rect 30900 -16770 31050 -16760
rect 30900 -16930 30910 -16770
rect 31040 -16930 31050 -16770
rect 30900 -16940 31050 -16930
rect 30910 -17800 31040 -16940
rect 31600 -17510 31700 -15850
rect 31860 -17070 31960 -15410
rect 32510 -16000 32640 -15990
rect 32510 -16680 32520 -16000
rect 32630 -16680 32640 -16000
rect 32510 -16770 32640 -16680
rect 32510 -16920 32520 -16770
rect 32630 -16920 32640 -16770
rect 31840 -17080 31980 -17070
rect 31840 -17200 31850 -17080
rect 31970 -17200 31980 -17080
rect 31840 -17210 31980 -17200
rect 31580 -17520 31720 -17510
rect 31580 -17640 31590 -17520
rect 31710 -17640 31720 -17520
rect 31580 -17650 31720 -17640
rect 30910 -18480 30920 -17800
rect 31030 -18480 31040 -17800
rect 30910 -18560 31040 -18480
rect 30900 -18570 31050 -18560
rect 30900 -18730 30910 -18570
rect 31040 -18730 31050 -18570
rect 30900 -18740 31050 -18730
rect 30910 -19600 31040 -18740
rect 31580 -18880 31720 -18870
rect 31580 -19000 31590 -18880
rect 31710 -19000 31720 -18880
rect 31580 -19010 31720 -19000
rect 30910 -20280 30920 -19600
rect 31030 -20280 31040 -19600
rect 30910 -20360 31040 -20280
rect 30900 -20370 31050 -20360
rect 30900 -20530 30910 -20370
rect 31040 -20530 31050 -20370
rect 30900 -20540 31050 -20530
rect 29310 -22080 29320 -21400
rect 29430 -22080 29440 -21400
rect 29310 -22160 29440 -22080
rect 30910 -21400 31040 -20540
rect 31600 -20670 31700 -19010
rect 31740 -19240 31820 -19230
rect 31740 -19520 31750 -19240
rect 31810 -19520 31820 -19240
rect 31740 -19530 31820 -19520
rect 31580 -20680 31720 -20670
rect 31580 -20800 31590 -20680
rect 31710 -20800 31720 -20680
rect 31580 -20810 31720 -20800
rect 30910 -22080 30920 -21400
rect 31030 -22080 31040 -21400
rect 30910 -22160 31040 -22080
rect 16500 -22170 16650 -22160
rect 16500 -22330 16510 -22170
rect 16640 -22330 16650 -22170
rect 16500 -22340 16650 -22330
rect 18100 -22170 18250 -22160
rect 18100 -22330 18110 -22170
rect 18240 -22330 18250 -22170
rect 18100 -22340 18250 -22330
rect 19700 -22170 19850 -22160
rect 19700 -22330 19710 -22170
rect 19840 -22330 19850 -22170
rect 19700 -22340 19850 -22330
rect 21300 -22170 21450 -22160
rect 21300 -22330 21310 -22170
rect 21440 -22330 21450 -22170
rect 21300 -22340 21450 -22330
rect 22900 -22170 23050 -22160
rect 22900 -22330 22910 -22170
rect 23040 -22330 23050 -22170
rect 22900 -22340 23050 -22330
rect 24500 -22170 24650 -22160
rect 24500 -22330 24510 -22170
rect 24640 -22330 24650 -22170
rect 24500 -22340 24650 -22330
rect 26100 -22170 26250 -22160
rect 26100 -22330 26110 -22170
rect 26240 -22330 26250 -22170
rect 26100 -22340 26250 -22330
rect 27700 -22170 27850 -22160
rect 27700 -22330 27710 -22170
rect 27840 -22330 27850 -22170
rect 27700 -22340 27850 -22330
rect 29300 -22170 29450 -22160
rect 29300 -22330 29310 -22170
rect 29440 -22330 29450 -22170
rect 29300 -22340 29450 -22330
rect 30900 -22170 31050 -22160
rect 30900 -22330 30910 -22170
rect 31040 -22330 31050 -22170
rect 30900 -22340 31050 -22330
rect 27710 -22740 27840 -22340
rect 27710 -22850 27720 -22740
rect 27830 -22850 27840 -22740
rect 27710 -22860 27840 -22850
rect 28140 -22730 28380 -22720
rect 28990 -22730 29230 -22720
rect 28140 -22870 28150 -22730
rect 28370 -22870 28380 -22730
rect 28140 -22880 28380 -22870
rect 28620 -22740 28750 -22730
rect 28620 -22870 28630 -22740
rect 28740 -22870 28750 -22740
rect 28620 -22880 28750 -22870
rect 28990 -22870 29000 -22730
rect 29220 -22870 29230 -22730
rect 29310 -22740 29440 -22340
rect 29310 -22850 29320 -22740
rect 29430 -22850 29440 -22740
rect 29310 -22860 29440 -22850
rect 30910 -22740 31040 -22340
rect 30910 -22850 30920 -22740
rect 31030 -22850 31040 -22740
rect 30910 -22860 31040 -22850
rect 28990 -22880 29230 -22870
rect 12410 -22980 12530 -22970
rect 12410 -23090 12420 -22980
rect 12520 -23090 12530 -22980
rect 12410 -23100 12530 -23090
rect 26520 -22980 26720 -22970
rect 26520 -23160 26530 -22980
rect 26710 -23160 26720 -22980
rect 1180 -23270 1360 -23260
rect 1180 -23450 1190 -23270
rect 1350 -23450 1360 -23270
rect 1180 -23460 1360 -23450
rect 2780 -23270 2960 -23260
rect 2780 -23450 2790 -23270
rect 2950 -23450 2960 -23270
rect 2780 -23460 2960 -23450
rect 4380 -23270 4560 -23260
rect 4380 -23450 4390 -23270
rect 4550 -23450 4560 -23270
rect 4380 -23460 4560 -23450
rect 5980 -23270 6160 -23260
rect 5980 -23450 5990 -23270
rect 6150 -23450 6160 -23270
rect 5980 -23460 6160 -23450
rect 7580 -23270 7760 -23260
rect 7580 -23450 7590 -23270
rect 7750 -23450 7760 -23270
rect 7580 -23460 7760 -23450
rect 9180 -23270 9360 -23260
rect 9180 -23450 9190 -23270
rect 9350 -23450 9360 -23270
rect 9180 -23460 9360 -23450
rect 23200 -23300 23400 -23290
rect 23200 -23480 23210 -23300
rect 23390 -23480 23400 -23300
rect 1620 -24070 1820 -24060
rect 1620 -24250 1630 -24070
rect 1810 -24250 1820 -24070
rect 1620 -24260 1820 -24250
rect 1280 -24470 1480 -24460
rect 1280 -24650 1290 -24470
rect 1470 -24650 1480 -24470
rect 1280 -24660 1480 -24650
rect 420 -26630 620 -26620
rect 420 -26710 430 -26630
rect 610 -26710 620 -26630
rect 420 -26720 620 -26710
rect 1420 -26860 1480 -24660
rect 1410 -26870 1490 -26860
rect 1410 -27020 1420 -26870
rect 1480 -27020 1490 -26870
rect 1410 -27030 1490 -27020
rect 420 -27430 620 -27420
rect 420 -27510 430 -27430
rect 610 -27510 620 -27430
rect 420 -27520 620 -27510
rect 420 -28230 620 -28220
rect 420 -28310 430 -28230
rect 610 -28310 620 -28230
rect 420 -28320 620 -28310
rect 420 -29030 620 -29020
rect 420 -29110 430 -29030
rect 610 -29110 620 -29030
rect 420 -29120 620 -29110
rect 1420 -29260 1480 -27030
rect 1620 -27660 1680 -24260
rect 2020 -25160 2080 -23820
rect 2240 -25160 2300 -23820
rect 2500 -25070 4020 -25060
rect 2500 -25130 2510 -25070
rect 4010 -25130 4020 -25070
rect 2500 -25140 4020 -25130
rect 4220 -25160 4280 -23820
rect 4440 -25160 4500 -23820
rect 4700 -25070 6220 -25060
rect 4700 -25130 4710 -25070
rect 6210 -25130 6220 -25070
rect 4700 -25140 6220 -25130
rect 6420 -25160 6480 -23820
rect 6640 -25160 6700 -23820
rect 6900 -25070 8420 -25060
rect 6900 -25130 6910 -25070
rect 8410 -25130 8420 -25070
rect 6900 -25140 8420 -25130
rect 8620 -25160 8680 -23820
rect 8840 -25160 8900 -23820
rect 9100 -25070 10620 -25060
rect 9100 -25130 9110 -25070
rect 10610 -25130 10620 -25070
rect 9100 -25140 10620 -25130
rect 10820 -25160 10880 -23820
rect 11040 -25160 11100 -23820
rect 11300 -25070 12820 -25060
rect 11300 -25130 11310 -25070
rect 12810 -25130 12820 -25070
rect 11300 -25140 12820 -25130
rect 13020 -25160 13080 -23820
rect 13240 -25160 13300 -23820
rect 13500 -25070 15020 -25060
rect 13500 -25130 13510 -25070
rect 15010 -25130 15020 -25070
rect 13500 -25140 15020 -25130
rect 15220 -25160 15280 -23820
rect 15440 -25160 15500 -23820
rect 15700 -25070 17220 -25060
rect 15700 -25130 15710 -25070
rect 17210 -25130 17220 -25070
rect 15700 -25140 17220 -25130
rect 17420 -25160 17480 -23820
rect 17640 -25160 17700 -23820
rect 17900 -25070 19420 -25060
rect 17900 -25130 17910 -25070
rect 19410 -25130 19420 -25070
rect 17900 -25140 19420 -25130
rect 19620 -25160 19680 -23820
rect 19840 -25160 19900 -23820
rect 20440 -24070 20640 -24060
rect 20440 -24250 20450 -24070
rect 20630 -24250 20640 -24070
rect 20440 -24260 20640 -24250
rect 20100 -24470 20300 -24460
rect 20100 -24650 20110 -24470
rect 20290 -24650 20300 -24470
rect 20100 -24660 20300 -24650
rect 2010 -25330 2090 -25160
rect 2230 -25260 2310 -25160
rect 2230 -25320 2240 -25260
rect 2300 -25320 2310 -25260
rect 2230 -25330 2310 -25320
rect 2020 -25960 2080 -25330
rect 2240 -25960 2300 -25330
rect 4210 -25350 4290 -25160
rect 4430 -25170 4510 -25160
rect 4430 -25230 4440 -25170
rect 4500 -25230 4510 -25170
rect 4430 -25280 4510 -25230
rect 4430 -25340 4440 -25280
rect 4500 -25340 4510 -25280
rect 4430 -25350 4510 -25340
rect 6410 -25280 6490 -25160
rect 6410 -25340 6420 -25280
rect 6480 -25340 6490 -25280
rect 6410 -25350 6490 -25340
rect 6630 -25170 6710 -25160
rect 6630 -25230 6640 -25170
rect 6700 -25230 6710 -25170
rect 6630 -25350 6710 -25230
rect 8610 -25170 8690 -25160
rect 8610 -25230 8620 -25170
rect 8680 -25230 8690 -25170
rect 8610 -25280 8690 -25230
rect 8610 -25340 8620 -25280
rect 8680 -25340 8690 -25280
rect 8610 -25350 8690 -25340
rect 8830 -25350 8910 -25160
rect 10810 -25170 10890 -25160
rect 10810 -25230 10820 -25170
rect 10880 -25230 10890 -25170
rect 10810 -25280 10890 -25230
rect 10810 -25340 10820 -25280
rect 10880 -25340 10890 -25280
rect 10810 -25350 10890 -25340
rect 11030 -25350 11110 -25160
rect 13010 -25170 13090 -25160
rect 13010 -25230 13020 -25170
rect 13080 -25230 13090 -25170
rect 13010 -25280 13090 -25230
rect 13010 -25340 13020 -25280
rect 13080 -25340 13090 -25280
rect 13010 -25350 13090 -25340
rect 13230 -25350 13310 -25160
rect 15210 -25170 15290 -25160
rect 15210 -25230 15220 -25170
rect 15280 -25230 15290 -25170
rect 15210 -25350 15290 -25230
rect 15430 -25280 15510 -25160
rect 15430 -25340 15440 -25280
rect 15500 -25340 15510 -25280
rect 15430 -25350 15510 -25340
rect 17410 -25350 17490 -25160
rect 17630 -25170 17710 -25160
rect 17630 -25230 17640 -25170
rect 17700 -25230 17710 -25170
rect 17630 -25280 17710 -25230
rect 17630 -25340 17640 -25280
rect 17700 -25340 17710 -25280
rect 17630 -25350 17710 -25340
rect 19610 -25350 19690 -25160
rect 19830 -25170 19910 -25160
rect 19830 -25230 19840 -25170
rect 19900 -25230 19910 -25170
rect 19830 -25350 19910 -25230
rect 2500 -25630 2700 -25550
rect 3160 -25630 3360 -25550
rect 3820 -25630 4020 -25550
rect 2500 -25700 2700 -25690
rect 2500 -25760 2510 -25700
rect 2690 -25760 2700 -25700
rect 2500 -25770 2700 -25760
rect 3160 -25700 3360 -25690
rect 3160 -25760 3170 -25700
rect 3350 -25760 3360 -25700
rect 3160 -25770 3360 -25760
rect 3820 -25700 4020 -25690
rect 3820 -25760 3830 -25700
rect 4010 -25760 4020 -25700
rect 3820 -25770 4020 -25760
rect 2500 -25870 4020 -25860
rect 2500 -25930 2510 -25870
rect 4010 -25930 4020 -25870
rect 2500 -25940 4020 -25930
rect 4220 -25960 4280 -25350
rect 4440 -25960 4500 -25350
rect 4700 -25630 4900 -25550
rect 5360 -25630 5560 -25550
rect 6020 -25630 6220 -25550
rect 4700 -25700 4900 -25690
rect 4700 -25760 4710 -25700
rect 4890 -25760 4900 -25700
rect 4700 -25770 4900 -25760
rect 5360 -25700 5560 -25690
rect 5360 -25760 5370 -25700
rect 5550 -25760 5560 -25700
rect 5360 -25770 5560 -25760
rect 6020 -25700 6220 -25690
rect 6020 -25760 6030 -25700
rect 6210 -25760 6220 -25700
rect 6020 -25770 6220 -25760
rect 4700 -25870 6220 -25860
rect 4700 -25930 4710 -25870
rect 6210 -25930 6220 -25870
rect 4700 -25940 6220 -25930
rect 6420 -25960 6480 -25350
rect 6640 -25960 6700 -25350
rect 6900 -25560 7100 -25550
rect 6900 -25620 6910 -25560
rect 7090 -25620 7100 -25560
rect 6900 -25630 7100 -25620
rect 7560 -25560 7760 -25550
rect 7560 -25620 7570 -25560
rect 7750 -25620 7760 -25560
rect 7560 -25630 7760 -25620
rect 8220 -25560 8420 -25550
rect 8220 -25620 8230 -25560
rect 8410 -25620 8420 -25560
rect 8220 -25630 8420 -25620
rect 6900 -25770 7100 -25690
rect 7560 -25770 7760 -25690
rect 8220 -25770 8420 -25690
rect 6900 -25870 8420 -25860
rect 6900 -25930 6910 -25870
rect 8410 -25930 8420 -25870
rect 6900 -25940 8420 -25930
rect 8620 -25960 8680 -25350
rect 8840 -25960 8900 -25350
rect 9100 -25560 9300 -25550
rect 9100 -25620 9110 -25560
rect 9290 -25620 9300 -25560
rect 9100 -25630 9300 -25620
rect 9760 -25560 9960 -25550
rect 9760 -25620 9770 -25560
rect 9950 -25620 9960 -25560
rect 9760 -25630 9960 -25620
rect 10420 -25560 10620 -25550
rect 10420 -25620 10430 -25560
rect 10610 -25620 10620 -25560
rect 10420 -25630 10620 -25620
rect 9100 -25770 9300 -25690
rect 9760 -25770 9960 -25690
rect 10420 -25770 10620 -25690
rect 9100 -25870 10620 -25860
rect 9100 -25930 9110 -25870
rect 10610 -25930 10620 -25870
rect 9100 -25940 10620 -25930
rect 10820 -25960 10880 -25350
rect 11040 -25960 11100 -25350
rect 11300 -25560 11500 -25550
rect 11300 -25620 11310 -25560
rect 11490 -25620 11500 -25560
rect 11300 -25630 11500 -25620
rect 11960 -25560 12160 -25550
rect 11960 -25620 11970 -25560
rect 12150 -25620 12160 -25560
rect 11960 -25630 12160 -25620
rect 12620 -25560 12820 -25550
rect 12620 -25620 12630 -25560
rect 12810 -25620 12820 -25560
rect 12620 -25630 12820 -25620
rect 11300 -25770 11500 -25690
rect 11960 -25770 12160 -25690
rect 12620 -25770 12820 -25690
rect 11300 -25870 12820 -25860
rect 11300 -25930 11310 -25870
rect 12810 -25930 12820 -25870
rect 11300 -25940 12820 -25930
rect 13020 -25960 13080 -25350
rect 13240 -25960 13300 -25350
rect 13500 -25560 13700 -25550
rect 13500 -25620 13510 -25560
rect 13690 -25620 13700 -25560
rect 13500 -25630 13700 -25620
rect 14160 -25560 14360 -25550
rect 14160 -25620 14170 -25560
rect 14350 -25620 14360 -25560
rect 14160 -25630 14360 -25620
rect 14820 -25560 15020 -25550
rect 14820 -25620 14830 -25560
rect 15010 -25620 15020 -25560
rect 14820 -25630 15020 -25620
rect 13500 -25770 13700 -25690
rect 14160 -25770 14360 -25690
rect 14820 -25770 15020 -25690
rect 13500 -25870 15020 -25860
rect 13500 -25930 13510 -25870
rect 15010 -25930 15020 -25870
rect 13500 -25940 15020 -25930
rect 15220 -25960 15280 -25350
rect 15440 -25960 15500 -25350
rect 15700 -25630 15900 -25550
rect 16360 -25630 16560 -25550
rect 17020 -25630 17220 -25550
rect 15700 -25700 15900 -25690
rect 15700 -25760 15710 -25700
rect 15890 -25760 15900 -25700
rect 15700 -25770 15900 -25760
rect 16360 -25700 16560 -25690
rect 16360 -25760 16370 -25700
rect 16550 -25760 16560 -25700
rect 16360 -25770 16560 -25760
rect 17020 -25700 17220 -25690
rect 17020 -25760 17030 -25700
rect 17210 -25760 17220 -25700
rect 17020 -25770 17220 -25760
rect 15700 -25870 17220 -25860
rect 15700 -25930 15710 -25870
rect 17210 -25930 17220 -25870
rect 15700 -25940 17220 -25930
rect 17420 -25960 17480 -25350
rect 17640 -25960 17700 -25350
rect 17900 -25630 18100 -25550
rect 18560 -25630 18760 -25550
rect 19220 -25630 19420 -25550
rect 17900 -25700 18100 -25690
rect 17900 -25760 17910 -25700
rect 18090 -25760 18100 -25700
rect 17900 -25770 18100 -25760
rect 18560 -25700 18760 -25690
rect 18560 -25760 18570 -25700
rect 18750 -25760 18760 -25700
rect 18560 -25770 18760 -25760
rect 19220 -25700 19420 -25690
rect 19220 -25760 19230 -25700
rect 19410 -25760 19420 -25700
rect 19220 -25770 19420 -25760
rect 17900 -25870 19420 -25860
rect 17900 -25930 17910 -25870
rect 19410 -25930 19420 -25870
rect 17900 -25940 19420 -25930
rect 19620 -25960 19680 -25350
rect 19840 -25960 19900 -25350
rect 2010 -26060 2090 -25960
rect 2010 -26120 2020 -26060
rect 2080 -26120 2090 -26060
rect 2010 -26130 2090 -26120
rect 2230 -26130 2310 -25960
rect 4210 -25970 4290 -25960
rect 4210 -26030 4220 -25970
rect 4280 -26030 4290 -25970
rect 4210 -26080 4290 -26030
rect 2020 -26760 2080 -26130
rect 2240 -26760 2300 -26130
rect 4210 -26140 4220 -26080
rect 4280 -26140 4290 -26080
rect 4210 -26150 4290 -26140
rect 4430 -26150 4510 -25960
rect 6410 -25970 6490 -25960
rect 6410 -26030 6420 -25970
rect 6480 -26030 6490 -25970
rect 6410 -26150 6490 -26030
rect 6630 -26080 6710 -25960
rect 6630 -26140 6640 -26080
rect 6700 -26140 6710 -26080
rect 6630 -26150 6710 -26140
rect 8610 -26150 8690 -25960
rect 8830 -25970 8910 -25960
rect 8830 -26030 8840 -25970
rect 8900 -26030 8910 -25970
rect 8830 -26080 8910 -26030
rect 8830 -26140 8840 -26080
rect 8900 -26140 8910 -26080
rect 8830 -26150 8910 -26140
rect 10810 -26150 10890 -25960
rect 11030 -25970 11110 -25960
rect 11030 -26030 11040 -25970
rect 11100 -26030 11110 -25970
rect 11030 -26080 11110 -26030
rect 11030 -26140 11040 -26080
rect 11100 -26140 11110 -26080
rect 11030 -26150 11110 -26140
rect 13010 -26150 13090 -25960
rect 13230 -25970 13310 -25960
rect 13230 -26030 13240 -25970
rect 13300 -26030 13310 -25970
rect 13230 -26080 13310 -26030
rect 13230 -26140 13240 -26080
rect 13300 -26140 13310 -26080
rect 13230 -26150 13310 -26140
rect 15210 -26080 15290 -25960
rect 15210 -26140 15220 -26080
rect 15280 -26140 15290 -26080
rect 15210 -26150 15290 -26140
rect 15430 -25970 15510 -25960
rect 15430 -26030 15440 -25970
rect 15500 -26030 15510 -25970
rect 15430 -26150 15510 -26030
rect 17410 -25970 17490 -25960
rect 17410 -26030 17420 -25970
rect 17480 -26030 17490 -25970
rect 17410 -26080 17490 -26030
rect 17410 -26140 17420 -26080
rect 17480 -26140 17490 -26080
rect 17410 -26150 17490 -26140
rect 17630 -26150 17710 -25960
rect 19610 -25970 19690 -25960
rect 19610 -26030 19620 -25970
rect 19680 -26030 19690 -25970
rect 19610 -26150 19690 -26030
rect 19830 -26150 19910 -25960
rect 2500 -26360 2700 -26350
rect 2500 -26420 2510 -26360
rect 2690 -26420 2700 -26360
rect 2500 -26430 2700 -26420
rect 3160 -26360 3360 -26350
rect 3160 -26420 3170 -26360
rect 3350 -26420 3360 -26360
rect 3160 -26430 3360 -26420
rect 3820 -26360 4020 -26350
rect 3820 -26420 3830 -26360
rect 4010 -26420 4020 -26360
rect 3820 -26430 4020 -26420
rect 2500 -26570 2700 -26490
rect 3160 -26570 3360 -26490
rect 3820 -26570 4020 -26490
rect 4220 -26760 4280 -26150
rect 4440 -26760 4500 -26150
rect 4700 -26360 4900 -26350
rect 4700 -26420 4710 -26360
rect 4890 -26420 4900 -26360
rect 4700 -26430 4900 -26420
rect 5360 -26360 5560 -26350
rect 5360 -26420 5370 -26360
rect 5550 -26420 5560 -26360
rect 5360 -26430 5560 -26420
rect 6020 -26360 6220 -26350
rect 6020 -26420 6030 -26360
rect 6210 -26420 6220 -26360
rect 6020 -26430 6220 -26420
rect 4700 -26570 4900 -26490
rect 5360 -26570 5560 -26490
rect 6020 -26570 6220 -26490
rect 4700 -26670 6220 -26660
rect 4700 -26730 4710 -26670
rect 6210 -26730 6220 -26670
rect 4700 -26740 6220 -26730
rect 6420 -26760 6480 -26150
rect 6640 -26760 6700 -26150
rect 6900 -26430 7100 -26350
rect 7560 -26430 7760 -26350
rect 8220 -26430 8420 -26350
rect 6900 -26500 7100 -26490
rect 6900 -26560 6910 -26500
rect 7090 -26560 7100 -26500
rect 6900 -26570 7100 -26560
rect 7560 -26500 7760 -26490
rect 7560 -26560 7570 -26500
rect 7750 -26560 7760 -26500
rect 7560 -26570 7760 -26560
rect 8220 -26500 8420 -26490
rect 8220 -26560 8230 -26500
rect 8410 -26560 8420 -26500
rect 8220 -26570 8420 -26560
rect 6900 -26670 8420 -26660
rect 6900 -26730 6910 -26670
rect 8410 -26730 8420 -26670
rect 6900 -26740 8420 -26730
rect 8620 -26760 8680 -26150
rect 8840 -26760 8900 -26150
rect 9100 -26430 9300 -26350
rect 9760 -26430 9960 -26350
rect 10420 -26430 10620 -26350
rect 9100 -26500 9300 -26490
rect 9100 -26560 9110 -26500
rect 9290 -26560 9300 -26500
rect 9100 -26570 9300 -26560
rect 9760 -26500 9960 -26490
rect 9760 -26560 9770 -26500
rect 9950 -26560 9960 -26500
rect 9760 -26570 9960 -26560
rect 10420 -26500 10620 -26490
rect 10420 -26560 10430 -26500
rect 10610 -26560 10620 -26500
rect 10420 -26570 10620 -26560
rect 9100 -26670 10620 -26660
rect 9100 -26730 9110 -26670
rect 10610 -26730 10620 -26670
rect 9100 -26740 10620 -26730
rect 10820 -26760 10880 -26150
rect 11040 -26760 11100 -26150
rect 11300 -26430 11500 -26350
rect 11960 -26430 12160 -26350
rect 12620 -26430 12820 -26350
rect 11300 -26500 11500 -26490
rect 11300 -26560 11310 -26500
rect 11490 -26560 11500 -26500
rect 11300 -26570 11500 -26560
rect 11960 -26500 12160 -26490
rect 11960 -26560 11970 -26500
rect 12150 -26560 12160 -26500
rect 11960 -26570 12160 -26560
rect 12620 -26500 12820 -26490
rect 12620 -26560 12630 -26500
rect 12810 -26560 12820 -26500
rect 12620 -26570 12820 -26560
rect 11300 -26670 12820 -26660
rect 11300 -26730 11310 -26670
rect 12810 -26730 12820 -26670
rect 11300 -26740 12820 -26730
rect 13020 -26760 13080 -26150
rect 13240 -26760 13300 -26150
rect 13500 -26430 13700 -26350
rect 14160 -26430 14360 -26350
rect 14820 -26430 15020 -26350
rect 13500 -26500 13700 -26490
rect 13500 -26560 13510 -26500
rect 13690 -26560 13700 -26500
rect 13500 -26570 13700 -26560
rect 14160 -26500 14360 -26490
rect 14160 -26560 14170 -26500
rect 14350 -26560 14360 -26500
rect 14160 -26570 14360 -26560
rect 14820 -26500 15020 -26490
rect 14820 -26560 14830 -26500
rect 15010 -26560 15020 -26500
rect 14820 -26570 15020 -26560
rect 13500 -26670 15020 -26660
rect 13500 -26730 13510 -26670
rect 15010 -26730 15020 -26670
rect 13500 -26740 15020 -26730
rect 15220 -26760 15280 -26150
rect 15440 -26760 15500 -26150
rect 15700 -26360 15900 -26350
rect 15700 -26420 15710 -26360
rect 15890 -26420 15900 -26360
rect 15700 -26430 15900 -26420
rect 16360 -26360 16560 -26350
rect 16360 -26420 16370 -26360
rect 16550 -26420 16560 -26360
rect 16360 -26430 16560 -26420
rect 17020 -26360 17220 -26350
rect 17020 -26420 17030 -26360
rect 17210 -26420 17220 -26360
rect 17020 -26430 17220 -26420
rect 15700 -26570 15900 -26490
rect 16360 -26570 16560 -26490
rect 17020 -26570 17220 -26490
rect 15700 -26670 17220 -26660
rect 15700 -26730 15710 -26670
rect 17210 -26730 17220 -26670
rect 15700 -26740 17220 -26730
rect 17420 -26760 17480 -26150
rect 17640 -26760 17700 -26150
rect 17900 -26360 18100 -26350
rect 17900 -26420 17910 -26360
rect 18090 -26420 18100 -26360
rect 17900 -26430 18100 -26420
rect 18560 -26360 18760 -26350
rect 18560 -26420 18570 -26360
rect 18750 -26420 18760 -26360
rect 18560 -26430 18760 -26420
rect 19220 -26360 19420 -26350
rect 19220 -26420 19230 -26360
rect 19410 -26420 19420 -26360
rect 19220 -26430 19420 -26420
rect 17900 -26570 18100 -26490
rect 18560 -26570 18760 -26490
rect 19220 -26570 19420 -26490
rect 19620 -26760 19680 -26150
rect 19840 -26760 19900 -26150
rect 2010 -26930 2090 -26760
rect 2230 -26930 2310 -26760
rect 2020 -27560 2080 -26930
rect 2240 -27560 2300 -26930
rect 4210 -26950 4290 -26760
rect 4430 -26880 4510 -26760
rect 4430 -26940 4440 -26880
rect 4500 -26940 4510 -26880
rect 4430 -26950 4510 -26940
rect 6410 -26880 6490 -26760
rect 6410 -26940 6420 -26880
rect 6480 -26940 6490 -26880
rect 6410 -26950 6490 -26940
rect 6630 -26770 6710 -26760
rect 6630 -26830 6640 -26770
rect 6700 -26830 6710 -26770
rect 6630 -26950 6710 -26830
rect 8610 -26770 8690 -26760
rect 8610 -26830 8620 -26770
rect 8680 -26830 8690 -26770
rect 8610 -26880 8690 -26830
rect 8610 -26940 8620 -26880
rect 8680 -26940 8690 -26880
rect 8610 -26950 8690 -26940
rect 8830 -26950 8910 -26760
rect 10810 -26770 10890 -26760
rect 10810 -26830 10820 -26770
rect 10880 -26830 10890 -26770
rect 10810 -26880 10890 -26830
rect 10810 -26940 10820 -26880
rect 10880 -26940 10890 -26880
rect 10810 -26950 10890 -26940
rect 11030 -26950 11110 -26760
rect 13010 -26770 13090 -26760
rect 13010 -26830 13020 -26770
rect 13080 -26830 13090 -26770
rect 13010 -26880 13090 -26830
rect 13010 -26940 13020 -26880
rect 13080 -26940 13090 -26880
rect 13010 -26950 13090 -26940
rect 13230 -26950 13310 -26760
rect 15210 -26770 15290 -26760
rect 15210 -26830 15220 -26770
rect 15280 -26830 15290 -26770
rect 15210 -26950 15290 -26830
rect 15430 -26880 15510 -26760
rect 15430 -26940 15440 -26880
rect 15500 -26940 15510 -26880
rect 15430 -26950 15510 -26940
rect 17410 -26950 17490 -26760
rect 17630 -26770 17710 -26760
rect 17630 -26830 17640 -26770
rect 17700 -26830 17710 -26770
rect 17630 -26950 17710 -26830
rect 19610 -26950 19690 -26760
rect 19830 -26950 19910 -26760
rect 20240 -26770 20300 -24660
rect 20230 -26780 20310 -26770
rect 20230 -26930 20240 -26780
rect 20300 -26930 20310 -26780
rect 20230 -26940 20310 -26930
rect 2500 -27230 2700 -27150
rect 3160 -27230 3360 -27150
rect 3820 -27230 4020 -27150
rect 2500 -27300 2700 -27290
rect 2500 -27360 2510 -27300
rect 2690 -27360 2700 -27300
rect 2500 -27370 2700 -27360
rect 3160 -27300 3360 -27290
rect 3160 -27360 3170 -27300
rect 3350 -27360 3360 -27300
rect 3160 -27370 3360 -27360
rect 3820 -27300 4020 -27290
rect 3820 -27360 3830 -27300
rect 4010 -27360 4020 -27300
rect 3820 -27370 4020 -27360
rect 4220 -27560 4280 -26950
rect 4440 -27560 4500 -26950
rect 4700 -27230 4900 -27150
rect 5360 -27230 5560 -27150
rect 6020 -27230 6220 -27150
rect 4700 -27300 4900 -27290
rect 4700 -27360 4710 -27300
rect 4890 -27360 4900 -27300
rect 4700 -27370 4900 -27360
rect 5360 -27300 5560 -27290
rect 5360 -27360 5370 -27300
rect 5550 -27360 5560 -27300
rect 5360 -27370 5560 -27360
rect 6020 -27300 6220 -27290
rect 6020 -27360 6030 -27300
rect 6210 -27360 6220 -27300
rect 6020 -27370 6220 -27360
rect 4700 -27470 6220 -27460
rect 4700 -27530 4710 -27470
rect 6210 -27530 6220 -27470
rect 4700 -27540 6220 -27530
rect 6420 -27560 6480 -26950
rect 6640 -27560 6700 -26950
rect 6900 -27160 7100 -27150
rect 6900 -27220 6910 -27160
rect 7090 -27220 7100 -27160
rect 6900 -27230 7100 -27220
rect 7560 -27160 7760 -27150
rect 7560 -27220 7570 -27160
rect 7750 -27220 7760 -27160
rect 7560 -27230 7760 -27220
rect 8220 -27160 8420 -27150
rect 8220 -27220 8230 -27160
rect 8410 -27220 8420 -27160
rect 8220 -27230 8420 -27220
rect 6900 -27370 7100 -27290
rect 7560 -27370 7760 -27290
rect 8220 -27370 8420 -27290
rect 6900 -27470 8420 -27460
rect 6900 -27530 6910 -27470
rect 8410 -27530 8420 -27470
rect 6900 -27540 8420 -27530
rect 8620 -27560 8680 -26950
rect 8840 -27560 8900 -26950
rect 9100 -27160 9300 -27150
rect 9100 -27220 9110 -27160
rect 9290 -27220 9300 -27160
rect 9100 -27230 9300 -27220
rect 9760 -27160 9960 -27150
rect 9760 -27220 9770 -27160
rect 9950 -27220 9960 -27160
rect 9760 -27230 9960 -27220
rect 10420 -27160 10620 -27150
rect 10420 -27220 10430 -27160
rect 10610 -27220 10620 -27160
rect 10420 -27230 10620 -27220
rect 9100 -27370 9300 -27290
rect 9760 -27370 9960 -27290
rect 10420 -27370 10620 -27290
rect 9100 -27470 10620 -27460
rect 9100 -27530 9110 -27470
rect 10610 -27530 10620 -27470
rect 9100 -27540 10620 -27530
rect 10820 -27560 10880 -26950
rect 11040 -27560 11100 -26950
rect 11300 -27160 11500 -27150
rect 11300 -27220 11310 -27160
rect 11490 -27220 11500 -27160
rect 11300 -27230 11500 -27220
rect 11960 -27160 12160 -27150
rect 11960 -27220 11970 -27160
rect 12150 -27220 12160 -27160
rect 11960 -27230 12160 -27220
rect 12620 -27160 12820 -27150
rect 12620 -27220 12630 -27160
rect 12810 -27220 12820 -27160
rect 12620 -27230 12820 -27220
rect 11300 -27370 11500 -27290
rect 11960 -27370 12160 -27290
rect 12620 -27370 12820 -27290
rect 11300 -27470 12820 -27460
rect 11300 -27530 11310 -27470
rect 12810 -27530 12820 -27470
rect 11300 -27540 12820 -27530
rect 13020 -27560 13080 -26950
rect 13240 -27560 13300 -26950
rect 13500 -27160 13700 -27150
rect 13500 -27220 13510 -27160
rect 13690 -27220 13700 -27160
rect 13500 -27230 13700 -27220
rect 14160 -27160 14360 -27150
rect 14160 -27220 14170 -27160
rect 14350 -27220 14360 -27160
rect 14160 -27230 14360 -27220
rect 14820 -27160 15020 -27150
rect 14820 -27220 14830 -27160
rect 15010 -27220 15020 -27160
rect 14820 -27230 15020 -27220
rect 13500 -27370 13700 -27290
rect 14160 -27370 14360 -27290
rect 14820 -27370 15020 -27290
rect 13500 -27470 15020 -27460
rect 13500 -27530 13510 -27470
rect 15010 -27530 15020 -27470
rect 13500 -27540 15020 -27530
rect 15220 -27560 15280 -26950
rect 15440 -27560 15500 -26950
rect 15700 -27230 15900 -27150
rect 16360 -27230 16560 -27150
rect 17020 -27230 17220 -27150
rect 15700 -27300 15900 -27290
rect 15700 -27360 15710 -27300
rect 15890 -27360 15900 -27300
rect 15700 -27370 15900 -27360
rect 16360 -27300 16560 -27290
rect 16360 -27360 16370 -27300
rect 16550 -27360 16560 -27300
rect 16360 -27370 16560 -27360
rect 17020 -27300 17220 -27290
rect 17020 -27360 17030 -27300
rect 17210 -27360 17220 -27300
rect 17020 -27370 17220 -27360
rect 15700 -27470 17220 -27460
rect 15700 -27530 15710 -27470
rect 17210 -27530 17220 -27470
rect 15700 -27540 17220 -27530
rect 17420 -27560 17480 -26950
rect 17640 -27560 17700 -26950
rect 17900 -27230 18100 -27150
rect 18560 -27230 18760 -27150
rect 19220 -27230 19420 -27150
rect 17900 -27300 18100 -27290
rect 17900 -27360 17910 -27300
rect 18090 -27360 18100 -27300
rect 17900 -27370 18100 -27360
rect 18560 -27300 18760 -27290
rect 18560 -27360 18570 -27300
rect 18750 -27360 18760 -27300
rect 18560 -27370 18760 -27360
rect 19220 -27300 19420 -27290
rect 19220 -27360 19230 -27300
rect 19410 -27360 19420 -27300
rect 19220 -27370 19420 -27360
rect 19620 -27560 19680 -26950
rect 19840 -27560 19900 -26950
rect 1610 -27670 1690 -27660
rect 1610 -27820 1620 -27670
rect 1680 -27820 1690 -27670
rect 2010 -27730 2090 -27560
rect 2230 -27730 2310 -27560
rect 4210 -27680 4290 -27560
rect 1610 -27830 1690 -27820
rect 1620 -28460 1680 -27830
rect 2020 -28360 2080 -27730
rect 2240 -28360 2300 -27730
rect 4210 -27740 4220 -27680
rect 4280 -27740 4290 -27680
rect 4210 -27750 4290 -27740
rect 4430 -27750 4510 -27560
rect 6410 -27570 6490 -27560
rect 6410 -27630 6420 -27570
rect 6480 -27630 6490 -27570
rect 6410 -27750 6490 -27630
rect 6630 -27680 6710 -27560
rect 6630 -27740 6640 -27680
rect 6700 -27740 6710 -27680
rect 6630 -27750 6710 -27740
rect 8610 -27750 8690 -27560
rect 8830 -27570 8910 -27560
rect 8830 -27630 8840 -27570
rect 8900 -27630 8910 -27570
rect 8830 -27680 8910 -27630
rect 8830 -27740 8840 -27680
rect 8900 -27740 8910 -27680
rect 8830 -27750 8910 -27740
rect 10810 -27750 10890 -27560
rect 11030 -27570 11110 -27560
rect 11030 -27630 11040 -27570
rect 11100 -27630 11110 -27570
rect 11030 -27680 11110 -27630
rect 11030 -27740 11040 -27680
rect 11100 -27740 11110 -27680
rect 11030 -27750 11110 -27740
rect 13010 -27750 13090 -27560
rect 13230 -27570 13310 -27560
rect 13230 -27630 13240 -27570
rect 13300 -27630 13310 -27570
rect 13230 -27680 13310 -27630
rect 13230 -27740 13240 -27680
rect 13300 -27740 13310 -27680
rect 13230 -27750 13310 -27740
rect 15210 -27680 15290 -27560
rect 15210 -27740 15220 -27680
rect 15280 -27740 15290 -27680
rect 15210 -27750 15290 -27740
rect 15430 -27570 15510 -27560
rect 15430 -27630 15440 -27570
rect 15500 -27630 15510 -27570
rect 15430 -27750 15510 -27630
rect 17410 -27570 17490 -27560
rect 17410 -27630 17420 -27570
rect 17480 -27630 17490 -27570
rect 17410 -27750 17490 -27630
rect 17630 -27750 17710 -27560
rect 19610 -27750 19690 -27560
rect 19830 -27750 19910 -27560
rect 2500 -27960 2700 -27950
rect 2500 -28020 2510 -27960
rect 2690 -28020 2700 -27960
rect 2500 -28030 2700 -28020
rect 3160 -27960 3360 -27950
rect 3160 -28020 3170 -27960
rect 3350 -28020 3360 -27960
rect 3160 -28030 3360 -28020
rect 3820 -27960 4020 -27950
rect 3820 -28020 3830 -27960
rect 4010 -28020 4020 -27960
rect 3820 -28030 4020 -28020
rect 2500 -28170 2700 -28090
rect 3160 -28170 3360 -28090
rect 3820 -28170 4020 -28090
rect 4220 -28360 4280 -27750
rect 4440 -28360 4500 -27750
rect 4700 -27960 4900 -27950
rect 4700 -28020 4710 -27960
rect 4890 -28020 4900 -27960
rect 4700 -28030 4900 -28020
rect 5360 -27960 5560 -27950
rect 5360 -28020 5370 -27960
rect 5550 -28020 5560 -27960
rect 5360 -28030 5560 -28020
rect 6020 -27960 6220 -27950
rect 6020 -28020 6030 -27960
rect 6210 -28020 6220 -27960
rect 6020 -28030 6220 -28020
rect 4700 -28170 4900 -28090
rect 5360 -28170 5560 -28090
rect 6020 -28170 6220 -28090
rect 4700 -28270 6220 -28260
rect 4700 -28330 4710 -28270
rect 6210 -28330 6220 -28270
rect 4700 -28340 6220 -28330
rect 6420 -28360 6480 -27750
rect 6640 -28360 6700 -27750
rect 6900 -28030 7100 -27950
rect 7560 -28030 7760 -27950
rect 8220 -28030 8420 -27950
rect 6900 -28100 7100 -28090
rect 6900 -28160 6910 -28100
rect 7090 -28160 7100 -28100
rect 6900 -28170 7100 -28160
rect 7560 -28100 7760 -28090
rect 7560 -28160 7570 -28100
rect 7750 -28160 7760 -28100
rect 7560 -28170 7760 -28160
rect 8220 -28100 8420 -28090
rect 8220 -28160 8230 -28100
rect 8410 -28160 8420 -28100
rect 8220 -28170 8420 -28160
rect 6900 -28270 8420 -28260
rect 6900 -28330 6910 -28270
rect 8410 -28330 8420 -28270
rect 6900 -28340 8420 -28330
rect 8620 -28360 8680 -27750
rect 8840 -28360 8900 -27750
rect 9100 -28030 9300 -27950
rect 9760 -28030 9960 -27950
rect 10420 -28030 10620 -27950
rect 9100 -28100 9300 -28090
rect 9100 -28160 9110 -28100
rect 9290 -28160 9300 -28100
rect 9100 -28170 9300 -28160
rect 9760 -28100 9960 -28090
rect 9760 -28160 9770 -28100
rect 9950 -28160 9960 -28100
rect 9760 -28170 9960 -28160
rect 10420 -28100 10620 -28090
rect 10420 -28160 10430 -28100
rect 10610 -28160 10620 -28100
rect 10420 -28170 10620 -28160
rect 9100 -28270 10620 -28260
rect 9100 -28330 9110 -28270
rect 10610 -28330 10620 -28270
rect 9100 -28340 10620 -28330
rect 10820 -28360 10880 -27750
rect 11040 -28360 11100 -27750
rect 11300 -28030 11500 -27950
rect 11960 -28030 12160 -27950
rect 12620 -28030 12820 -27950
rect 11300 -28100 11500 -28090
rect 11300 -28160 11310 -28100
rect 11490 -28160 11500 -28100
rect 11300 -28170 11500 -28160
rect 11960 -28100 12160 -28090
rect 11960 -28160 11970 -28100
rect 12150 -28160 12160 -28100
rect 11960 -28170 12160 -28160
rect 12620 -28100 12820 -28090
rect 12620 -28160 12630 -28100
rect 12810 -28160 12820 -28100
rect 12620 -28170 12820 -28160
rect 11300 -28270 12820 -28260
rect 11300 -28330 11310 -28270
rect 12810 -28330 12820 -28270
rect 11300 -28340 12820 -28330
rect 13020 -28360 13080 -27750
rect 13240 -28360 13300 -27750
rect 13500 -28030 13700 -27950
rect 14160 -28030 14360 -27950
rect 14820 -28030 15020 -27950
rect 13500 -28100 13700 -28090
rect 13500 -28160 13510 -28100
rect 13690 -28160 13700 -28100
rect 13500 -28170 13700 -28160
rect 14160 -28100 14360 -28090
rect 14160 -28160 14170 -28100
rect 14350 -28160 14360 -28100
rect 14160 -28170 14360 -28160
rect 14820 -28100 15020 -28090
rect 14820 -28160 14830 -28100
rect 15010 -28160 15020 -28100
rect 14820 -28170 15020 -28160
rect 13500 -28270 15020 -28260
rect 13500 -28330 13510 -28270
rect 15010 -28330 15020 -28270
rect 13500 -28340 15020 -28330
rect 15220 -28360 15280 -27750
rect 15440 -28360 15500 -27750
rect 15700 -27960 15900 -27950
rect 15700 -28020 15710 -27960
rect 15890 -28020 15900 -27960
rect 15700 -28030 15900 -28020
rect 16360 -27960 16560 -27950
rect 16360 -28020 16370 -27960
rect 16550 -28020 16560 -27960
rect 16360 -28030 16560 -28020
rect 17020 -27960 17220 -27950
rect 17020 -28020 17030 -27960
rect 17210 -28020 17220 -27960
rect 17020 -28030 17220 -28020
rect 15700 -28170 15900 -28090
rect 16360 -28170 16560 -28090
rect 17020 -28170 17220 -28090
rect 15700 -28270 17220 -28260
rect 15700 -28330 15710 -28270
rect 17210 -28330 17220 -28270
rect 15700 -28340 17220 -28330
rect 17420 -28360 17480 -27750
rect 17640 -28360 17700 -27750
rect 17900 -27960 18100 -27950
rect 17900 -28020 17910 -27960
rect 18090 -28020 18100 -27960
rect 17900 -28030 18100 -28020
rect 18560 -27960 18760 -27950
rect 18560 -28020 18570 -27960
rect 18750 -28020 18760 -27960
rect 18560 -28030 18760 -28020
rect 19220 -27960 19420 -27950
rect 19220 -28020 19230 -27960
rect 19410 -28020 19420 -27960
rect 19220 -28030 19420 -28020
rect 17900 -28170 18100 -28090
rect 18560 -28170 18760 -28090
rect 19220 -28170 19420 -28090
rect 19620 -28360 19680 -27750
rect 19840 -28360 19900 -27750
rect 1610 -28470 1690 -28460
rect 1610 -28620 1620 -28470
rect 1680 -28620 1690 -28470
rect 2010 -28530 2090 -28360
rect 2230 -28530 2310 -28360
rect 4210 -28480 4290 -28360
rect 1610 -28630 1690 -28620
rect 1410 -29270 1490 -29260
rect 1410 -29420 1420 -29270
rect 1480 -29420 1490 -29270
rect 1410 -29430 1490 -29420
rect 1620 -29430 1680 -28630
rect 2020 -29160 2080 -28530
rect 2240 -29160 2300 -28530
rect 4210 -28540 4220 -28480
rect 4280 -28540 4290 -28480
rect 4210 -28550 4290 -28540
rect 4430 -28550 4510 -28360
rect 6410 -28370 6490 -28360
rect 6410 -28430 6420 -28370
rect 6480 -28430 6490 -28370
rect 6410 -28550 6490 -28430
rect 6630 -28480 6710 -28360
rect 6630 -28540 6640 -28480
rect 6700 -28540 6710 -28480
rect 6630 -28550 6710 -28540
rect 8610 -28550 8690 -28360
rect 8830 -28370 8910 -28360
rect 8830 -28430 8840 -28370
rect 8900 -28430 8910 -28370
rect 8830 -28480 8910 -28430
rect 8830 -28540 8840 -28480
rect 8900 -28540 8910 -28480
rect 8830 -28550 8910 -28540
rect 10810 -28550 10890 -28360
rect 11030 -28370 11110 -28360
rect 11030 -28430 11040 -28370
rect 11100 -28430 11110 -28370
rect 11030 -28480 11110 -28430
rect 11030 -28540 11040 -28480
rect 11100 -28540 11110 -28480
rect 11030 -28550 11110 -28540
rect 13010 -28550 13090 -28360
rect 13230 -28370 13310 -28360
rect 13230 -28430 13240 -28370
rect 13300 -28430 13310 -28370
rect 13230 -28480 13310 -28430
rect 13230 -28540 13240 -28480
rect 13300 -28540 13310 -28480
rect 13230 -28550 13310 -28540
rect 15210 -28480 15290 -28360
rect 15210 -28540 15220 -28480
rect 15280 -28540 15290 -28480
rect 15210 -28550 15290 -28540
rect 15430 -28370 15510 -28360
rect 15430 -28430 15440 -28370
rect 15500 -28430 15510 -28370
rect 15430 -28550 15510 -28430
rect 17410 -28370 17490 -28360
rect 17410 -28430 17420 -28370
rect 17480 -28430 17490 -28370
rect 17410 -28550 17490 -28430
rect 17630 -28550 17710 -28360
rect 19610 -28550 19690 -28360
rect 19830 -28550 19910 -28360
rect 2500 -28760 2700 -28750
rect 2500 -28820 2510 -28760
rect 2690 -28820 2700 -28760
rect 2500 -28830 2700 -28820
rect 3160 -28760 3360 -28750
rect 3160 -28820 3170 -28760
rect 3350 -28820 3360 -28760
rect 3160 -28830 3360 -28820
rect 3820 -28760 4020 -28750
rect 3820 -28820 3830 -28760
rect 4010 -28820 4020 -28760
rect 3820 -28830 4020 -28820
rect 2500 -28970 2700 -28890
rect 3160 -28970 3360 -28890
rect 3820 -28970 4020 -28890
rect 4220 -29160 4280 -28550
rect 4440 -29160 4500 -28550
rect 4700 -28760 4900 -28750
rect 4700 -28820 4710 -28760
rect 4890 -28820 4900 -28760
rect 4700 -28830 4900 -28820
rect 5360 -28760 5560 -28750
rect 5360 -28820 5370 -28760
rect 5550 -28820 5560 -28760
rect 5360 -28830 5560 -28820
rect 6020 -28760 6220 -28750
rect 6020 -28820 6030 -28760
rect 6210 -28820 6220 -28760
rect 6020 -28830 6220 -28820
rect 4700 -28970 4900 -28890
rect 5360 -28970 5560 -28890
rect 6020 -28970 6220 -28890
rect 4700 -29070 6220 -29060
rect 4700 -29130 4710 -29070
rect 6210 -29130 6220 -29070
rect 4700 -29140 6220 -29130
rect 6420 -29160 6480 -28550
rect 6640 -29160 6700 -28550
rect 6900 -28830 7100 -28750
rect 7560 -28830 7760 -28750
rect 8220 -28830 8420 -28750
rect 6900 -28900 7100 -28890
rect 6900 -28960 6910 -28900
rect 7090 -28960 7100 -28900
rect 6900 -28970 7100 -28960
rect 7560 -28900 7760 -28890
rect 7560 -28960 7570 -28900
rect 7750 -28960 7760 -28900
rect 7560 -28970 7760 -28960
rect 8220 -28900 8420 -28890
rect 8220 -28960 8230 -28900
rect 8410 -28960 8420 -28900
rect 8220 -28970 8420 -28960
rect 6900 -29070 8420 -29060
rect 6900 -29130 6910 -29070
rect 8410 -29130 8420 -29070
rect 6900 -29140 8420 -29130
rect 8620 -29160 8680 -28550
rect 8840 -29160 8900 -28550
rect 9100 -28830 9300 -28750
rect 9760 -28830 9960 -28750
rect 10420 -28830 10620 -28750
rect 9100 -28900 9300 -28890
rect 9100 -28960 9110 -28900
rect 9290 -28960 9300 -28900
rect 9100 -28970 9300 -28960
rect 9760 -28900 9960 -28890
rect 9760 -28960 9770 -28900
rect 9950 -28960 9960 -28900
rect 9760 -28970 9960 -28960
rect 10420 -28900 10620 -28890
rect 10420 -28960 10430 -28900
rect 10610 -28960 10620 -28900
rect 10420 -28970 10620 -28960
rect 9100 -29070 10620 -29060
rect 9100 -29130 9110 -29070
rect 10610 -29130 10620 -29070
rect 9100 -29140 10620 -29130
rect 10820 -29160 10880 -28550
rect 11040 -29160 11100 -28550
rect 11300 -28830 11500 -28750
rect 11960 -28830 12160 -28750
rect 12620 -28830 12820 -28750
rect 11300 -28900 11500 -28890
rect 11300 -28960 11310 -28900
rect 11490 -28960 11500 -28900
rect 11300 -28970 11500 -28960
rect 11960 -28900 12160 -28890
rect 11960 -28960 11970 -28900
rect 12150 -28960 12160 -28900
rect 11960 -28970 12160 -28960
rect 12620 -28900 12820 -28890
rect 12620 -28960 12630 -28900
rect 12810 -28960 12820 -28900
rect 12620 -28970 12820 -28960
rect 11300 -29070 12820 -29060
rect 11300 -29130 11310 -29070
rect 12810 -29130 12820 -29070
rect 11300 -29140 12820 -29130
rect 13020 -29160 13080 -28550
rect 13240 -29160 13300 -28550
rect 13500 -28830 13700 -28750
rect 14160 -28830 14360 -28750
rect 14820 -28830 15020 -28750
rect 13500 -28900 13700 -28890
rect 13500 -28960 13510 -28900
rect 13690 -28960 13700 -28900
rect 13500 -28970 13700 -28960
rect 14160 -28900 14360 -28890
rect 14160 -28960 14170 -28900
rect 14350 -28960 14360 -28900
rect 14160 -28970 14360 -28960
rect 14820 -28900 15020 -28890
rect 14820 -28960 14830 -28900
rect 15010 -28960 15020 -28900
rect 14820 -28970 15020 -28960
rect 13500 -29070 15020 -29060
rect 13500 -29130 13510 -29070
rect 15010 -29130 15020 -29070
rect 13500 -29140 15020 -29130
rect 15220 -29160 15280 -28550
rect 15440 -29160 15500 -28550
rect 15700 -28760 15900 -28750
rect 15700 -28820 15710 -28760
rect 15890 -28820 15900 -28760
rect 15700 -28830 15900 -28820
rect 16360 -28760 16560 -28750
rect 16360 -28820 16370 -28760
rect 16550 -28820 16560 -28760
rect 16360 -28830 16560 -28820
rect 17020 -28760 17220 -28750
rect 17020 -28820 17030 -28760
rect 17210 -28820 17220 -28760
rect 17020 -28830 17220 -28820
rect 15700 -28970 15900 -28890
rect 16360 -28970 16560 -28890
rect 17020 -28970 17220 -28890
rect 15700 -29070 17220 -29060
rect 15700 -29130 15710 -29070
rect 17210 -29130 17220 -29070
rect 15700 -29140 17220 -29130
rect 17420 -29160 17480 -28550
rect 17640 -29160 17700 -28550
rect 17900 -28760 18100 -28750
rect 17900 -28820 17910 -28760
rect 18090 -28820 18100 -28760
rect 17900 -28830 18100 -28820
rect 18560 -28760 18760 -28750
rect 18560 -28820 18570 -28760
rect 18750 -28820 18760 -28760
rect 18560 -28830 18760 -28820
rect 19220 -28760 19420 -28750
rect 19220 -28820 19230 -28760
rect 19410 -28820 19420 -28760
rect 19220 -28830 19420 -28820
rect 17900 -28970 18100 -28890
rect 18560 -28970 18760 -28890
rect 19220 -28970 19420 -28890
rect 19620 -29160 19680 -28550
rect 19840 -29160 19900 -28550
rect 2010 -29330 2090 -29160
rect 2230 -29330 2310 -29160
rect 2020 -29960 2080 -29330
rect 2240 -29960 2300 -29330
rect 4210 -29350 4290 -29160
rect 4430 -29280 4510 -29160
rect 4430 -29340 4440 -29280
rect 4500 -29340 4510 -29280
rect 4430 -29350 4510 -29340
rect 6410 -29280 6490 -29160
rect 6410 -29340 6420 -29280
rect 6480 -29340 6490 -29280
rect 6410 -29350 6490 -29340
rect 6630 -29170 6710 -29160
rect 6630 -29230 6640 -29170
rect 6700 -29230 6710 -29170
rect 6630 -29350 6710 -29230
rect 8610 -29170 8690 -29160
rect 8610 -29230 8620 -29170
rect 8680 -29230 8690 -29170
rect 8610 -29280 8690 -29230
rect 8610 -29340 8620 -29280
rect 8680 -29340 8690 -29280
rect 8610 -29350 8690 -29340
rect 8830 -29350 8910 -29160
rect 10810 -29170 10890 -29160
rect 10810 -29230 10820 -29170
rect 10880 -29230 10890 -29170
rect 10810 -29280 10890 -29230
rect 10810 -29340 10820 -29280
rect 10880 -29340 10890 -29280
rect 10810 -29350 10890 -29340
rect 11030 -29350 11110 -29160
rect 13010 -29170 13090 -29160
rect 13010 -29230 13020 -29170
rect 13080 -29230 13090 -29170
rect 13010 -29280 13090 -29230
rect 13010 -29340 13020 -29280
rect 13080 -29340 13090 -29280
rect 13010 -29350 13090 -29340
rect 13230 -29350 13310 -29160
rect 15210 -29170 15290 -29160
rect 15210 -29230 15220 -29170
rect 15280 -29230 15290 -29170
rect 15210 -29350 15290 -29230
rect 15430 -29280 15510 -29160
rect 15430 -29340 15440 -29280
rect 15500 -29340 15510 -29280
rect 15430 -29350 15510 -29340
rect 17410 -29350 17490 -29160
rect 17630 -29170 17710 -29160
rect 17630 -29230 17640 -29170
rect 17700 -29230 17710 -29170
rect 17630 -29350 17710 -29230
rect 19610 -29350 19690 -29160
rect 19830 -29350 19910 -29160
rect 20240 -29170 20300 -26940
rect 20440 -27570 20500 -24260
rect 23200 -24680 23400 -23480
rect 23030 -24690 23570 -24680
rect 23030 -25070 23040 -24690
rect 23560 -25070 23570 -24690
rect 23030 -25080 23570 -25070
rect 26520 -25500 26720 -23160
rect 31600 -23290 31700 -20810
rect 31750 -21030 31810 -19530
rect 31740 -21040 31820 -21030
rect 31740 -21320 31750 -21040
rect 31810 -21320 31820 -21040
rect 31740 -21330 31820 -21320
rect 31550 -23300 31750 -23290
rect 31550 -23480 31560 -23300
rect 31740 -23480 31750 -23300
rect 31550 -23490 31750 -23480
rect 29740 -23520 29890 -23510
rect 29740 -23590 29750 -23520
rect 29880 -23590 29890 -23520
rect 29740 -23600 29890 -23590
rect 28490 -24040 28670 -24030
rect 27620 -24070 27820 -24060
rect 27620 -24250 27630 -24070
rect 27810 -24250 27820 -24070
rect 28490 -24200 28500 -24040
rect 28660 -24050 28670 -24040
rect 28660 -24110 29740 -24050
rect 28660 -24200 28670 -24110
rect 28490 -24210 28670 -24200
rect 27620 -24260 27820 -24250
rect 27390 -24470 27590 -24460
rect 27390 -24650 27400 -24470
rect 27580 -24650 27590 -24470
rect 27390 -24660 27590 -24650
rect 27240 -24890 27440 -24880
rect 27240 -25070 27250 -24890
rect 27430 -25070 27440 -24890
rect 27240 -25080 27440 -25070
rect 26520 -25510 27330 -25500
rect 26520 -25600 27260 -25510
rect 27320 -25600 27330 -25510
rect 26520 -25610 27330 -25600
rect 26520 -25630 27320 -25610
rect 21300 -26630 21500 -26620
rect 21300 -26710 21310 -26630
rect 21490 -26710 21500 -26630
rect 21300 -26720 21500 -26710
rect 21300 -27430 21500 -27420
rect 21300 -27510 21310 -27430
rect 21490 -27510 21500 -27430
rect 21300 -27520 21500 -27510
rect 20430 -27580 20510 -27570
rect 20430 -27730 20440 -27580
rect 20500 -27730 20510 -27580
rect 20430 -27740 20510 -27730
rect 20440 -28370 20500 -27740
rect 21300 -28230 21500 -28220
rect 21300 -28310 21310 -28230
rect 21490 -28310 21500 -28230
rect 21300 -28320 21500 -28310
rect 20430 -28380 20510 -28370
rect 20430 -28530 20440 -28380
rect 20500 -28530 20510 -28380
rect 20430 -28540 20510 -28530
rect 20230 -29180 20310 -29170
rect 20230 -29330 20240 -29180
rect 20300 -29330 20310 -29180
rect 20230 -29340 20310 -29330
rect 20440 -29340 20500 -28540
rect 21300 -29030 21500 -29020
rect 21300 -29110 21310 -29030
rect 21490 -29110 21500 -29030
rect 21300 -29120 21500 -29110
rect 2500 -29630 2700 -29550
rect 3160 -29630 3360 -29550
rect 3820 -29630 4020 -29550
rect 2500 -29700 2700 -29690
rect 2500 -29760 2510 -29700
rect 2690 -29760 2700 -29700
rect 2500 -29770 2700 -29760
rect 3160 -29700 3360 -29690
rect 3160 -29760 3170 -29700
rect 3350 -29760 3360 -29700
rect 3160 -29770 3360 -29760
rect 3820 -29700 4020 -29690
rect 3820 -29760 3830 -29700
rect 4010 -29760 4020 -29700
rect 3820 -29770 4020 -29760
rect 2500 -29870 4020 -29860
rect 2500 -29930 2510 -29870
rect 4010 -29930 4020 -29870
rect 2500 -29940 4020 -29930
rect 4220 -29960 4280 -29350
rect 4440 -29960 4500 -29350
rect 4700 -29630 4900 -29550
rect 5360 -29630 5560 -29550
rect 6020 -29630 6220 -29550
rect 4700 -29700 4900 -29690
rect 4700 -29760 4710 -29700
rect 4890 -29760 4900 -29700
rect 4700 -29770 4900 -29760
rect 5360 -29700 5560 -29690
rect 5360 -29760 5370 -29700
rect 5550 -29760 5560 -29700
rect 5360 -29770 5560 -29760
rect 6020 -29700 6220 -29690
rect 6020 -29760 6030 -29700
rect 6210 -29760 6220 -29700
rect 6020 -29770 6220 -29760
rect 4700 -29870 6220 -29860
rect 4700 -29930 4710 -29870
rect 6210 -29930 6220 -29870
rect 4700 -29940 6220 -29930
rect 6420 -29960 6480 -29350
rect 6640 -29960 6700 -29350
rect 6900 -29560 7100 -29550
rect 6900 -29620 6910 -29560
rect 7090 -29620 7100 -29560
rect 6900 -29630 7100 -29620
rect 7560 -29560 7760 -29550
rect 7560 -29620 7570 -29560
rect 7750 -29620 7760 -29560
rect 7560 -29630 7760 -29620
rect 8220 -29560 8420 -29550
rect 8220 -29620 8230 -29560
rect 8410 -29620 8420 -29560
rect 8220 -29630 8420 -29620
rect 6900 -29770 7100 -29690
rect 7560 -29770 7760 -29690
rect 8220 -29770 8420 -29690
rect 6900 -29870 8420 -29860
rect 6900 -29930 6910 -29870
rect 8410 -29930 8420 -29870
rect 6900 -29940 8420 -29930
rect 8620 -29960 8680 -29350
rect 8840 -29960 8900 -29350
rect 9100 -29560 9300 -29550
rect 9100 -29620 9110 -29560
rect 9290 -29620 9300 -29560
rect 9100 -29630 9300 -29620
rect 9760 -29560 9960 -29550
rect 9760 -29620 9770 -29560
rect 9950 -29620 9960 -29560
rect 9760 -29630 9960 -29620
rect 10420 -29560 10620 -29550
rect 10420 -29620 10430 -29560
rect 10610 -29620 10620 -29560
rect 10420 -29630 10620 -29620
rect 9100 -29770 9300 -29690
rect 9760 -29770 9960 -29690
rect 10420 -29770 10620 -29690
rect 9100 -29870 10620 -29860
rect 9100 -29930 9110 -29870
rect 10610 -29930 10620 -29870
rect 9100 -29940 10620 -29930
rect 10820 -29960 10880 -29350
rect 11040 -29960 11100 -29350
rect 11300 -29560 11500 -29550
rect 11300 -29620 11310 -29560
rect 11490 -29620 11500 -29560
rect 11300 -29630 11500 -29620
rect 11960 -29560 12160 -29550
rect 11960 -29620 11970 -29560
rect 12150 -29620 12160 -29560
rect 11960 -29630 12160 -29620
rect 12620 -29560 12820 -29550
rect 12620 -29620 12630 -29560
rect 12810 -29620 12820 -29560
rect 12620 -29630 12820 -29620
rect 11300 -29770 11500 -29690
rect 11960 -29770 12160 -29690
rect 12620 -29770 12820 -29690
rect 11300 -29870 12820 -29860
rect 11300 -29930 11310 -29870
rect 12810 -29930 12820 -29870
rect 11300 -29940 12820 -29930
rect 13020 -29960 13080 -29350
rect 13240 -29960 13300 -29350
rect 13500 -29560 13700 -29550
rect 13500 -29620 13510 -29560
rect 13690 -29620 13700 -29560
rect 13500 -29630 13700 -29620
rect 14160 -29560 14360 -29550
rect 14160 -29620 14170 -29560
rect 14350 -29620 14360 -29560
rect 14160 -29630 14360 -29620
rect 14820 -29560 15020 -29550
rect 14820 -29620 14830 -29560
rect 15010 -29620 15020 -29560
rect 14820 -29630 15020 -29620
rect 13500 -29770 13700 -29690
rect 14160 -29770 14360 -29690
rect 14820 -29770 15020 -29690
rect 13500 -29870 15020 -29860
rect 13500 -29930 13510 -29870
rect 15010 -29930 15020 -29870
rect 13500 -29940 15020 -29930
rect 15220 -29960 15280 -29350
rect 15440 -29960 15500 -29350
rect 15700 -29630 15900 -29550
rect 16360 -29630 16560 -29550
rect 17020 -29630 17220 -29550
rect 15700 -29700 15900 -29690
rect 15700 -29760 15710 -29700
rect 15890 -29760 15900 -29700
rect 15700 -29770 15900 -29760
rect 16360 -29700 16560 -29690
rect 16360 -29760 16370 -29700
rect 16550 -29760 16560 -29700
rect 16360 -29770 16560 -29760
rect 17020 -29700 17220 -29690
rect 17020 -29760 17030 -29700
rect 17210 -29760 17220 -29700
rect 17020 -29770 17220 -29760
rect 15700 -29870 17220 -29860
rect 15700 -29930 15710 -29870
rect 17210 -29930 17220 -29870
rect 15700 -29940 17220 -29930
rect 17420 -29960 17480 -29350
rect 17640 -29960 17700 -29350
rect 17900 -29630 18100 -29550
rect 18560 -29630 18760 -29550
rect 19220 -29630 19420 -29550
rect 17900 -29700 18100 -29690
rect 17900 -29760 17910 -29700
rect 18090 -29760 18100 -29700
rect 17900 -29770 18100 -29760
rect 18560 -29700 18760 -29690
rect 18560 -29760 18570 -29700
rect 18750 -29760 18760 -29700
rect 18560 -29770 18760 -29760
rect 19220 -29700 19420 -29690
rect 19220 -29760 19230 -29700
rect 19410 -29760 19420 -29700
rect 19220 -29770 19420 -29760
rect 17900 -29870 19420 -29860
rect 17900 -29930 17910 -29870
rect 19410 -29930 19420 -29870
rect 17900 -29940 19420 -29930
rect 19620 -29960 19680 -29350
rect 19840 -29960 19900 -29350
rect 2010 -30060 2090 -29960
rect 2010 -30120 2020 -30060
rect 2080 -30120 2090 -30060
rect 2010 -30130 2090 -30120
rect 2230 -30130 2310 -29960
rect 4210 -29970 4290 -29960
rect 4210 -30030 4220 -29970
rect 4280 -30030 4290 -29970
rect 4210 -30080 4290 -30030
rect 2020 -30760 2080 -30130
rect 2240 -30760 2300 -30130
rect 4210 -30140 4220 -30080
rect 4280 -30140 4290 -30080
rect 4210 -30150 4290 -30140
rect 4430 -30150 4510 -29960
rect 6410 -29970 6490 -29960
rect 6410 -30030 6420 -29970
rect 6480 -30030 6490 -29970
rect 6410 -30150 6490 -30030
rect 6630 -30080 6710 -29960
rect 6630 -30140 6640 -30080
rect 6700 -30140 6710 -30080
rect 6630 -30150 6710 -30140
rect 8610 -30150 8690 -29960
rect 8830 -29970 8910 -29960
rect 8830 -30030 8840 -29970
rect 8900 -30030 8910 -29970
rect 8830 -30080 8910 -30030
rect 8830 -30140 8840 -30080
rect 8900 -30140 8910 -30080
rect 8830 -30150 8910 -30140
rect 10810 -30150 10890 -29960
rect 11030 -29970 11110 -29960
rect 11030 -30030 11040 -29970
rect 11100 -30030 11110 -29970
rect 11030 -30080 11110 -30030
rect 11030 -30140 11040 -30080
rect 11100 -30140 11110 -30080
rect 11030 -30150 11110 -30140
rect 13010 -30150 13090 -29960
rect 13230 -29970 13310 -29960
rect 13230 -30030 13240 -29970
rect 13300 -30030 13310 -29970
rect 13230 -30080 13310 -30030
rect 13230 -30140 13240 -30080
rect 13300 -30140 13310 -30080
rect 13230 -30150 13310 -30140
rect 15210 -30080 15290 -29960
rect 15210 -30140 15220 -30080
rect 15280 -30140 15290 -30080
rect 15210 -30150 15290 -30140
rect 15430 -29970 15510 -29960
rect 15430 -30030 15440 -29970
rect 15500 -30030 15510 -29970
rect 15430 -30150 15510 -30030
rect 17410 -29970 17490 -29960
rect 17410 -30030 17420 -29970
rect 17480 -30030 17490 -29970
rect 17410 -30080 17490 -30030
rect 17410 -30140 17420 -30080
rect 17480 -30140 17490 -30080
rect 17410 -30150 17490 -30140
rect 17630 -30150 17710 -29960
rect 19610 -29970 19690 -29960
rect 19610 -30030 19620 -29970
rect 19680 -30030 19690 -29970
rect 19610 -30150 19690 -30030
rect 19830 -30150 19910 -29960
rect 2500 -30360 2700 -30350
rect 2500 -30420 2510 -30360
rect 2690 -30420 2700 -30360
rect 2500 -30430 2700 -30420
rect 3160 -30360 3360 -30350
rect 3160 -30420 3170 -30360
rect 3350 -30420 3360 -30360
rect 3160 -30430 3360 -30420
rect 3820 -30360 4020 -30350
rect 3820 -30420 3830 -30360
rect 4010 -30420 4020 -30360
rect 3820 -30430 4020 -30420
rect 2500 -30570 2700 -30490
rect 3160 -30570 3360 -30490
rect 3820 -30570 4020 -30490
rect 2500 -30670 4020 -30660
rect 2500 -30730 2510 -30670
rect 4010 -30730 4020 -30670
rect 2500 -30740 4020 -30730
rect 4220 -30760 4280 -30150
rect 4440 -30760 4500 -30150
rect 4700 -30360 4900 -30350
rect 4700 -30420 4710 -30360
rect 4890 -30420 4900 -30360
rect 4700 -30430 4900 -30420
rect 5360 -30360 5560 -30350
rect 5360 -30420 5370 -30360
rect 5550 -30420 5560 -30360
rect 5360 -30430 5560 -30420
rect 6020 -30360 6220 -30350
rect 6020 -30420 6030 -30360
rect 6210 -30420 6220 -30360
rect 6020 -30430 6220 -30420
rect 4700 -30570 4900 -30490
rect 5360 -30570 5560 -30490
rect 6020 -30570 6220 -30490
rect 4700 -30670 6220 -30660
rect 4700 -30730 4710 -30670
rect 6210 -30730 6220 -30670
rect 4700 -30740 6220 -30730
rect 6420 -30760 6480 -30150
rect 6640 -30760 6700 -30150
rect 6900 -30430 7100 -30350
rect 7560 -30430 7760 -30350
rect 8220 -30430 8420 -30350
rect 6900 -30500 7100 -30490
rect 6900 -30560 6910 -30500
rect 7090 -30560 7100 -30500
rect 6900 -30570 7100 -30560
rect 7560 -30500 7760 -30490
rect 7560 -30560 7570 -30500
rect 7750 -30560 7760 -30500
rect 7560 -30570 7760 -30560
rect 8220 -30500 8420 -30490
rect 8220 -30560 8230 -30500
rect 8410 -30560 8420 -30500
rect 8220 -30570 8420 -30560
rect 6900 -30670 8420 -30660
rect 6900 -30730 6910 -30670
rect 8410 -30730 8420 -30670
rect 6900 -30740 8420 -30730
rect 8620 -30760 8680 -30150
rect 8840 -30760 8900 -30150
rect 9100 -30430 9300 -30350
rect 9760 -30430 9960 -30350
rect 10420 -30430 10620 -30350
rect 9100 -30500 9300 -30490
rect 9100 -30560 9110 -30500
rect 9290 -30560 9300 -30500
rect 9100 -30570 9300 -30560
rect 9760 -30500 9960 -30490
rect 9760 -30560 9770 -30500
rect 9950 -30560 9960 -30500
rect 9760 -30570 9960 -30560
rect 10420 -30500 10620 -30490
rect 10420 -30560 10430 -30500
rect 10610 -30560 10620 -30500
rect 10420 -30570 10620 -30560
rect 9100 -30670 10620 -30660
rect 9100 -30730 9110 -30670
rect 10610 -30730 10620 -30670
rect 9100 -30740 10620 -30730
rect 10820 -30760 10880 -30150
rect 11040 -30760 11100 -30150
rect 11300 -30430 11500 -30350
rect 11960 -30430 12160 -30350
rect 12620 -30430 12820 -30350
rect 11300 -30500 11500 -30490
rect 11300 -30560 11310 -30500
rect 11490 -30560 11500 -30500
rect 11300 -30570 11500 -30560
rect 11960 -30500 12160 -30490
rect 11960 -30560 11970 -30500
rect 12150 -30560 12160 -30500
rect 11960 -30570 12160 -30560
rect 12620 -30500 12820 -30490
rect 12620 -30560 12630 -30500
rect 12810 -30560 12820 -30500
rect 12620 -30570 12820 -30560
rect 11300 -30670 12820 -30660
rect 11300 -30730 11310 -30670
rect 12810 -30730 12820 -30670
rect 11300 -30740 12820 -30730
rect 13020 -30760 13080 -30150
rect 13240 -30760 13300 -30150
rect 13500 -30430 13700 -30350
rect 14160 -30430 14360 -30350
rect 14820 -30430 15020 -30350
rect 13500 -30500 13700 -30490
rect 13500 -30560 13510 -30500
rect 13690 -30560 13700 -30500
rect 13500 -30570 13700 -30560
rect 14160 -30500 14360 -30490
rect 14160 -30560 14170 -30500
rect 14350 -30560 14360 -30500
rect 14160 -30570 14360 -30560
rect 14820 -30500 15020 -30490
rect 14820 -30560 14830 -30500
rect 15010 -30560 15020 -30500
rect 14820 -30570 15020 -30560
rect 13500 -30670 15020 -30660
rect 13500 -30730 13510 -30670
rect 15010 -30730 15020 -30670
rect 13500 -30740 15020 -30730
rect 15220 -30760 15280 -30150
rect 15440 -30760 15500 -30150
rect 15700 -30360 15900 -30350
rect 15700 -30420 15710 -30360
rect 15890 -30420 15900 -30360
rect 15700 -30430 15900 -30420
rect 16360 -30360 16560 -30350
rect 16360 -30420 16370 -30360
rect 16550 -30420 16560 -30360
rect 16360 -30430 16560 -30420
rect 17020 -30360 17220 -30350
rect 17020 -30420 17030 -30360
rect 17210 -30420 17220 -30360
rect 17020 -30430 17220 -30420
rect 15700 -30570 15900 -30490
rect 16360 -30570 16560 -30490
rect 17020 -30570 17220 -30490
rect 15700 -30670 17220 -30660
rect 15700 -30730 15710 -30670
rect 17210 -30730 17220 -30670
rect 15700 -30740 17220 -30730
rect 17420 -30760 17480 -30150
rect 17640 -30760 17700 -30150
rect 17900 -30360 18100 -30350
rect 17900 -30420 17910 -30360
rect 18090 -30420 18100 -30360
rect 17900 -30430 18100 -30420
rect 18560 -30360 18760 -30350
rect 18560 -30420 18570 -30360
rect 18750 -30420 18760 -30360
rect 18560 -30430 18760 -30420
rect 19220 -30360 19420 -30350
rect 19220 -30420 19230 -30360
rect 19410 -30420 19420 -30360
rect 19220 -30430 19420 -30420
rect 17900 -30570 18100 -30490
rect 18560 -30570 18760 -30490
rect 19220 -30570 19420 -30490
rect 17900 -30670 19420 -30660
rect 17900 -30730 17910 -30670
rect 19410 -30730 19420 -30670
rect 17900 -30740 19420 -30730
rect 19620 -30760 19680 -30150
rect 19840 -30760 19900 -30150
rect 2010 -30930 2090 -30760
rect 2230 -30860 2310 -30760
rect 2230 -30920 2240 -30860
rect 2300 -30920 2310 -30860
rect 2230 -30930 2310 -30920
rect 2020 -31700 2080 -30930
rect 80 -32110 90 -31730
rect 270 -32110 280 -31730
rect 1980 -31710 2120 -31700
rect 1980 -31830 1990 -31710
rect 2110 -31830 2120 -31710
rect 1980 -31840 2120 -31830
rect 80 -32120 280 -32110
rect 2020 -32140 2080 -31840
rect 2240 -32000 2300 -30930
rect 4210 -30950 4290 -30760
rect 4430 -30770 4510 -30760
rect 4430 -30830 4440 -30770
rect 4500 -30830 4510 -30770
rect 4430 -30880 4510 -30830
rect 4430 -30940 4440 -30880
rect 4500 -30940 4510 -30880
rect 4430 -30950 4510 -30940
rect 6410 -30880 6490 -30760
rect 6410 -30940 6420 -30880
rect 6480 -30940 6490 -30880
rect 6410 -30950 6490 -30940
rect 6630 -30770 6710 -30760
rect 6630 -30830 6640 -30770
rect 6700 -30830 6710 -30770
rect 6630 -30950 6710 -30830
rect 8610 -30770 8690 -30760
rect 8610 -30830 8620 -30770
rect 8680 -30830 8690 -30770
rect 8610 -30880 8690 -30830
rect 8610 -30940 8620 -30880
rect 8680 -30940 8690 -30880
rect 8610 -30950 8690 -30940
rect 8830 -30950 8910 -30760
rect 10810 -30770 10890 -30760
rect 10810 -30830 10820 -30770
rect 10880 -30830 10890 -30770
rect 10810 -30880 10890 -30830
rect 10810 -30940 10820 -30880
rect 10880 -30940 10890 -30880
rect 10810 -30950 10890 -30940
rect 11030 -30950 11110 -30760
rect 13010 -30770 13090 -30760
rect 13010 -30830 13020 -30770
rect 13080 -30830 13090 -30770
rect 13010 -30880 13090 -30830
rect 13010 -30940 13020 -30880
rect 13080 -30940 13090 -30880
rect 13010 -30950 13090 -30940
rect 13230 -30950 13310 -30760
rect 15210 -30770 15290 -30760
rect 15210 -30830 15220 -30770
rect 15280 -30830 15290 -30770
rect 15210 -30950 15290 -30830
rect 15430 -30880 15510 -30760
rect 15430 -30940 15440 -30880
rect 15500 -30940 15510 -30880
rect 15430 -30950 15510 -30940
rect 17410 -30950 17490 -30760
rect 17630 -30770 17710 -30760
rect 17630 -30830 17640 -30770
rect 17700 -30830 17710 -30770
rect 17630 -30880 17710 -30830
rect 17630 -30940 17640 -30880
rect 17700 -30940 17710 -30880
rect 17630 -30950 17710 -30940
rect 19610 -30950 19690 -30760
rect 19830 -30770 19910 -30760
rect 19830 -30830 19840 -30770
rect 19900 -30830 19910 -30770
rect 19830 -30950 19910 -30830
rect 2500 -31230 2700 -31150
rect 3160 -31230 3360 -31150
rect 3820 -31230 4020 -31150
rect 2500 -31300 2700 -31290
rect 2500 -31360 2510 -31300
rect 2690 -31360 2700 -31300
rect 2500 -31370 2700 -31360
rect 3160 -31300 3360 -31290
rect 3160 -31360 3170 -31300
rect 3350 -31360 3360 -31300
rect 3160 -31370 3360 -31360
rect 3820 -31300 4020 -31290
rect 3820 -31360 3830 -31300
rect 4010 -31360 4020 -31300
rect 3820 -31370 4020 -31360
rect 4220 -31700 4280 -30950
rect 4180 -31710 4320 -31700
rect 4180 -31830 4190 -31710
rect 4310 -31830 4320 -31710
rect 4180 -31840 4320 -31830
rect 2200 -32010 2340 -32000
rect 2200 -32130 2210 -32010
rect 2330 -32130 2340 -32010
rect 2200 -32140 2340 -32130
rect 4220 -32140 4280 -31840
rect 4440 -32000 4500 -30950
rect 4700 -31230 4900 -31150
rect 5360 -31230 5560 -31150
rect 6020 -31230 6220 -31150
rect 4700 -31300 4900 -31290
rect 4700 -31360 4710 -31300
rect 4890 -31360 4900 -31300
rect 4700 -31370 4900 -31360
rect 5360 -31300 5560 -31290
rect 5360 -31360 5370 -31300
rect 5550 -31360 5560 -31300
rect 5360 -31370 5560 -31360
rect 6020 -31300 6220 -31290
rect 6020 -31360 6030 -31300
rect 6210 -31360 6220 -31300
rect 6020 -31370 6220 -31360
rect 6420 -31700 6480 -30950
rect 6380 -31710 6520 -31700
rect 6380 -31830 6390 -31710
rect 6510 -31830 6520 -31710
rect 6380 -31840 6520 -31830
rect 4400 -32010 4540 -32000
rect 4400 -32130 4410 -32010
rect 4530 -32130 4540 -32010
rect 4400 -32140 4540 -32130
rect 6420 -32140 6480 -31840
rect 6640 -32000 6700 -30950
rect 6900 -31160 7100 -31150
rect 6900 -31220 6910 -31160
rect 7090 -31220 7100 -31160
rect 6900 -31230 7100 -31220
rect 7560 -31160 7760 -31150
rect 7560 -31220 7570 -31160
rect 7750 -31220 7760 -31160
rect 7560 -31230 7760 -31220
rect 8220 -31160 8420 -31150
rect 8220 -31220 8230 -31160
rect 8410 -31220 8420 -31160
rect 8220 -31230 8420 -31220
rect 6900 -31370 7100 -31290
rect 7560 -31370 7760 -31290
rect 8220 -31370 8420 -31290
rect 8620 -31700 8680 -30950
rect 8580 -31710 8720 -31700
rect 8580 -31830 8590 -31710
rect 8710 -31830 8720 -31710
rect 8580 -31840 8720 -31830
rect 6600 -32010 6740 -32000
rect 6600 -32130 6610 -32010
rect 6730 -32130 6740 -32010
rect 6600 -32140 6740 -32130
rect 8620 -32140 8680 -31840
rect 8840 -32000 8900 -30950
rect 9100 -31160 9300 -31150
rect 9100 -31220 9110 -31160
rect 9290 -31220 9300 -31160
rect 9100 -31230 9300 -31220
rect 9760 -31160 9960 -31150
rect 9760 -31220 9770 -31160
rect 9950 -31220 9960 -31160
rect 9760 -31230 9960 -31220
rect 10420 -31160 10620 -31150
rect 10420 -31220 10430 -31160
rect 10610 -31220 10620 -31160
rect 10420 -31230 10620 -31220
rect 9100 -31370 9300 -31290
rect 9760 -31370 9960 -31290
rect 10420 -31370 10620 -31290
rect 10820 -31700 10880 -30950
rect 10780 -31710 10920 -31700
rect 10780 -31830 10790 -31710
rect 10910 -31830 10920 -31710
rect 10780 -31840 10920 -31830
rect 8800 -32010 8940 -32000
rect 8800 -32130 8810 -32010
rect 8930 -32130 8940 -32010
rect 8800 -32140 8940 -32130
rect 10820 -32140 10880 -31840
rect 11040 -32000 11100 -30950
rect 11300 -31160 11500 -31150
rect 11300 -31220 11310 -31160
rect 11490 -31220 11500 -31160
rect 11300 -31230 11500 -31220
rect 11960 -31160 12160 -31150
rect 11960 -31220 11970 -31160
rect 12150 -31220 12160 -31160
rect 11960 -31230 12160 -31220
rect 12620 -31160 12820 -31150
rect 12620 -31220 12630 -31160
rect 12810 -31220 12820 -31160
rect 12620 -31230 12820 -31220
rect 11300 -31370 11500 -31290
rect 11960 -31370 12160 -31290
rect 12620 -31370 12820 -31290
rect 13020 -31700 13080 -30950
rect 12980 -31710 13120 -31700
rect 12980 -31830 12990 -31710
rect 13110 -31830 13120 -31710
rect 12980 -31840 13120 -31830
rect 11000 -32010 11140 -32000
rect 11000 -32130 11010 -32010
rect 11130 -32130 11140 -32010
rect 11000 -32140 11140 -32130
rect 13020 -32140 13080 -31840
rect 13240 -32000 13300 -30950
rect 13500 -31160 13700 -31150
rect 13500 -31220 13510 -31160
rect 13690 -31220 13700 -31160
rect 13500 -31230 13700 -31220
rect 14160 -31160 14360 -31150
rect 14160 -31220 14170 -31160
rect 14350 -31220 14360 -31160
rect 14160 -31230 14360 -31220
rect 14820 -31160 15020 -31150
rect 14820 -31220 14830 -31160
rect 15010 -31220 15020 -31160
rect 14820 -31230 15020 -31220
rect 13500 -31370 13700 -31290
rect 14160 -31370 14360 -31290
rect 14820 -31370 15020 -31290
rect 15220 -31700 15280 -30950
rect 15180 -31710 15320 -31700
rect 15180 -31830 15190 -31710
rect 15310 -31830 15320 -31710
rect 15180 -31840 15320 -31830
rect 13200 -32010 13340 -32000
rect 13200 -32130 13210 -32010
rect 13330 -32130 13340 -32010
rect 13200 -32140 13340 -32130
rect 15220 -32140 15280 -31840
rect 15440 -32000 15500 -30950
rect 15700 -31230 15900 -31150
rect 16360 -31230 16560 -31150
rect 17020 -31230 17220 -31150
rect 15700 -31300 15900 -31290
rect 15700 -31360 15710 -31300
rect 15890 -31360 15900 -31300
rect 15700 -31370 15900 -31360
rect 16360 -31300 16560 -31290
rect 16360 -31360 16370 -31300
rect 16550 -31360 16560 -31300
rect 16360 -31370 16560 -31360
rect 17020 -31300 17220 -31290
rect 17020 -31360 17030 -31300
rect 17210 -31360 17220 -31300
rect 17020 -31370 17220 -31360
rect 17420 -31700 17480 -30950
rect 17380 -31710 17520 -31700
rect 17380 -31830 17390 -31710
rect 17510 -31830 17520 -31710
rect 17380 -31840 17520 -31830
rect 15400 -32010 15540 -32000
rect 15400 -32130 15410 -32010
rect 15530 -32130 15540 -32010
rect 15400 -32140 15540 -32130
rect 17420 -32140 17480 -31840
rect 17640 -32000 17700 -30950
rect 17900 -31230 18100 -31150
rect 18560 -31230 18760 -31150
rect 19220 -31230 19420 -31150
rect 17900 -31300 18100 -31290
rect 17900 -31360 17910 -31300
rect 18090 -31360 18100 -31300
rect 17900 -31370 18100 -31360
rect 18560 -31300 18760 -31290
rect 18560 -31360 18570 -31300
rect 18750 -31360 18760 -31300
rect 18560 -31370 18760 -31360
rect 19220 -31300 19420 -31290
rect 19220 -31360 19230 -31300
rect 19410 -31360 19420 -31300
rect 19220 -31370 19420 -31360
rect 19620 -31700 19680 -30950
rect 19580 -31710 19720 -31700
rect 19580 -31830 19590 -31710
rect 19710 -31830 19720 -31710
rect 19580 -31840 19720 -31830
rect 17600 -32010 17740 -32000
rect 17600 -32130 17610 -32010
rect 17730 -32130 17740 -32010
rect 17600 -32140 17740 -32130
rect 19620 -32140 19680 -31840
rect 19840 -32000 19900 -30950
rect 25690 -31510 26230 -31500
rect 25690 -31880 25700 -31510
rect 26220 -31600 26230 -31510
rect 26520 -31600 26720 -25630
rect 27260 -25820 27320 -25630
rect 27250 -25830 27330 -25820
rect 27250 -25920 27260 -25830
rect 27320 -25920 27330 -25830
rect 27250 -25930 27330 -25920
rect 27260 -26135 27320 -25930
rect 27250 -26145 27330 -26135
rect 27250 -26235 27260 -26145
rect 27320 -26235 27330 -26145
rect 27250 -26245 27330 -26235
rect 27260 -27585 27320 -26245
rect 27380 -26700 27440 -25080
rect 27370 -26710 27450 -26700
rect 27370 -26800 27380 -26710
rect 27440 -26800 27450 -26710
rect 27370 -26810 27450 -26800
rect 27380 -27015 27440 -26810
rect 27370 -27025 27450 -27015
rect 27370 -27115 27380 -27025
rect 27440 -27115 27450 -27025
rect 27370 -27125 27450 -27115
rect 27250 -27595 27330 -27585
rect 27250 -27685 27260 -27595
rect 27320 -27685 27330 -27595
rect 27250 -27695 27330 -27685
rect 27260 -27900 27320 -27695
rect 27250 -27910 27330 -27900
rect 27250 -28000 27260 -27910
rect 27320 -28000 27330 -27910
rect 27250 -28010 27330 -28000
rect 27260 -28215 27320 -28010
rect 27250 -28225 27330 -28215
rect 27250 -28315 27260 -28225
rect 27320 -28315 27330 -28225
rect 27250 -28325 27330 -28315
rect 27260 -28620 27320 -28325
rect 27250 -28630 27330 -28620
rect 27250 -28720 27260 -28630
rect 27320 -28720 27330 -28630
rect 27250 -28730 27330 -28720
rect 27260 -28940 27320 -28730
rect 27250 -28950 27330 -28940
rect 27250 -29040 27260 -28950
rect 27320 -29040 27330 -28950
rect 27250 -29050 27330 -29040
rect 27260 -29250 27320 -29050
rect 27250 -29260 27330 -29250
rect 27250 -29350 27260 -29260
rect 27320 -29350 27330 -29260
rect 27250 -29360 27330 -29350
rect 27260 -31600 27320 -29360
rect 27380 -29660 27440 -27125
rect 27500 -27740 27560 -24660
rect 27490 -27750 27570 -27740
rect 27490 -27840 27500 -27750
rect 27560 -27840 27570 -27750
rect 27490 -27850 27570 -27840
rect 27500 -28055 27560 -27850
rect 27490 -28065 27570 -28055
rect 27490 -28155 27500 -28065
rect 27560 -28155 27570 -28065
rect 27490 -28165 27570 -28155
rect 27370 -29670 27450 -29660
rect 27370 -29760 27380 -29670
rect 27440 -29760 27450 -29670
rect 27370 -29770 27450 -29760
rect 27380 -29975 27440 -29770
rect 27370 -29985 27450 -29975
rect 27370 -30075 27380 -29985
rect 27440 -30075 27450 -29985
rect 27370 -30085 27450 -30075
rect 27380 -30290 27440 -30085
rect 27370 -30300 27450 -30290
rect 27370 -30390 27380 -30300
rect 27440 -30390 27450 -30300
rect 27370 -30400 27450 -30390
rect 27380 -30700 27440 -30400
rect 27370 -30710 27450 -30700
rect 27370 -30800 27380 -30710
rect 27440 -30800 27450 -30710
rect 27370 -30810 27450 -30800
rect 27380 -31015 27440 -30810
rect 27500 -30860 27560 -28165
rect 27620 -28780 27680 -24260
rect 29370 -24490 29450 -24480
rect 29370 -24720 29380 -24490
rect 29440 -24720 29450 -24490
rect 29370 -24730 29450 -24720
rect 29520 -24640 29600 -24630
rect 27730 -25670 27810 -25660
rect 27730 -25760 27740 -25670
rect 27800 -25760 27810 -25670
rect 29380 -25760 29440 -24730
rect 29520 -24870 29530 -24640
rect 29590 -24870 29600 -24640
rect 29520 -24880 29600 -24870
rect 27730 -25770 27810 -25760
rect 29370 -25770 29450 -25760
rect 27740 -25975 27800 -25770
rect 29370 -25970 29380 -25770
rect 29440 -25970 29450 -25770
rect 27730 -25985 27810 -25975
rect 29370 -25980 29450 -25970
rect 27730 -26075 27740 -25985
rect 27800 -26075 27810 -25985
rect 27730 -26085 27810 -26075
rect 27740 -26540 27800 -26085
rect 27730 -26550 27810 -26540
rect 27730 -26640 27740 -26550
rect 27800 -26640 27810 -26550
rect 27730 -26650 27810 -26640
rect 27740 -26860 27800 -26650
rect 27730 -26870 27810 -26860
rect 27730 -26960 27740 -26870
rect 27800 -26960 27810 -26870
rect 27730 -26970 27810 -26960
rect 27740 -27175 27800 -26970
rect 27730 -27185 27810 -27175
rect 27730 -27275 27740 -27185
rect 27800 -27275 27810 -27185
rect 27730 -27285 27810 -27275
rect 29070 -27850 29150 -27840
rect 29070 -28050 29080 -27850
rect 29140 -28050 29150 -27850
rect 29070 -28060 29150 -28050
rect 27610 -28790 27690 -28780
rect 27610 -28880 27620 -28790
rect 27680 -28880 27690 -28790
rect 27610 -28890 27690 -28880
rect 27620 -29100 27680 -28890
rect 27610 -29110 27690 -29100
rect 27610 -29200 27620 -29110
rect 27680 -29200 27690 -29110
rect 27610 -29210 27690 -29200
rect 27620 -29820 27680 -29210
rect 27610 -29830 27690 -29820
rect 27610 -29920 27620 -29830
rect 27680 -29920 27690 -29830
rect 29080 -29920 29140 -28060
rect 29220 -28890 29300 -28880
rect 29220 -29090 29230 -28890
rect 29290 -29090 29300 -28890
rect 29220 -29100 29300 -29090
rect 27610 -29930 27690 -29920
rect 29070 -29930 29150 -29920
rect 27620 -30135 27680 -29930
rect 29070 -30130 29080 -29930
rect 29140 -30130 29150 -29930
rect 27610 -30145 27690 -30135
rect 29070 -30140 29150 -30130
rect 27610 -30235 27620 -30145
rect 27680 -30235 27690 -30145
rect 27610 -30245 27690 -30235
rect 27490 -30870 27570 -30860
rect 27490 -30960 27500 -30870
rect 27560 -30960 27570 -30870
rect 27490 -30970 27570 -30960
rect 27370 -31025 27450 -31015
rect 27370 -31115 27380 -31025
rect 27440 -31115 27450 -31025
rect 27370 -31125 27450 -31115
rect 27380 -31330 27440 -31125
rect 27500 -31175 27560 -30970
rect 27490 -31185 27570 -31175
rect 27490 -31275 27500 -31185
rect 27560 -31275 27570 -31185
rect 27490 -31285 27570 -31275
rect 27370 -31340 27450 -31330
rect 27370 -31430 27380 -31340
rect 27440 -31430 27450 -31340
rect 27370 -31440 27450 -31430
rect 27380 -31600 27440 -31440
rect 27500 -31600 27560 -31285
rect 27620 -31600 27680 -30245
rect 29080 -30800 29140 -30140
rect 28930 -30810 29170 -30800
rect 28930 -30880 28940 -30810
rect 29160 -30880 29170 -30810
rect 28930 -30890 29170 -30880
rect 29230 -30950 29290 -29100
rect 29060 -30960 29300 -30950
rect 29060 -31030 29070 -30960
rect 29290 -31030 29300 -30960
rect 29060 -31040 29300 -31030
rect 29380 -31100 29440 -25980
rect 29530 -26800 29590 -24880
rect 29520 -26810 29600 -26800
rect 29520 -27010 29530 -26810
rect 29590 -27010 29600 -26810
rect 29520 -27020 29600 -27010
rect 29210 -31110 29450 -31100
rect 29210 -31180 29220 -31110
rect 29440 -31180 29450 -31110
rect 29210 -31190 29450 -31180
rect 29530 -31250 29590 -27020
rect 29680 -28710 29740 -24110
rect 29670 -28720 29750 -28710
rect 29670 -28940 29680 -28720
rect 29740 -28940 29750 -28720
rect 29830 -28860 29890 -23600
rect 31860 -23660 31960 -17210
rect 32510 -17800 32640 -16920
rect 32510 -18480 32520 -17800
rect 32630 -18480 32640 -17800
rect 32510 -18490 32640 -18480
rect 32510 -19600 32640 -19590
rect 32510 -20280 32520 -19600
rect 32630 -20280 32640 -19600
rect 32510 -20360 32640 -20280
rect 33180 -20340 33320 -20330
rect 32500 -20370 32650 -20360
rect 32500 -20530 32510 -20370
rect 32640 -20530 32650 -20370
rect 33180 -20460 33190 -20340
rect 33310 -20460 33320 -20340
rect 33180 -20470 33320 -20460
rect 32500 -20540 32650 -20530
rect 32510 -21400 32640 -20540
rect 32510 -22080 32520 -21400
rect 32630 -22080 32640 -21400
rect 32510 -22090 32640 -22080
rect 33200 -22140 33300 -20470
rect 33200 -22240 33210 -22140
rect 33290 -22240 33300 -22140
rect 33200 -22420 33300 -22240
rect 32620 -22430 33310 -22420
rect 32620 -22490 32630 -22430
rect 33300 -22490 33310 -22430
rect 32620 -22500 33310 -22490
rect 32690 -23070 33240 -23060
rect 32690 -23150 32700 -23070
rect 32910 -23150 33020 -23070
rect 33230 -23150 33240 -23070
rect 32690 -23160 33240 -23150
rect 31810 -23670 32010 -23660
rect 31810 -23850 31820 -23670
rect 32000 -23850 32010 -23670
rect 31810 -23860 32010 -23850
rect 29970 -24140 30050 -24130
rect 29970 -24370 29980 -24140
rect 30040 -24370 30050 -24140
rect 29970 -24380 30050 -24370
rect 29670 -28950 29750 -28940
rect 29820 -28870 29900 -28860
rect 29820 -29090 29830 -28870
rect 29890 -29090 29900 -28870
rect 29980 -29010 30040 -24380
rect 32880 -24470 32940 -23160
rect 33440 -23550 33540 -9640
rect 34100 -9570 34250 -9560
rect 34100 -9730 34110 -9570
rect 34240 -9730 34250 -9570
rect 34100 -9740 34250 -9730
rect 34110 -10600 34240 -9740
rect 34820 -9860 34920 -8200
rect 35710 -8800 35840 -8790
rect 35710 -9360 35720 -8800
rect 35830 -9360 35840 -8800
rect 35710 -9560 35840 -9360
rect 35700 -9570 35850 -9560
rect 35700 -9730 35710 -9570
rect 35840 -9730 35850 -9570
rect 35700 -9740 35850 -9730
rect 34800 -9870 34940 -9860
rect 34800 -9990 34810 -9870
rect 34930 -9990 34940 -9870
rect 34800 -10000 34940 -9990
rect 34110 -11110 34120 -10600
rect 34230 -11110 34240 -10600
rect 34110 -11360 34240 -11110
rect 34100 -11370 34250 -11360
rect 34100 -11530 34110 -11370
rect 34240 -11530 34250 -11370
rect 34100 -11540 34250 -11530
rect 34110 -12400 34240 -11540
rect 34820 -11660 34920 -10000
rect 35710 -10600 35840 -9740
rect 35710 -11110 35720 -10600
rect 35830 -11110 35840 -10600
rect 35000 -11310 35140 -11300
rect 35000 -11430 35010 -11310
rect 35130 -11430 35140 -11310
rect 35710 -11360 35840 -11110
rect 35000 -11440 35140 -11430
rect 34800 -11670 34940 -11660
rect 34800 -11790 34810 -11670
rect 34930 -11790 34940 -11670
rect 34800 -11800 34940 -11790
rect 34110 -12910 34120 -12400
rect 34230 -12910 34240 -12400
rect 34110 -13160 34240 -12910
rect 34100 -13170 34250 -13160
rect 34100 -13330 34110 -13170
rect 34240 -13330 34250 -13170
rect 34100 -13340 34250 -13330
rect 34110 -14200 34240 -13340
rect 34820 -13460 34920 -11800
rect 35040 -13100 35140 -11440
rect 35700 -11370 35850 -11360
rect 35700 -11530 35710 -11370
rect 35840 -11530 35850 -11370
rect 35700 -11540 35850 -11530
rect 35000 -13110 35140 -13100
rect 35000 -13230 35010 -13110
rect 35130 -13230 35140 -13110
rect 35710 -12400 35840 -11540
rect 35710 -12910 35720 -12400
rect 35830 -12910 35840 -12400
rect 35710 -13160 35840 -12910
rect 35000 -13240 35140 -13230
rect 34800 -13470 34940 -13460
rect 34800 -13590 34810 -13470
rect 34930 -13590 34940 -13470
rect 34800 -13600 34940 -13590
rect 34110 -14710 34120 -14200
rect 34230 -14710 34240 -14200
rect 34110 -14890 34240 -14710
rect 34110 -16000 34240 -15990
rect 34110 -16680 34120 -16000
rect 34230 -16680 34240 -16000
rect 34110 -16770 34240 -16680
rect 34110 -16920 34120 -16770
rect 34230 -16920 34240 -16770
rect 34110 -17800 34240 -16920
rect 34110 -18480 34120 -17800
rect 34230 -18480 34240 -17800
rect 34110 -18490 34240 -18480
rect 34110 -19600 34240 -19590
rect 34110 -20280 34120 -19600
rect 34230 -20280 34240 -19600
rect 34110 -20360 34240 -20280
rect 34100 -20370 34250 -20360
rect 34100 -20530 34110 -20370
rect 34240 -20530 34250 -20370
rect 34100 -20540 34250 -20530
rect 34110 -21400 34240 -20540
rect 34110 -22080 34120 -21400
rect 34230 -22080 34240 -21400
rect 34110 -22090 34240 -22080
rect 34010 -22170 34370 -22160
rect 34010 -22240 34020 -22170
rect 34360 -22240 34370 -22170
rect 34010 -22250 34370 -22240
rect 34030 -22430 34320 -22250
rect 34030 -22490 34040 -22430
rect 34310 -22490 34320 -22430
rect 34030 -22500 34320 -22490
rect 34060 -23100 34310 -23090
rect 34060 -23160 34070 -23100
rect 34300 -23160 34310 -23100
rect 34060 -23170 34310 -23160
rect 33400 -23560 33920 -23550
rect 33400 -23620 33410 -23560
rect 33910 -23620 33920 -23560
rect 33400 -23630 33920 -23620
rect 33160 -24220 34150 -24210
rect 33160 -24280 33170 -24220
rect 33280 -24280 33410 -24220
rect 33600 -24280 33730 -24220
rect 33920 -24280 34040 -24220
rect 34140 -24280 34150 -24220
rect 33160 -24290 34150 -24280
rect 32790 -24480 33040 -24470
rect 32790 -24550 32800 -24480
rect 33030 -24550 33040 -24480
rect 32790 -24560 33040 -24550
rect 33640 -24770 33700 -24290
rect 34200 -24620 34260 -23170
rect 34820 -23460 34920 -13600
rect 35040 -14900 35140 -13240
rect 35700 -13170 35850 -13160
rect 35700 -13330 35710 -13170
rect 35840 -13330 35850 -13170
rect 35700 -13340 35850 -13330
rect 35710 -14200 35840 -13340
rect 35710 -14710 35720 -14200
rect 35830 -14710 35840 -14200
rect 35710 -14890 35840 -14710
rect 35000 -14910 35140 -14900
rect 35000 -15030 35010 -14910
rect 35130 -15030 35140 -14910
rect 35000 -15040 35140 -15030
rect 34610 -24220 34780 -24210
rect 34610 -24280 34620 -24220
rect 34770 -24280 34780 -24220
rect 34610 -24290 34780 -24280
rect 34840 -24480 34900 -23460
rect 35040 -23550 35140 -15040
rect 35710 -16000 35840 -15990
rect 35710 -16680 35720 -16000
rect 35830 -16680 35840 -16000
rect 35710 -16770 35840 -16680
rect 35710 -16920 35720 -16770
rect 35830 -16920 35840 -16770
rect 35710 -17800 35840 -16920
rect 35710 -18480 35720 -17800
rect 35830 -18480 35840 -17800
rect 35710 -18490 35840 -18480
rect 35710 -19600 35840 -19590
rect 35710 -20280 35720 -19600
rect 35830 -20280 35840 -19600
rect 35710 -20360 35840 -20280
rect 35700 -20370 35850 -20360
rect 35700 -20530 35710 -20370
rect 35840 -20530 35850 -20370
rect 35700 -20540 35850 -20530
rect 35710 -21400 35840 -20540
rect 35710 -22080 35720 -21400
rect 35830 -22080 35840 -21400
rect 35710 -22090 35840 -22080
rect 35000 -23560 37030 -23550
rect 37020 -23620 37030 -23560
rect 35000 -23630 37030 -23620
rect 34980 -24220 37030 -24210
rect 34980 -24280 34990 -24220
rect 37020 -24280 37030 -24220
rect 34980 -24290 37030 -24280
rect 34800 -24490 34940 -24480
rect 34800 -24610 34810 -24490
rect 34930 -24610 34940 -24490
rect 34800 -24620 34940 -24610
rect 34110 -24630 34360 -24620
rect 34110 -24700 34120 -24630
rect 34350 -24700 34360 -24630
rect 37120 -24640 37290 -24630
rect 34110 -24710 34360 -24700
rect 34800 -24660 34910 -24650
rect 30280 -24780 30520 -24770
rect 30280 -24850 30290 -24780
rect 30510 -24850 30520 -24780
rect 30280 -24860 30520 -24850
rect 33550 -24780 33800 -24770
rect 33550 -24850 33560 -24780
rect 33790 -24850 33800 -24780
rect 33550 -24860 33800 -24850
rect 34800 -24860 34810 -24660
rect 34900 -24860 34910 -24660
rect 37120 -24780 37130 -24640
rect 37270 -24780 37290 -24640
rect 37120 -24790 37290 -24780
rect 30120 -24940 30200 -24930
rect 30120 -25170 30130 -24940
rect 30190 -25170 30200 -24940
rect 30120 -25180 30200 -25170
rect 29820 -29100 29900 -29090
rect 29970 -29020 30050 -29010
rect 29970 -29240 29980 -29020
rect 30040 -29240 30050 -29020
rect 30130 -29160 30190 -25180
rect 29970 -29250 30050 -29240
rect 30120 -29170 30200 -29160
rect 30120 -29390 30130 -29170
rect 30190 -29390 30200 -29170
rect 30280 -29310 30340 -24860
rect 34800 -24940 34910 -24860
rect 34800 -25010 34810 -24940
rect 34900 -25010 34910 -24940
rect 30420 -25090 30500 -25080
rect 30420 -25320 30430 -25090
rect 30490 -25320 30500 -25090
rect 30420 -25330 30500 -25320
rect 34800 -25200 34910 -25010
rect 34800 -25270 34810 -25200
rect 34900 -25270 34910 -25200
rect 30120 -29400 30200 -29390
rect 30270 -29320 30350 -29310
rect 30270 -29540 30280 -29320
rect 30340 -29540 30350 -29320
rect 30430 -29460 30490 -25330
rect 34800 -25460 34910 -25270
rect 34800 -25530 34810 -25460
rect 34900 -25530 34910 -25460
rect 34800 -25720 34910 -25530
rect 34800 -25790 34810 -25720
rect 34900 -25790 34910 -25720
rect 34800 -25980 34910 -25790
rect 34800 -26050 34810 -25980
rect 34900 -26050 34910 -25980
rect 34800 -26240 34910 -26050
rect 34800 -26310 34810 -26240
rect 34900 -26310 34910 -26240
rect 34800 -26500 34910 -26310
rect 34800 -26570 34810 -26500
rect 34900 -26570 34910 -26500
rect 34800 -26760 34910 -26570
rect 34800 -26830 34810 -26760
rect 34900 -26830 34910 -26760
rect 34800 -26840 34910 -26830
rect 37180 -24940 37290 -24790
rect 37180 -25010 37190 -24940
rect 37280 -25010 37290 -24940
rect 37180 -25200 37290 -25010
rect 37180 -25270 37190 -25200
rect 37280 -25270 37290 -25200
rect 37180 -25460 37290 -25270
rect 37180 -25530 37190 -25460
rect 37280 -25530 37290 -25460
rect 37180 -25720 37290 -25530
rect 37180 -25790 37190 -25720
rect 37280 -25790 37290 -25720
rect 37180 -25980 37290 -25790
rect 37180 -26050 37190 -25980
rect 37280 -26050 37290 -25980
rect 37180 -26240 37290 -26050
rect 37180 -26310 37190 -26240
rect 37280 -26310 37290 -26240
rect 37180 -26500 37290 -26310
rect 37180 -26570 37190 -26500
rect 37280 -26570 37290 -26500
rect 37180 -26760 37290 -26570
rect 37180 -26830 37190 -26760
rect 37280 -26830 37290 -26760
rect 37180 -26840 37290 -26830
rect 36020 -27010 36420 -27000
rect 36020 -27140 36030 -27010
rect 36410 -27140 36420 -27010
rect 36020 -27150 36420 -27140
rect 36520 -27010 36920 -27000
rect 36520 -27140 36530 -27010
rect 36910 -27140 36920 -27010
rect 36520 -27150 36920 -27140
rect 33420 -27640 33600 -27620
rect 33420 -27780 33440 -27640
rect 33580 -27780 33600 -27640
rect 33420 -27800 33600 -27780
rect 31810 -28050 33170 -28040
rect 31810 -28290 31820 -28050
rect 33160 -28290 33170 -28050
rect 31810 -28300 33170 -28290
rect 31988 -28528 32058 -28522
rect 31988 -28700 31994 -28528
rect 31790 -28710 31994 -28700
rect 32052 -28700 32058 -28528
rect 32200 -28528 32270 -28522
rect 31790 -28780 31800 -28710
rect 31790 -28790 31994 -28780
rect 31988 -28914 31994 -28790
rect 32052 -28790 32060 -28700
rect 32052 -28914 32058 -28790
rect 32200 -28850 32206 -28528
rect 30270 -29550 30350 -29540
rect 30420 -29470 30500 -29460
rect 30420 -29690 30430 -29470
rect 30490 -29690 30500 -29470
rect 30420 -29700 30500 -29690
rect 31988 -29548 32058 -28914
rect 32190 -28860 32206 -28850
rect 32264 -28850 32270 -28528
rect 32264 -28860 32460 -28850
rect 32190 -28930 32200 -28860
rect 32450 -28930 32460 -28860
rect 32190 -28940 32460 -28930
rect 31988 -29734 31994 -29548
rect 32052 -29734 32058 -29548
rect 31988 -29740 32058 -29734
rect 32200 -29550 32270 -28940
rect 33460 -29200 33560 -27800
rect 35620 -27840 35800 -27820
rect 35620 -27980 35640 -27840
rect 35780 -27980 35800 -27840
rect 35620 -28000 35800 -27980
rect 34188 -28528 34258 -28522
rect 34188 -28914 34194 -28528
rect 34252 -28914 34258 -28528
rect 34188 -29000 34258 -28914
rect 34400 -28528 34470 -28522
rect 34400 -28914 34406 -28528
rect 34464 -28914 34470 -28528
rect 33990 -29010 34260 -29000
rect 33990 -29080 34000 -29010
rect 34250 -29080 34260 -29010
rect 33990 -29090 34260 -29080
rect 33350 -29210 33570 -29200
rect 32328 -29276 33172 -29270
rect 32328 -29334 32334 -29276
rect 32472 -29334 33004 -29276
rect 33142 -29334 33172 -29276
rect 33350 -29290 33360 -29210
rect 33560 -29290 33570 -29210
rect 33350 -29300 33570 -29290
rect 32328 -29340 33172 -29334
rect 32200 -29736 32206 -29550
rect 32264 -29736 32270 -29550
rect 32200 -29742 32270 -29736
rect 33072 -29376 33172 -29340
rect 33072 -29378 33594 -29376
rect 33072 -29430 33454 -29378
rect 33588 -29430 33594 -29378
rect 33072 -29432 33594 -29430
rect 33072 -29546 33172 -29432
rect 33072 -29736 33078 -29546
rect 33166 -29736 33172 -29546
rect 33072 -29742 33172 -29736
rect 34188 -29548 34258 -29090
rect 34188 -29734 34194 -29548
rect 34252 -29734 34258 -29548
rect 34188 -29740 34258 -29734
rect 34400 -29140 34470 -28914
rect 34400 -29150 34670 -29140
rect 34400 -29220 34410 -29150
rect 34660 -29220 34670 -29150
rect 35660 -29200 35760 -28000
rect 37720 -28040 37900 -28020
rect 37720 -28180 37740 -28040
rect 37880 -28180 37900 -28040
rect 37720 -28200 37900 -28180
rect 36388 -28528 36458 -28522
rect 36388 -28914 36394 -28528
rect 36452 -28914 36458 -28528
rect 34400 -29230 34670 -29220
rect 35550 -29210 35770 -29200
rect 34400 -29550 34470 -29230
rect 34528 -29276 35372 -29270
rect 34528 -29334 34534 -29276
rect 34672 -29334 35204 -29276
rect 35342 -29334 35372 -29276
rect 35550 -29290 35560 -29210
rect 35760 -29290 35770 -29210
rect 35550 -29300 35770 -29290
rect 36388 -29300 36458 -28914
rect 36600 -28528 36670 -28522
rect 36600 -28914 36606 -28528
rect 36664 -28914 36670 -28528
rect 34528 -29340 35372 -29334
rect 34400 -29736 34406 -29550
rect 34464 -29736 34470 -29550
rect 34400 -29742 34470 -29736
rect 35272 -29376 35372 -29340
rect 36190 -29310 36460 -29300
rect 35272 -29378 35794 -29376
rect 35272 -29430 35654 -29378
rect 35788 -29430 35794 -29378
rect 36190 -29380 36200 -29310
rect 36450 -29380 36460 -29310
rect 36190 -29390 36460 -29380
rect 35272 -29432 35794 -29430
rect 35272 -29546 35372 -29432
rect 35272 -29736 35278 -29546
rect 35366 -29736 35372 -29546
rect 35272 -29742 35372 -29736
rect 36388 -29548 36458 -29390
rect 36600 -29450 36670 -28914
rect 37760 -29200 37860 -28200
rect 37750 -29210 37970 -29200
rect 36728 -29276 37572 -29270
rect 36728 -29334 36734 -29276
rect 36872 -29334 37404 -29276
rect 37542 -29334 37572 -29276
rect 37750 -29290 37760 -29210
rect 37960 -29290 37970 -29210
rect 37750 -29300 37970 -29290
rect 36728 -29340 37572 -29334
rect 37472 -29376 37572 -29340
rect 37472 -29378 37994 -29376
rect 37472 -29430 37854 -29378
rect 37988 -29430 37994 -29378
rect 37472 -29432 37994 -29430
rect 36590 -29460 36860 -29450
rect 36590 -29530 36600 -29460
rect 36850 -29530 36860 -29460
rect 36590 -29540 36860 -29530
rect 36388 -29734 36394 -29548
rect 36452 -29734 36458 -29548
rect 36388 -29740 36458 -29734
rect 36600 -29550 36670 -29540
rect 36600 -29736 36606 -29550
rect 36664 -29736 36670 -29550
rect 36600 -29742 36670 -29736
rect 37472 -29546 37572 -29432
rect 37472 -29736 37478 -29546
rect 37566 -29736 37572 -29546
rect 37472 -29742 37572 -29736
rect 37240 -29920 37700 -29910
rect 37240 -30110 37250 -29920
rect 37690 -30110 37700 -29920
rect 37240 -30120 37700 -30110
rect 32250 -30288 32350 -30282
rect 32250 -30478 32256 -30288
rect 32344 -30478 32350 -30288
rect 32250 -30592 32350 -30478
rect 31828 -30594 32350 -30592
rect 31828 -30646 31834 -30594
rect 31968 -30646 32350 -30594
rect 31828 -30648 32350 -30646
rect 32250 -30684 32350 -30648
rect 33152 -30288 33222 -30282
rect 33152 -30474 33158 -30288
rect 33216 -30474 33222 -30288
rect 32250 -30690 33094 -30684
rect 31840 -30730 32060 -30720
rect 31840 -30810 31850 -30730
rect 32050 -30810 32060 -30730
rect 32250 -30748 32280 -30690
rect 32418 -30748 32950 -30690
rect 33088 -30748 33094 -30690
rect 32250 -30754 33094 -30748
rect 33152 -30800 33222 -30474
rect 31840 -30820 32060 -30810
rect 32950 -30810 33222 -30800
rect 29360 -31260 29600 -31250
rect 29360 -31330 29370 -31260
rect 29590 -31330 29600 -31260
rect 29360 -31340 29600 -31330
rect 26220 -31800 27320 -31600
rect 26220 -31880 26230 -31800
rect 31880 -31880 31980 -30820
rect 32950 -30880 32960 -30810
rect 33210 -30880 33222 -30810
rect 32950 -30890 33222 -30880
rect 33152 -31110 33222 -30890
rect 33364 -30290 33434 -30284
rect 33364 -30476 33370 -30290
rect 33428 -30476 33434 -30290
rect 33364 -30950 33434 -30476
rect 34450 -30288 34550 -30282
rect 34450 -30478 34456 -30288
rect 34544 -30478 34550 -30288
rect 34450 -30592 34550 -30478
rect 34028 -30594 34550 -30592
rect 34028 -30646 34034 -30594
rect 34168 -30646 34550 -30594
rect 34028 -30648 34550 -30646
rect 34450 -30684 34550 -30648
rect 35352 -30288 35422 -30282
rect 35352 -30474 35358 -30288
rect 35416 -30474 35422 -30288
rect 34450 -30690 35294 -30684
rect 34050 -30730 34270 -30720
rect 34050 -30810 34060 -30730
rect 34260 -30810 34270 -30730
rect 34450 -30748 34480 -30690
rect 34618 -30748 35150 -30690
rect 35288 -30748 35294 -30690
rect 34450 -30754 35294 -30748
rect 34050 -30820 34270 -30810
rect 33320 -30960 33590 -30950
rect 33320 -31030 33330 -30960
rect 33580 -31030 33590 -30960
rect 33320 -31040 33590 -31030
rect 33152 -31496 33158 -31110
rect 33216 -31496 33222 -31110
rect 33152 -31502 33222 -31496
rect 33364 -31110 33434 -31040
rect 33364 -31496 33370 -31110
rect 33428 -31496 33434 -31110
rect 33364 -31502 33434 -31496
rect 32530 -31730 33700 -31720
rect 25690 -31890 26230 -31880
rect 32530 -31950 32540 -31730
rect 33690 -31950 33700 -31730
rect 34080 -31880 34180 -30820
rect 35352 -31110 35422 -30474
rect 35564 -30290 35634 -30284
rect 35564 -30476 35570 -30290
rect 35628 -30476 35634 -30290
rect 35564 -31100 35634 -30476
rect 36650 -30288 36750 -30282
rect 36650 -30478 36656 -30288
rect 36744 -30478 36750 -30288
rect 36650 -30592 36750 -30478
rect 36228 -30594 36750 -30592
rect 36228 -30646 36234 -30594
rect 36368 -30646 36750 -30594
rect 36228 -30648 36750 -30646
rect 36650 -30684 36750 -30648
rect 37552 -30288 37622 -30282
rect 37552 -30474 37558 -30288
rect 37616 -30474 37622 -30288
rect 36650 -30690 37494 -30684
rect 36250 -30740 36470 -30730
rect 36250 -30820 36260 -30740
rect 36460 -30820 36470 -30740
rect 36650 -30748 36680 -30690
rect 36818 -30748 37350 -30690
rect 37488 -30748 37494 -30690
rect 36650 -30754 37494 -30748
rect 36250 -30830 36470 -30820
rect 35352 -31496 35358 -31110
rect 35416 -31496 35422 -31110
rect 35550 -31110 35820 -31100
rect 35550 -31180 35560 -31110
rect 35810 -31180 35820 -31110
rect 35550 -31190 35570 -31180
rect 35352 -31502 35422 -31496
rect 35564 -31496 35570 -31190
rect 35628 -31190 35820 -31180
rect 35628 -31496 35634 -31190
rect 35564 -31502 35634 -31496
rect 36280 -31880 36380 -30830
rect 37552 -31110 37622 -30474
rect 37552 -31496 37558 -31110
rect 37616 -31496 37622 -31110
rect 37764 -30290 37834 -30284
rect 37764 -30476 37770 -30290
rect 37828 -30476 37834 -30290
rect 37764 -31110 37834 -30476
rect 37764 -31250 37770 -31110
rect 37700 -31260 37770 -31250
rect 37828 -31250 37834 -31110
rect 37828 -31260 37970 -31250
rect 37700 -31330 37710 -31260
rect 37960 -31330 37970 -31260
rect 37700 -31340 37770 -31330
rect 37552 -31502 37622 -31496
rect 37764 -31496 37770 -31340
rect 37828 -31340 37970 -31330
rect 37828 -31496 37834 -31340
rect 37764 -31502 37834 -31496
rect 32530 -31960 33700 -31950
rect 19800 -32010 19940 -32000
rect 19800 -32130 19810 -32010
rect 19930 -32130 19940 -32010
rect 19800 -32140 19940 -32130
<< via2 >>
rect -350 11610 -170 11990
rect 2210 11890 2330 12010
rect 90 11310 270 11690
rect 1990 11590 2110 11710
rect -70 10870 -10 10930
rect -70 10070 -10 10130
rect -70 9270 -10 9330
rect -70 8470 -10 8530
rect -70 7670 -10 7730
rect -70 6870 -10 6930
rect -70 6070 -10 6130
rect -70 5270 -10 5330
rect -350 -31830 -170 -31450
rect 2130 10870 2190 10930
rect 4410 11890 4530 12010
rect 4190 11590 4310 11710
rect 2510 11180 2690 11240
rect 3170 11180 3350 11240
rect 3830 11180 4010 11240
rect 4330 10870 4390 10930
rect 6610 11890 6730 12010
rect 6390 11590 6510 11710
rect 4710 11180 4890 11240
rect 5370 11180 5550 11240
rect 6030 11180 6210 11240
rect 6530 10870 6590 10930
rect 8810 11890 8930 12010
rect 8590 11590 8710 11710
rect 6910 11040 7090 11100
rect 7570 11040 7750 11100
rect 8230 11040 8410 11100
rect 8730 10870 8790 10930
rect 11010 11890 11130 12010
rect 10790 11590 10910 11710
rect 9110 11040 9290 11100
rect 9770 11040 9950 11100
rect 10430 11040 10610 11100
rect 10930 10870 10990 10930
rect 13210 11890 13330 12010
rect 12990 11590 13110 11710
rect 11310 11040 11490 11100
rect 11970 11040 12150 11100
rect 12630 11040 12810 11100
rect 13130 10870 13190 10930
rect 15410 11890 15530 12010
rect 15190 11590 15310 11710
rect 13510 11040 13690 11100
rect 14170 11040 14350 11100
rect 14830 11040 15010 11100
rect 15330 10870 15390 10930
rect 17610 11890 17730 12010
rect 17390 11590 17510 11710
rect 15710 11180 15890 11240
rect 16370 11180 16550 11240
rect 17030 11180 17210 11240
rect 17530 10870 17590 10930
rect 19810 11890 19930 12010
rect 19590 11590 19710 11710
rect 17910 11180 18090 11240
rect 18570 11180 18750 11240
rect 19230 11180 19410 11240
rect 19730 10870 19790 10930
rect 21930 10870 21990 10930
rect 2130 10070 2190 10130
rect 2510 10550 4010 10610
rect 2510 10240 2690 10300
rect 3170 10240 3350 10300
rect 3830 10240 4010 10300
rect 4330 10070 4390 10130
rect 4710 10550 6210 10610
rect 4710 10240 4890 10300
rect 5370 10240 5550 10300
rect 6030 10240 6210 10300
rect 6530 10070 6590 10130
rect 6910 10550 8410 10610
rect 6910 10380 7090 10440
rect 7570 10380 7750 10440
rect 8230 10380 8410 10440
rect 8730 10070 8790 10130
rect 9110 10550 10610 10610
rect 9110 10380 9290 10440
rect 9770 10380 9950 10440
rect 10430 10380 10610 10440
rect 10930 10070 10990 10130
rect 11310 10550 12810 10610
rect 11310 10380 11490 10440
rect 11970 10380 12150 10440
rect 12630 10380 12810 10440
rect 13130 10070 13190 10130
rect 13510 10550 15010 10610
rect 13510 10380 13690 10440
rect 14170 10380 14350 10440
rect 14830 10380 15010 10440
rect 15330 10070 15390 10130
rect 15710 10550 17210 10610
rect 15710 10240 15890 10300
rect 16370 10240 16550 10300
rect 17030 10240 17210 10300
rect 17530 10070 17590 10130
rect 17910 10550 19410 10610
rect 17910 10240 18090 10300
rect 18570 10240 18750 10300
rect 19230 10240 19410 10300
rect 19730 10070 19790 10130
rect 21930 10070 21990 10130
rect 2130 9270 2190 9330
rect 2510 9750 4010 9810
rect 2510 9580 2690 9640
rect 3170 9580 3350 9640
rect 3830 9580 4010 9640
rect 4330 9270 4390 9330
rect 4710 9750 6210 9810
rect 4710 9580 4890 9640
rect 5370 9580 5550 9640
rect 6030 9580 6210 9640
rect 6530 9270 6590 9330
rect 6910 9750 8410 9810
rect 6910 9440 7090 9500
rect 7570 9440 7750 9500
rect 8230 9440 8410 9500
rect 8730 9270 8790 9330
rect 9110 9750 10610 9810
rect 9110 9440 9290 9500
rect 9770 9440 9950 9500
rect 10430 9440 10610 9500
rect 10930 9270 10990 9330
rect 11310 9750 12810 9810
rect 11310 9440 11490 9500
rect 11970 9440 12150 9500
rect 12630 9440 12810 9500
rect 13130 9270 13190 9330
rect 13510 9750 15010 9810
rect 13510 9440 13690 9500
rect 14170 9440 14350 9500
rect 14830 9440 15010 9500
rect 15330 9270 15390 9330
rect 15710 9750 17210 9810
rect 15710 9580 15890 9640
rect 16370 9580 16550 9640
rect 17030 9580 17210 9640
rect 17530 9270 17590 9330
rect 17910 9750 19410 9810
rect 17910 9580 18090 9640
rect 18570 9580 18750 9640
rect 19230 9580 19410 9640
rect 430 8910 610 8990
rect 430 8110 610 8190
rect 430 7310 610 7390
rect 19730 9270 19790 9330
rect 2130 8470 2190 8530
rect 2510 8640 2690 8700
rect 3170 8640 3350 8700
rect 3830 8640 4010 8700
rect 4330 8470 4390 8530
rect 4710 8950 6210 9010
rect 4710 8640 4890 8700
rect 5370 8640 5550 8700
rect 6030 8640 6210 8700
rect 6530 8470 6590 8530
rect 6910 8950 8410 9010
rect 6910 8780 7090 8840
rect 7570 8780 7750 8840
rect 8230 8780 8410 8840
rect 8730 8470 8790 8530
rect 9110 8950 10610 9010
rect 9110 8780 9290 8840
rect 9770 8780 9950 8840
rect 10430 8780 10610 8840
rect 10930 8470 10990 8530
rect 11310 8950 12810 9010
rect 11310 8780 11490 8840
rect 11970 8780 12150 8840
rect 12630 8780 12810 8840
rect 13130 8470 13190 8530
rect 13510 8950 15010 9010
rect 13510 8780 13690 8840
rect 14170 8780 14350 8840
rect 14830 8780 15010 8840
rect 15330 8470 15390 8530
rect 15710 8950 17210 9010
rect 15710 8640 15890 8700
rect 16370 8640 16550 8700
rect 17030 8640 17210 8700
rect 17530 8470 17590 8530
rect 17910 8640 18090 8700
rect 18570 8640 18750 8700
rect 19230 8640 19410 8700
rect 19730 8470 19790 8530
rect 2130 7670 2190 7730
rect 2510 7840 2690 7900
rect 3170 7840 3350 7900
rect 3830 7840 4010 7900
rect 4330 7670 4390 7730
rect 4710 8150 6210 8210
rect 4710 7840 4890 7900
rect 5370 7840 5550 7900
rect 6030 7840 6210 7900
rect 6530 7670 6590 7730
rect 6910 8150 8410 8210
rect 6910 7980 7090 8040
rect 7570 7980 7750 8040
rect 8230 7980 8410 8040
rect 8730 7670 8790 7730
rect 9110 8150 10610 8210
rect 9110 7980 9290 8040
rect 9770 7980 9950 8040
rect 10430 7980 10610 8040
rect 10930 7670 10990 7730
rect 11310 8150 12810 8210
rect 11310 7980 11490 8040
rect 11970 7980 12150 8040
rect 12630 7980 12810 8040
rect 13130 7670 13190 7730
rect 13510 8150 15010 8210
rect 13510 7980 13690 8040
rect 14170 7980 14350 8040
rect 14830 7980 15010 8040
rect 15330 7670 15390 7730
rect 15710 8150 17210 8210
rect 15710 7840 15890 7900
rect 16370 7840 16550 7900
rect 17030 7840 17210 7900
rect 17530 7670 17590 7730
rect 17910 7840 18090 7900
rect 18570 7840 18750 7900
rect 19230 7840 19410 7900
rect 430 6510 610 6590
rect 1290 4350 1470 4530
rect 19730 7670 19790 7730
rect 2130 6870 2190 6930
rect 2510 7180 2690 7240
rect 3170 7180 3350 7240
rect 3830 7180 4010 7240
rect 4330 6870 4390 6930
rect 4710 7350 6210 7410
rect 4710 7180 4890 7240
rect 5370 7180 5550 7240
rect 6030 7180 6210 7240
rect 6530 6870 6590 6930
rect 6910 7350 8410 7410
rect 6910 7040 7090 7100
rect 7570 7040 7750 7100
rect 8230 7040 8410 7100
rect 8730 6870 8790 6930
rect 9110 7350 10610 7410
rect 9110 7040 9290 7100
rect 9770 7040 9950 7100
rect 10430 7040 10610 7100
rect 10930 6870 10990 6930
rect 11310 7350 12810 7410
rect 11310 7040 11490 7100
rect 11970 7040 12150 7100
rect 12630 7040 12810 7100
rect 13130 6870 13190 6930
rect 13510 7350 15010 7410
rect 13510 7040 13690 7100
rect 14170 7040 14350 7100
rect 14830 7040 15010 7100
rect 15330 6870 15390 6930
rect 15710 7350 17210 7410
rect 15710 7180 15890 7240
rect 16370 7180 16550 7240
rect 17030 7180 17210 7240
rect 17530 6870 17590 6930
rect 17910 7180 18090 7240
rect 18570 7180 18750 7240
rect 19230 7180 19410 7240
rect 19730 6870 19790 6930
rect 21930 9270 21990 9330
rect 21310 8910 21490 8990
rect 21930 8470 21990 8530
rect 21310 8110 21490 8190
rect 21930 7670 21990 7730
rect 2130 6070 2190 6130
rect 2510 6240 2690 6300
rect 3170 6240 3350 6300
rect 3830 6240 4010 6300
rect 4330 6070 4390 6130
rect 4710 6550 6210 6610
rect 4710 6240 4890 6300
rect 5370 6240 5550 6300
rect 6030 6240 6210 6300
rect 6530 6070 6590 6130
rect 6910 6550 8410 6610
rect 6910 6380 7090 6440
rect 7570 6380 7750 6440
rect 8230 6380 8410 6440
rect 8730 6070 8790 6130
rect 9110 6550 10610 6610
rect 9110 6380 9290 6440
rect 9770 6380 9950 6440
rect 10430 6380 10610 6440
rect 10930 6070 10990 6130
rect 11310 6550 12810 6610
rect 11310 6380 11490 6440
rect 11970 6380 12150 6440
rect 12630 6380 12810 6440
rect 13130 6070 13190 6130
rect 13510 6550 15010 6610
rect 13510 6380 13690 6440
rect 14170 6380 14350 6440
rect 14830 6380 15010 6440
rect 15330 6070 15390 6130
rect 15710 6550 17210 6610
rect 15710 6240 15890 6300
rect 16370 6240 16550 6300
rect 17030 6240 17210 6300
rect 17530 6070 17590 6130
rect 17910 6240 18090 6300
rect 18570 6240 18750 6300
rect 19230 6240 19410 6300
rect 19730 6070 19790 6130
rect 2130 5270 2190 5330
rect 2510 5750 4010 5810
rect 2510 5580 2690 5640
rect 3170 5580 3350 5640
rect 3830 5580 4010 5640
rect 4330 5270 4390 5330
rect 4710 5750 6210 5810
rect 4710 5580 4890 5640
rect 5370 5580 5550 5640
rect 6030 5580 6210 5640
rect 6530 5270 6590 5330
rect 6910 5750 8410 5810
rect 6910 5440 7090 5500
rect 7570 5440 7750 5500
rect 8230 5440 8410 5500
rect 8730 5270 8790 5330
rect 9110 5750 10610 5810
rect 9110 5440 9290 5500
rect 9770 5440 9950 5500
rect 10430 5440 10610 5500
rect 10930 5270 10990 5330
rect 11310 5750 12810 5810
rect 11310 5440 11490 5500
rect 11970 5440 12150 5500
rect 12630 5440 12810 5500
rect 13130 5270 13190 5330
rect 13510 5750 15010 5810
rect 13510 5440 13690 5500
rect 14170 5440 14350 5500
rect 14830 5440 15010 5500
rect 15330 5270 15390 5330
rect 15710 5750 17210 5810
rect 15710 5580 15890 5640
rect 16370 5580 16550 5640
rect 17030 5580 17210 5640
rect 17530 5270 17590 5330
rect 17910 5750 19410 5810
rect 17910 5580 18090 5640
rect 18570 5580 18750 5640
rect 19230 5580 19410 5640
rect 19730 5270 19790 5330
rect 2510 4950 4010 5010
rect 4710 4950 6210 5010
rect 6910 4950 8410 5010
rect 1630 3950 1810 4130
rect 1170 3150 1330 3330
rect 2770 3150 2930 3330
rect 4370 3150 4530 3330
rect 5970 3150 6130 3330
rect 7570 3150 7730 3330
rect 480 -4780 660 2220
rect 2110 2090 2230 2250
rect 3710 2090 3830 2250
rect 2110 290 2230 450
rect 5310 2090 5430 2250
rect 3710 290 3830 450
rect 2110 -1510 2230 -1350
rect 6910 2090 7030 2250
rect 5310 290 5430 450
rect 3710 -1510 3830 -1350
rect 2110 -3310 2230 -3150
rect 9110 4950 10610 5010
rect 11310 4950 12810 5010
rect 13510 4950 15010 5010
rect 15710 4950 17210 5010
rect 17910 4950 19410 5010
rect 20110 4350 20290 4530
rect 21310 7310 21490 7390
rect 21930 6870 21990 6930
rect 21310 6510 21490 6590
rect 21930 6070 21990 6130
rect 21930 5270 21990 5330
rect 23050 4710 23580 4970
rect 20450 3950 20630 4130
rect 9170 3150 9330 3330
rect 7810 2810 7930 2930
rect 8510 2090 8630 2250
rect 6910 290 7030 450
rect 5310 -1510 5430 -1350
rect 3710 -3310 3830 -3150
rect 28780 11040 28840 11260
rect 29280 11120 29510 11190
rect 28960 10970 29190 11040
rect 28870 10710 28930 10880
rect 29020 10570 29080 10740
rect 27250 4750 27430 4930
rect 27370 4350 27550 4530
rect 29140 4290 29200 4520
rect 31290 11110 31530 11200
rect 30300 10080 30400 10180
rect 33490 10970 33730 11060
rect 32380 9900 32480 10000
rect 35700 10900 35940 10920
rect 35700 10830 35878 10900
rect 35878 10830 35936 10900
rect 35936 10830 35940 10900
rect 36480 11510 36810 11980
rect 36090 10650 36148 10740
rect 36148 10650 36330 10740
rect 34560 9720 34660 9820
rect 31460 9220 31670 9410
rect 31450 8780 31680 8990
rect 30040 5070 30320 5170
rect 29770 4640 30550 4710
rect 29280 4190 29510 4260
rect 27630 3950 27810 4130
rect 30080 3860 30260 4040
rect 31680 3860 31860 4040
rect 34750 7960 34890 8180
rect 35170 7760 35310 7980
rect 36230 6080 36410 6260
rect 36530 6080 36710 6260
rect 32560 5280 32620 5510
rect 33330 5020 33630 5290
rect 36300 5300 36390 5370
rect 36300 5110 36390 5300
rect 36300 5040 36390 5110
rect 32410 4650 32470 4880
rect 32500 4340 32640 4480
rect 34090 4340 34230 4480
rect 31530 3550 31690 3730
rect 32080 3610 32210 3740
rect 26620 3220 26760 3360
rect 10890 2870 11030 3010
rect 14190 2870 14350 3030
rect 18060 2870 18200 3010
rect 23220 2910 23400 3090
rect 11700 2620 11840 2770
rect 11000 2400 11140 2540
rect 10110 2090 10230 2250
rect 12600 2400 12740 2540
rect 13980 2400 14120 2540
rect 11710 2090 11830 2250
rect 8510 290 8630 450
rect 6910 -1510 7030 -1350
rect 5310 -3310 5430 -3150
rect 13310 2090 13430 2250
rect 10110 290 10230 450
rect 8510 -1510 8630 -1350
rect 6910 -3310 7030 -3150
rect 11710 290 11830 450
rect 10110 -1510 10230 -1350
rect 8510 -3310 8630 -3150
rect 13310 290 13430 450
rect 11710 -1510 11830 -1350
rect 10110 -3310 10230 -3150
rect 12880 -1260 13240 -1110
rect 13310 -1510 13430 -1350
rect 11710 -3310 11830 -3150
rect 16910 2640 17130 2780
rect 17380 2640 17490 2780
rect 17740 2640 17960 2780
rect 16510 2090 16630 2250
rect 14910 1320 15030 1980
rect 18110 2090 18230 2250
rect 19710 2090 19830 2250
rect 21310 2090 21430 2250
rect 22910 2090 23030 2250
rect 24510 2090 24630 2250
rect 26110 2090 26230 2250
rect 27710 2070 27830 2250
rect 29310 2070 29430 2250
rect 14910 -1510 15030 -1350
rect 15250 -1510 15370 -1350
rect 13310 -3310 13430 -3150
rect 16510 290 16630 450
rect 7810 -7990 7930 -7870
rect 490 -22380 670 -8090
rect 2130 -9750 2230 -9590
rect 2130 -11550 2230 -11390
rect 3730 -9750 3830 -9590
rect 2130 -13350 2230 -13190
rect 3730 -11550 3830 -11390
rect 2130 -15150 2230 -14990
rect 5330 -9750 5430 -9590
rect 3730 -13350 3830 -13190
rect 2130 -16950 2230 -16790
rect 5330 -11550 5430 -11390
rect 3730 -15150 3830 -14990
rect 2130 -18750 2230 -18590
rect 6930 -9750 7030 -9590
rect 5330 -13350 5430 -13190
rect 3730 -16950 3830 -16790
rect 2130 -20550 2230 -20390
rect 6930 -11550 7030 -11390
rect 5330 -15150 5430 -14990
rect 3730 -18750 3830 -18590
rect 2130 -22350 2230 -22190
rect 8530 -9750 8630 -9590
rect 6930 -13350 7030 -13190
rect 5330 -16950 5430 -16790
rect 3730 -20550 3830 -20390
rect 10810 -8380 10930 -8260
rect 8530 -11550 8630 -11390
rect 6930 -15150 7030 -14990
rect 5330 -18750 5430 -18590
rect 3730 -22350 3830 -22190
rect 10130 -9750 10230 -9590
rect 8530 -13350 8630 -13190
rect 6930 -16950 7030 -16790
rect 5330 -20550 5430 -20390
rect 10130 -11550 10230 -11390
rect 8530 -15150 8630 -14990
rect 6930 -18750 7030 -18590
rect 5330 -22350 5430 -22190
rect 10130 -13350 10230 -13190
rect 8530 -16950 8630 -16790
rect 6930 -20550 7030 -20390
rect 10130 -15150 10230 -14990
rect 8530 -18750 8630 -18590
rect 6930 -22350 7030 -22190
rect 10130 -16950 10230 -16790
rect 8530 -20550 8630 -20390
rect 10130 -18750 10230 -18590
rect 8530 -22350 8630 -22190
rect 10130 -20550 10230 -20390
rect 12950 -6990 13110 -6830
rect 14910 -3310 15030 -3150
rect 16510 -1510 16630 -1350
rect 13310 -8380 13440 -8260
rect 13290 -13330 13460 -13170
rect 18110 290 18230 450
rect 16510 -3310 16630 -3150
rect 15570 -5350 15730 -5170
rect 15570 -5750 15730 -5570
rect 14910 -6610 15030 -6490
rect 13290 -15130 13460 -14970
rect 13300 -16950 13450 -16790
rect 13300 -18750 13450 -18590
rect 15790 -6150 15950 -5970
rect 18110 -1510 18230 -1350
rect 19710 290 19830 450
rect 18110 -3310 18230 -3150
rect 19710 -1510 19830 -1350
rect 21310 290 21430 450
rect 19710 -3310 19830 -3150
rect 21310 -1510 21430 -1350
rect 18770 -5350 18930 -5170
rect 18770 -5750 18930 -5570
rect 17390 -6950 17550 -6770
rect 17170 -7350 17330 -7170
rect 17170 -7750 17330 -7570
rect 16510 -8380 16640 -8260
rect 16510 -9730 16640 -9570
rect 18990 -6150 19150 -5970
rect 22910 290 23030 450
rect 21310 -3310 21430 -3150
rect 22910 -1510 23030 -1350
rect 24510 290 24630 450
rect 22910 -3310 23030 -3150
rect 24510 -1510 24630 -1350
rect 21970 -5350 22130 -5170
rect 21970 -5750 22130 -5570
rect 20590 -6950 20750 -6770
rect 20370 -7350 20530 -7170
rect 20370 -7750 20530 -7570
rect 18110 -9730 18240 -9570
rect 16510 -11530 16640 -11370
rect 14890 -13330 15060 -13170
rect 19710 -9730 19840 -9570
rect 18110 -11530 18240 -11370
rect 16510 -13330 16640 -13170
rect 14890 -15130 15060 -14970
rect 22190 -6150 22350 -5970
rect 24510 -3310 24630 -3150
rect 26110 290 26230 450
rect 26110 -1510 26230 -1350
rect 27710 270 27830 450
rect 26110 -3310 26230 -3150
rect 27710 -1530 27830 -1350
rect 25170 -5350 25330 -5170
rect 25170 -5750 25330 -5570
rect 23790 -6950 23950 -6770
rect 23570 -7350 23730 -7170
rect 23570 -7750 23730 -7570
rect 21310 -9730 21440 -9570
rect 19710 -11530 19840 -11370
rect 18110 -13330 18240 -13170
rect 16510 -15130 16640 -14970
rect 14900 -16950 15050 -16790
rect 22910 -9730 23040 -9570
rect 21310 -11530 21440 -11370
rect 19710 -13330 19840 -13170
rect 18110 -15130 18240 -14970
rect 16510 -16930 16640 -16770
rect 14900 -18750 15050 -18590
rect 25390 -6150 25550 -5970
rect 29310 270 29430 450
rect 27710 -3330 27830 -3150
rect 29310 -1530 29430 -1350
rect 30910 2070 31030 2250
rect 30910 270 31030 450
rect 33130 4070 33290 4110
rect 33130 4010 33290 4070
rect 31830 2910 31990 3090
rect 33180 2390 33330 2550
rect 32510 1030 32630 1150
rect 33180 280 33330 440
rect 32510 -490 32630 190
rect 30910 -1530 31030 -1350
rect 35700 4150 35840 4290
rect 34870 4010 35190 4090
rect 34780 2620 34930 2780
rect 34110 1030 34230 1150
rect 34790 1030 34920 1150
rect 34110 -490 34230 190
rect 29310 -3330 29430 -3150
rect 28370 -5350 28530 -5170
rect 28370 -5750 28530 -5570
rect 27690 -6150 27850 -5970
rect 26990 -6950 27150 -6770
rect 26770 -7350 26930 -7170
rect 26770 -7750 26930 -7570
rect 24510 -9730 24640 -9570
rect 22910 -11530 23040 -11370
rect 21310 -13330 21440 -13170
rect 19710 -15130 19840 -14970
rect 18110 -16930 18240 -16770
rect 16510 -18730 16640 -18570
rect 10130 -22350 10230 -22190
rect 10110 -22590 10250 -22450
rect 11050 -22850 11150 -22740
rect 11720 -22850 11820 -22740
rect 26110 -9730 26240 -9570
rect 24510 -11530 24640 -11370
rect 22910 -13330 23040 -13170
rect 21310 -15130 21440 -14970
rect 19710 -16930 19840 -16770
rect 18110 -18730 18240 -18570
rect 16510 -20530 16640 -20370
rect 28590 -6150 28750 -5970
rect 29290 -6150 29450 -5970
rect 30910 -3330 31030 -3150
rect 32510 -2570 32630 -2450
rect 37680 5300 37770 5370
rect 37680 5110 37770 5300
rect 37680 5040 37770 5110
rect 37880 3580 38010 3710
rect 35710 1030 35830 1150
rect 35710 -490 35830 190
rect 34110 -2570 34230 -2450
rect 34790 -2570 34920 -2450
rect 35710 -2570 35830 -2450
rect 36590 3220 36730 3360
rect 37310 1030 37430 1150
rect 30890 -6150 31050 -5970
rect 30190 -6950 30350 -6770
rect 29970 -7350 30130 -7170
rect 29970 -7750 30130 -7570
rect 27710 -9730 27840 -9570
rect 26110 -11530 26240 -11370
rect 24510 -13330 24640 -13170
rect 22910 -15130 23040 -14970
rect 21310 -16930 21440 -16770
rect 19710 -18730 19840 -18570
rect 18110 -20530 18240 -20370
rect 29310 -9730 29440 -9570
rect 27710 -11530 27840 -11370
rect 26110 -13330 26240 -13170
rect 24510 -15130 24640 -14970
rect 22910 -16930 23040 -16770
rect 21310 -18730 21440 -18570
rect 19710 -20530 19840 -20370
rect 30910 -9730 31040 -9570
rect 29310 -11530 29440 -11370
rect 27710 -13330 27840 -13170
rect 26110 -15130 26240 -14970
rect 32510 -9730 32640 -9570
rect 30910 -11530 31040 -11370
rect 29310 -13330 29440 -13170
rect 27710 -15130 27840 -14970
rect 24510 -16930 24640 -16770
rect 26110 -16930 26240 -16770
rect 22910 -18730 23040 -18570
rect 21310 -20530 21440 -20370
rect 32510 -11530 32640 -11370
rect 30910 -13330 31040 -13170
rect 29310 -15130 29440 -14970
rect 27710 -16930 27840 -16770
rect 24510 -18730 24640 -18570
rect 26110 -18730 26240 -18570
rect 22910 -20530 23040 -20370
rect 29310 -16930 29440 -16770
rect 27710 -18730 27840 -18570
rect 24510 -20530 24640 -20370
rect 26110 -20530 26240 -20370
rect 29310 -18730 29440 -18570
rect 27710 -20530 27840 -20370
rect 29310 -20530 29440 -20370
rect 32510 -13330 32640 -13170
rect 30910 -15130 31040 -14970
rect 30910 -16930 31040 -16770
rect 32520 -16920 32630 -16770
rect 30910 -18730 31040 -18570
rect 30910 -20530 31040 -20370
rect 16510 -22330 16640 -22170
rect 18110 -22330 18240 -22170
rect 19710 -22330 19840 -22170
rect 21310 -22330 21440 -22170
rect 22910 -22330 23040 -22170
rect 24510 -22330 24640 -22170
rect 26110 -22330 26240 -22170
rect 27710 -22330 27840 -22170
rect 29310 -22330 29440 -22170
rect 30910 -22330 31040 -22170
rect 27720 -22850 27830 -22740
rect 28150 -22870 28370 -22730
rect 28630 -22870 28740 -22740
rect 29000 -22870 29220 -22730
rect 29320 -22850 29430 -22740
rect 30920 -22850 31030 -22740
rect 12420 -23090 12520 -22980
rect 26530 -23160 26710 -22980
rect 1190 -23450 1350 -23270
rect 2790 -23450 2950 -23270
rect 4390 -23450 4550 -23270
rect 5990 -23450 6150 -23270
rect 7590 -23450 7750 -23270
rect 9190 -23450 9350 -23270
rect 23210 -23480 23390 -23300
rect 1630 -24250 1810 -24070
rect 1290 -24650 1470 -24470
rect 430 -26710 610 -26630
rect 430 -27510 610 -27430
rect 430 -28310 610 -28230
rect 430 -29110 610 -29030
rect 2510 -25130 4010 -25070
rect 4710 -25130 6210 -25070
rect 6910 -25130 8410 -25070
rect 9110 -25130 10610 -25070
rect 11310 -25130 12810 -25070
rect 13510 -25130 15010 -25070
rect 15710 -25130 17210 -25070
rect 17910 -25130 19410 -25070
rect 20450 -24250 20630 -24070
rect 20110 -24650 20290 -24470
rect 2510 -25760 2690 -25700
rect 3170 -25760 3350 -25700
rect 3830 -25760 4010 -25700
rect 2510 -25930 4010 -25870
rect 4710 -25760 4890 -25700
rect 5370 -25760 5550 -25700
rect 6030 -25760 6210 -25700
rect 4710 -25930 6210 -25870
rect 6910 -25620 7090 -25560
rect 7570 -25620 7750 -25560
rect 8230 -25620 8410 -25560
rect 6910 -25930 8410 -25870
rect 9110 -25620 9290 -25560
rect 9770 -25620 9950 -25560
rect 10430 -25620 10610 -25560
rect 9110 -25930 10610 -25870
rect 11310 -25620 11490 -25560
rect 11970 -25620 12150 -25560
rect 12630 -25620 12810 -25560
rect 11310 -25930 12810 -25870
rect 13510 -25620 13690 -25560
rect 14170 -25620 14350 -25560
rect 14830 -25620 15010 -25560
rect 13510 -25930 15010 -25870
rect 15710 -25760 15890 -25700
rect 16370 -25760 16550 -25700
rect 17030 -25760 17210 -25700
rect 15710 -25930 17210 -25870
rect 17910 -25760 18090 -25700
rect 18570 -25760 18750 -25700
rect 19230 -25760 19410 -25700
rect 17910 -25930 19410 -25870
rect 2510 -26420 2690 -26360
rect 3170 -26420 3350 -26360
rect 3830 -26420 4010 -26360
rect 4710 -26420 4890 -26360
rect 5370 -26420 5550 -26360
rect 6030 -26420 6210 -26360
rect 4710 -26730 6210 -26670
rect 6910 -26560 7090 -26500
rect 7570 -26560 7750 -26500
rect 8230 -26560 8410 -26500
rect 6910 -26730 8410 -26670
rect 9110 -26560 9290 -26500
rect 9770 -26560 9950 -26500
rect 10430 -26560 10610 -26500
rect 9110 -26730 10610 -26670
rect 11310 -26560 11490 -26500
rect 11970 -26560 12150 -26500
rect 12630 -26560 12810 -26500
rect 11310 -26730 12810 -26670
rect 13510 -26560 13690 -26500
rect 14170 -26560 14350 -26500
rect 14830 -26560 15010 -26500
rect 13510 -26730 15010 -26670
rect 15710 -26420 15890 -26360
rect 16370 -26420 16550 -26360
rect 17030 -26420 17210 -26360
rect 15710 -26730 17210 -26670
rect 17910 -26420 18090 -26360
rect 18570 -26420 18750 -26360
rect 19230 -26420 19410 -26360
rect 2510 -27360 2690 -27300
rect 3170 -27360 3350 -27300
rect 3830 -27360 4010 -27300
rect 4710 -27360 4890 -27300
rect 5370 -27360 5550 -27300
rect 6030 -27360 6210 -27300
rect 4710 -27530 6210 -27470
rect 6910 -27220 7090 -27160
rect 7570 -27220 7750 -27160
rect 8230 -27220 8410 -27160
rect 6910 -27530 8410 -27470
rect 9110 -27220 9290 -27160
rect 9770 -27220 9950 -27160
rect 10430 -27220 10610 -27160
rect 9110 -27530 10610 -27470
rect 11310 -27220 11490 -27160
rect 11970 -27220 12150 -27160
rect 12630 -27220 12810 -27160
rect 11310 -27530 12810 -27470
rect 13510 -27220 13690 -27160
rect 14170 -27220 14350 -27160
rect 14830 -27220 15010 -27160
rect 13510 -27530 15010 -27470
rect 15710 -27360 15890 -27300
rect 16370 -27360 16550 -27300
rect 17030 -27360 17210 -27300
rect 15710 -27530 17210 -27470
rect 17910 -27360 18090 -27300
rect 18570 -27360 18750 -27300
rect 19230 -27360 19410 -27300
rect 2510 -28020 2690 -27960
rect 3170 -28020 3350 -27960
rect 3830 -28020 4010 -27960
rect 4710 -28020 4890 -27960
rect 5370 -28020 5550 -27960
rect 6030 -28020 6210 -27960
rect 4710 -28330 6210 -28270
rect 6910 -28160 7090 -28100
rect 7570 -28160 7750 -28100
rect 8230 -28160 8410 -28100
rect 6910 -28330 8410 -28270
rect 9110 -28160 9290 -28100
rect 9770 -28160 9950 -28100
rect 10430 -28160 10610 -28100
rect 9110 -28330 10610 -28270
rect 11310 -28160 11490 -28100
rect 11970 -28160 12150 -28100
rect 12630 -28160 12810 -28100
rect 11310 -28330 12810 -28270
rect 13510 -28160 13690 -28100
rect 14170 -28160 14350 -28100
rect 14830 -28160 15010 -28100
rect 13510 -28330 15010 -28270
rect 15710 -28020 15890 -27960
rect 16370 -28020 16550 -27960
rect 17030 -28020 17210 -27960
rect 15710 -28330 17210 -28270
rect 17910 -28020 18090 -27960
rect 18570 -28020 18750 -27960
rect 19230 -28020 19410 -27960
rect 2510 -28820 2690 -28760
rect 3170 -28820 3350 -28760
rect 3830 -28820 4010 -28760
rect 4710 -28820 4890 -28760
rect 5370 -28820 5550 -28760
rect 6030 -28820 6210 -28760
rect 4710 -29130 6210 -29070
rect 6910 -28960 7090 -28900
rect 7570 -28960 7750 -28900
rect 8230 -28960 8410 -28900
rect 6910 -29130 8410 -29070
rect 9110 -28960 9290 -28900
rect 9770 -28960 9950 -28900
rect 10430 -28960 10610 -28900
rect 9110 -29130 10610 -29070
rect 11310 -28960 11490 -28900
rect 11970 -28960 12150 -28900
rect 12630 -28960 12810 -28900
rect 11310 -29130 12810 -29070
rect 13510 -28960 13690 -28900
rect 14170 -28960 14350 -28900
rect 14830 -28960 15010 -28900
rect 13510 -29130 15010 -29070
rect 15710 -28820 15890 -28760
rect 16370 -28820 16550 -28760
rect 17030 -28820 17210 -28760
rect 15710 -29130 17210 -29070
rect 17910 -28820 18090 -28760
rect 18570 -28820 18750 -28760
rect 19230 -28820 19410 -28760
rect 23040 -25070 23560 -24820
rect 31560 -23480 31740 -23300
rect 27630 -24250 27810 -24070
rect 28500 -24200 28660 -24040
rect 27400 -24650 27580 -24470
rect 27250 -25070 27430 -24890
rect 21310 -26710 21490 -26630
rect 21310 -27510 21490 -27430
rect 21310 -28310 21490 -28230
rect 21310 -29110 21490 -29030
rect 2510 -29760 2690 -29700
rect 3170 -29760 3350 -29700
rect 3830 -29760 4010 -29700
rect 2510 -29930 4010 -29870
rect 4710 -29760 4890 -29700
rect 5370 -29760 5550 -29700
rect 6030 -29760 6210 -29700
rect 4710 -29930 6210 -29870
rect 6910 -29620 7090 -29560
rect 7570 -29620 7750 -29560
rect 8230 -29620 8410 -29560
rect 6910 -29930 8410 -29870
rect 9110 -29620 9290 -29560
rect 9770 -29620 9950 -29560
rect 10430 -29620 10610 -29560
rect 9110 -29930 10610 -29870
rect 11310 -29620 11490 -29560
rect 11970 -29620 12150 -29560
rect 12630 -29620 12810 -29560
rect 11310 -29930 12810 -29870
rect 13510 -29620 13690 -29560
rect 14170 -29620 14350 -29560
rect 14830 -29620 15010 -29560
rect 13510 -29930 15010 -29870
rect 15710 -29760 15890 -29700
rect 16370 -29760 16550 -29700
rect 17030 -29760 17210 -29700
rect 15710 -29930 17210 -29870
rect 17910 -29760 18090 -29700
rect 18570 -29760 18750 -29700
rect 19230 -29760 19410 -29700
rect 17910 -29930 19410 -29870
rect 2510 -30420 2690 -30360
rect 3170 -30420 3350 -30360
rect 3830 -30420 4010 -30360
rect 2510 -30730 4010 -30670
rect 4710 -30420 4890 -30360
rect 5370 -30420 5550 -30360
rect 6030 -30420 6210 -30360
rect 4710 -30730 6210 -30670
rect 6910 -30560 7090 -30500
rect 7570 -30560 7750 -30500
rect 8230 -30560 8410 -30500
rect 6910 -30730 8410 -30670
rect 9110 -30560 9290 -30500
rect 9770 -30560 9950 -30500
rect 10430 -30560 10610 -30500
rect 9110 -30730 10610 -30670
rect 11310 -30560 11490 -30500
rect 11970 -30560 12150 -30500
rect 12630 -30560 12810 -30500
rect 11310 -30730 12810 -30670
rect 13510 -30560 13690 -30500
rect 14170 -30560 14350 -30500
rect 14830 -30560 15010 -30500
rect 13510 -30730 15010 -30670
rect 15710 -30420 15890 -30360
rect 16370 -30420 16550 -30360
rect 17030 -30420 17210 -30360
rect 15710 -30730 17210 -30670
rect 17910 -30420 18090 -30360
rect 18570 -30420 18750 -30360
rect 19230 -30420 19410 -30360
rect 17910 -30730 19410 -30670
rect 90 -32110 270 -31730
rect 1990 -31830 2110 -31710
rect 2510 -31360 2690 -31300
rect 3170 -31360 3350 -31300
rect 3830 -31360 4010 -31300
rect 4190 -31830 4310 -31710
rect 2210 -32130 2330 -32010
rect 4710 -31360 4890 -31300
rect 5370 -31360 5550 -31300
rect 6030 -31360 6210 -31300
rect 6390 -31830 6510 -31710
rect 4410 -32130 4530 -32010
rect 6910 -31220 7090 -31160
rect 7570 -31220 7750 -31160
rect 8230 -31220 8410 -31160
rect 8590 -31830 8710 -31710
rect 6610 -32130 6730 -32010
rect 9110 -31220 9290 -31160
rect 9770 -31220 9950 -31160
rect 10430 -31220 10610 -31160
rect 10790 -31830 10910 -31710
rect 8810 -32130 8930 -32010
rect 11310 -31220 11490 -31160
rect 11970 -31220 12150 -31160
rect 12630 -31220 12810 -31160
rect 12990 -31830 13110 -31710
rect 11010 -32130 11130 -32010
rect 13510 -31220 13690 -31160
rect 14170 -31220 14350 -31160
rect 14830 -31220 15010 -31160
rect 15190 -31830 15310 -31710
rect 13210 -32130 13330 -32010
rect 15710 -31360 15890 -31300
rect 16370 -31360 16550 -31300
rect 17030 -31360 17210 -31300
rect 17390 -31830 17510 -31710
rect 15410 -32130 15530 -32010
rect 17910 -31360 18090 -31300
rect 18570 -31360 18750 -31300
rect 19230 -31360 19410 -31300
rect 19590 -31830 19710 -31710
rect 17610 -32130 17730 -32010
rect 29380 -24720 29440 -24490
rect 29530 -24870 29590 -24640
rect 28940 -30880 29160 -30810
rect 29070 -31030 29290 -30960
rect 29220 -31180 29440 -31110
rect 29680 -28940 29740 -28720
rect 32510 -20530 32640 -20370
rect 31820 -23850 32000 -23670
rect 29980 -24370 30040 -24140
rect 29830 -29090 29890 -28870
rect 34110 -9730 34240 -9570
rect 35710 -9730 35840 -9570
rect 34110 -11530 34240 -11370
rect 34110 -13330 34240 -13170
rect 35710 -11530 35840 -11370
rect 34120 -16920 34230 -16770
rect 34110 -20530 34240 -20370
rect 32800 -24550 33030 -24480
rect 35710 -13330 35840 -13170
rect 34620 -24280 34770 -24220
rect 35720 -16920 35830 -16770
rect 35710 -20530 35840 -20370
rect 34990 -24280 35130 -24220
rect 35130 -24280 35260 -24220
rect 35260 -24280 35450 -24220
rect 35450 -24280 35570 -24220
rect 35570 -24280 35760 -24220
rect 35760 -24280 35890 -24220
rect 35890 -24280 36080 -24220
rect 36080 -24280 36200 -24220
rect 36200 -24280 36390 -24220
rect 36390 -24280 36520 -24220
rect 36520 -24280 36710 -24220
rect 36710 -24280 36830 -24220
rect 36830 -24280 37020 -24220
rect 34120 -24700 34350 -24630
rect 30290 -24850 30510 -24780
rect 33560 -24850 33790 -24780
rect 34810 -24860 34900 -24660
rect 37130 -24780 37270 -24640
rect 30130 -25170 30190 -24940
rect 29980 -29240 30040 -29020
rect 30130 -29390 30190 -29170
rect 30430 -25320 30490 -25090
rect 30280 -29540 30340 -29320
rect 36030 -27140 36410 -27010
rect 36530 -27140 36910 -27010
rect 33440 -27780 33580 -27640
rect 31820 -28290 33160 -28050
rect 31800 -28780 31994 -28710
rect 31994 -28780 32050 -28710
rect 30430 -29690 30490 -29470
rect 32200 -28914 32206 -28860
rect 32206 -28914 32264 -28860
rect 32264 -28914 32450 -28860
rect 32200 -28930 32450 -28914
rect 35640 -27980 35780 -27840
rect 34000 -29080 34250 -29010
rect 34410 -29220 34660 -29150
rect 37740 -28180 37880 -28040
rect 36200 -29380 36450 -29310
rect 36600 -29530 36850 -29460
rect 37250 -30110 37690 -29920
rect 29370 -31330 29590 -31260
rect 32960 -30880 33210 -30810
rect 33330 -31030 33580 -30960
rect 32540 -31950 33690 -31730
rect 35560 -31180 35570 -31110
rect 35570 -31180 35628 -31110
rect 35628 -31180 35810 -31110
rect 37710 -31330 37770 -31260
rect 37770 -31330 37828 -31260
rect 37828 -31330 37960 -31260
rect 19810 -32130 19930 -32010
<< metal3 >>
rect 2200 12010 2340 12020
rect 2200 12000 2210 12010
rect -360 11990 2210 12000
rect -360 11610 -350 11990
rect -170 11900 2210 11990
rect -170 11610 -160 11900
rect 2200 11890 2210 11900
rect 2330 12000 2340 12010
rect 4400 12010 4540 12020
rect 4400 12000 4410 12010
rect 2330 11900 4410 12000
rect 2330 11890 2340 11900
rect 2200 11880 2340 11890
rect 4400 11890 4410 11900
rect 4530 12000 4540 12010
rect 6600 12010 6740 12020
rect 6600 12000 6610 12010
rect 4530 11900 6610 12000
rect 4530 11890 4540 11900
rect 4400 11880 4540 11890
rect 6600 11890 6610 11900
rect 6730 12000 6740 12010
rect 8800 12010 8940 12020
rect 8800 12000 8810 12010
rect 6730 11900 8810 12000
rect 6730 11890 6740 11900
rect 6600 11880 6740 11890
rect 8800 11890 8810 11900
rect 8930 12000 8940 12010
rect 11000 12010 11140 12020
rect 11000 12000 11010 12010
rect 8930 11900 11010 12000
rect 8930 11890 8940 11900
rect 8800 11880 8940 11890
rect 11000 11890 11010 11900
rect 11130 12000 11140 12010
rect 13200 12010 13340 12020
rect 13200 12000 13210 12010
rect 11130 11900 13210 12000
rect 11130 11890 11140 11900
rect 11000 11880 11140 11890
rect 13200 11890 13210 11900
rect 13330 12000 13340 12010
rect 15400 12010 15540 12020
rect 15400 12000 15410 12010
rect 13330 11900 15410 12000
rect 13330 11890 13340 11900
rect 13200 11880 13340 11890
rect 15400 11890 15410 11900
rect 15530 12000 15540 12010
rect 17600 12010 17740 12020
rect 17600 12000 17610 12010
rect 15530 11900 17610 12000
rect 15530 11890 15540 11900
rect 15400 11880 15540 11890
rect 17600 11890 17610 11900
rect 17730 12000 17740 12010
rect 19800 12010 19940 12020
rect 19800 12000 19810 12010
rect 17730 11900 19810 12000
rect 17730 11890 17740 11900
rect 17600 11880 17740 11890
rect 19800 11890 19810 11900
rect 19930 12000 19940 12010
rect 19930 11900 22160 12000
rect 36470 11980 36820 11990
rect 19930 11890 19940 11900
rect 19800 11880 19940 11890
rect 1980 11710 2120 11720
rect 1980 11700 1990 11710
rect -360 11600 -160 11610
rect 80 11690 1990 11700
rect 80 11310 90 11690
rect 270 11600 1990 11690
rect 270 11310 280 11600
rect 1980 11590 1990 11600
rect 2110 11700 2120 11710
rect 4180 11710 4320 11720
rect 4180 11700 4190 11710
rect 2110 11600 4190 11700
rect 2110 11590 2120 11600
rect 1980 11580 2120 11590
rect 4180 11590 4190 11600
rect 4310 11700 4320 11710
rect 6380 11710 6520 11720
rect 6380 11700 6390 11710
rect 4310 11600 6390 11700
rect 4310 11590 4320 11600
rect 4180 11580 4320 11590
rect 6380 11590 6390 11600
rect 6510 11700 6520 11710
rect 8580 11710 8720 11720
rect 8580 11700 8590 11710
rect 6510 11600 8590 11700
rect 6510 11590 6520 11600
rect 6380 11580 6520 11590
rect 8580 11590 8590 11600
rect 8710 11700 8720 11710
rect 10780 11710 10920 11720
rect 10780 11700 10790 11710
rect 8710 11600 10790 11700
rect 8710 11590 8720 11600
rect 8580 11580 8720 11590
rect 10780 11590 10790 11600
rect 10910 11700 10920 11710
rect 12980 11710 13120 11720
rect 12980 11700 12990 11710
rect 10910 11600 12990 11700
rect 10910 11590 10920 11600
rect 10780 11580 10920 11590
rect 12980 11590 12990 11600
rect 13110 11700 13120 11710
rect 15180 11710 15320 11720
rect 15180 11700 15190 11710
rect 13110 11600 15190 11700
rect 13110 11590 13120 11600
rect 12980 11580 13120 11590
rect 15180 11590 15190 11600
rect 15310 11700 15320 11710
rect 17380 11710 17520 11720
rect 17380 11700 17390 11710
rect 15310 11600 17390 11700
rect 15310 11590 15320 11600
rect 15180 11580 15320 11590
rect 17380 11590 17390 11600
rect 17510 11700 17520 11710
rect 19580 11710 19720 11720
rect 19580 11700 19590 11710
rect 17510 11600 19590 11700
rect 17510 11590 17520 11600
rect 17380 11580 17520 11590
rect 19580 11590 19590 11600
rect 19710 11700 19720 11710
rect 19710 11600 22160 11700
rect 19710 11590 19720 11600
rect 19580 11580 19720 11590
rect 36470 11510 36480 11980
rect 36810 11510 36820 11980
rect 36470 11500 36820 11510
rect 80 11300 280 11310
rect 28770 11260 28850 11270
rect 820 11250 1020 11260
rect 20500 11250 20700 11260
rect 820 11240 830 11250
rect -220 11180 830 11240
rect 820 11170 830 11180
rect 1010 11240 1020 11250
rect 2500 11240 2700 11250
rect 3160 11240 3360 11250
rect 3820 11240 4020 11250
rect 4700 11240 4900 11250
rect 5360 11240 5560 11250
rect 6020 11240 6220 11250
rect 6900 11240 7100 11250
rect 7560 11240 7760 11250
rect 8220 11240 8420 11250
rect 9100 11240 9300 11250
rect 9760 11240 9960 11250
rect 10420 11240 10620 11250
rect 11300 11240 11500 11250
rect 11960 11240 12160 11250
rect 12620 11240 12820 11250
rect 13500 11240 13700 11250
rect 14160 11240 14360 11250
rect 14820 11240 15020 11250
rect 15700 11240 15900 11250
rect 16360 11240 16560 11250
rect 17020 11240 17220 11250
rect 17900 11240 18100 11250
rect 18560 11240 18760 11250
rect 19220 11240 19420 11250
rect 20500 11240 20510 11250
rect 1010 11180 2510 11240
rect 2690 11180 3170 11240
rect 3350 11180 3830 11240
rect 4010 11180 4710 11240
rect 4890 11180 5370 11240
rect 5550 11180 6030 11240
rect 6210 11180 15710 11240
rect 15890 11180 16370 11240
rect 16550 11180 17030 11240
rect 17210 11180 17910 11240
rect 18090 11180 18570 11240
rect 18750 11180 19230 11240
rect 19410 11180 20510 11240
rect 1010 11170 1020 11180
rect 2500 11170 2700 11180
rect 3160 11170 3360 11180
rect 3820 11170 4020 11180
rect 4700 11170 4900 11180
rect 5360 11170 5560 11180
rect 6020 11170 6220 11180
rect 6900 11170 7100 11180
rect 7560 11170 7760 11180
rect 8220 11170 8420 11180
rect 9100 11170 9300 11180
rect 9760 11170 9960 11180
rect 10420 11170 10620 11180
rect 11300 11170 11500 11180
rect 11960 11170 12160 11180
rect 12620 11170 12820 11180
rect 13500 11170 13700 11180
rect 14160 11170 14360 11180
rect 14820 11170 15020 11180
rect 15700 11170 15900 11180
rect 16360 11170 16560 11180
rect 17020 11170 17220 11180
rect 17900 11170 18100 11180
rect 18560 11170 18760 11180
rect 19220 11170 19420 11180
rect 20500 11170 20510 11180
rect 20690 11240 20700 11250
rect 20690 11180 22180 11240
rect 20690 11170 20700 11180
rect 820 11160 1020 11170
rect 20500 11160 20700 11170
rect 1220 11110 1420 11120
rect 20900 11110 21100 11120
rect 1220 11100 1230 11110
rect -220 11040 1230 11100
rect 1220 11030 1230 11040
rect 1410 11100 1420 11110
rect 2500 11100 2700 11110
rect 3160 11100 3360 11110
rect 3820 11100 4020 11110
rect 4700 11100 4900 11110
rect 5360 11100 5560 11110
rect 6020 11100 6220 11110
rect 6900 11100 7100 11110
rect 7560 11100 7760 11110
rect 8220 11100 8420 11110
rect 9100 11100 9300 11110
rect 9760 11100 9960 11110
rect 10420 11100 10620 11110
rect 11300 11100 11500 11110
rect 11960 11100 12160 11110
rect 12620 11100 12820 11110
rect 13500 11100 13700 11110
rect 14160 11100 14360 11110
rect 14820 11100 15020 11110
rect 15700 11100 15900 11110
rect 16360 11100 16560 11110
rect 17020 11100 17220 11110
rect 17900 11100 18100 11110
rect 18560 11100 18760 11110
rect 19220 11100 19420 11110
rect 20900 11100 20910 11110
rect 1410 11040 6910 11100
rect 7090 11040 7570 11100
rect 7750 11040 8230 11100
rect 8410 11040 9110 11100
rect 9290 11040 9770 11100
rect 9950 11040 10430 11100
rect 10610 11040 11310 11100
rect 11490 11040 11970 11100
rect 12150 11040 12630 11100
rect 12810 11040 13510 11100
rect 13690 11040 14170 11100
rect 14350 11040 14830 11100
rect 15010 11040 20910 11100
rect 1410 11030 1420 11040
rect 2500 11030 2700 11040
rect 3160 11030 3360 11040
rect 3820 11030 4020 11040
rect 4700 11030 4900 11040
rect 5360 11030 5560 11040
rect 6020 11030 6220 11040
rect 6900 11030 7100 11040
rect 7560 11030 7760 11040
rect 8220 11030 8420 11040
rect 9100 11030 9300 11040
rect 9760 11030 9960 11040
rect 10420 11030 10620 11040
rect 11300 11030 11500 11040
rect 11960 11030 12160 11040
rect 12620 11030 12820 11040
rect 13500 11030 13700 11040
rect 14160 11030 14360 11040
rect 14820 11030 15020 11040
rect 15700 11030 15900 11040
rect 16360 11030 16560 11040
rect 17020 11030 17220 11040
rect 17900 11030 18100 11040
rect 18560 11030 18760 11040
rect 19220 11030 19420 11040
rect 20900 11030 20910 11040
rect 21090 11100 21100 11110
rect 21090 11040 22180 11100
rect 28770 11040 28780 11260
rect 28840 11190 28850 11260
rect 31280 11200 31540 11210
rect 29270 11190 29520 11200
rect 31280 11190 31290 11200
rect 28840 11120 29280 11190
rect 29510 11120 31290 11190
rect 28840 11040 28850 11120
rect 29270 11110 29520 11120
rect 31280 11110 31290 11120
rect 31530 11110 31540 11200
rect 31280 11100 31540 11110
rect 33480 11060 33740 11070
rect 21090 11030 21100 11040
rect 28770 11030 28850 11040
rect 28950 11040 29200 11050
rect 1220 11020 1420 11030
rect 20900 11020 21100 11030
rect 28950 10970 28960 11040
rect 29190 11030 29200 11040
rect 33480 11030 33490 11060
rect 29190 10970 33490 11030
rect 33730 10970 33740 11060
rect 28950 10960 33740 10970
rect -110 10940 30 10960
rect -110 10690 -80 10940
rect 0 10690 30 10940
rect -110 10660 30 10690
rect 2090 10940 2230 10960
rect 2090 10690 2120 10940
rect 2200 10690 2230 10940
rect 2090 10660 2230 10690
rect 4290 10940 4430 10960
rect 4290 10690 4320 10940
rect 4400 10690 4430 10940
rect 4290 10660 4430 10690
rect 6490 10940 6630 10960
rect 6490 10690 6520 10940
rect 6600 10690 6630 10940
rect 6490 10660 6630 10690
rect 8690 10940 8830 10960
rect 8690 10690 8720 10940
rect 8800 10690 8830 10940
rect 8690 10660 8830 10690
rect 10890 10940 11030 10960
rect 10890 10690 10920 10940
rect 11000 10690 11030 10940
rect 10890 10660 11030 10690
rect 13090 10940 13230 10960
rect 13090 10690 13120 10940
rect 13200 10690 13230 10940
rect 13090 10660 13230 10690
rect 15290 10940 15430 10960
rect 15290 10690 15320 10940
rect 15400 10690 15430 10940
rect 15290 10660 15430 10690
rect 17490 10940 17630 10960
rect 17490 10690 17520 10940
rect 17600 10690 17630 10940
rect 17490 10660 17630 10690
rect 19690 10940 19830 10960
rect 19690 10690 19720 10940
rect 19800 10690 19830 10940
rect 19690 10660 19830 10690
rect 21890 10940 22030 10960
rect 21890 10690 21920 10940
rect 22000 10690 22030 10940
rect 35690 10920 35950 10930
rect 35690 10890 35700 10920
rect 28860 10880 35700 10890
rect 28860 10710 28870 10880
rect 28930 10830 35700 10880
rect 35940 10830 35950 10920
rect 28930 10820 35950 10830
rect 28930 10710 28940 10820
rect 28860 10700 28940 10710
rect 29010 10740 36340 10750
rect 21890 10660 22030 10690
rect 2500 10610 4020 10620
rect 1620 10590 1820 10600
rect 1620 10580 1630 10590
rect 1600 10520 1630 10580
rect 1620 10510 1630 10520
rect 1810 10580 1820 10590
rect 2500 10580 2510 10610
rect 1810 10550 2510 10580
rect 4010 10580 4020 10610
rect 4700 10610 6220 10620
rect 4700 10580 4710 10610
rect 4010 10550 4710 10580
rect 6210 10580 6220 10610
rect 6900 10610 8420 10620
rect 6900 10580 6910 10610
rect 6210 10550 6910 10580
rect 8410 10580 8420 10610
rect 9100 10610 10620 10620
rect 9100 10580 9110 10610
rect 8410 10550 9110 10580
rect 10610 10580 10620 10610
rect 11300 10610 12820 10620
rect 11300 10580 11310 10610
rect 10610 10550 11310 10580
rect 12810 10580 12820 10610
rect 13500 10610 15020 10620
rect 13500 10580 13510 10610
rect 12810 10550 13510 10580
rect 15010 10580 15020 10610
rect 15700 10610 17220 10620
rect 15700 10580 15710 10610
rect 15010 10550 15710 10580
rect 17210 10580 17220 10610
rect 17900 10610 19420 10620
rect 17900 10580 17910 10610
rect 17210 10550 17910 10580
rect 19410 10580 19420 10610
rect 20100 10590 20300 10600
rect 20100 10580 20110 10590
rect 19410 10550 20110 10580
rect 1810 10520 20110 10550
rect 1810 10510 1820 10520
rect 1620 10500 1820 10510
rect 20100 10510 20110 10520
rect 20290 10580 20300 10590
rect 20290 10520 20320 10580
rect 29010 10570 29020 10740
rect 29080 10680 36090 10740
rect 29080 10570 29090 10680
rect 36080 10650 36090 10680
rect 36330 10650 36340 10740
rect 36080 10640 36340 10650
rect 29010 10560 29090 10570
rect 20290 10510 20300 10520
rect 20100 10500 20300 10510
rect 820 10450 1020 10460
rect 20500 10450 20700 10460
rect 820 10440 830 10450
rect -220 10380 830 10440
rect 820 10370 830 10380
rect 1010 10440 1020 10450
rect 2500 10440 2700 10450
rect 3160 10440 3360 10450
rect 3820 10440 4020 10450
rect 4700 10440 4900 10450
rect 5360 10440 5560 10450
rect 6020 10440 6220 10450
rect 6900 10440 7100 10450
rect 7560 10440 7760 10450
rect 8220 10440 8420 10450
rect 9100 10440 9300 10450
rect 9760 10440 9960 10450
rect 10420 10440 10620 10450
rect 11300 10440 11500 10450
rect 11960 10440 12160 10450
rect 12620 10440 12820 10450
rect 13500 10440 13700 10450
rect 14160 10440 14360 10450
rect 14820 10440 15020 10450
rect 15700 10440 15900 10450
rect 16360 10440 16560 10450
rect 17020 10440 17220 10450
rect 17900 10440 18100 10450
rect 18560 10440 18760 10450
rect 19220 10440 19420 10450
rect 20500 10440 20510 10450
rect 1010 10380 6910 10440
rect 7090 10380 7570 10440
rect 7750 10380 8230 10440
rect 8410 10380 9110 10440
rect 9290 10380 9770 10440
rect 9950 10380 10430 10440
rect 10610 10380 11310 10440
rect 11490 10380 11970 10440
rect 12150 10380 12630 10440
rect 12810 10380 13510 10440
rect 13690 10380 14170 10440
rect 14350 10380 14830 10440
rect 15010 10380 20510 10440
rect 1010 10370 1020 10380
rect 2500 10370 2700 10380
rect 3160 10370 3360 10380
rect 3820 10370 4020 10380
rect 4700 10370 4900 10380
rect 5360 10370 5560 10380
rect 6020 10370 6220 10380
rect 6900 10370 7100 10380
rect 7560 10370 7760 10380
rect 8220 10370 8420 10380
rect 9100 10370 9300 10380
rect 9760 10370 9960 10380
rect 10420 10370 10620 10380
rect 11300 10370 11500 10380
rect 11960 10370 12160 10380
rect 12620 10370 12820 10380
rect 13500 10370 13700 10380
rect 14160 10370 14360 10380
rect 14820 10370 15020 10380
rect 15700 10370 15900 10380
rect 16360 10370 16560 10380
rect 17020 10370 17220 10380
rect 17900 10370 18100 10380
rect 18560 10370 18760 10380
rect 19220 10370 19420 10380
rect 20500 10370 20510 10380
rect 20690 10440 20700 10450
rect 20690 10380 22180 10440
rect 20690 10370 20700 10380
rect 820 10360 1020 10370
rect 20500 10360 20700 10370
rect 1220 10310 1420 10320
rect 20900 10310 21100 10320
rect 1220 10300 1230 10310
rect -220 10240 1230 10300
rect 1220 10230 1230 10240
rect 1410 10300 1420 10310
rect 2500 10300 2700 10310
rect 3160 10300 3360 10310
rect 3820 10300 4020 10310
rect 4700 10300 4900 10310
rect 5360 10300 5560 10310
rect 6020 10300 6220 10310
rect 6900 10300 7100 10310
rect 7560 10300 7760 10310
rect 8220 10300 8420 10310
rect 9100 10300 9300 10310
rect 9760 10300 9960 10310
rect 10420 10300 10620 10310
rect 11300 10300 11500 10310
rect 11960 10300 12160 10310
rect 12620 10300 12820 10310
rect 13500 10300 13700 10310
rect 14160 10300 14360 10310
rect 14820 10300 15020 10310
rect 15700 10300 15900 10310
rect 16360 10300 16560 10310
rect 17020 10300 17220 10310
rect 17900 10300 18100 10310
rect 18560 10300 18760 10310
rect 19220 10300 19420 10310
rect 20900 10300 20910 10310
rect 1410 10240 2510 10300
rect 2690 10240 3170 10300
rect 3350 10240 3830 10300
rect 4010 10240 4710 10300
rect 4890 10240 5370 10300
rect 5550 10240 6030 10300
rect 6210 10240 15710 10300
rect 15890 10240 16370 10300
rect 16550 10240 17030 10300
rect 17210 10240 17910 10300
rect 18090 10240 18570 10300
rect 18750 10240 19230 10300
rect 19410 10240 20910 10300
rect 1410 10230 1420 10240
rect 2500 10230 2700 10240
rect 3160 10230 3360 10240
rect 3820 10230 4020 10240
rect 4700 10230 4900 10240
rect 5360 10230 5560 10240
rect 6020 10230 6220 10240
rect 6900 10230 7100 10240
rect 7560 10230 7760 10240
rect 8220 10230 8420 10240
rect 9100 10230 9300 10240
rect 9760 10230 9960 10240
rect 10420 10230 10620 10240
rect 11300 10230 11500 10240
rect 11960 10230 12160 10240
rect 12620 10230 12820 10240
rect 13500 10230 13700 10240
rect 14160 10230 14360 10240
rect 14820 10230 15020 10240
rect 15700 10230 15900 10240
rect 16360 10230 16560 10240
rect 17020 10230 17220 10240
rect 17900 10230 18100 10240
rect 18560 10230 18760 10240
rect 19220 10230 19420 10240
rect 20900 10230 20910 10240
rect 21090 10300 21100 10310
rect 21090 10240 22180 10300
rect 21090 10230 21100 10240
rect 1220 10220 1420 10230
rect 20900 10220 21100 10230
rect 30290 10180 30410 10190
rect -110 10140 30 10160
rect -110 9890 -80 10140
rect 0 9890 30 10140
rect -110 9860 30 9890
rect 2090 10140 2230 10160
rect 2090 9890 2120 10140
rect 2200 9890 2230 10140
rect 2090 9860 2230 9890
rect 4290 10140 4430 10160
rect 4290 9890 4320 10140
rect 4400 9890 4430 10140
rect 4290 9860 4430 9890
rect 6490 10140 6630 10160
rect 6490 9890 6520 10140
rect 6600 9890 6630 10140
rect 6490 9860 6630 9890
rect 8690 10140 8830 10160
rect 8690 9890 8720 10140
rect 8800 9890 8830 10140
rect 8690 9860 8830 9890
rect 10890 10140 11030 10160
rect 10890 9890 10920 10140
rect 11000 9890 11030 10140
rect 10890 9860 11030 9890
rect 13090 10140 13230 10160
rect 13090 9890 13120 10140
rect 13200 9890 13230 10140
rect 13090 9860 13230 9890
rect 15290 10140 15430 10160
rect 15290 9890 15320 10140
rect 15400 9890 15430 10140
rect 15290 9860 15430 9890
rect 17490 10140 17630 10160
rect 17490 9890 17520 10140
rect 17600 9890 17630 10140
rect 17490 9860 17630 9890
rect 19690 10140 19830 10160
rect 19690 9890 19720 10140
rect 19800 9890 19830 10140
rect 19690 9860 19830 9890
rect 21890 10140 22030 10160
rect 21890 9890 21920 10140
rect 22000 9890 22030 10140
rect 30290 10080 30300 10180
rect 30400 10170 30410 10180
rect 30400 10090 37470 10170
rect 30400 10080 30410 10090
rect 30290 10070 30410 10080
rect 32370 10000 32490 10010
rect 32370 9900 32380 10000
rect 32480 9990 32490 10000
rect 32480 9910 37470 9990
rect 32480 9900 32490 9910
rect 32370 9890 32490 9900
rect 21890 9860 22030 9890
rect 34550 9820 34670 9830
rect 2500 9810 4020 9820
rect 1620 9790 1820 9800
rect 1620 9780 1630 9790
rect 1600 9720 1630 9780
rect 1620 9710 1630 9720
rect 1810 9780 1820 9790
rect 2500 9780 2510 9810
rect 1810 9750 2510 9780
rect 4010 9780 4020 9810
rect 4700 9810 6220 9820
rect 4700 9780 4710 9810
rect 4010 9750 4710 9780
rect 6210 9780 6220 9810
rect 6900 9810 8420 9820
rect 6900 9780 6910 9810
rect 6210 9750 6910 9780
rect 8410 9780 8420 9810
rect 9100 9810 10620 9820
rect 9100 9780 9110 9810
rect 8410 9750 9110 9780
rect 10610 9780 10620 9810
rect 11300 9810 12820 9820
rect 11300 9780 11310 9810
rect 10610 9750 11310 9780
rect 12810 9780 12820 9810
rect 13500 9810 15020 9820
rect 13500 9780 13510 9810
rect 12810 9750 13510 9780
rect 15010 9780 15020 9810
rect 15700 9810 17220 9820
rect 15700 9780 15710 9810
rect 15010 9750 15710 9780
rect 17210 9780 17220 9810
rect 17900 9810 19420 9820
rect 17900 9780 17910 9810
rect 17210 9750 17910 9780
rect 19410 9780 19420 9810
rect 20100 9790 20300 9800
rect 20100 9780 20110 9790
rect 19410 9750 20110 9780
rect 1810 9720 20110 9750
rect 1810 9710 1820 9720
rect 1620 9700 1820 9710
rect 20100 9710 20110 9720
rect 20290 9780 20300 9790
rect 20290 9720 20320 9780
rect 34550 9720 34560 9820
rect 34660 9810 34670 9820
rect 34660 9730 37470 9810
rect 34660 9720 34670 9730
rect 20290 9710 20300 9720
rect 34550 9710 34670 9720
rect 20100 9700 20300 9710
rect 820 9650 1020 9660
rect 20500 9650 20700 9660
rect 820 9640 830 9650
rect -220 9580 830 9640
rect 820 9570 830 9580
rect 1010 9640 1020 9650
rect 2500 9640 2700 9650
rect 3160 9640 3360 9650
rect 3820 9640 4020 9650
rect 4700 9640 4900 9650
rect 5360 9640 5560 9650
rect 6020 9640 6220 9650
rect 6900 9640 7100 9650
rect 7560 9640 7760 9650
rect 8220 9640 8420 9650
rect 9100 9640 9300 9650
rect 9760 9640 9960 9650
rect 10420 9640 10620 9650
rect 11300 9640 11500 9650
rect 11960 9640 12160 9650
rect 12620 9640 12820 9650
rect 13500 9640 13700 9650
rect 14160 9640 14360 9650
rect 14820 9640 15020 9650
rect 15700 9640 15900 9650
rect 16360 9640 16560 9650
rect 17020 9640 17220 9650
rect 17900 9640 18100 9650
rect 18560 9640 18760 9650
rect 19220 9640 19420 9650
rect 20500 9640 20510 9650
rect 1010 9580 2510 9640
rect 2690 9580 3170 9640
rect 3350 9580 3830 9640
rect 4010 9580 4710 9640
rect 4890 9580 5370 9640
rect 5550 9580 6030 9640
rect 6210 9580 15710 9640
rect 15890 9580 16370 9640
rect 16550 9580 17030 9640
rect 17210 9580 17910 9640
rect 18090 9580 18570 9640
rect 18750 9580 19230 9640
rect 19410 9580 20510 9640
rect 1010 9570 1020 9580
rect 2500 9570 2700 9580
rect 3160 9570 3360 9580
rect 3820 9570 4020 9580
rect 4700 9570 4900 9580
rect 5360 9570 5560 9580
rect 6020 9570 6220 9580
rect 6900 9570 7100 9580
rect 7560 9570 7760 9580
rect 8220 9570 8420 9580
rect 9100 9570 9300 9580
rect 9760 9570 9960 9580
rect 10420 9570 10620 9580
rect 11300 9570 11500 9580
rect 11960 9570 12160 9580
rect 12620 9570 12820 9580
rect 13500 9570 13700 9580
rect 14160 9570 14360 9580
rect 14820 9570 15020 9580
rect 15700 9570 15900 9580
rect 16360 9570 16560 9580
rect 17020 9570 17220 9580
rect 17900 9570 18100 9580
rect 18560 9570 18760 9580
rect 19220 9570 19420 9580
rect 20500 9570 20510 9580
rect 20690 9640 20700 9650
rect 20690 9580 22180 9640
rect 20690 9570 20700 9580
rect 820 9560 1020 9570
rect 20500 9560 20700 9570
rect 1220 9510 1420 9520
rect 20900 9510 21100 9520
rect 1220 9500 1230 9510
rect -220 9440 1230 9500
rect 1220 9430 1230 9440
rect 1410 9500 1420 9510
rect 2500 9500 2700 9510
rect 3160 9500 3360 9510
rect 3820 9500 4020 9510
rect 4700 9500 4900 9510
rect 5360 9500 5560 9510
rect 6020 9500 6220 9510
rect 6900 9500 7100 9510
rect 7560 9500 7760 9510
rect 8220 9500 8420 9510
rect 9100 9500 9300 9510
rect 9760 9500 9960 9510
rect 10420 9500 10620 9510
rect 11300 9500 11500 9510
rect 11960 9500 12160 9510
rect 12620 9500 12820 9510
rect 13500 9500 13700 9510
rect 14160 9500 14360 9510
rect 14820 9500 15020 9510
rect 15700 9500 15900 9510
rect 16360 9500 16560 9510
rect 17020 9500 17220 9510
rect 17900 9500 18100 9510
rect 18560 9500 18760 9510
rect 19220 9500 19420 9510
rect 20900 9500 20910 9510
rect 1410 9440 6910 9500
rect 7090 9440 7570 9500
rect 7750 9440 8230 9500
rect 8410 9440 9110 9500
rect 9290 9440 9770 9500
rect 9950 9440 10430 9500
rect 10610 9440 11310 9500
rect 11490 9440 11970 9500
rect 12150 9440 12630 9500
rect 12810 9440 13510 9500
rect 13690 9440 14170 9500
rect 14350 9440 14830 9500
rect 15010 9440 20910 9500
rect 1410 9430 1420 9440
rect 2500 9430 2700 9440
rect 3160 9430 3360 9440
rect 3820 9430 4020 9440
rect 4700 9430 4900 9440
rect 5360 9430 5560 9440
rect 6020 9430 6220 9440
rect 6900 9430 7100 9440
rect 7560 9430 7760 9440
rect 8220 9430 8420 9440
rect 9100 9430 9300 9440
rect 9760 9430 9960 9440
rect 10420 9430 10620 9440
rect 11300 9430 11500 9440
rect 11960 9430 12160 9440
rect 12620 9430 12820 9440
rect 13500 9430 13700 9440
rect 14160 9430 14360 9440
rect 14820 9430 15020 9440
rect 15700 9430 15900 9440
rect 16360 9430 16560 9440
rect 17020 9430 17220 9440
rect 17900 9430 18100 9440
rect 18560 9430 18760 9440
rect 19220 9430 19420 9440
rect 20900 9430 20910 9440
rect 21090 9500 21100 9510
rect 21090 9440 22180 9500
rect 21090 9430 21100 9440
rect 1220 9420 1420 9430
rect 20900 9420 21100 9430
rect 31450 9410 31680 9420
rect 31450 9390 31460 9410
rect -110 9340 30 9360
rect -110 9090 -80 9340
rect 0 9090 30 9340
rect -110 9060 30 9090
rect 2090 9340 2230 9360
rect 2090 9090 2120 9340
rect 2200 9090 2230 9340
rect 2090 9060 2230 9090
rect 4290 9340 4430 9360
rect 4290 9090 4320 9340
rect 4400 9090 4430 9340
rect 4290 9060 4430 9090
rect 6490 9340 6630 9360
rect 6490 9090 6520 9340
rect 6600 9090 6630 9340
rect 6490 9060 6630 9090
rect 8690 9340 8830 9360
rect 8690 9090 8720 9340
rect 8800 9090 8830 9340
rect 8690 9060 8830 9090
rect 10890 9340 11030 9360
rect 10890 9090 10920 9340
rect 11000 9090 11030 9340
rect 10890 9060 11030 9090
rect 13090 9340 13230 9360
rect 13090 9090 13120 9340
rect 13200 9090 13230 9340
rect 13090 9060 13230 9090
rect 15290 9340 15430 9360
rect 15290 9090 15320 9340
rect 15400 9090 15430 9340
rect 15290 9060 15430 9090
rect 17490 9340 17630 9360
rect 17490 9090 17520 9340
rect 17600 9090 17630 9340
rect 17490 9060 17630 9090
rect 19690 9340 19830 9360
rect 19690 9090 19720 9340
rect 19800 9090 19830 9340
rect 19690 9060 19830 9090
rect 21890 9340 22030 9360
rect 21890 9090 21920 9340
rect 22000 9090 22030 9340
rect 21890 9060 22030 9090
rect 31440 9220 31460 9390
rect 31670 9390 31680 9410
rect 31670 9380 38100 9390
rect 31670 9220 37910 9380
rect 31440 9200 37910 9220
rect 38090 9200 38100 9380
rect 31440 9190 38100 9200
rect 4700 9010 6220 9020
rect 420 8990 620 9000
rect 420 8910 430 8990
rect 610 8910 620 8990
rect 1620 8990 1820 9000
rect 1620 8980 1630 8990
rect 1600 8920 1630 8980
rect 420 8900 620 8910
rect 1620 8910 1630 8920
rect 1810 8980 1820 8990
rect 4700 8980 4710 9010
rect 1810 8950 4710 8980
rect 6210 8980 6220 9010
rect 6900 9010 8420 9020
rect 6900 8980 6910 9010
rect 6210 8950 6910 8980
rect 8410 8980 8420 9010
rect 9100 9010 10620 9020
rect 9100 8980 9110 9010
rect 8410 8950 9110 8980
rect 10610 8980 10620 9010
rect 11300 9010 12820 9020
rect 11300 8980 11310 9010
rect 10610 8950 11310 8980
rect 12810 8980 12820 9010
rect 13500 9010 15020 9020
rect 13500 8980 13510 9010
rect 12810 8950 13510 8980
rect 15010 8980 15020 9010
rect 15700 9010 17220 9020
rect 15700 8980 15710 9010
rect 15010 8950 15710 8980
rect 17210 8980 17220 9010
rect 20100 8990 20300 9000
rect 20100 8980 20110 8990
rect 17210 8950 20110 8980
rect 1810 8920 20110 8950
rect 1810 8910 1820 8920
rect 1620 8900 1820 8910
rect 20100 8910 20110 8920
rect 20290 8980 20300 8990
rect 21300 8990 21500 9000
rect 20290 8920 20320 8980
rect 20290 8910 20300 8920
rect 20100 8900 20300 8910
rect 21300 8910 21310 8990
rect 21490 8910 21500 8990
rect 21300 8900 21500 8910
rect 31440 8990 31690 9190
rect 820 8850 1020 8860
rect 20500 8850 20700 8860
rect 820 8840 830 8850
rect -220 8780 830 8840
rect 820 8770 830 8780
rect 1010 8840 1020 8850
rect 2500 8840 2700 8850
rect 3160 8840 3360 8850
rect 3820 8840 4020 8850
rect 4700 8840 4900 8850
rect 5360 8840 5560 8850
rect 6020 8840 6220 8850
rect 6900 8840 7100 8850
rect 7560 8840 7760 8850
rect 8220 8840 8420 8850
rect 9100 8840 9300 8850
rect 9760 8840 9960 8850
rect 10420 8840 10620 8850
rect 11300 8840 11500 8850
rect 11960 8840 12160 8850
rect 12620 8840 12820 8850
rect 13500 8840 13700 8850
rect 14160 8840 14360 8850
rect 14820 8840 15020 8850
rect 15700 8840 15900 8850
rect 16360 8840 16560 8850
rect 17020 8840 17220 8850
rect 17900 8840 18100 8850
rect 18560 8840 18760 8850
rect 19220 8840 19420 8850
rect 20500 8840 20510 8850
rect 1010 8780 6910 8840
rect 7090 8780 7570 8840
rect 7750 8780 8230 8840
rect 8410 8780 9110 8840
rect 9290 8780 9770 8840
rect 9950 8780 10430 8840
rect 10610 8780 11310 8840
rect 11490 8780 11970 8840
rect 12150 8780 12630 8840
rect 12810 8780 13510 8840
rect 13690 8780 14170 8840
rect 14350 8780 14830 8840
rect 15010 8780 20510 8840
rect 1010 8770 1020 8780
rect 2500 8770 2700 8780
rect 3160 8770 3360 8780
rect 3820 8770 4020 8780
rect 4700 8770 4900 8780
rect 5360 8770 5560 8780
rect 6020 8770 6220 8780
rect 6900 8770 7100 8780
rect 7560 8770 7760 8780
rect 8220 8770 8420 8780
rect 9100 8770 9300 8780
rect 9760 8770 9960 8780
rect 10420 8770 10620 8780
rect 11300 8770 11500 8780
rect 11960 8770 12160 8780
rect 12620 8770 12820 8780
rect 13500 8770 13700 8780
rect 14160 8770 14360 8780
rect 14820 8770 15020 8780
rect 15700 8770 15900 8780
rect 16360 8770 16560 8780
rect 17020 8770 17220 8780
rect 17900 8770 18100 8780
rect 18560 8770 18760 8780
rect 19220 8770 19420 8780
rect 20500 8770 20510 8780
rect 20690 8840 20700 8850
rect 20690 8780 22180 8840
rect 31440 8780 31450 8990
rect 31680 8780 31690 8990
rect 20690 8770 20700 8780
rect 31440 8770 31690 8780
rect 820 8760 1020 8770
rect 20500 8760 20700 8770
rect 1220 8710 1420 8720
rect 20900 8710 21100 8720
rect 1220 8700 1230 8710
rect -220 8640 1230 8700
rect 1220 8630 1230 8640
rect 1410 8700 1420 8710
rect 2500 8700 2700 8710
rect 3160 8700 3360 8710
rect 3820 8700 4020 8710
rect 4700 8700 4900 8710
rect 5360 8700 5560 8710
rect 6020 8700 6220 8710
rect 6900 8700 7100 8710
rect 7560 8700 7760 8710
rect 8220 8700 8420 8710
rect 9100 8700 9300 8710
rect 9760 8700 9960 8710
rect 10420 8700 10620 8710
rect 11300 8700 11500 8710
rect 11960 8700 12160 8710
rect 12620 8700 12820 8710
rect 13500 8700 13700 8710
rect 14160 8700 14360 8710
rect 14820 8700 15020 8710
rect 15700 8700 15900 8710
rect 16360 8700 16560 8710
rect 17020 8700 17220 8710
rect 17900 8700 18100 8710
rect 18560 8700 18760 8710
rect 19220 8700 19420 8710
rect 20900 8700 20910 8710
rect 1410 8640 2510 8700
rect 2690 8640 3170 8700
rect 3350 8640 3830 8700
rect 4010 8640 4710 8700
rect 4890 8640 5370 8700
rect 5550 8640 6030 8700
rect 6210 8640 15710 8700
rect 15890 8640 16370 8700
rect 16550 8640 17030 8700
rect 17210 8640 17910 8700
rect 18090 8640 18570 8700
rect 18750 8640 19230 8700
rect 19410 8640 20910 8700
rect 1410 8630 1420 8640
rect 2500 8630 2700 8640
rect 3160 8630 3360 8640
rect 3820 8630 4020 8640
rect 4700 8630 4900 8640
rect 5360 8630 5560 8640
rect 6020 8630 6220 8640
rect 6900 8630 7100 8640
rect 7560 8630 7760 8640
rect 8220 8630 8420 8640
rect 9100 8630 9300 8640
rect 9760 8630 9960 8640
rect 10420 8630 10620 8640
rect 11300 8630 11500 8640
rect 11960 8630 12160 8640
rect 12620 8630 12820 8640
rect 13500 8630 13700 8640
rect 14160 8630 14360 8640
rect 14820 8630 15020 8640
rect 15700 8630 15900 8640
rect 16360 8630 16560 8640
rect 17020 8630 17220 8640
rect 17900 8630 18100 8640
rect 18560 8630 18760 8640
rect 19220 8630 19420 8640
rect 20900 8630 20910 8640
rect 21090 8700 21100 8710
rect 21090 8640 22180 8700
rect 21090 8630 21100 8640
rect 1220 8620 1420 8630
rect 20900 8620 21100 8630
rect -110 8540 30 8560
rect -110 8290 -80 8540
rect 0 8290 30 8540
rect -110 8260 30 8290
rect 2090 8540 2230 8560
rect 2090 8290 2120 8540
rect 2200 8290 2230 8540
rect 2090 8260 2230 8290
rect 4290 8540 4430 8560
rect 4290 8290 4320 8540
rect 4400 8290 4430 8540
rect 4290 8260 4430 8290
rect 6490 8540 6630 8560
rect 6490 8290 6520 8540
rect 6600 8290 6630 8540
rect 6490 8260 6630 8290
rect 8690 8540 8830 8560
rect 8690 8290 8720 8540
rect 8800 8290 8830 8540
rect 8690 8260 8830 8290
rect 10890 8540 11030 8560
rect 10890 8290 10920 8540
rect 11000 8290 11030 8540
rect 10890 8260 11030 8290
rect 13090 8540 13230 8560
rect 13090 8290 13120 8540
rect 13200 8290 13230 8540
rect 13090 8260 13230 8290
rect 15290 8540 15430 8560
rect 15290 8290 15320 8540
rect 15400 8290 15430 8540
rect 15290 8260 15430 8290
rect 17490 8540 17630 8560
rect 17490 8290 17520 8540
rect 17600 8290 17630 8540
rect 17490 8260 17630 8290
rect 19690 8540 19830 8560
rect 19690 8290 19720 8540
rect 19800 8290 19830 8540
rect 19690 8260 19830 8290
rect 21890 8540 22030 8560
rect 21890 8290 21920 8540
rect 22000 8290 22030 8540
rect 21890 8260 22030 8290
rect 4700 8210 6220 8220
rect 420 8190 620 8200
rect 420 8110 430 8190
rect 610 8110 620 8190
rect 1620 8190 1820 8200
rect 1620 8180 1630 8190
rect 1600 8120 1630 8180
rect 420 8100 620 8110
rect 1620 8110 1630 8120
rect 1810 8180 1820 8190
rect 4700 8180 4710 8210
rect 1810 8150 4710 8180
rect 6210 8180 6220 8210
rect 6900 8210 8420 8220
rect 6900 8180 6910 8210
rect 6210 8150 6910 8180
rect 8410 8180 8420 8210
rect 9100 8210 10620 8220
rect 9100 8180 9110 8210
rect 8410 8150 9110 8180
rect 10610 8180 10620 8210
rect 11300 8210 12820 8220
rect 11300 8180 11310 8210
rect 10610 8150 11310 8180
rect 12810 8180 12820 8210
rect 13500 8210 15020 8220
rect 13500 8180 13510 8210
rect 12810 8150 13510 8180
rect 15010 8180 15020 8210
rect 15700 8210 17220 8220
rect 15700 8180 15710 8210
rect 15010 8150 15710 8180
rect 17210 8180 17220 8210
rect 20100 8190 20300 8200
rect 20100 8180 20110 8190
rect 17210 8150 20110 8180
rect 1810 8120 20110 8150
rect 1810 8110 1820 8120
rect 1620 8100 1820 8110
rect 20100 8110 20110 8120
rect 20290 8180 20300 8190
rect 21300 8190 21500 8200
rect 20290 8120 20320 8180
rect 20290 8110 20300 8120
rect 20100 8100 20300 8110
rect 21300 8110 21310 8190
rect 21490 8110 21500 8190
rect 21300 8100 21500 8110
rect 34740 8180 34900 8190
rect 820 8050 1020 8060
rect 20500 8050 20700 8060
rect 820 8040 830 8050
rect -220 7980 830 8040
rect 820 7970 830 7980
rect 1010 8040 1020 8050
rect 2500 8040 2700 8050
rect 3160 8040 3360 8050
rect 3820 8040 4020 8050
rect 4700 8040 4900 8050
rect 5360 8040 5560 8050
rect 6020 8040 6220 8050
rect 6900 8040 7100 8050
rect 7560 8040 7760 8050
rect 8220 8040 8420 8050
rect 9100 8040 9300 8050
rect 9760 8040 9960 8050
rect 10420 8040 10620 8050
rect 11300 8040 11500 8050
rect 11960 8040 12160 8050
rect 12620 8040 12820 8050
rect 13500 8040 13700 8050
rect 14160 8040 14360 8050
rect 14820 8040 15020 8050
rect 15700 8040 15900 8050
rect 16360 8040 16560 8050
rect 17020 8040 17220 8050
rect 17900 8040 18100 8050
rect 18560 8040 18760 8050
rect 19220 8040 19420 8050
rect 20500 8040 20510 8050
rect 1010 7980 6910 8040
rect 7090 7980 7570 8040
rect 7750 7980 8230 8040
rect 8410 7980 9110 8040
rect 9290 7980 9770 8040
rect 9950 7980 10430 8040
rect 10610 7980 11310 8040
rect 11490 7980 11970 8040
rect 12150 7980 12630 8040
rect 12810 7980 13510 8040
rect 13690 7980 14170 8040
rect 14350 7980 14830 8040
rect 15010 7980 20510 8040
rect 1010 7970 1020 7980
rect 2500 7970 2700 7980
rect 3160 7970 3360 7980
rect 3820 7970 4020 7980
rect 4700 7970 4900 7980
rect 5360 7970 5560 7980
rect 6020 7970 6220 7980
rect 6900 7970 7100 7980
rect 7560 7970 7760 7980
rect 8220 7970 8420 7980
rect 9100 7970 9300 7980
rect 9760 7970 9960 7980
rect 10420 7970 10620 7980
rect 11300 7970 11500 7980
rect 11960 7970 12160 7980
rect 12620 7970 12820 7980
rect 13500 7970 13700 7980
rect 14160 7970 14360 7980
rect 14820 7970 15020 7980
rect 15700 7970 15900 7980
rect 16360 7970 16560 7980
rect 17020 7970 17220 7980
rect 17900 7970 18100 7980
rect 18560 7970 18760 7980
rect 19220 7970 19420 7980
rect 20500 7970 20510 7980
rect 20690 8040 20700 8050
rect 20690 7980 22180 8040
rect 20690 7970 20700 7980
rect 820 7960 1020 7970
rect 20500 7960 20700 7970
rect 34740 7960 34750 8180
rect 34890 8130 34900 8180
rect 36780 8170 37020 8180
rect 36780 8130 36790 8170
rect 34890 8070 36790 8130
rect 34890 7960 34900 8070
rect 36780 8030 36790 8070
rect 37010 8030 37020 8170
rect 36780 8020 37020 8030
rect 34740 7950 34900 7960
rect 35160 7980 35320 7990
rect 1220 7910 1420 7920
rect 20900 7910 21100 7920
rect 1220 7900 1230 7910
rect -220 7840 1230 7900
rect 1220 7830 1230 7840
rect 1410 7900 1420 7910
rect 2500 7900 2700 7910
rect 3160 7900 3360 7910
rect 3820 7900 4020 7910
rect 4700 7900 4900 7910
rect 5360 7900 5560 7910
rect 6020 7900 6220 7910
rect 6900 7900 7100 7910
rect 7560 7900 7760 7910
rect 8220 7900 8420 7910
rect 9100 7900 9300 7910
rect 9760 7900 9960 7910
rect 10420 7900 10620 7910
rect 11300 7900 11500 7910
rect 11960 7900 12160 7910
rect 12620 7900 12820 7910
rect 13500 7900 13700 7910
rect 14160 7900 14360 7910
rect 14820 7900 15020 7910
rect 15700 7900 15900 7910
rect 16360 7900 16560 7910
rect 17020 7900 17220 7910
rect 17900 7900 18100 7910
rect 18560 7900 18760 7910
rect 19220 7900 19420 7910
rect 20900 7900 20910 7910
rect 1410 7840 2510 7900
rect 2690 7840 3170 7900
rect 3350 7840 3830 7900
rect 4010 7840 4710 7900
rect 4890 7840 5370 7900
rect 5550 7840 6030 7900
rect 6210 7840 15710 7900
rect 15890 7840 16370 7900
rect 16550 7840 17030 7900
rect 17210 7840 17910 7900
rect 18090 7840 18570 7900
rect 18750 7840 19230 7900
rect 19410 7840 20910 7900
rect 1410 7830 1420 7840
rect 2500 7830 2700 7840
rect 3160 7830 3360 7840
rect 3820 7830 4020 7840
rect 4700 7830 4900 7840
rect 5360 7830 5560 7840
rect 6020 7830 6220 7840
rect 6900 7830 7100 7840
rect 7560 7830 7760 7840
rect 8220 7830 8420 7840
rect 9100 7830 9300 7840
rect 9760 7830 9960 7840
rect 10420 7830 10620 7840
rect 11300 7830 11500 7840
rect 11960 7830 12160 7840
rect 12620 7830 12820 7840
rect 13500 7830 13700 7840
rect 14160 7830 14360 7840
rect 14820 7830 15020 7840
rect 15700 7830 15900 7840
rect 16360 7830 16560 7840
rect 17020 7830 17220 7840
rect 17900 7830 18100 7840
rect 18560 7830 18760 7840
rect 19220 7830 19420 7840
rect 20900 7830 20910 7840
rect 21090 7900 21100 7910
rect 21090 7840 22180 7900
rect 21090 7830 21100 7840
rect 1220 7820 1420 7830
rect 20900 7820 21100 7830
rect 35160 7760 35170 7980
rect 35310 7930 35320 7980
rect 37120 7970 37360 7980
rect 37120 7930 37130 7970
rect 35310 7870 37130 7930
rect 35310 7760 35320 7870
rect 37120 7830 37130 7870
rect 37350 7830 37360 7970
rect 37120 7820 37360 7830
rect -110 7740 30 7760
rect -110 7490 -80 7740
rect 0 7490 30 7740
rect -110 7460 30 7490
rect 2090 7740 2230 7760
rect 2090 7490 2120 7740
rect 2200 7490 2230 7740
rect 2090 7460 2230 7490
rect 4290 7740 4430 7760
rect 4290 7490 4320 7740
rect 4400 7490 4430 7740
rect 4290 7460 4430 7490
rect 6490 7740 6630 7760
rect 6490 7490 6520 7740
rect 6600 7490 6630 7740
rect 6490 7460 6630 7490
rect 8690 7740 8830 7760
rect 8690 7490 8720 7740
rect 8800 7490 8830 7740
rect 8690 7460 8830 7490
rect 10890 7740 11030 7760
rect 10890 7490 10920 7740
rect 11000 7490 11030 7740
rect 10890 7460 11030 7490
rect 13090 7740 13230 7760
rect 13090 7490 13120 7740
rect 13200 7490 13230 7740
rect 13090 7460 13230 7490
rect 15290 7740 15430 7760
rect 15290 7490 15320 7740
rect 15400 7490 15430 7740
rect 15290 7460 15430 7490
rect 17490 7740 17630 7760
rect 17490 7490 17520 7740
rect 17600 7490 17630 7740
rect 17490 7460 17630 7490
rect 19690 7740 19830 7760
rect 19690 7490 19720 7740
rect 19800 7490 19830 7740
rect 19690 7460 19830 7490
rect 21890 7740 22030 7760
rect 35160 7750 35320 7760
rect 21890 7490 21920 7740
rect 22000 7490 22030 7740
rect 21890 7460 22030 7490
rect 4700 7410 6220 7420
rect 420 7390 620 7400
rect 420 7310 430 7390
rect 610 7310 620 7390
rect 1620 7390 1820 7400
rect 1620 7380 1630 7390
rect 1600 7320 1630 7380
rect 420 7300 620 7310
rect 1620 7310 1630 7320
rect 1810 7380 1820 7390
rect 4700 7380 4710 7410
rect 1810 7350 4710 7380
rect 6210 7380 6220 7410
rect 6900 7410 8420 7420
rect 6900 7380 6910 7410
rect 6210 7350 6910 7380
rect 8410 7380 8420 7410
rect 9100 7410 10620 7420
rect 9100 7380 9110 7410
rect 8410 7350 9110 7380
rect 10610 7380 10620 7410
rect 11300 7410 12820 7420
rect 11300 7380 11310 7410
rect 10610 7350 11310 7380
rect 12810 7380 12820 7410
rect 13500 7410 15020 7420
rect 13500 7380 13510 7410
rect 12810 7350 13510 7380
rect 15010 7380 15020 7410
rect 15700 7410 17220 7420
rect 15700 7380 15710 7410
rect 15010 7350 15710 7380
rect 17210 7380 17220 7410
rect 20100 7390 20300 7400
rect 20100 7380 20110 7390
rect 17210 7350 20110 7380
rect 1810 7320 20110 7350
rect 1810 7310 1820 7320
rect 1620 7300 1820 7310
rect 20100 7310 20110 7320
rect 20290 7380 20300 7390
rect 21300 7390 21500 7400
rect 20290 7320 20320 7380
rect 20290 7310 20300 7320
rect 20100 7300 20300 7310
rect 21300 7310 21310 7390
rect 21490 7310 21500 7390
rect 21300 7300 21500 7310
rect 820 7250 1020 7260
rect 20500 7250 20700 7260
rect 820 7240 830 7250
rect -220 7180 830 7240
rect 820 7170 830 7180
rect 1010 7240 1020 7250
rect 2500 7240 2700 7250
rect 3160 7240 3360 7250
rect 3820 7240 4020 7250
rect 4700 7240 4900 7250
rect 5360 7240 5560 7250
rect 6020 7240 6220 7250
rect 6900 7240 7100 7250
rect 7560 7240 7760 7250
rect 8220 7240 8420 7250
rect 9100 7240 9300 7250
rect 9760 7240 9960 7250
rect 10420 7240 10620 7250
rect 11300 7240 11500 7250
rect 11960 7240 12160 7250
rect 12620 7240 12820 7250
rect 13500 7240 13700 7250
rect 14160 7240 14360 7250
rect 14820 7240 15020 7250
rect 15700 7240 15900 7250
rect 16360 7240 16560 7250
rect 17020 7240 17220 7250
rect 17900 7240 18100 7250
rect 18560 7240 18760 7250
rect 19220 7240 19420 7250
rect 20500 7240 20510 7250
rect 1010 7180 2510 7240
rect 2690 7180 3170 7240
rect 3350 7180 3830 7240
rect 4010 7180 4710 7240
rect 4890 7180 5370 7240
rect 5550 7180 6030 7240
rect 6210 7180 15710 7240
rect 15890 7180 16370 7240
rect 16550 7180 17030 7240
rect 17210 7180 17910 7240
rect 18090 7180 18570 7240
rect 18750 7180 19230 7240
rect 19410 7180 20510 7240
rect 1010 7170 1020 7180
rect 2500 7170 2700 7180
rect 3160 7170 3360 7180
rect 3820 7170 4020 7180
rect 4700 7170 4900 7180
rect 5360 7170 5560 7180
rect 6020 7170 6220 7180
rect 6900 7170 7100 7180
rect 7560 7170 7760 7180
rect 8220 7170 8420 7180
rect 9100 7170 9300 7180
rect 9760 7170 9960 7180
rect 10420 7170 10620 7180
rect 11300 7170 11500 7180
rect 11960 7170 12160 7180
rect 12620 7170 12820 7180
rect 13500 7170 13700 7180
rect 14160 7170 14360 7180
rect 14820 7170 15020 7180
rect 15700 7170 15900 7180
rect 16360 7170 16560 7180
rect 17020 7170 17220 7180
rect 17900 7170 18100 7180
rect 18560 7170 18760 7180
rect 19220 7170 19420 7180
rect 20500 7170 20510 7180
rect 20690 7240 20700 7250
rect 20690 7180 22180 7240
rect 20690 7170 20700 7180
rect 820 7160 1020 7170
rect 20500 7160 20700 7170
rect 1220 7110 1420 7120
rect 20900 7110 21100 7120
rect 1220 7100 1230 7110
rect -220 7040 1230 7100
rect 1220 7030 1230 7040
rect 1410 7100 1420 7110
rect 2500 7100 2700 7110
rect 3160 7100 3360 7110
rect 3820 7100 4020 7110
rect 4700 7100 4900 7110
rect 5360 7100 5560 7110
rect 6020 7100 6220 7110
rect 6900 7100 7100 7110
rect 7560 7100 7760 7110
rect 8220 7100 8420 7110
rect 9100 7100 9300 7110
rect 9760 7100 9960 7110
rect 10420 7100 10620 7110
rect 11300 7100 11500 7110
rect 11960 7100 12160 7110
rect 12620 7100 12820 7110
rect 13500 7100 13700 7110
rect 14160 7100 14360 7110
rect 14820 7100 15020 7110
rect 15700 7100 15900 7110
rect 16360 7100 16560 7110
rect 17020 7100 17220 7110
rect 17900 7100 18100 7110
rect 18560 7100 18760 7110
rect 19220 7100 19420 7110
rect 20900 7100 20910 7110
rect 1410 7040 6910 7100
rect 7090 7040 7570 7100
rect 7750 7040 8230 7100
rect 8410 7040 9110 7100
rect 9290 7040 9770 7100
rect 9950 7040 10430 7100
rect 10610 7040 11310 7100
rect 11490 7040 11970 7100
rect 12150 7040 12630 7100
rect 12810 7040 13510 7100
rect 13690 7040 14170 7100
rect 14350 7040 14830 7100
rect 15010 7040 20910 7100
rect 1410 7030 1420 7040
rect 2500 7030 2700 7040
rect 3160 7030 3360 7040
rect 3820 7030 4020 7040
rect 4700 7030 4900 7040
rect 5360 7030 5560 7040
rect 6020 7030 6220 7040
rect 6900 7030 7100 7040
rect 7560 7030 7760 7040
rect 8220 7030 8420 7040
rect 9100 7030 9300 7040
rect 9760 7030 9960 7040
rect 10420 7030 10620 7040
rect 11300 7030 11500 7040
rect 11960 7030 12160 7040
rect 12620 7030 12820 7040
rect 13500 7030 13700 7040
rect 14160 7030 14360 7040
rect 14820 7030 15020 7040
rect 15700 7030 15900 7040
rect 16360 7030 16560 7040
rect 17020 7030 17220 7040
rect 17900 7030 18100 7040
rect 18560 7030 18760 7040
rect 19220 7030 19420 7040
rect 20900 7030 20910 7040
rect 21090 7100 21100 7110
rect 21090 7040 22180 7100
rect 21090 7030 21100 7040
rect 1220 7020 1420 7030
rect 20900 7020 21100 7030
rect -110 6940 30 6960
rect -110 6690 -80 6940
rect 0 6690 30 6940
rect -110 6660 30 6690
rect 2090 6940 2230 6960
rect 2090 6690 2120 6940
rect 2200 6690 2230 6940
rect 2090 6660 2230 6690
rect 4290 6940 4430 6960
rect 4290 6690 4320 6940
rect 4400 6690 4430 6940
rect 4290 6660 4430 6690
rect 6490 6940 6630 6960
rect 6490 6690 6520 6940
rect 6600 6690 6630 6940
rect 6490 6660 6630 6690
rect 8690 6940 8830 6960
rect 8690 6690 8720 6940
rect 8800 6690 8830 6940
rect 8690 6660 8830 6690
rect 10890 6940 11030 6960
rect 10890 6690 10920 6940
rect 11000 6690 11030 6940
rect 10890 6660 11030 6690
rect 13090 6940 13230 6960
rect 13090 6690 13120 6940
rect 13200 6690 13230 6940
rect 13090 6660 13230 6690
rect 15290 6940 15430 6960
rect 15290 6690 15320 6940
rect 15400 6690 15430 6940
rect 15290 6660 15430 6690
rect 17490 6940 17630 6960
rect 17490 6690 17520 6940
rect 17600 6690 17630 6940
rect 17490 6660 17630 6690
rect 19690 6940 19830 6960
rect 19690 6690 19720 6940
rect 19800 6690 19830 6940
rect 19690 6660 19830 6690
rect 21890 6940 22030 6960
rect 21890 6690 21920 6940
rect 22000 6690 22030 6940
rect 21890 6660 22030 6690
rect 4700 6610 6220 6620
rect 420 6590 620 6600
rect 420 6510 430 6590
rect 610 6510 620 6590
rect 1620 6590 1820 6600
rect 1620 6580 1630 6590
rect 1600 6520 1630 6580
rect 420 6500 620 6510
rect 1620 6510 1630 6520
rect 1810 6580 1820 6590
rect 4700 6580 4710 6610
rect 1810 6550 4710 6580
rect 6210 6580 6220 6610
rect 6900 6610 8420 6620
rect 6900 6580 6910 6610
rect 6210 6550 6910 6580
rect 8410 6580 8420 6610
rect 9100 6610 10620 6620
rect 9100 6580 9110 6610
rect 8410 6550 9110 6580
rect 10610 6580 10620 6610
rect 11300 6610 12820 6620
rect 11300 6580 11310 6610
rect 10610 6550 11310 6580
rect 12810 6580 12820 6610
rect 13500 6610 15020 6620
rect 13500 6580 13510 6610
rect 12810 6550 13510 6580
rect 15010 6580 15020 6610
rect 15700 6610 17220 6620
rect 15700 6580 15710 6610
rect 15010 6550 15710 6580
rect 17210 6580 17220 6610
rect 20100 6590 20300 6600
rect 20100 6580 20110 6590
rect 17210 6550 20110 6580
rect 1810 6520 20110 6550
rect 1810 6510 1820 6520
rect 1620 6500 1820 6510
rect 20100 6510 20110 6520
rect 20290 6580 20300 6590
rect 21300 6590 21500 6600
rect 20290 6520 20320 6580
rect 20290 6510 20300 6520
rect 20100 6500 20300 6510
rect 21300 6510 21310 6590
rect 21490 6510 21500 6590
rect 21300 6500 21500 6510
rect 820 6450 1020 6460
rect 20500 6450 20700 6460
rect 820 6440 830 6450
rect -220 6380 830 6440
rect 820 6370 830 6380
rect 1010 6440 1020 6450
rect 2500 6440 2700 6450
rect 3160 6440 3360 6450
rect 3820 6440 4020 6450
rect 4700 6440 4900 6450
rect 5360 6440 5560 6450
rect 6020 6440 6220 6450
rect 6900 6440 7100 6450
rect 7560 6440 7760 6450
rect 8220 6440 8420 6450
rect 9100 6440 9300 6450
rect 9760 6440 9960 6450
rect 10420 6440 10620 6450
rect 11300 6440 11500 6450
rect 11960 6440 12160 6450
rect 12620 6440 12820 6450
rect 13500 6440 13700 6450
rect 14160 6440 14360 6450
rect 14820 6440 15020 6450
rect 15700 6440 15900 6450
rect 16360 6440 16560 6450
rect 17020 6440 17220 6450
rect 17900 6440 18100 6450
rect 18560 6440 18760 6450
rect 19220 6440 19420 6450
rect 20500 6440 20510 6450
rect 1010 6380 6910 6440
rect 7090 6380 7570 6440
rect 7750 6380 8230 6440
rect 8410 6380 9110 6440
rect 9290 6380 9770 6440
rect 9950 6380 10430 6440
rect 10610 6380 11310 6440
rect 11490 6380 11970 6440
rect 12150 6380 12630 6440
rect 12810 6380 13510 6440
rect 13690 6380 14170 6440
rect 14350 6380 14830 6440
rect 15010 6380 20510 6440
rect 1010 6370 1020 6380
rect 2500 6370 2700 6380
rect 3160 6370 3360 6380
rect 3820 6370 4020 6380
rect 4700 6370 4900 6380
rect 5360 6370 5560 6380
rect 6020 6370 6220 6380
rect 6900 6370 7100 6380
rect 7560 6370 7760 6380
rect 8220 6370 8420 6380
rect 9100 6370 9300 6380
rect 9760 6370 9960 6380
rect 10420 6370 10620 6380
rect 11300 6370 11500 6380
rect 11960 6370 12160 6380
rect 12620 6370 12820 6380
rect 13500 6370 13700 6380
rect 14160 6370 14360 6380
rect 14820 6370 15020 6380
rect 15700 6370 15900 6380
rect 16360 6370 16560 6380
rect 17020 6370 17220 6380
rect 17900 6370 18100 6380
rect 18560 6370 18760 6380
rect 19220 6370 19420 6380
rect 20500 6370 20510 6380
rect 20690 6440 20700 6450
rect 20690 6380 22180 6440
rect 20690 6370 20700 6380
rect 820 6360 1020 6370
rect 20500 6360 20700 6370
rect 1220 6310 1420 6320
rect 20900 6310 21100 6320
rect 1220 6300 1230 6310
rect -220 6240 1230 6300
rect 1220 6230 1230 6240
rect 1410 6300 1420 6310
rect 2500 6300 2700 6310
rect 3160 6300 3360 6310
rect 3820 6300 4020 6310
rect 4700 6300 4900 6310
rect 5360 6300 5560 6310
rect 6020 6300 6220 6310
rect 6900 6300 7100 6310
rect 7560 6300 7760 6310
rect 8220 6300 8420 6310
rect 9100 6300 9300 6310
rect 9760 6300 9960 6310
rect 10420 6300 10620 6310
rect 11300 6300 11500 6310
rect 11960 6300 12160 6310
rect 12620 6300 12820 6310
rect 13500 6300 13700 6310
rect 14160 6300 14360 6310
rect 14820 6300 15020 6310
rect 15700 6300 15900 6310
rect 16360 6300 16560 6310
rect 17020 6300 17220 6310
rect 17900 6300 18100 6310
rect 18560 6300 18760 6310
rect 19220 6300 19420 6310
rect 20900 6300 20910 6310
rect 1410 6240 2510 6300
rect 2690 6240 3170 6300
rect 3350 6240 3830 6300
rect 4010 6240 4710 6300
rect 4890 6240 5370 6300
rect 5550 6240 6030 6300
rect 6210 6240 15710 6300
rect 15890 6240 16370 6300
rect 16550 6240 17030 6300
rect 17210 6240 17910 6300
rect 18090 6240 18570 6300
rect 18750 6240 19230 6300
rect 19410 6240 20910 6300
rect 1410 6230 1420 6240
rect 2500 6230 2700 6240
rect 3160 6230 3360 6240
rect 3820 6230 4020 6240
rect 4700 6230 4900 6240
rect 5360 6230 5560 6240
rect 6020 6230 6220 6240
rect 6900 6230 7100 6240
rect 7560 6230 7760 6240
rect 8220 6230 8420 6240
rect 9100 6230 9300 6240
rect 9760 6230 9960 6240
rect 10420 6230 10620 6240
rect 11300 6230 11500 6240
rect 11960 6230 12160 6240
rect 12620 6230 12820 6240
rect 13500 6230 13700 6240
rect 14160 6230 14360 6240
rect 14820 6230 15020 6240
rect 15700 6230 15900 6240
rect 16360 6230 16560 6240
rect 17020 6230 17220 6240
rect 17900 6230 18100 6240
rect 18560 6230 18760 6240
rect 19220 6230 19420 6240
rect 20900 6230 20910 6240
rect 21090 6300 21100 6310
rect 21090 6240 22180 6300
rect 36220 6260 36420 6270
rect 21090 6230 21100 6240
rect 1220 6220 1420 6230
rect 20900 6220 21100 6230
rect -110 6140 30 6160
rect -110 5890 -80 6140
rect 0 5890 30 6140
rect -110 5860 30 5890
rect 2090 6140 2230 6160
rect 2090 5890 2120 6140
rect 2200 5890 2230 6140
rect 2090 5860 2230 5890
rect 4290 6140 4430 6160
rect 4290 5890 4320 6140
rect 4400 5890 4430 6140
rect 4290 5860 4430 5890
rect 6490 6140 6630 6160
rect 6490 5890 6520 6140
rect 6600 5890 6630 6140
rect 6490 5860 6630 5890
rect 8690 6140 8830 6160
rect 8690 5890 8720 6140
rect 8800 5890 8830 6140
rect 8690 5860 8830 5890
rect 10890 6140 11030 6160
rect 10890 5890 10920 6140
rect 11000 5890 11030 6140
rect 10890 5860 11030 5890
rect 13090 6140 13230 6160
rect 13090 5890 13120 6140
rect 13200 5890 13230 6140
rect 13090 5860 13230 5890
rect 15290 6140 15430 6160
rect 15290 5890 15320 6140
rect 15400 5890 15430 6140
rect 15290 5860 15430 5890
rect 17490 6140 17630 6160
rect 17490 5890 17520 6140
rect 17600 5890 17630 6140
rect 17490 5860 17630 5890
rect 19690 6140 19830 6160
rect 19690 5890 19720 6140
rect 19800 5890 19830 6140
rect 19690 5860 19830 5890
rect 21890 6140 22030 6160
rect 21890 5890 21920 6140
rect 22000 5890 22030 6140
rect 36220 6080 36230 6260
rect 36410 6080 36420 6260
rect 36220 6070 36420 6080
rect 36520 6260 36720 6270
rect 36520 6080 36530 6260
rect 36710 6080 36720 6260
rect 36520 6070 36720 6080
rect 21890 5860 22030 5890
rect 2500 5810 4020 5820
rect 1620 5790 1820 5800
rect 1620 5780 1630 5790
rect 1600 5720 1630 5780
rect 1620 5710 1630 5720
rect 1810 5780 1820 5790
rect 2500 5780 2510 5810
rect 1810 5750 2510 5780
rect 4010 5780 4020 5810
rect 4700 5810 6220 5820
rect 4700 5780 4710 5810
rect 4010 5750 4710 5780
rect 6210 5780 6220 5810
rect 6900 5810 8420 5820
rect 6900 5780 6910 5810
rect 6210 5750 6910 5780
rect 8410 5780 8420 5810
rect 9100 5810 10620 5820
rect 9100 5780 9110 5810
rect 8410 5750 9110 5780
rect 10610 5780 10620 5810
rect 11300 5810 12820 5820
rect 11300 5780 11310 5810
rect 10610 5750 11310 5780
rect 12810 5780 12820 5810
rect 13500 5810 15020 5820
rect 13500 5780 13510 5810
rect 12810 5750 13510 5780
rect 15010 5780 15020 5810
rect 15700 5810 17220 5820
rect 15700 5780 15710 5810
rect 15010 5750 15710 5780
rect 17210 5780 17220 5810
rect 17900 5810 19420 5820
rect 17900 5780 17910 5810
rect 17210 5750 17910 5780
rect 19410 5780 19420 5810
rect 20100 5790 20300 5800
rect 20100 5780 20110 5790
rect 19410 5750 20110 5780
rect 1810 5720 20110 5750
rect 1810 5710 1820 5720
rect 1620 5700 1820 5710
rect 20100 5710 20110 5720
rect 20290 5780 20300 5790
rect 20290 5720 20320 5780
rect 20290 5710 20300 5720
rect 20100 5700 20300 5710
rect 820 5650 1020 5660
rect 20500 5650 20700 5660
rect 820 5640 830 5650
rect -220 5580 830 5640
rect 820 5570 830 5580
rect 1010 5640 1020 5650
rect 2500 5640 2700 5650
rect 3160 5640 3360 5650
rect 3820 5640 4020 5650
rect 4700 5640 4900 5650
rect 5360 5640 5560 5650
rect 6020 5640 6220 5650
rect 6900 5640 7100 5650
rect 7560 5640 7760 5650
rect 8220 5640 8420 5650
rect 9100 5640 9300 5650
rect 9760 5640 9960 5650
rect 10420 5640 10620 5650
rect 11300 5640 11500 5650
rect 11960 5640 12160 5650
rect 12620 5640 12820 5650
rect 13500 5640 13700 5650
rect 14160 5640 14360 5650
rect 14820 5640 15020 5650
rect 15700 5640 15900 5650
rect 16360 5640 16560 5650
rect 17020 5640 17220 5650
rect 17900 5640 18100 5650
rect 18560 5640 18760 5650
rect 19220 5640 19420 5650
rect 20500 5640 20510 5650
rect 1010 5580 2510 5640
rect 2690 5580 3170 5640
rect 3350 5580 3830 5640
rect 4010 5580 4710 5640
rect 4890 5580 5370 5640
rect 5550 5580 6030 5640
rect 6210 5580 15710 5640
rect 15890 5580 16370 5640
rect 16550 5580 17030 5640
rect 17210 5580 17910 5640
rect 18090 5580 18570 5640
rect 18750 5580 19230 5640
rect 19410 5580 20510 5640
rect 1010 5570 1020 5580
rect 2500 5570 2700 5580
rect 3160 5570 3360 5580
rect 3820 5570 4020 5580
rect 4700 5570 4900 5580
rect 5360 5570 5560 5580
rect 6020 5570 6220 5580
rect 6900 5570 7100 5580
rect 7560 5570 7760 5580
rect 8220 5570 8420 5580
rect 9100 5570 9300 5580
rect 9760 5570 9960 5580
rect 10420 5570 10620 5580
rect 11300 5570 11500 5580
rect 11960 5570 12160 5580
rect 12620 5570 12820 5580
rect 13500 5570 13700 5580
rect 14160 5570 14360 5580
rect 14820 5570 15020 5580
rect 15700 5570 15900 5580
rect 16360 5570 16560 5580
rect 17020 5570 17220 5580
rect 17900 5570 18100 5580
rect 18560 5570 18760 5580
rect 19220 5570 19420 5580
rect 20500 5570 20510 5580
rect 20690 5640 20700 5650
rect 20690 5580 22180 5640
rect 20690 5570 20700 5580
rect 820 5560 1020 5570
rect 20500 5560 20700 5570
rect 1220 5510 1420 5520
rect 20900 5510 21100 5520
rect 1220 5500 1230 5510
rect -220 5440 1230 5500
rect 1220 5430 1230 5440
rect 1410 5500 1420 5510
rect 2500 5500 2700 5510
rect 3160 5500 3360 5510
rect 3820 5500 4020 5510
rect 4700 5500 4900 5510
rect 5360 5500 5560 5510
rect 6020 5500 6220 5510
rect 6900 5500 7100 5510
rect 7560 5500 7760 5510
rect 8220 5500 8420 5510
rect 9100 5500 9300 5510
rect 9760 5500 9960 5510
rect 10420 5500 10620 5510
rect 11300 5500 11500 5510
rect 11960 5500 12160 5510
rect 12620 5500 12820 5510
rect 13500 5500 13700 5510
rect 14160 5500 14360 5510
rect 14820 5500 15020 5510
rect 15700 5500 15900 5510
rect 16360 5500 16560 5510
rect 17020 5500 17220 5510
rect 17900 5500 18100 5510
rect 18560 5500 18760 5510
rect 19220 5500 19420 5510
rect 20900 5500 20910 5510
rect 1410 5440 6910 5500
rect 7090 5440 7570 5500
rect 7750 5440 8230 5500
rect 8410 5440 9110 5500
rect 9290 5440 9770 5500
rect 9950 5440 10430 5500
rect 10610 5440 11310 5500
rect 11490 5440 11970 5500
rect 12150 5440 12630 5500
rect 12810 5440 13510 5500
rect 13690 5440 14170 5500
rect 14350 5440 14830 5500
rect 15010 5440 20910 5500
rect 1410 5430 1420 5440
rect 2500 5430 2700 5440
rect 3160 5430 3360 5440
rect 3820 5430 4020 5440
rect 4700 5430 4900 5440
rect 5360 5430 5560 5440
rect 6020 5430 6220 5440
rect 6900 5430 7100 5440
rect 7560 5430 7760 5440
rect 8220 5430 8420 5440
rect 9100 5430 9300 5440
rect 9760 5430 9960 5440
rect 10420 5430 10620 5440
rect 11300 5430 11500 5440
rect 11960 5430 12160 5440
rect 12620 5430 12820 5440
rect 13500 5430 13700 5440
rect 14160 5430 14360 5440
rect 14820 5430 15020 5440
rect 15700 5430 15900 5440
rect 16360 5430 16560 5440
rect 17020 5430 17220 5440
rect 17900 5430 18100 5440
rect 18560 5430 18760 5440
rect 19220 5430 19420 5440
rect 20900 5430 20910 5440
rect 21090 5500 21100 5510
rect 32550 5510 32630 5520
rect 21090 5440 22180 5500
rect 21090 5430 21100 5440
rect 1220 5420 1420 5430
rect 20900 5420 21100 5430
rect 28490 5400 28670 5410
rect -110 5340 30 5360
rect -110 5090 -80 5340
rect 0 5090 30 5340
rect -110 5060 30 5090
rect 2090 5340 2230 5360
rect 2090 5090 2120 5340
rect 2200 5090 2230 5340
rect 2090 5060 2230 5090
rect 4290 5340 4430 5360
rect 4290 5090 4320 5340
rect 4400 5090 4430 5340
rect 4290 5060 4430 5090
rect 6490 5340 6630 5360
rect 6490 5090 6520 5340
rect 6600 5090 6630 5340
rect 6490 5060 6630 5090
rect 8690 5340 8830 5360
rect 8690 5090 8720 5340
rect 8800 5090 8830 5340
rect 8690 5060 8830 5090
rect 10890 5340 11030 5360
rect 10890 5090 10920 5340
rect 11000 5090 11030 5340
rect 10890 5060 11030 5090
rect 13090 5340 13230 5360
rect 13090 5090 13120 5340
rect 13200 5090 13230 5340
rect 13090 5060 13230 5090
rect 15290 5340 15430 5360
rect 15290 5090 15320 5340
rect 15400 5090 15430 5340
rect 15290 5060 15430 5090
rect 17490 5340 17630 5360
rect 17490 5090 17520 5340
rect 17600 5090 17630 5340
rect 17490 5060 17630 5090
rect 19690 5340 19830 5360
rect 19690 5090 19720 5340
rect 19800 5090 19830 5340
rect 19690 5060 19830 5090
rect 21890 5340 22030 5360
rect 21890 5090 21920 5340
rect 22000 5090 22030 5340
rect 28490 5240 28500 5400
rect 28660 5370 28670 5400
rect 32550 5370 32560 5510
rect 28660 5280 32560 5370
rect 32620 5280 32630 5510
rect 36290 5370 36400 5380
rect 28660 5270 32630 5280
rect 33320 5290 33640 5300
rect 28660 5240 28670 5270
rect 28490 5230 28670 5240
rect 21890 5060 22030 5090
rect 30030 5170 30330 5180
rect 33320 5170 33330 5290
rect 30030 5070 30040 5170
rect 30320 5070 33330 5170
rect 30030 5060 33330 5070
rect 33320 5020 33330 5060
rect 33630 5020 33640 5290
rect 36290 5040 36300 5370
rect 36390 5250 36400 5370
rect 37670 5370 37780 5380
rect 36860 5320 37020 5330
rect 36860 5250 36870 5320
rect 36390 5170 36870 5250
rect 36390 5040 36400 5170
rect 36860 5100 36870 5170
rect 37010 5100 37020 5320
rect 36860 5090 37020 5100
rect 37120 5320 37280 5330
rect 37120 5100 37130 5320
rect 37270 5250 37280 5320
rect 37670 5250 37680 5370
rect 37270 5170 37680 5250
rect 37270 5100 37280 5170
rect 37120 5090 37280 5100
rect 36290 5030 36400 5040
rect 37670 5040 37680 5170
rect 37770 5040 37780 5370
rect 37670 5030 37780 5040
rect 2500 5010 4020 5020
rect 1620 4990 1820 5000
rect 1620 4980 1630 4990
rect 1600 4920 1630 4980
rect 1620 4910 1630 4920
rect 1810 4980 1820 4990
rect 2500 4980 2510 5010
rect 1810 4950 2510 4980
rect 4010 4980 4020 5010
rect 4700 5010 6220 5020
rect 4700 4980 4710 5010
rect 4010 4950 4710 4980
rect 6210 4980 6220 5010
rect 6900 5010 8420 5020
rect 6900 4980 6910 5010
rect 6210 4950 6910 4980
rect 8410 4980 8420 5010
rect 9100 5010 10620 5020
rect 9100 4980 9110 5010
rect 8410 4950 9110 4980
rect 10610 4980 10620 5010
rect 11300 5010 12820 5020
rect 11300 4980 11310 5010
rect 10610 4950 11310 4980
rect 12810 4980 12820 5010
rect 13500 5010 15020 5020
rect 13500 4980 13510 5010
rect 12810 4950 13510 4980
rect 15010 4980 15020 5010
rect 15700 5010 17220 5020
rect 15700 4980 15710 5010
rect 15010 4950 15710 4980
rect 17210 4980 17220 5010
rect 17900 5010 19420 5020
rect 33320 5010 33640 5020
rect 17900 4980 17910 5010
rect 17210 4950 17910 4980
rect 19410 4980 19420 5010
rect 20100 4990 20300 5000
rect 20100 4980 20110 4990
rect 19410 4950 20110 4980
rect 1810 4920 20110 4950
rect 1810 4910 1820 4920
rect 1620 4900 1820 4910
rect 20100 4910 20110 4920
rect 20290 4980 20300 4990
rect 20290 4920 20320 4980
rect 23040 4970 23590 4980
rect 20290 4910 20300 4920
rect 20100 4900 20300 4910
rect 23040 4710 23050 4970
rect 23580 4940 23590 4970
rect 23580 4930 27440 4940
rect 23580 4750 27250 4930
rect 27430 4750 27440 4930
rect 23580 4710 23590 4750
rect 27240 4740 27440 4750
rect 32400 4880 32480 4890
rect 23040 4700 23590 4710
rect 29760 4710 30560 4720
rect 32400 4710 32410 4880
rect 29760 4640 29770 4710
rect 30550 4650 32410 4710
rect 32470 4650 32480 4880
rect 30550 4640 32480 4650
rect 29760 4630 30560 4640
rect -300 4530 27560 4540
rect -300 4350 1290 4530
rect 1470 4350 20110 4530
rect 20290 4350 27370 4530
rect 27550 4350 27560 4530
rect -300 4340 27560 4350
rect 29130 4520 29210 4530
rect 29130 4290 29140 4520
rect 29200 4410 29210 4520
rect 32490 4480 32650 4490
rect 32490 4410 32500 4480
rect 29200 4340 32500 4410
rect 32640 4410 32650 4480
rect 34080 4480 34240 4490
rect 34080 4410 34090 4480
rect 32640 4340 34090 4410
rect 34230 4340 34240 4480
rect 29200 4290 29210 4340
rect 32490 4330 32650 4340
rect 34080 4330 34240 4340
rect 29130 4280 29210 4290
rect 35690 4290 35850 4300
rect 29270 4260 29520 4270
rect 35690 4260 35700 4290
rect 29270 4190 29280 4260
rect 29510 4190 35700 4260
rect 29270 4180 29520 4190
rect 35690 4150 35700 4190
rect 35840 4150 35850 4290
rect 35690 4140 35850 4150
rect -300 4130 27820 4140
rect -300 3950 1630 4130
rect 1810 3950 20450 4130
rect 20630 3950 27630 4130
rect 27810 3950 27820 4130
rect 33120 4110 33300 4120
rect -300 3940 27820 3950
rect 30070 4040 30270 4050
rect 30070 3860 30080 4040
rect 30260 3860 30270 4040
rect 30070 3850 30270 3860
rect 31670 4040 31870 4050
rect 31670 3860 31680 4040
rect 31860 3860 31870 4040
rect 33120 4010 33130 4110
rect 33290 4010 33300 4110
rect 33120 4000 33300 4010
rect 34860 4090 35200 4100
rect 34860 4010 34870 4090
rect 35190 4010 35200 4090
rect 34860 4000 35200 4010
rect 31670 3850 31870 3860
rect 32070 3740 32220 3750
rect -300 3730 31700 3740
rect -300 3550 430 3730
rect 610 3550 21310 3730
rect 21490 3550 31530 3730
rect 31690 3550 31700 3730
rect 32070 3610 32080 3740
rect 32210 3720 32220 3740
rect 32210 3710 38020 3720
rect 32210 3620 37880 3710
rect 32210 3610 32220 3620
rect 32070 3600 32220 3610
rect 37870 3580 37880 3620
rect 38010 3580 38020 3710
rect 37870 3570 38020 3580
rect -300 3540 31700 3550
rect 26200 3400 26380 3410
rect 26200 3370 26210 3400
rect 1160 3330 20300 3340
rect 1160 3150 1170 3330
rect 1330 3150 1630 3330
rect 1810 3150 2770 3330
rect 2930 3150 4370 3330
rect 4530 3150 5970 3330
rect 6130 3150 7570 3330
rect 7730 3150 9170 3330
rect 9330 3150 20110 3330
rect 20290 3150 20300 3330
rect 1160 3140 20300 3150
rect 20700 3270 26210 3370
rect 14180 3030 14360 3040
rect 10880 3010 11040 3020
rect 7800 2930 7940 2940
rect 7800 2810 7810 2930
rect 7930 2810 7940 2930
rect 10880 2870 10890 3010
rect 11030 3000 11040 3010
rect 14180 3000 14190 3030
rect 11030 2880 14190 3000
rect 11030 2870 11040 2880
rect 10880 2860 11040 2870
rect 14180 2870 14190 2880
rect 14350 2870 14360 3030
rect 14180 2860 14360 2870
rect 18050 3010 18210 3020
rect 18050 2870 18060 3010
rect 18200 2990 18210 3010
rect 20700 2990 20800 3270
rect 26200 3240 26210 3270
rect 26370 3370 26380 3400
rect 26370 3270 26410 3370
rect 26610 3360 26770 3370
rect 26370 3240 26380 3270
rect 26200 3230 26380 3240
rect 26610 3220 26620 3360
rect 26760 3340 26770 3360
rect 36580 3360 36740 3370
rect 36580 3340 36590 3360
rect 26760 3240 36590 3340
rect 26760 3220 26770 3240
rect 26610 3210 26770 3220
rect 36580 3220 36590 3240
rect 36730 3220 36740 3360
rect 36580 3210 36740 3220
rect 18200 2890 20800 2990
rect 23210 3090 32000 3100
rect 23210 2910 23220 3090
rect 23400 2910 31830 3090
rect 31990 2910 32000 3090
rect 23210 2900 32000 2910
rect 18200 2870 18210 2890
rect 18050 2860 18210 2870
rect 7800 2790 7940 2810
rect 16900 2780 17140 2790
rect 11690 2770 11850 2780
rect 11690 2620 11700 2770
rect 11840 2760 11850 2770
rect 16900 2760 16910 2780
rect 11840 2640 16910 2760
rect 17130 2760 17140 2780
rect 17370 2780 17500 2790
rect 17370 2760 17380 2780
rect 17130 2640 17380 2760
rect 17490 2760 17500 2780
rect 17730 2780 17970 2790
rect 17730 2760 17740 2780
rect 17490 2640 17740 2760
rect 17960 2760 17970 2780
rect 34770 2780 34940 2790
rect 34770 2760 34780 2780
rect 17960 2640 34780 2760
rect 11840 2630 34780 2640
rect 11840 2620 11850 2630
rect 11690 2610 11850 2620
rect 34770 2620 34780 2630
rect 34930 2620 34940 2780
rect 34770 2610 34940 2620
rect 33170 2550 33340 2560
rect 10990 2540 11150 2550
rect 10990 2530 11000 2540
rect 530 2400 11000 2530
rect 11140 2530 11150 2540
rect 12590 2540 12750 2550
rect 12590 2530 12600 2540
rect 11140 2400 12600 2530
rect 12740 2530 12750 2540
rect 13970 2540 14130 2550
rect 13970 2530 13980 2540
rect 12740 2400 13980 2530
rect 14120 2400 14130 2540
rect 33170 2530 33180 2550
rect 10990 2390 11150 2400
rect 12590 2390 12750 2400
rect 13970 2390 14130 2400
rect 14900 2400 33180 2530
rect 2090 2250 13440 2260
rect 470 2220 670 2240
rect 470 -4780 480 2220
rect 660 -4780 670 2220
rect 2090 2090 2110 2250
rect 2230 2090 3710 2250
rect 3830 2090 5310 2250
rect 5430 2090 6910 2250
rect 7030 2090 8510 2250
rect 8630 2090 10110 2250
rect 10230 2090 11710 2250
rect 11830 2090 13310 2250
rect 13430 2090 13440 2250
rect 2090 2080 13440 2090
rect 14900 1980 15040 2400
rect 33170 2390 33180 2400
rect 33330 2390 33340 2550
rect 33170 2380 33340 2390
rect 16500 2250 26240 2260
rect 16500 2090 16510 2250
rect 16630 2090 18110 2250
rect 18230 2090 19710 2250
rect 19830 2090 21310 2250
rect 21430 2090 22910 2250
rect 23030 2090 24510 2250
rect 24630 2090 26110 2250
rect 26230 2090 26240 2250
rect 16500 2080 26240 2090
rect 27700 2250 31040 2260
rect 27700 2070 27710 2250
rect 27830 2070 29310 2250
rect 29430 2070 30910 2250
rect 31030 2070 31040 2250
rect 27700 2060 31040 2070
rect 14900 1320 14910 1980
rect 15030 1320 15040 1980
rect 14900 1290 15040 1320
rect 32500 1150 32640 1160
rect 34100 1150 34240 1160
rect 34780 1150 34930 1160
rect 35700 1150 37440 1160
rect 32500 1030 32510 1150
rect 32630 1030 34110 1150
rect 34230 1030 34790 1150
rect 34920 1030 35710 1150
rect 35830 1030 37310 1150
rect 37430 1030 37440 1150
rect 32500 1020 32640 1030
rect 34100 1020 34240 1030
rect 34780 1020 34930 1030
rect 35700 1020 37440 1030
rect 2090 450 13440 460
rect 2090 290 2110 450
rect 2230 290 3710 450
rect 3830 290 5310 450
rect 5430 290 6910 450
rect 7030 290 8510 450
rect 8630 290 10110 450
rect 10230 290 11710 450
rect 11830 290 13310 450
rect 13430 290 13440 450
rect 2090 280 13440 290
rect 16500 450 26240 460
rect 16500 290 16510 450
rect 16630 290 18110 450
rect 18230 290 19710 450
rect 19830 290 21310 450
rect 21430 290 22910 450
rect 23030 290 24510 450
rect 24630 290 26110 450
rect 26230 290 26240 450
rect 16500 280 26240 290
rect 27700 450 31040 460
rect 27700 270 27710 450
rect 27830 270 29310 450
rect 29430 270 30910 450
rect 31030 270 31040 450
rect 27700 260 31040 270
rect 32500 440 35840 450
rect 32500 280 33180 440
rect 33330 280 35840 440
rect 32500 270 35840 280
rect 32500 190 32640 270
rect 32500 -490 32510 190
rect 32630 -490 32640 190
rect 32500 -500 32640 -490
rect 34100 190 34240 270
rect 34100 -490 34110 190
rect 34230 -490 34240 190
rect 34100 -500 34240 -490
rect 35700 190 35840 270
rect 35700 -490 35710 190
rect 35830 -490 35840 190
rect 35700 -500 35840 -490
rect 12870 -1110 13250 -1100
rect 12870 -1260 12880 -1110
rect 13240 -1260 13250 -1110
rect 12870 -1270 13250 -1260
rect 2090 -1350 15040 -1340
rect 2090 -1510 2110 -1350
rect 2230 -1510 3710 -1350
rect 3830 -1510 5310 -1350
rect 5430 -1510 6910 -1350
rect 7030 -1510 8510 -1350
rect 8630 -1510 10110 -1350
rect 10230 -1510 11710 -1350
rect 11830 -1510 13310 -1350
rect 13430 -1510 14910 -1350
rect 15030 -1510 15040 -1350
rect 2090 -1520 15040 -1510
rect 15240 -1350 26270 -1340
rect 15240 -1510 15250 -1350
rect 15370 -1510 16510 -1350
rect 16630 -1510 18110 -1350
rect 18230 -1510 19710 -1350
rect 19830 -1510 21310 -1350
rect 21430 -1510 22910 -1350
rect 23030 -1510 24510 -1350
rect 24630 -1510 26110 -1350
rect 26230 -1510 26270 -1350
rect 15240 -1520 26270 -1510
rect 27700 -1350 31040 -1340
rect 27700 -1530 27710 -1350
rect 27830 -1530 29310 -1350
rect 29430 -1530 30910 -1350
rect 31030 -1530 31040 -1350
rect 27700 -1540 31040 -1530
rect 32500 -2450 32640 -2440
rect 34100 -2450 34240 -2440
rect 34780 -2450 34930 -2440
rect 35700 -2450 35840 -2440
rect 32500 -2570 32510 -2450
rect 32630 -2570 34110 -2450
rect 34230 -2570 34790 -2450
rect 34920 -2570 35710 -2450
rect 35830 -2570 35840 -2450
rect 32500 -2580 32640 -2570
rect 34100 -2580 34240 -2570
rect 34780 -2580 34930 -2570
rect 35700 -2580 35840 -2570
rect 2090 -3150 15040 -3140
rect 2090 -3310 2110 -3150
rect 2230 -3310 3710 -3150
rect 3830 -3310 5310 -3150
rect 5430 -3310 6910 -3150
rect 7030 -3310 8510 -3150
rect 8630 -3310 10110 -3150
rect 10230 -3310 11710 -3150
rect 11830 -3310 13310 -3150
rect 13430 -3310 14910 -3150
rect 15030 -3310 15040 -3150
rect 2090 -3320 15040 -3310
rect 16500 -3150 26240 -3140
rect 16500 -3310 16510 -3150
rect 16630 -3310 18110 -3150
rect 18230 -3310 19710 -3150
rect 19830 -3310 21310 -3150
rect 21430 -3310 22910 -3150
rect 23030 -3310 24510 -3150
rect 24630 -3310 26110 -3150
rect 26230 -3310 26240 -3150
rect 16500 -3320 26240 -3310
rect 27700 -3150 31040 -3140
rect 27700 -3330 27710 -3150
rect 27830 -3330 29310 -3150
rect 29430 -3330 30910 -3150
rect 31030 -3330 31040 -3150
rect 27700 -3340 31040 -3330
rect 470 -4800 670 -4780
rect 680 -5170 37760 -5160
rect 680 -5350 2810 -5170
rect 2990 -5350 15570 -5170
rect 15730 -5350 18770 -5170
rect 18930 -5350 21280 -5170
rect 21460 -5350 21970 -5170
rect 22130 -5350 25170 -5170
rect 25330 -5350 28370 -5170
rect 28530 -5350 36030 -5170
rect 36210 -5350 37760 -5170
rect 680 -5360 37760 -5350
rect 680 -5570 37760 -5560
rect 680 -5750 1270 -5570
rect 1450 -5750 15570 -5570
rect 15730 -5750 18770 -5570
rect 18930 -5750 20510 -5570
rect 20690 -5750 21970 -5570
rect 22130 -5750 25170 -5570
rect 25330 -5750 28370 -5570
rect 28530 -5750 36230 -5570
rect 36410 -5750 37760 -5570
rect 680 -5760 37760 -5750
rect 15780 -5970 31990 -5960
rect 15780 -6150 15790 -5970
rect 15950 -6150 18990 -5970
rect 19150 -6150 22190 -5970
rect 22350 -6150 25390 -5970
rect 25550 -6150 27690 -5970
rect 27850 -6150 28590 -5970
rect 28750 -6150 29290 -5970
rect 29450 -6150 30890 -5970
rect 31050 -6150 31680 -5970
rect 31860 -6150 31990 -5970
rect 15780 -6160 31990 -6150
rect 14900 -6490 15040 -6480
rect 14900 -6610 14910 -6490
rect 15030 -6610 15040 -6490
rect 14900 -6620 15040 -6610
rect 17380 -6770 31990 -6760
rect 12940 -6830 13120 -6820
rect 12940 -6990 12950 -6830
rect 13110 -6990 13120 -6830
rect 17380 -6950 17390 -6770
rect 17550 -6950 20590 -6770
rect 20750 -6950 23790 -6770
rect 23950 -6950 26990 -6770
rect 27150 -6950 30080 -6770
rect 30350 -6950 31990 -6770
rect 17380 -6960 31990 -6950
rect 12940 -7000 13120 -6990
rect 680 -7170 37760 -7160
rect 680 -7350 1260 -7170
rect 1440 -7350 17170 -7170
rect 17330 -7350 20370 -7170
rect 20690 -7350 23570 -7170
rect 23730 -7350 26770 -7170
rect 26930 -7350 29970 -7170
rect 30130 -7350 36530 -7170
rect 36710 -7350 37760 -7170
rect 680 -7360 37760 -7350
rect 680 -7570 37760 -7560
rect 680 -7750 2080 -7570
rect 2260 -7750 17170 -7570
rect 17330 -7750 20370 -7570
rect 20530 -7750 22070 -7570
rect 22250 -7750 23570 -7570
rect 23730 -7750 26770 -7570
rect 26930 -7750 29970 -7570
rect 30130 -7750 36230 -7570
rect 36410 -7750 37760 -7570
rect 680 -7760 37760 -7750
rect 7800 -7870 7940 -7860
rect 7800 -7990 7810 -7870
rect 7930 -7990 7940 -7870
rect 7800 -8000 7940 -7990
rect 480 -8090 680 -8080
rect 480 -22380 490 -8090
rect 670 -22380 680 -8090
rect 10800 -8260 16650 -8250
rect 10800 -8380 10810 -8260
rect 10930 -8380 13310 -8260
rect 13440 -8380 16510 -8260
rect 16640 -8380 16650 -8260
rect 10800 -8390 16650 -8380
rect 16500 -9570 26250 -9560
rect 2120 -9590 10240 -9580
rect 2120 -9750 2130 -9590
rect 2230 -9750 3730 -9590
rect 3830 -9750 5330 -9590
rect 5430 -9750 6930 -9590
rect 7030 -9750 8530 -9590
rect 8630 -9750 10130 -9590
rect 10230 -9750 10240 -9590
rect 16500 -9730 16510 -9570
rect 16640 -9730 18110 -9570
rect 18240 -9730 19710 -9570
rect 19840 -9730 21310 -9570
rect 21440 -9730 22910 -9570
rect 23040 -9730 24510 -9570
rect 24640 -9730 26110 -9570
rect 26240 -9730 26250 -9570
rect 16500 -9740 26250 -9730
rect 27700 -9570 35850 -9560
rect 27700 -9730 27710 -9570
rect 27840 -9730 29310 -9570
rect 29440 -9730 30910 -9570
rect 31040 -9730 32510 -9570
rect 32640 -9730 34110 -9570
rect 34240 -9730 35710 -9570
rect 35840 -9730 35850 -9570
rect 27700 -9740 35850 -9730
rect 2120 -9760 10240 -9750
rect 16500 -11370 26250 -11360
rect 2120 -11390 10240 -11380
rect 2120 -11550 2130 -11390
rect 2230 -11550 3730 -11390
rect 3830 -11550 5330 -11390
rect 5430 -11550 6930 -11390
rect 7030 -11550 8530 -11390
rect 8630 -11550 10130 -11390
rect 10230 -11550 10240 -11390
rect 16500 -11530 16510 -11370
rect 16640 -11530 18110 -11370
rect 18240 -11530 19710 -11370
rect 19840 -11530 21310 -11370
rect 21440 -11530 22910 -11370
rect 23040 -11530 24510 -11370
rect 24640 -11530 26110 -11370
rect 26240 -11530 26250 -11370
rect 16500 -11540 26250 -11530
rect 27700 -11370 35850 -11360
rect 27700 -11530 27710 -11370
rect 27840 -11530 29310 -11370
rect 29440 -11530 30910 -11370
rect 31040 -11530 32510 -11370
rect 32640 -11530 34110 -11370
rect 34240 -11530 35710 -11370
rect 35840 -11530 35850 -11370
rect 27700 -11540 35850 -11530
rect 2120 -11560 10240 -11550
rect 13280 -13170 26250 -13160
rect 2120 -13190 10240 -13180
rect 2120 -13350 2130 -13190
rect 2230 -13350 3730 -13190
rect 3830 -13350 5330 -13190
rect 5430 -13350 6930 -13190
rect 7030 -13350 8530 -13190
rect 8630 -13350 10130 -13190
rect 10230 -13350 10240 -13190
rect 2120 -13360 10240 -13350
rect 13280 -13330 13290 -13170
rect 13460 -13330 14890 -13170
rect 15060 -13330 16510 -13170
rect 16640 -13330 18110 -13170
rect 18240 -13330 19710 -13170
rect 19840 -13330 21310 -13170
rect 21440 -13330 22910 -13170
rect 23040 -13330 24510 -13170
rect 24640 -13330 26110 -13170
rect 26240 -13330 26250 -13170
rect 13280 -13340 26250 -13330
rect 27700 -13170 35850 -13160
rect 27700 -13330 27710 -13170
rect 27840 -13330 29310 -13170
rect 29440 -13330 30910 -13170
rect 31040 -13330 32510 -13170
rect 32640 -13330 34110 -13170
rect 34240 -13330 35710 -13170
rect 35840 -13330 35850 -13170
rect 27700 -13340 35850 -13330
rect 13280 -13360 15070 -13340
rect 13280 -14970 26250 -14960
rect 2120 -14990 10240 -14980
rect 2120 -15150 2130 -14990
rect 2230 -15150 3730 -14990
rect 3830 -15150 5330 -14990
rect 5430 -15150 6930 -14990
rect 7030 -15150 8530 -14990
rect 8630 -15150 10130 -14990
rect 10230 -15150 10240 -14990
rect 2120 -15160 10240 -15150
rect 13280 -15130 13290 -14970
rect 13460 -15130 14890 -14970
rect 15060 -15130 16510 -14970
rect 16640 -15130 18110 -14970
rect 18240 -15130 19710 -14970
rect 19840 -15130 21310 -14970
rect 21440 -15130 22910 -14970
rect 23040 -15130 24510 -14970
rect 24640 -15130 26110 -14970
rect 26240 -15130 26250 -14970
rect 13280 -15140 26250 -15130
rect 27700 -14970 31050 -14960
rect 27700 -15130 27710 -14970
rect 27840 -15130 29310 -14970
rect 29440 -15130 30910 -14970
rect 31040 -15130 31050 -14970
rect 27700 -15140 31050 -15130
rect 13280 -15160 15070 -15140
rect 16500 -16770 26250 -16760
rect 2120 -16790 15090 -16780
rect 2120 -16950 2130 -16790
rect 2230 -16950 3730 -16790
rect 3830 -16950 5330 -16790
rect 5430 -16950 6930 -16790
rect 7030 -16950 8530 -16790
rect 8630 -16950 10130 -16790
rect 10230 -16950 13300 -16790
rect 13450 -16950 14900 -16790
rect 15050 -16950 15090 -16790
rect 16500 -16930 16510 -16770
rect 16640 -16930 18110 -16770
rect 18240 -16930 19710 -16770
rect 19840 -16930 21310 -16770
rect 21440 -16930 22910 -16770
rect 23040 -16930 24510 -16770
rect 24640 -16930 26110 -16770
rect 26240 -16930 26250 -16770
rect 16500 -16940 26250 -16930
rect 27700 -16770 31050 -16760
rect 27700 -16930 27710 -16770
rect 27840 -16930 29310 -16770
rect 29440 -16930 30910 -16770
rect 31040 -16930 31050 -16770
rect 32510 -16770 35840 -16760
rect 32510 -16920 32520 -16770
rect 32630 -16920 34120 -16770
rect 34230 -16920 34910 -16770
rect 35050 -16920 35720 -16770
rect 35830 -16920 35840 -16770
rect 32510 -16930 35840 -16920
rect 27700 -16940 31050 -16930
rect 2120 -16960 15090 -16950
rect 16500 -18570 26250 -18560
rect 2120 -18590 15060 -18580
rect 2120 -18750 2130 -18590
rect 2230 -18750 3730 -18590
rect 3830 -18750 5330 -18590
rect 5430 -18750 6930 -18590
rect 7030 -18750 8530 -18590
rect 8630 -18750 10130 -18590
rect 10230 -18750 13300 -18590
rect 13450 -18750 14900 -18590
rect 15050 -18750 15060 -18590
rect 16500 -18730 16510 -18570
rect 16640 -18730 18110 -18570
rect 18240 -18730 19710 -18570
rect 19840 -18730 21310 -18570
rect 21440 -18730 22910 -18570
rect 23040 -18730 24510 -18570
rect 24640 -18730 26110 -18570
rect 26240 -18730 26250 -18570
rect 16500 -18740 26250 -18730
rect 27700 -18570 31050 -18560
rect 27700 -18730 27710 -18570
rect 27840 -18730 29310 -18570
rect 29440 -18730 30910 -18570
rect 31040 -18730 31050 -18570
rect 27700 -18740 31050 -18730
rect 2120 -18760 15060 -18750
rect 16500 -20370 26250 -20360
rect 2120 -20390 10240 -20380
rect 2120 -20550 2130 -20390
rect 2230 -20550 3730 -20390
rect 3830 -20550 5330 -20390
rect 5430 -20550 6930 -20390
rect 7030 -20550 8530 -20390
rect 8630 -20550 10130 -20390
rect 10230 -20550 10240 -20390
rect 16500 -20530 16510 -20370
rect 16640 -20530 18110 -20370
rect 18240 -20530 19710 -20370
rect 19840 -20530 21310 -20370
rect 21440 -20530 22910 -20370
rect 23040 -20530 24510 -20370
rect 24640 -20530 26110 -20370
rect 26240 -20530 26250 -20370
rect 16500 -20540 26250 -20530
rect 27700 -20370 35860 -20360
rect 27700 -20530 27710 -20370
rect 27840 -20530 29310 -20370
rect 29440 -20530 30910 -20370
rect 31040 -20530 32510 -20370
rect 32640 -20530 34110 -20370
rect 34240 -20530 35710 -20370
rect 35840 -20530 35860 -20370
rect 27700 -20540 35860 -20530
rect 2120 -20560 10240 -20550
rect 16500 -22170 26250 -22160
rect 2120 -22190 10240 -22180
rect 2120 -22350 2130 -22190
rect 2230 -22350 3730 -22190
rect 3830 -22350 5330 -22190
rect 5430 -22350 6930 -22190
rect 7030 -22350 8530 -22190
rect 8630 -22350 10130 -22190
rect 10230 -22350 10240 -22190
rect 16500 -22330 16510 -22170
rect 16640 -22330 18110 -22170
rect 18240 -22330 19710 -22170
rect 19840 -22330 21310 -22170
rect 21440 -22330 22910 -22170
rect 23040 -22330 24510 -22170
rect 24640 -22330 26110 -22170
rect 26240 -22330 26250 -22170
rect 16500 -22340 26250 -22330
rect 27700 -22170 31050 -22160
rect 27700 -22330 27710 -22170
rect 27840 -22330 29310 -22170
rect 29440 -22330 30910 -22170
rect 31040 -22330 31050 -22170
rect 27700 -22340 31050 -22330
rect 2120 -22360 10240 -22350
rect 480 -22400 680 -22380
rect 10120 -22440 10240 -22360
rect 10100 -22450 10260 -22440
rect 10100 -22590 10110 -22450
rect 10250 -22460 10260 -22450
rect 10250 -22470 35120 -22460
rect 10250 -22590 34910 -22470
rect 10100 -22600 10260 -22590
rect 34900 -22610 34910 -22590
rect 35050 -22590 35120 -22470
rect 35050 -22610 35060 -22590
rect 34900 -22620 35060 -22610
rect 28140 -22730 28380 -22720
rect 28990 -22730 29230 -22720
rect 11040 -22740 28150 -22730
rect 11040 -22850 11050 -22740
rect 11150 -22850 11720 -22740
rect 11820 -22850 27720 -22740
rect 27830 -22850 28150 -22740
rect 11040 -22860 28150 -22850
rect 28140 -22870 28150 -22860
rect 28370 -22740 29000 -22730
rect 28370 -22860 28630 -22740
rect 28370 -22870 28380 -22860
rect 28140 -22880 28380 -22870
rect 28620 -22870 28630 -22860
rect 28740 -22860 29000 -22740
rect 28740 -22870 28750 -22860
rect 28620 -22880 28750 -22870
rect 28990 -22870 29000 -22860
rect 29220 -22740 31040 -22730
rect 29220 -22850 29320 -22740
rect 29430 -22850 30920 -22740
rect 31030 -22850 31040 -22740
rect 29220 -22860 31040 -22850
rect 29220 -22870 29230 -22860
rect 28990 -22880 29230 -22870
rect 12410 -22980 26720 -22970
rect 12410 -23090 12420 -22980
rect 12520 -23090 26530 -22980
rect 12410 -23100 26530 -23090
rect 26520 -23160 26530 -23100
rect 26710 -23160 26720 -22980
rect 26520 -23170 26720 -23160
rect -300 -23270 20300 -23260
rect -300 -23450 1190 -23270
rect 1350 -23450 1630 -23270
rect 1810 -23450 2790 -23270
rect 2950 -23450 4390 -23270
rect 4550 -23450 5990 -23270
rect 6150 -23450 7590 -23270
rect 7750 -23450 9190 -23270
rect 9350 -23450 20110 -23270
rect 20290 -23450 20300 -23270
rect -300 -23460 20300 -23450
rect 23200 -23300 23400 -23290
rect 23200 -23480 23210 -23300
rect 23390 -23330 23400 -23300
rect 31550 -23300 31750 -23290
rect 31550 -23330 31560 -23300
rect 23390 -23460 31560 -23330
rect 23390 -23480 23400 -23460
rect 23200 -23490 23400 -23480
rect 31550 -23480 31560 -23460
rect 31740 -23480 31750 -23300
rect 31550 -23490 31750 -23480
rect -300 -23670 32010 -23660
rect -300 -23850 430 -23670
rect 610 -23850 21310 -23670
rect 21490 -23850 31820 -23670
rect 32000 -23850 32010 -23670
rect -300 -23860 32010 -23850
rect 28490 -24040 28670 -24030
rect -300 -24070 27820 -24060
rect -300 -24250 1630 -24070
rect 1810 -24250 20450 -24070
rect 20630 -24250 27630 -24070
rect 27810 -24250 27820 -24070
rect 28490 -24200 28500 -24040
rect 28660 -24200 28670 -24040
rect 28490 -24210 28670 -24200
rect 29970 -24140 30050 -24130
rect -300 -24260 27820 -24250
rect 29970 -24370 29980 -24140
rect 30040 -24210 30050 -24140
rect 30040 -24220 37030 -24210
rect 30040 -24280 34620 -24220
rect 34770 -24280 34990 -24220
rect 37020 -24280 37030 -24220
rect 30040 -24370 30050 -24280
rect 34610 -24290 37030 -24280
rect 29970 -24380 30050 -24370
rect -300 -24470 27590 -24460
rect -300 -24650 1290 -24470
rect 1470 -24650 20110 -24470
rect 20290 -24650 27400 -24470
rect 27580 -24650 27590 -24470
rect 32790 -24480 33040 -24470
rect -300 -24660 27590 -24650
rect 29370 -24490 32800 -24480
rect 29370 -24720 29380 -24490
rect 29440 -24550 32800 -24490
rect 33030 -24550 33040 -24480
rect 29440 -24720 29450 -24550
rect 32790 -24560 33040 -24550
rect 34110 -24630 34360 -24620
rect 29370 -24730 29450 -24720
rect 29520 -24640 34120 -24630
rect 23030 -24820 23570 -24810
rect 1620 -25030 1820 -25020
rect 1620 -25040 1630 -25030
rect 1600 -25100 1630 -25040
rect 1620 -25110 1630 -25100
rect 1810 -25040 1820 -25030
rect 20100 -25030 20300 -25020
rect 20100 -25040 20110 -25030
rect 1810 -25070 20110 -25040
rect 1810 -25100 2510 -25070
rect 1810 -25110 1820 -25100
rect 1620 -25120 1820 -25110
rect 2500 -25130 2510 -25100
rect 4010 -25100 4710 -25070
rect 4010 -25130 4020 -25100
rect 2500 -25140 4020 -25130
rect 4700 -25130 4710 -25100
rect 6210 -25100 6910 -25070
rect 6210 -25130 6220 -25100
rect 4700 -25140 6220 -25130
rect 6900 -25130 6910 -25100
rect 8410 -25100 9110 -25070
rect 8410 -25130 8420 -25100
rect 6900 -25140 8420 -25130
rect 9100 -25130 9110 -25100
rect 10610 -25100 11310 -25070
rect 10610 -25130 10620 -25100
rect 9100 -25140 10620 -25130
rect 11300 -25130 11310 -25100
rect 12810 -25100 13510 -25070
rect 12810 -25130 12820 -25100
rect 11300 -25140 12820 -25130
rect 13500 -25130 13510 -25100
rect 15010 -25100 15710 -25070
rect 15010 -25130 15020 -25100
rect 13500 -25140 15020 -25130
rect 15700 -25130 15710 -25100
rect 17210 -25100 17910 -25070
rect 17210 -25130 17220 -25100
rect 15700 -25140 17220 -25130
rect 17900 -25130 17910 -25100
rect 19410 -25100 20110 -25070
rect 19410 -25130 19420 -25100
rect 20100 -25110 20110 -25100
rect 20290 -25040 20300 -25030
rect 20290 -25100 20320 -25040
rect 23030 -25070 23040 -24820
rect 23560 -24880 23570 -24820
rect 29520 -24870 29530 -24640
rect 29590 -24700 34120 -24640
rect 34350 -24700 34360 -24630
rect 36860 -24640 37020 -24630
rect 36860 -24650 36870 -24640
rect 29590 -24870 29600 -24700
rect 34110 -24710 34360 -24700
rect 34800 -24660 36870 -24650
rect 30280 -24780 30520 -24770
rect 33550 -24780 33800 -24770
rect 30280 -24850 30290 -24780
rect 30510 -24850 33560 -24780
rect 33790 -24850 33800 -24780
rect 30280 -24860 30520 -24850
rect 33550 -24860 33800 -24850
rect 34800 -24860 34810 -24660
rect 34900 -24780 36870 -24660
rect 37010 -24780 37020 -24640
rect 34900 -24790 37020 -24780
rect 37120 -24640 37280 -24630
rect 37120 -24780 37130 -24640
rect 37270 -24780 37280 -24640
rect 37120 -24790 37280 -24780
rect 34900 -24860 34910 -24790
rect 34800 -24870 34910 -24860
rect 29520 -24880 29600 -24870
rect 23560 -24890 27440 -24880
rect 23560 -25070 27250 -24890
rect 27430 -25070 27440 -24890
rect 33020 -24930 33300 -24920
rect 23030 -25080 27440 -25070
rect 30120 -24940 33030 -24930
rect 20290 -25110 20300 -25100
rect 20100 -25120 20300 -25110
rect 17900 -25140 19420 -25130
rect 30120 -25170 30130 -24940
rect 30190 -25000 33030 -24940
rect 33290 -25000 33300 -24930
rect 30190 -25170 30200 -25000
rect 33020 -25010 33300 -25000
rect 33220 -25080 33500 -25070
rect 30120 -25180 30200 -25170
rect 30420 -25090 33230 -25080
rect 30420 -25320 30430 -25090
rect 30490 -25150 33230 -25090
rect 33490 -25150 33500 -25080
rect 30490 -25320 30500 -25150
rect 33220 -25160 33500 -25150
rect 30420 -25330 30500 -25320
rect 820 -25550 1020 -25540
rect 20500 -25550 20700 -25540
rect 820 -25560 830 -25550
rect -260 -25620 830 -25560
rect 820 -25630 830 -25620
rect 1010 -25560 1020 -25550
rect 2500 -25560 2700 -25550
rect 3160 -25560 3360 -25550
rect 3820 -25560 4020 -25550
rect 4700 -25560 4900 -25550
rect 5360 -25560 5560 -25550
rect 6020 -25560 6220 -25550
rect 6900 -25560 7100 -25550
rect 7560 -25560 7760 -25550
rect 8220 -25560 8420 -25550
rect 9100 -25560 9300 -25550
rect 9760 -25560 9960 -25550
rect 10420 -25560 10620 -25550
rect 11300 -25560 11500 -25550
rect 11960 -25560 12160 -25550
rect 12620 -25560 12820 -25550
rect 13500 -25560 13700 -25550
rect 14160 -25560 14360 -25550
rect 14820 -25560 15020 -25550
rect 15700 -25560 15900 -25550
rect 16360 -25560 16560 -25550
rect 17020 -25560 17220 -25550
rect 17900 -25560 18100 -25550
rect 18560 -25560 18760 -25550
rect 19220 -25560 19420 -25550
rect 20500 -25560 20510 -25550
rect 1010 -25620 6910 -25560
rect 7090 -25620 7570 -25560
rect 7750 -25620 8230 -25560
rect 8410 -25620 9110 -25560
rect 9290 -25620 9770 -25560
rect 9950 -25620 10430 -25560
rect 10610 -25620 11310 -25560
rect 11490 -25620 11970 -25560
rect 12150 -25620 12630 -25560
rect 12810 -25620 13510 -25560
rect 13690 -25620 14170 -25560
rect 14350 -25620 14830 -25560
rect 15010 -25620 20510 -25560
rect 1010 -25630 1020 -25620
rect 2500 -25630 2700 -25620
rect 3160 -25630 3360 -25620
rect 3820 -25630 4020 -25620
rect 4700 -25630 4900 -25620
rect 5360 -25630 5560 -25620
rect 6020 -25630 6220 -25620
rect 6900 -25630 7100 -25620
rect 7560 -25630 7760 -25620
rect 8220 -25630 8420 -25620
rect 9100 -25630 9300 -25620
rect 9760 -25630 9960 -25620
rect 10420 -25630 10620 -25620
rect 11300 -25630 11500 -25620
rect 11960 -25630 12160 -25620
rect 12620 -25630 12820 -25620
rect 13500 -25630 13700 -25620
rect 14160 -25630 14360 -25620
rect 14820 -25630 15020 -25620
rect 15700 -25630 15900 -25620
rect 16360 -25630 16560 -25620
rect 17020 -25630 17220 -25620
rect 17900 -25630 18100 -25620
rect 18560 -25630 18760 -25620
rect 19220 -25630 19420 -25620
rect 20500 -25630 20510 -25620
rect 20690 -25560 20700 -25550
rect 20690 -25620 22140 -25560
rect 20690 -25630 20700 -25620
rect 820 -25640 1020 -25630
rect 20500 -25640 20700 -25630
rect 1220 -25690 1420 -25680
rect 20900 -25690 21100 -25680
rect 1220 -25700 1230 -25690
rect -260 -25760 1230 -25700
rect 1220 -25770 1230 -25760
rect 1410 -25700 1420 -25690
rect 2500 -25700 2700 -25690
rect 3160 -25700 3360 -25690
rect 3820 -25700 4020 -25690
rect 4700 -25700 4900 -25690
rect 5360 -25700 5560 -25690
rect 6020 -25700 6220 -25690
rect 6900 -25700 7100 -25690
rect 7560 -25700 7760 -25690
rect 8220 -25700 8420 -25690
rect 9100 -25700 9300 -25690
rect 9760 -25700 9960 -25690
rect 10420 -25700 10620 -25690
rect 11300 -25700 11500 -25690
rect 11960 -25700 12160 -25690
rect 12620 -25700 12820 -25690
rect 13500 -25700 13700 -25690
rect 14160 -25700 14360 -25690
rect 14820 -25700 15020 -25690
rect 15700 -25700 15900 -25690
rect 16360 -25700 16560 -25690
rect 17020 -25700 17220 -25690
rect 17900 -25700 18100 -25690
rect 18560 -25700 18760 -25690
rect 19220 -25700 19420 -25690
rect 20900 -25700 20910 -25690
rect 1410 -25760 2510 -25700
rect 2690 -25760 3170 -25700
rect 3350 -25760 3830 -25700
rect 4010 -25760 4710 -25700
rect 4890 -25760 5370 -25700
rect 5550 -25760 6030 -25700
rect 6210 -25760 15710 -25700
rect 15890 -25760 16370 -25700
rect 16550 -25760 17030 -25700
rect 17210 -25760 17910 -25700
rect 18090 -25760 18570 -25700
rect 18750 -25760 19230 -25700
rect 19410 -25760 20910 -25700
rect 1410 -25770 1420 -25760
rect 2500 -25770 2700 -25760
rect 3160 -25770 3360 -25760
rect 3820 -25770 4020 -25760
rect 4700 -25770 4900 -25760
rect 5360 -25770 5560 -25760
rect 6020 -25770 6220 -25760
rect 6900 -25770 7100 -25760
rect 7560 -25770 7760 -25760
rect 8220 -25770 8420 -25760
rect 9100 -25770 9300 -25760
rect 9760 -25770 9960 -25760
rect 10420 -25770 10620 -25760
rect 11300 -25770 11500 -25760
rect 11960 -25770 12160 -25760
rect 12620 -25770 12820 -25760
rect 13500 -25770 13700 -25760
rect 14160 -25770 14360 -25760
rect 14820 -25770 15020 -25760
rect 15700 -25770 15900 -25760
rect 16360 -25770 16560 -25760
rect 17020 -25770 17220 -25760
rect 17900 -25770 18100 -25760
rect 18560 -25770 18760 -25760
rect 19220 -25770 19420 -25760
rect 20900 -25770 20910 -25760
rect 21090 -25700 21100 -25690
rect 21090 -25760 22140 -25700
rect 21090 -25770 21100 -25760
rect 1220 -25780 1420 -25770
rect 20900 -25780 21100 -25770
rect 1620 -25830 1820 -25820
rect 1620 -25840 1630 -25830
rect 1600 -25900 1630 -25840
rect 1620 -25910 1630 -25900
rect 1810 -25840 1820 -25830
rect 20100 -25830 20300 -25820
rect 20100 -25840 20110 -25830
rect 1810 -25870 20110 -25840
rect 1810 -25900 2510 -25870
rect 1810 -25910 1820 -25900
rect 1620 -25920 1820 -25910
rect 2500 -25930 2510 -25900
rect 4010 -25900 4710 -25870
rect 4010 -25930 4020 -25900
rect 2500 -25940 4020 -25930
rect 4700 -25930 4710 -25900
rect 6210 -25900 6910 -25870
rect 6210 -25930 6220 -25900
rect 4700 -25940 6220 -25930
rect 6900 -25930 6910 -25900
rect 8410 -25900 9110 -25870
rect 8410 -25930 8420 -25900
rect 6900 -25940 8420 -25930
rect 9100 -25930 9110 -25900
rect 10610 -25900 11310 -25870
rect 10610 -25930 10620 -25900
rect 9100 -25940 10620 -25930
rect 11300 -25930 11310 -25900
rect 12810 -25900 13510 -25870
rect 12810 -25930 12820 -25900
rect 11300 -25940 12820 -25930
rect 13500 -25930 13510 -25900
rect 15010 -25900 15710 -25870
rect 15010 -25930 15020 -25900
rect 13500 -25940 15020 -25930
rect 15700 -25930 15710 -25900
rect 17210 -25900 17910 -25870
rect 17210 -25930 17220 -25900
rect 15700 -25940 17220 -25930
rect 17900 -25930 17910 -25900
rect 19410 -25900 20110 -25870
rect 19410 -25930 19420 -25900
rect 20100 -25910 20110 -25900
rect 20290 -25840 20300 -25830
rect 20290 -25900 20320 -25840
rect 20290 -25910 20300 -25900
rect 20100 -25920 20300 -25910
rect 17900 -25940 19420 -25930
rect 820 -26350 1020 -26340
rect 20500 -26350 20700 -26340
rect 820 -26360 830 -26350
rect -260 -26420 830 -26360
rect 820 -26430 830 -26420
rect 1010 -26360 1020 -26350
rect 2500 -26360 2700 -26350
rect 3160 -26360 3360 -26350
rect 3820 -26360 4020 -26350
rect 4700 -26360 4900 -26350
rect 5360 -26360 5560 -26350
rect 6020 -26360 6220 -26350
rect 6900 -26360 7100 -26350
rect 7560 -26360 7760 -26350
rect 8220 -26360 8420 -26350
rect 9100 -26360 9300 -26350
rect 9760 -26360 9960 -26350
rect 10420 -26360 10620 -26350
rect 11300 -26360 11500 -26350
rect 11960 -26360 12160 -26350
rect 12620 -26360 12820 -26350
rect 13500 -26360 13700 -26350
rect 14160 -26360 14360 -26350
rect 14820 -26360 15020 -26350
rect 15700 -26360 15900 -26350
rect 16360 -26360 16560 -26350
rect 17020 -26360 17220 -26350
rect 17900 -26360 18100 -26350
rect 18560 -26360 18760 -26350
rect 19220 -26360 19420 -26350
rect 20500 -26360 20510 -26350
rect 1010 -26420 2510 -26360
rect 2690 -26420 3170 -26360
rect 3350 -26420 3830 -26360
rect 4010 -26420 4710 -26360
rect 4890 -26420 5370 -26360
rect 5550 -26420 6030 -26360
rect 6210 -26420 15710 -26360
rect 15890 -26420 16370 -26360
rect 16550 -26420 17030 -26360
rect 17210 -26420 17910 -26360
rect 18090 -26420 18570 -26360
rect 18750 -26420 19230 -26360
rect 19410 -26420 20510 -26360
rect 1010 -26430 1020 -26420
rect 2500 -26430 2700 -26420
rect 3160 -26430 3360 -26420
rect 3820 -26430 4020 -26420
rect 4700 -26430 4900 -26420
rect 5360 -26430 5560 -26420
rect 6020 -26430 6220 -26420
rect 6900 -26430 7100 -26420
rect 7560 -26430 7760 -26420
rect 8220 -26430 8420 -26420
rect 9100 -26430 9300 -26420
rect 9760 -26430 9960 -26420
rect 10420 -26430 10620 -26420
rect 11300 -26430 11500 -26420
rect 11960 -26430 12160 -26420
rect 12620 -26430 12820 -26420
rect 13500 -26430 13700 -26420
rect 14160 -26430 14360 -26420
rect 14820 -26430 15020 -26420
rect 15700 -26430 15900 -26420
rect 16360 -26430 16560 -26420
rect 17020 -26430 17220 -26420
rect 17900 -26430 18100 -26420
rect 18560 -26430 18760 -26420
rect 19220 -26430 19420 -26420
rect 20500 -26430 20510 -26420
rect 20690 -26360 20700 -26350
rect 20690 -26420 22140 -26360
rect 20690 -26430 20700 -26420
rect 820 -26440 1020 -26430
rect 20500 -26440 20700 -26430
rect 1220 -26490 1420 -26480
rect 20900 -26490 21100 -26480
rect 1220 -26500 1230 -26490
rect -260 -26560 1230 -26500
rect 1220 -26570 1230 -26560
rect 1410 -26500 1420 -26490
rect 2500 -26500 2700 -26490
rect 3160 -26500 3360 -26490
rect 3820 -26500 4020 -26490
rect 4700 -26500 4900 -26490
rect 5360 -26500 5560 -26490
rect 6020 -26500 6220 -26490
rect 6900 -26500 7100 -26490
rect 7560 -26500 7760 -26490
rect 8220 -26500 8420 -26490
rect 9100 -26500 9300 -26490
rect 9760 -26500 9960 -26490
rect 10420 -26500 10620 -26490
rect 11300 -26500 11500 -26490
rect 11960 -26500 12160 -26490
rect 12620 -26500 12820 -26490
rect 13500 -26500 13700 -26490
rect 14160 -26500 14360 -26490
rect 14820 -26500 15020 -26490
rect 15700 -26500 15900 -26490
rect 16360 -26500 16560 -26490
rect 17020 -26500 17220 -26490
rect 17900 -26500 18100 -26490
rect 18560 -26500 18760 -26490
rect 19220 -26500 19420 -26490
rect 20900 -26500 20910 -26490
rect 1410 -26560 6910 -26500
rect 7090 -26560 7570 -26500
rect 7750 -26560 8230 -26500
rect 8410 -26560 9110 -26500
rect 9290 -26560 9770 -26500
rect 9950 -26560 10430 -26500
rect 10610 -26560 11310 -26500
rect 11490 -26560 11970 -26500
rect 12150 -26560 12630 -26500
rect 12810 -26560 13510 -26500
rect 13690 -26560 14170 -26500
rect 14350 -26560 14830 -26500
rect 15010 -26560 20910 -26500
rect 1410 -26570 1420 -26560
rect 2500 -26570 2700 -26560
rect 3160 -26570 3360 -26560
rect 3820 -26570 4020 -26560
rect 4700 -26570 4900 -26560
rect 5360 -26570 5560 -26560
rect 6020 -26570 6220 -26560
rect 6900 -26570 7100 -26560
rect 7560 -26570 7760 -26560
rect 8220 -26570 8420 -26560
rect 9100 -26570 9300 -26560
rect 9760 -26570 9960 -26560
rect 10420 -26570 10620 -26560
rect 11300 -26570 11500 -26560
rect 11960 -26570 12160 -26560
rect 12620 -26570 12820 -26560
rect 13500 -26570 13700 -26560
rect 14160 -26570 14360 -26560
rect 14820 -26570 15020 -26560
rect 15700 -26570 15900 -26560
rect 16360 -26570 16560 -26560
rect 17020 -26570 17220 -26560
rect 17900 -26570 18100 -26560
rect 18560 -26570 18760 -26560
rect 19220 -26570 19420 -26560
rect 20900 -26570 20910 -26560
rect 21090 -26500 21100 -26490
rect 21090 -26560 22140 -26500
rect 21090 -26570 21100 -26560
rect 1220 -26580 1420 -26570
rect 20900 -26580 21100 -26570
rect 420 -26630 620 -26620
rect 420 -26710 430 -26630
rect 610 -26710 620 -26630
rect 1620 -26630 1820 -26620
rect 1620 -26640 1630 -26630
rect 1600 -26700 1630 -26640
rect 420 -26720 620 -26710
rect 1620 -26710 1630 -26700
rect 1810 -26640 1820 -26630
rect 20100 -26630 20300 -26620
rect 20100 -26640 20110 -26630
rect 1810 -26670 20110 -26640
rect 1810 -26700 4710 -26670
rect 1810 -26710 1820 -26700
rect 1620 -26720 1820 -26710
rect 4700 -26730 4710 -26700
rect 6210 -26700 6910 -26670
rect 6210 -26730 6220 -26700
rect 4700 -26740 6220 -26730
rect 6900 -26730 6910 -26700
rect 8410 -26700 9110 -26670
rect 8410 -26730 8420 -26700
rect 6900 -26740 8420 -26730
rect 9100 -26730 9110 -26700
rect 10610 -26700 11310 -26670
rect 10610 -26730 10620 -26700
rect 9100 -26740 10620 -26730
rect 11300 -26730 11310 -26700
rect 12810 -26700 13510 -26670
rect 12810 -26730 12820 -26700
rect 11300 -26740 12820 -26730
rect 13500 -26730 13510 -26700
rect 15010 -26700 15710 -26670
rect 15010 -26730 15020 -26700
rect 13500 -26740 15020 -26730
rect 15700 -26730 15710 -26700
rect 17210 -26700 20110 -26670
rect 17210 -26730 17220 -26700
rect 20100 -26710 20110 -26700
rect 20290 -26640 20300 -26630
rect 21300 -26630 21500 -26620
rect 20290 -26700 20320 -26640
rect 20290 -26710 20300 -26700
rect 20100 -26720 20300 -26710
rect 21300 -26710 21310 -26630
rect 21490 -26710 21500 -26630
rect 21300 -26720 21500 -26710
rect 15700 -26740 17220 -26730
rect 36020 -27010 36420 -27000
rect 36020 -27140 36030 -27010
rect 36410 -27140 36420 -27010
rect 820 -27150 1020 -27140
rect 20500 -27150 20700 -27140
rect 36020 -27150 36420 -27140
rect 36520 -27010 36920 -27000
rect 36520 -27140 36530 -27010
rect 36910 -27140 36920 -27010
rect 36520 -27150 36920 -27140
rect 820 -27160 830 -27150
rect -260 -27220 830 -27160
rect 820 -27230 830 -27220
rect 1010 -27160 1020 -27150
rect 2500 -27160 2700 -27150
rect 3160 -27160 3360 -27150
rect 3820 -27160 4020 -27150
rect 4700 -27160 4900 -27150
rect 5360 -27160 5560 -27150
rect 6020 -27160 6220 -27150
rect 6900 -27160 7100 -27150
rect 7560 -27160 7760 -27150
rect 8220 -27160 8420 -27150
rect 9100 -27160 9300 -27150
rect 9760 -27160 9960 -27150
rect 10420 -27160 10620 -27150
rect 11300 -27160 11500 -27150
rect 11960 -27160 12160 -27150
rect 12620 -27160 12820 -27150
rect 13500 -27160 13700 -27150
rect 14160 -27160 14360 -27150
rect 14820 -27160 15020 -27150
rect 15700 -27160 15900 -27150
rect 16360 -27160 16560 -27150
rect 17020 -27160 17220 -27150
rect 17900 -27160 18100 -27150
rect 18560 -27160 18760 -27150
rect 19220 -27160 19420 -27150
rect 20500 -27160 20510 -27150
rect 1010 -27220 6910 -27160
rect 7090 -27220 7570 -27160
rect 7750 -27220 8230 -27160
rect 8410 -27220 9110 -27160
rect 9290 -27220 9770 -27160
rect 9950 -27220 10430 -27160
rect 10610 -27220 11310 -27160
rect 11490 -27220 11970 -27160
rect 12150 -27220 12630 -27160
rect 12810 -27220 13510 -27160
rect 13690 -27220 14170 -27160
rect 14350 -27220 14830 -27160
rect 15010 -27220 20510 -27160
rect 1010 -27230 1020 -27220
rect 2500 -27230 2700 -27220
rect 3160 -27230 3360 -27220
rect 3820 -27230 4020 -27220
rect 4700 -27230 4900 -27220
rect 5360 -27230 5560 -27220
rect 6020 -27230 6220 -27220
rect 6900 -27230 7100 -27220
rect 7560 -27230 7760 -27220
rect 8220 -27230 8420 -27220
rect 9100 -27230 9300 -27220
rect 9760 -27230 9960 -27220
rect 10420 -27230 10620 -27220
rect 11300 -27230 11500 -27220
rect 11960 -27230 12160 -27220
rect 12620 -27230 12820 -27220
rect 13500 -27230 13700 -27220
rect 14160 -27230 14360 -27220
rect 14820 -27230 15020 -27220
rect 15700 -27230 15900 -27220
rect 16360 -27230 16560 -27220
rect 17020 -27230 17220 -27220
rect 17900 -27230 18100 -27220
rect 18560 -27230 18760 -27220
rect 19220 -27230 19420 -27220
rect 20500 -27230 20510 -27220
rect 20690 -27160 20700 -27150
rect 20690 -27220 22140 -27160
rect 20690 -27230 20700 -27220
rect 820 -27240 1020 -27230
rect 20500 -27240 20700 -27230
rect 1220 -27290 1420 -27280
rect 20900 -27290 21100 -27280
rect 1220 -27300 1230 -27290
rect -260 -27360 1230 -27300
rect 1220 -27370 1230 -27360
rect 1410 -27300 1420 -27290
rect 2500 -27300 2700 -27290
rect 3160 -27300 3360 -27290
rect 3820 -27300 4020 -27290
rect 4700 -27300 4900 -27290
rect 5360 -27300 5560 -27290
rect 6020 -27300 6220 -27290
rect 6900 -27300 7100 -27290
rect 7560 -27300 7760 -27290
rect 8220 -27300 8420 -27290
rect 9100 -27300 9300 -27290
rect 9760 -27300 9960 -27290
rect 10420 -27300 10620 -27290
rect 11300 -27300 11500 -27290
rect 11960 -27300 12160 -27290
rect 12620 -27300 12820 -27290
rect 13500 -27300 13700 -27290
rect 14160 -27300 14360 -27290
rect 14820 -27300 15020 -27290
rect 15700 -27300 15900 -27290
rect 16360 -27300 16560 -27290
rect 17020 -27300 17220 -27290
rect 17900 -27300 18100 -27290
rect 18560 -27300 18760 -27290
rect 19220 -27300 19420 -27290
rect 20900 -27300 20910 -27290
rect 1410 -27360 2510 -27300
rect 2690 -27360 3170 -27300
rect 3350 -27360 3830 -27300
rect 4010 -27360 4710 -27300
rect 4890 -27360 5370 -27300
rect 5550 -27360 6030 -27300
rect 6210 -27360 15710 -27300
rect 15890 -27360 16370 -27300
rect 16550 -27360 17030 -27300
rect 17210 -27360 17910 -27300
rect 18090 -27360 18570 -27300
rect 18750 -27360 19230 -27300
rect 19410 -27360 20910 -27300
rect 1410 -27370 1420 -27360
rect 2500 -27370 2700 -27360
rect 3160 -27370 3360 -27360
rect 3820 -27370 4020 -27360
rect 4700 -27370 4900 -27360
rect 5360 -27370 5560 -27360
rect 6020 -27370 6220 -27360
rect 6900 -27370 7100 -27360
rect 7560 -27370 7760 -27360
rect 8220 -27370 8420 -27360
rect 9100 -27370 9300 -27360
rect 9760 -27370 9960 -27360
rect 10420 -27370 10620 -27360
rect 11300 -27370 11500 -27360
rect 11960 -27370 12160 -27360
rect 12620 -27370 12820 -27360
rect 13500 -27370 13700 -27360
rect 14160 -27370 14360 -27360
rect 14820 -27370 15020 -27360
rect 15700 -27370 15900 -27360
rect 16360 -27370 16560 -27360
rect 17020 -27370 17220 -27360
rect 17900 -27370 18100 -27360
rect 18560 -27370 18760 -27360
rect 19220 -27370 19420 -27360
rect 20900 -27370 20910 -27360
rect 21090 -27300 21100 -27290
rect 21090 -27360 22140 -27300
rect 21090 -27370 21100 -27360
rect 1220 -27380 1420 -27370
rect 20900 -27380 21100 -27370
rect 420 -27430 620 -27420
rect 420 -27510 430 -27430
rect 610 -27510 620 -27430
rect 1620 -27430 1820 -27420
rect 1620 -27440 1630 -27430
rect 1600 -27500 1630 -27440
rect 420 -27520 620 -27510
rect 1620 -27510 1630 -27500
rect 1810 -27440 1820 -27430
rect 20100 -27430 20300 -27420
rect 20100 -27440 20110 -27430
rect 1810 -27470 20110 -27440
rect 1810 -27500 4710 -27470
rect 1810 -27510 1820 -27500
rect 1620 -27520 1820 -27510
rect 4700 -27530 4710 -27500
rect 6210 -27500 6910 -27470
rect 6210 -27530 6220 -27500
rect 4700 -27540 6220 -27530
rect 6900 -27530 6910 -27500
rect 8410 -27500 9110 -27470
rect 8410 -27530 8420 -27500
rect 6900 -27540 8420 -27530
rect 9100 -27530 9110 -27500
rect 10610 -27500 11310 -27470
rect 10610 -27530 10620 -27500
rect 9100 -27540 10620 -27530
rect 11300 -27530 11310 -27500
rect 12810 -27500 13510 -27470
rect 12810 -27530 12820 -27500
rect 11300 -27540 12820 -27530
rect 13500 -27530 13510 -27500
rect 15010 -27500 15710 -27470
rect 15010 -27530 15020 -27500
rect 13500 -27540 15020 -27530
rect 15700 -27530 15710 -27500
rect 17210 -27500 20110 -27470
rect 17210 -27530 17220 -27500
rect 20100 -27510 20110 -27500
rect 20290 -27440 20300 -27430
rect 21300 -27430 21500 -27420
rect 20290 -27500 20320 -27440
rect 20290 -27510 20300 -27500
rect 20100 -27520 20300 -27510
rect 21300 -27510 21310 -27430
rect 21490 -27510 21500 -27430
rect 21300 -27520 21500 -27510
rect 15700 -27540 17220 -27530
rect 33420 -27640 33600 -27620
rect 33420 -27780 33440 -27640
rect 33580 -27660 33600 -27640
rect 33580 -27760 38080 -27660
rect 33580 -27780 33600 -27760
rect 33420 -27800 33600 -27780
rect 35620 -27840 35800 -27820
rect 820 -27950 1020 -27940
rect 20500 -27950 20700 -27940
rect 820 -27960 830 -27950
rect -260 -28020 830 -27960
rect 820 -28030 830 -28020
rect 1010 -27960 1020 -27950
rect 2500 -27960 2700 -27950
rect 3160 -27960 3360 -27950
rect 3820 -27960 4020 -27950
rect 4700 -27960 4900 -27950
rect 5360 -27960 5560 -27950
rect 6020 -27960 6220 -27950
rect 6900 -27960 7100 -27950
rect 7560 -27960 7760 -27950
rect 8220 -27960 8420 -27950
rect 9100 -27960 9300 -27950
rect 9760 -27960 9960 -27950
rect 10420 -27960 10620 -27950
rect 11300 -27960 11500 -27950
rect 11960 -27960 12160 -27950
rect 12620 -27960 12820 -27950
rect 13500 -27960 13700 -27950
rect 14160 -27960 14360 -27950
rect 14820 -27960 15020 -27950
rect 15700 -27960 15900 -27950
rect 16360 -27960 16560 -27950
rect 17020 -27960 17220 -27950
rect 17900 -27960 18100 -27950
rect 18560 -27960 18760 -27950
rect 19220 -27960 19420 -27950
rect 20500 -27960 20510 -27950
rect 1010 -28020 2510 -27960
rect 2690 -28020 3170 -27960
rect 3350 -28020 3830 -27960
rect 4010 -28020 4710 -27960
rect 4890 -28020 5370 -27960
rect 5550 -28020 6030 -27960
rect 6210 -28020 15710 -27960
rect 15890 -28020 16370 -27960
rect 16550 -28020 17030 -27960
rect 17210 -28020 17910 -27960
rect 18090 -28020 18570 -27960
rect 18750 -28020 19230 -27960
rect 19410 -28020 20510 -27960
rect 1010 -28030 1020 -28020
rect 2500 -28030 2700 -28020
rect 3160 -28030 3360 -28020
rect 3820 -28030 4020 -28020
rect 4700 -28030 4900 -28020
rect 5360 -28030 5560 -28020
rect 6020 -28030 6220 -28020
rect 6900 -28030 7100 -28020
rect 7560 -28030 7760 -28020
rect 8220 -28030 8420 -28020
rect 9100 -28030 9300 -28020
rect 9760 -28030 9960 -28020
rect 10420 -28030 10620 -28020
rect 11300 -28030 11500 -28020
rect 11960 -28030 12160 -28020
rect 12620 -28030 12820 -28020
rect 13500 -28030 13700 -28020
rect 14160 -28030 14360 -28020
rect 14820 -28030 15020 -28020
rect 15700 -28030 15900 -28020
rect 16360 -28030 16560 -28020
rect 17020 -28030 17220 -28020
rect 17900 -28030 18100 -28020
rect 18560 -28030 18760 -28020
rect 19220 -28030 19420 -28020
rect 20500 -28030 20510 -28020
rect 20690 -27960 20700 -27950
rect 20690 -28020 22140 -27960
rect 35620 -27980 35640 -27840
rect 35780 -27860 35800 -27840
rect 35780 -27960 38080 -27860
rect 35780 -27980 35800 -27960
rect 35620 -28000 35800 -27980
rect 20690 -28030 20700 -28020
rect 820 -28040 1020 -28030
rect 20500 -28040 20700 -28030
rect 37720 -28040 37900 -28020
rect 31810 -28050 33170 -28040
rect 1220 -28090 1420 -28080
rect 20900 -28090 21100 -28080
rect 1220 -28100 1230 -28090
rect -260 -28160 1230 -28100
rect 1220 -28170 1230 -28160
rect 1410 -28100 1420 -28090
rect 2500 -28100 2700 -28090
rect 3160 -28100 3360 -28090
rect 3820 -28100 4020 -28090
rect 4700 -28100 4900 -28090
rect 5360 -28100 5560 -28090
rect 6020 -28100 6220 -28090
rect 6900 -28100 7100 -28090
rect 7560 -28100 7760 -28090
rect 8220 -28100 8420 -28090
rect 9100 -28100 9300 -28090
rect 9760 -28100 9960 -28090
rect 10420 -28100 10620 -28090
rect 11300 -28100 11500 -28090
rect 11960 -28100 12160 -28090
rect 12620 -28100 12820 -28090
rect 13500 -28100 13700 -28090
rect 14160 -28100 14360 -28090
rect 14820 -28100 15020 -28090
rect 15700 -28100 15900 -28090
rect 16360 -28100 16560 -28090
rect 17020 -28100 17220 -28090
rect 17900 -28100 18100 -28090
rect 18560 -28100 18760 -28090
rect 19220 -28100 19420 -28090
rect 20900 -28100 20910 -28090
rect 1410 -28160 6910 -28100
rect 7090 -28160 7570 -28100
rect 7750 -28160 8230 -28100
rect 8410 -28160 9110 -28100
rect 9290 -28160 9770 -28100
rect 9950 -28160 10430 -28100
rect 10610 -28160 11310 -28100
rect 11490 -28160 11970 -28100
rect 12150 -28160 12630 -28100
rect 12810 -28160 13510 -28100
rect 13690 -28160 14170 -28100
rect 14350 -28160 14830 -28100
rect 15010 -28160 20910 -28100
rect 1410 -28170 1420 -28160
rect 2500 -28170 2700 -28160
rect 3160 -28170 3360 -28160
rect 3820 -28170 4020 -28160
rect 4700 -28170 4900 -28160
rect 5360 -28170 5560 -28160
rect 6020 -28170 6220 -28160
rect 6900 -28170 7100 -28160
rect 7560 -28170 7760 -28160
rect 8220 -28170 8420 -28160
rect 9100 -28170 9300 -28160
rect 9760 -28170 9960 -28160
rect 10420 -28170 10620 -28160
rect 11300 -28170 11500 -28160
rect 11960 -28170 12160 -28160
rect 12620 -28170 12820 -28160
rect 13500 -28170 13700 -28160
rect 14160 -28170 14360 -28160
rect 14820 -28170 15020 -28160
rect 15700 -28170 15900 -28160
rect 16360 -28170 16560 -28160
rect 17020 -28170 17220 -28160
rect 17900 -28170 18100 -28160
rect 18560 -28170 18760 -28160
rect 19220 -28170 19420 -28160
rect 20900 -28170 20910 -28160
rect 21090 -28100 21100 -28090
rect 21090 -28160 22140 -28100
rect 21090 -28170 21100 -28160
rect 1220 -28180 1420 -28170
rect 20900 -28180 21100 -28170
rect 420 -28230 620 -28220
rect 420 -28310 430 -28230
rect 610 -28310 620 -28230
rect 1620 -28230 1820 -28220
rect 1620 -28240 1630 -28230
rect 1600 -28300 1630 -28240
rect 420 -28320 620 -28310
rect 1620 -28310 1630 -28300
rect 1810 -28240 1820 -28230
rect 20100 -28230 20300 -28220
rect 20100 -28240 20110 -28230
rect 1810 -28270 20110 -28240
rect 1810 -28300 4710 -28270
rect 1810 -28310 1820 -28300
rect 1620 -28320 1820 -28310
rect 4700 -28330 4710 -28300
rect 6210 -28300 6910 -28270
rect 6210 -28330 6220 -28300
rect 4700 -28340 6220 -28330
rect 6900 -28330 6910 -28300
rect 8410 -28300 9110 -28270
rect 8410 -28330 8420 -28300
rect 6900 -28340 8420 -28330
rect 9100 -28330 9110 -28300
rect 10610 -28300 11310 -28270
rect 10610 -28330 10620 -28300
rect 9100 -28340 10620 -28330
rect 11300 -28330 11310 -28300
rect 12810 -28300 13510 -28270
rect 12810 -28330 12820 -28300
rect 11300 -28340 12820 -28330
rect 13500 -28330 13510 -28300
rect 15010 -28300 15710 -28270
rect 15010 -28330 15020 -28300
rect 13500 -28340 15020 -28330
rect 15700 -28330 15710 -28300
rect 17210 -28300 20110 -28270
rect 17210 -28330 17220 -28300
rect 20100 -28310 20110 -28300
rect 20290 -28240 20300 -28230
rect 21300 -28230 21500 -28220
rect 20290 -28300 20320 -28240
rect 20290 -28310 20300 -28300
rect 20100 -28320 20300 -28310
rect 21300 -28310 21310 -28230
rect 21490 -28310 21500 -28230
rect 31810 -28290 31820 -28050
rect 33160 -28290 33170 -28050
rect 37720 -28180 37740 -28040
rect 37880 -28060 37900 -28040
rect 37880 -28160 38080 -28060
rect 37880 -28180 37900 -28160
rect 37720 -28200 37900 -28180
rect 31810 -28300 33170 -28290
rect 21300 -28320 21500 -28310
rect 15700 -28340 17220 -28330
rect 31790 -28710 32060 -28700
rect 29670 -28720 31800 -28710
rect 820 -28750 1020 -28740
rect 20500 -28750 20700 -28740
rect 820 -28760 830 -28750
rect -260 -28820 830 -28760
rect 820 -28830 830 -28820
rect 1010 -28760 1020 -28750
rect 2500 -28760 2700 -28750
rect 3160 -28760 3360 -28750
rect 3820 -28760 4020 -28750
rect 4700 -28760 4900 -28750
rect 5360 -28760 5560 -28750
rect 6020 -28760 6220 -28750
rect 6900 -28760 7100 -28750
rect 7560 -28760 7760 -28750
rect 8220 -28760 8420 -28750
rect 9100 -28760 9300 -28750
rect 9760 -28760 9960 -28750
rect 10420 -28760 10620 -28750
rect 11300 -28760 11500 -28750
rect 11960 -28760 12160 -28750
rect 12620 -28760 12820 -28750
rect 13500 -28760 13700 -28750
rect 14160 -28760 14360 -28750
rect 14820 -28760 15020 -28750
rect 15700 -28760 15900 -28750
rect 16360 -28760 16560 -28750
rect 17020 -28760 17220 -28750
rect 17900 -28760 18100 -28750
rect 18560 -28760 18760 -28750
rect 19220 -28760 19420 -28750
rect 20500 -28760 20510 -28750
rect 1010 -28820 2510 -28760
rect 2690 -28820 3170 -28760
rect 3350 -28820 3830 -28760
rect 4010 -28820 4710 -28760
rect 4890 -28820 5370 -28760
rect 5550 -28820 6030 -28760
rect 6210 -28820 15710 -28760
rect 15890 -28820 16370 -28760
rect 16550 -28820 17030 -28760
rect 17210 -28820 17910 -28760
rect 18090 -28820 18570 -28760
rect 18750 -28820 19230 -28760
rect 19410 -28820 20510 -28760
rect 1010 -28830 1020 -28820
rect 2500 -28830 2700 -28820
rect 3160 -28830 3360 -28820
rect 3820 -28830 4020 -28820
rect 4700 -28830 4900 -28820
rect 5360 -28830 5560 -28820
rect 6020 -28830 6220 -28820
rect 6900 -28830 7100 -28820
rect 7560 -28830 7760 -28820
rect 8220 -28830 8420 -28820
rect 9100 -28830 9300 -28820
rect 9760 -28830 9960 -28820
rect 10420 -28830 10620 -28820
rect 11300 -28830 11500 -28820
rect 11960 -28830 12160 -28820
rect 12620 -28830 12820 -28820
rect 13500 -28830 13700 -28820
rect 14160 -28830 14360 -28820
rect 14820 -28830 15020 -28820
rect 15700 -28830 15900 -28820
rect 16360 -28830 16560 -28820
rect 17020 -28830 17220 -28820
rect 17900 -28830 18100 -28820
rect 18560 -28830 18760 -28820
rect 19220 -28830 19420 -28820
rect 20500 -28830 20510 -28820
rect 20690 -28760 20700 -28750
rect 20690 -28820 22140 -28760
rect 20690 -28830 20700 -28820
rect 820 -28840 1020 -28830
rect 20500 -28840 20700 -28830
rect 1220 -28890 1420 -28880
rect 20900 -28890 21100 -28880
rect 1220 -28900 1230 -28890
rect -260 -28960 1230 -28900
rect 1220 -28970 1230 -28960
rect 1410 -28900 1420 -28890
rect 2500 -28900 2700 -28890
rect 3160 -28900 3360 -28890
rect 3820 -28900 4020 -28890
rect 4700 -28900 4900 -28890
rect 5360 -28900 5560 -28890
rect 6020 -28900 6220 -28890
rect 6900 -28900 7100 -28890
rect 7560 -28900 7760 -28890
rect 8220 -28900 8420 -28890
rect 9100 -28900 9300 -28890
rect 9760 -28900 9960 -28890
rect 10420 -28900 10620 -28890
rect 11300 -28900 11500 -28890
rect 11960 -28900 12160 -28890
rect 12620 -28900 12820 -28890
rect 13500 -28900 13700 -28890
rect 14160 -28900 14360 -28890
rect 14820 -28900 15020 -28890
rect 15700 -28900 15900 -28890
rect 16360 -28900 16560 -28890
rect 17020 -28900 17220 -28890
rect 17900 -28900 18100 -28890
rect 18560 -28900 18760 -28890
rect 19220 -28900 19420 -28890
rect 20900 -28900 20910 -28890
rect 1410 -28960 6910 -28900
rect 7090 -28960 7570 -28900
rect 7750 -28960 8230 -28900
rect 8410 -28960 9110 -28900
rect 9290 -28960 9770 -28900
rect 9950 -28960 10430 -28900
rect 10610 -28960 11310 -28900
rect 11490 -28960 11970 -28900
rect 12150 -28960 12630 -28900
rect 12810 -28960 13510 -28900
rect 13690 -28960 14170 -28900
rect 14350 -28960 14830 -28900
rect 15010 -28960 20910 -28900
rect 1410 -28970 1420 -28960
rect 2500 -28970 2700 -28960
rect 3160 -28970 3360 -28960
rect 3820 -28970 4020 -28960
rect 4700 -28970 4900 -28960
rect 5360 -28970 5560 -28960
rect 6020 -28970 6220 -28960
rect 6900 -28970 7100 -28960
rect 7560 -28970 7760 -28960
rect 8220 -28970 8420 -28960
rect 9100 -28970 9300 -28960
rect 9760 -28970 9960 -28960
rect 10420 -28970 10620 -28960
rect 11300 -28970 11500 -28960
rect 11960 -28970 12160 -28960
rect 12620 -28970 12820 -28960
rect 13500 -28970 13700 -28960
rect 14160 -28970 14360 -28960
rect 14820 -28970 15020 -28960
rect 15700 -28970 15900 -28960
rect 16360 -28970 16560 -28960
rect 17020 -28970 17220 -28960
rect 17900 -28970 18100 -28960
rect 18560 -28970 18760 -28960
rect 19220 -28970 19420 -28960
rect 20900 -28970 20910 -28960
rect 21090 -28900 21100 -28890
rect 21090 -28960 22140 -28900
rect 29670 -28940 29680 -28720
rect 29740 -28780 31800 -28720
rect 32050 -28780 32060 -28710
rect 29740 -28940 29750 -28780
rect 31790 -28790 32060 -28780
rect 32190 -28860 32460 -28850
rect 29670 -28950 29750 -28940
rect 29820 -28870 32200 -28860
rect 21090 -28970 21100 -28960
rect 1220 -28980 1420 -28970
rect 20900 -28980 21100 -28970
rect 420 -29030 620 -29020
rect 420 -29110 430 -29030
rect 610 -29110 620 -29030
rect 1620 -29030 1820 -29020
rect 1620 -29040 1630 -29030
rect 1600 -29100 1630 -29040
rect 420 -29120 620 -29110
rect 1620 -29110 1630 -29100
rect 1810 -29040 1820 -29030
rect 20100 -29030 20300 -29020
rect 20100 -29040 20110 -29030
rect 1810 -29070 20110 -29040
rect 1810 -29100 4710 -29070
rect 1810 -29110 1820 -29100
rect 1620 -29120 1820 -29110
rect 4700 -29130 4710 -29100
rect 6210 -29100 6910 -29070
rect 6210 -29130 6220 -29100
rect 4700 -29140 6220 -29130
rect 6900 -29130 6910 -29100
rect 8410 -29100 9110 -29070
rect 8410 -29130 8420 -29100
rect 6900 -29140 8420 -29130
rect 9100 -29130 9110 -29100
rect 10610 -29100 11310 -29070
rect 10610 -29130 10620 -29100
rect 9100 -29140 10620 -29130
rect 11300 -29130 11310 -29100
rect 12810 -29100 13510 -29070
rect 12810 -29130 12820 -29100
rect 11300 -29140 12820 -29130
rect 13500 -29130 13510 -29100
rect 15010 -29100 15710 -29070
rect 15010 -29130 15020 -29100
rect 13500 -29140 15020 -29130
rect 15700 -29130 15710 -29100
rect 17210 -29100 20110 -29070
rect 17210 -29130 17220 -29100
rect 20100 -29110 20110 -29100
rect 20290 -29040 20300 -29030
rect 21300 -29030 21500 -29020
rect 20290 -29100 20320 -29040
rect 20290 -29110 20300 -29100
rect 20100 -29120 20300 -29110
rect 21300 -29110 21310 -29030
rect 21490 -29110 21500 -29030
rect 29820 -29090 29830 -28870
rect 29890 -28930 32200 -28870
rect 32450 -28930 32460 -28860
rect 29890 -29090 29900 -28930
rect 32190 -28940 32460 -28930
rect 33990 -29010 34260 -29000
rect 29820 -29100 29900 -29090
rect 29970 -29020 34000 -29010
rect 21300 -29120 21500 -29110
rect 15700 -29140 17220 -29130
rect 29970 -29240 29980 -29020
rect 30040 -29080 34000 -29020
rect 34250 -29080 34260 -29010
rect 30040 -29240 30050 -29080
rect 33990 -29090 34260 -29080
rect 34400 -29150 34670 -29140
rect 34400 -29160 34410 -29150
rect 29970 -29250 30050 -29240
rect 30120 -29170 34410 -29160
rect 30120 -29390 30130 -29170
rect 30190 -29220 34410 -29170
rect 34660 -29220 34670 -29150
rect 30190 -29230 34670 -29220
rect 30190 -29390 30200 -29230
rect 36190 -29310 36460 -29300
rect 30120 -29400 30200 -29390
rect 30270 -29320 36200 -29310
rect 30270 -29540 30280 -29320
rect 30340 -29380 36200 -29320
rect 36450 -29380 36460 -29310
rect 30340 -29540 30350 -29380
rect 36190 -29390 36460 -29380
rect 36590 -29460 36860 -29450
rect 820 -29550 1020 -29540
rect 20500 -29550 20700 -29540
rect 30270 -29550 30350 -29540
rect 30420 -29470 36600 -29460
rect 820 -29560 830 -29550
rect -260 -29620 830 -29560
rect 820 -29630 830 -29620
rect 1010 -29560 1020 -29550
rect 2500 -29560 2700 -29550
rect 3160 -29560 3360 -29550
rect 3820 -29560 4020 -29550
rect 4700 -29560 4900 -29550
rect 5360 -29560 5560 -29550
rect 6020 -29560 6220 -29550
rect 6900 -29560 7100 -29550
rect 7560 -29560 7760 -29550
rect 8220 -29560 8420 -29550
rect 9100 -29560 9300 -29550
rect 9760 -29560 9960 -29550
rect 10420 -29560 10620 -29550
rect 11300 -29560 11500 -29550
rect 11960 -29560 12160 -29550
rect 12620 -29560 12820 -29550
rect 13500 -29560 13700 -29550
rect 14160 -29560 14360 -29550
rect 14820 -29560 15020 -29550
rect 15700 -29560 15900 -29550
rect 16360 -29560 16560 -29550
rect 17020 -29560 17220 -29550
rect 17900 -29560 18100 -29550
rect 18560 -29560 18760 -29550
rect 19220 -29560 19420 -29550
rect 20500 -29560 20510 -29550
rect 1010 -29620 6910 -29560
rect 7090 -29620 7570 -29560
rect 7750 -29620 8230 -29560
rect 8410 -29620 9110 -29560
rect 9290 -29620 9770 -29560
rect 9950 -29620 10430 -29560
rect 10610 -29620 11310 -29560
rect 11490 -29620 11970 -29560
rect 12150 -29620 12630 -29560
rect 12810 -29620 13510 -29560
rect 13690 -29620 14170 -29560
rect 14350 -29620 14830 -29560
rect 15010 -29620 20510 -29560
rect 1010 -29630 1020 -29620
rect 2500 -29630 2700 -29620
rect 3160 -29630 3360 -29620
rect 3820 -29630 4020 -29620
rect 4700 -29630 4900 -29620
rect 5360 -29630 5560 -29620
rect 6020 -29630 6220 -29620
rect 6900 -29630 7100 -29620
rect 7560 -29630 7760 -29620
rect 8220 -29630 8420 -29620
rect 9100 -29630 9300 -29620
rect 9760 -29630 9960 -29620
rect 10420 -29630 10620 -29620
rect 11300 -29630 11500 -29620
rect 11960 -29630 12160 -29620
rect 12620 -29630 12820 -29620
rect 13500 -29630 13700 -29620
rect 14160 -29630 14360 -29620
rect 14820 -29630 15020 -29620
rect 15700 -29630 15900 -29620
rect 16360 -29630 16560 -29620
rect 17020 -29630 17220 -29620
rect 17900 -29630 18100 -29620
rect 18560 -29630 18760 -29620
rect 19220 -29630 19420 -29620
rect 20500 -29630 20510 -29620
rect 20690 -29560 20700 -29550
rect 20690 -29620 22140 -29560
rect 20690 -29630 20700 -29620
rect 820 -29640 1020 -29630
rect 20500 -29640 20700 -29630
rect 1220 -29690 1420 -29680
rect 20900 -29690 21100 -29680
rect 1220 -29700 1230 -29690
rect -260 -29760 1230 -29700
rect 1220 -29770 1230 -29760
rect 1410 -29700 1420 -29690
rect 2500 -29700 2700 -29690
rect 3160 -29700 3360 -29690
rect 3820 -29700 4020 -29690
rect 4700 -29700 4900 -29690
rect 5360 -29700 5560 -29690
rect 6020 -29700 6220 -29690
rect 6900 -29700 7100 -29690
rect 7560 -29700 7760 -29690
rect 8220 -29700 8420 -29690
rect 9100 -29700 9300 -29690
rect 9760 -29700 9960 -29690
rect 10420 -29700 10620 -29690
rect 11300 -29700 11500 -29690
rect 11960 -29700 12160 -29690
rect 12620 -29700 12820 -29690
rect 13500 -29700 13700 -29690
rect 14160 -29700 14360 -29690
rect 14820 -29700 15020 -29690
rect 15700 -29700 15900 -29690
rect 16360 -29700 16560 -29690
rect 17020 -29700 17220 -29690
rect 17900 -29700 18100 -29690
rect 18560 -29700 18760 -29690
rect 19220 -29700 19420 -29690
rect 20900 -29700 20910 -29690
rect 1410 -29760 2510 -29700
rect 2690 -29760 3170 -29700
rect 3350 -29760 3830 -29700
rect 4010 -29760 4710 -29700
rect 4890 -29760 5370 -29700
rect 5550 -29760 6030 -29700
rect 6210 -29760 15710 -29700
rect 15890 -29760 16370 -29700
rect 16550 -29760 17030 -29700
rect 17210 -29760 17910 -29700
rect 18090 -29760 18570 -29700
rect 18750 -29760 19230 -29700
rect 19410 -29760 20910 -29700
rect 1410 -29770 1420 -29760
rect 2500 -29770 2700 -29760
rect 3160 -29770 3360 -29760
rect 3820 -29770 4020 -29760
rect 4700 -29770 4900 -29760
rect 5360 -29770 5560 -29760
rect 6020 -29770 6220 -29760
rect 6900 -29770 7100 -29760
rect 7560 -29770 7760 -29760
rect 8220 -29770 8420 -29760
rect 9100 -29770 9300 -29760
rect 9760 -29770 9960 -29760
rect 10420 -29770 10620 -29760
rect 11300 -29770 11500 -29760
rect 11960 -29770 12160 -29760
rect 12620 -29770 12820 -29760
rect 13500 -29770 13700 -29760
rect 14160 -29770 14360 -29760
rect 14820 -29770 15020 -29760
rect 15700 -29770 15900 -29760
rect 16360 -29770 16560 -29760
rect 17020 -29770 17220 -29760
rect 17900 -29770 18100 -29760
rect 18560 -29770 18760 -29760
rect 19220 -29770 19420 -29760
rect 20900 -29770 20910 -29760
rect 21090 -29700 21100 -29690
rect 30420 -29690 30430 -29470
rect 30490 -29530 36600 -29470
rect 36850 -29530 36860 -29460
rect 30490 -29690 30500 -29530
rect 36590 -29540 36860 -29530
rect 30420 -29700 30500 -29690
rect 21090 -29760 22140 -29700
rect 21090 -29770 21100 -29760
rect 1220 -29780 1420 -29770
rect 20900 -29780 21100 -29770
rect 1620 -29830 1820 -29820
rect 1620 -29840 1630 -29830
rect 1600 -29900 1630 -29840
rect 1620 -29910 1630 -29900
rect 1810 -29840 1820 -29830
rect 20100 -29830 20300 -29820
rect 20100 -29840 20110 -29830
rect 1810 -29870 20110 -29840
rect 1810 -29900 2510 -29870
rect 1810 -29910 1820 -29900
rect 1620 -29920 1820 -29910
rect 2500 -29930 2510 -29900
rect 4010 -29900 4710 -29870
rect 4010 -29930 4020 -29900
rect 2500 -29940 4020 -29930
rect 4700 -29930 4710 -29900
rect 6210 -29900 6910 -29870
rect 6210 -29930 6220 -29900
rect 4700 -29940 6220 -29930
rect 6900 -29930 6910 -29900
rect 8410 -29900 9110 -29870
rect 8410 -29930 8420 -29900
rect 6900 -29940 8420 -29930
rect 9100 -29930 9110 -29900
rect 10610 -29900 11310 -29870
rect 10610 -29930 10620 -29900
rect 9100 -29940 10620 -29930
rect 11300 -29930 11310 -29900
rect 12810 -29900 13510 -29870
rect 12810 -29930 12820 -29900
rect 11300 -29940 12820 -29930
rect 13500 -29930 13510 -29900
rect 15010 -29900 15710 -29870
rect 15010 -29930 15020 -29900
rect 13500 -29940 15020 -29930
rect 15700 -29930 15710 -29900
rect 17210 -29900 17910 -29870
rect 17210 -29930 17220 -29900
rect 15700 -29940 17220 -29930
rect 17900 -29930 17910 -29900
rect 19410 -29900 20110 -29870
rect 19410 -29930 19420 -29900
rect 20100 -29910 20110 -29900
rect 20290 -29840 20300 -29830
rect 20290 -29900 20320 -29840
rect 20290 -29910 20300 -29900
rect 20100 -29920 20300 -29910
rect 37240 -29920 37700 -29910
rect 17900 -29940 19420 -29930
rect 37240 -30110 37250 -29920
rect 37690 -30110 37700 -29920
rect 37240 -30120 37700 -30110
rect 820 -30350 1020 -30340
rect 20500 -30350 20700 -30340
rect 820 -30360 830 -30350
rect -260 -30420 830 -30360
rect 820 -30430 830 -30420
rect 1010 -30360 1020 -30350
rect 2500 -30360 2700 -30350
rect 3160 -30360 3360 -30350
rect 3820 -30360 4020 -30350
rect 4700 -30360 4900 -30350
rect 5360 -30360 5560 -30350
rect 6020 -30360 6220 -30350
rect 6900 -30360 7100 -30350
rect 7560 -30360 7760 -30350
rect 8220 -30360 8420 -30350
rect 9100 -30360 9300 -30350
rect 9760 -30360 9960 -30350
rect 10420 -30360 10620 -30350
rect 11300 -30360 11500 -30350
rect 11960 -30360 12160 -30350
rect 12620 -30360 12820 -30350
rect 13500 -30360 13700 -30350
rect 14160 -30360 14360 -30350
rect 14820 -30360 15020 -30350
rect 15700 -30360 15900 -30350
rect 16360 -30360 16560 -30350
rect 17020 -30360 17220 -30350
rect 17900 -30360 18100 -30350
rect 18560 -30360 18760 -30350
rect 19220 -30360 19420 -30350
rect 20500 -30360 20510 -30350
rect 1010 -30420 2510 -30360
rect 2690 -30420 3170 -30360
rect 3350 -30420 3830 -30360
rect 4010 -30420 4710 -30360
rect 4890 -30420 5370 -30360
rect 5550 -30420 6030 -30360
rect 6210 -30420 15710 -30360
rect 15890 -30420 16370 -30360
rect 16550 -30420 17030 -30360
rect 17210 -30420 17910 -30360
rect 18090 -30420 18570 -30360
rect 18750 -30420 19230 -30360
rect 19410 -30420 20510 -30360
rect 1010 -30430 1020 -30420
rect 2500 -30430 2700 -30420
rect 3160 -30430 3360 -30420
rect 3820 -30430 4020 -30420
rect 4700 -30430 4900 -30420
rect 5360 -30430 5560 -30420
rect 6020 -30430 6220 -30420
rect 6900 -30430 7100 -30420
rect 7560 -30430 7760 -30420
rect 8220 -30430 8420 -30420
rect 9100 -30430 9300 -30420
rect 9760 -30430 9960 -30420
rect 10420 -30430 10620 -30420
rect 11300 -30430 11500 -30420
rect 11960 -30430 12160 -30420
rect 12620 -30430 12820 -30420
rect 13500 -30430 13700 -30420
rect 14160 -30430 14360 -30420
rect 14820 -30430 15020 -30420
rect 15700 -30430 15900 -30420
rect 16360 -30430 16560 -30420
rect 17020 -30430 17220 -30420
rect 17900 -30430 18100 -30420
rect 18560 -30430 18760 -30420
rect 19220 -30430 19420 -30420
rect 20500 -30430 20510 -30420
rect 20690 -30360 20700 -30350
rect 20690 -30420 22140 -30360
rect 20690 -30430 20700 -30420
rect 820 -30440 1020 -30430
rect 20500 -30440 20700 -30430
rect 1220 -30490 1420 -30480
rect 20900 -30490 21100 -30480
rect 1220 -30500 1230 -30490
rect -260 -30560 1230 -30500
rect 1220 -30570 1230 -30560
rect 1410 -30500 1420 -30490
rect 2500 -30500 2700 -30490
rect 3160 -30500 3360 -30490
rect 3820 -30500 4020 -30490
rect 4700 -30500 4900 -30490
rect 5360 -30500 5560 -30490
rect 6020 -30500 6220 -30490
rect 6900 -30500 7100 -30490
rect 7560 -30500 7760 -30490
rect 8220 -30500 8420 -30490
rect 9100 -30500 9300 -30490
rect 9760 -30500 9960 -30490
rect 10420 -30500 10620 -30490
rect 11300 -30500 11500 -30490
rect 11960 -30500 12160 -30490
rect 12620 -30500 12820 -30490
rect 13500 -30500 13700 -30490
rect 14160 -30500 14360 -30490
rect 14820 -30500 15020 -30490
rect 15700 -30500 15900 -30490
rect 16360 -30500 16560 -30490
rect 17020 -30500 17220 -30490
rect 17900 -30500 18100 -30490
rect 18560 -30500 18760 -30490
rect 19220 -30500 19420 -30490
rect 20900 -30500 20910 -30490
rect 1410 -30560 6910 -30500
rect 7090 -30560 7570 -30500
rect 7750 -30560 8230 -30500
rect 8410 -30560 9110 -30500
rect 9290 -30560 9770 -30500
rect 9950 -30560 10430 -30500
rect 10610 -30560 11310 -30500
rect 11490 -30560 11970 -30500
rect 12150 -30560 12630 -30500
rect 12810 -30560 13510 -30500
rect 13690 -30560 14170 -30500
rect 14350 -30560 14830 -30500
rect 15010 -30560 20910 -30500
rect 1410 -30570 1420 -30560
rect 2500 -30570 2700 -30560
rect 3160 -30570 3360 -30560
rect 3820 -30570 4020 -30560
rect 4700 -30570 4900 -30560
rect 5360 -30570 5560 -30560
rect 6020 -30570 6220 -30560
rect 6900 -30570 7100 -30560
rect 7560 -30570 7760 -30560
rect 8220 -30570 8420 -30560
rect 9100 -30570 9300 -30560
rect 9760 -30570 9960 -30560
rect 10420 -30570 10620 -30560
rect 11300 -30570 11500 -30560
rect 11960 -30570 12160 -30560
rect 12620 -30570 12820 -30560
rect 13500 -30570 13700 -30560
rect 14160 -30570 14360 -30560
rect 14820 -30570 15020 -30560
rect 15700 -30570 15900 -30560
rect 16360 -30570 16560 -30560
rect 17020 -30570 17220 -30560
rect 17900 -30570 18100 -30560
rect 18560 -30570 18760 -30560
rect 19220 -30570 19420 -30560
rect 20900 -30570 20910 -30560
rect 21090 -30500 21100 -30490
rect 21090 -30560 22140 -30500
rect 21090 -30570 21100 -30560
rect 1220 -30580 1420 -30570
rect 20900 -30580 21100 -30570
rect 1620 -30630 1820 -30620
rect 1620 -30640 1630 -30630
rect 1600 -30700 1630 -30640
rect 1620 -30710 1630 -30700
rect 1810 -30640 1820 -30630
rect 20100 -30630 20300 -30620
rect 20100 -30640 20110 -30630
rect 1810 -30670 20110 -30640
rect 1810 -30700 2510 -30670
rect 1810 -30710 1820 -30700
rect 1620 -30720 1820 -30710
rect 2500 -30730 2510 -30700
rect 4010 -30700 4710 -30670
rect 4010 -30730 4020 -30700
rect 2500 -30740 4020 -30730
rect 4700 -30730 4710 -30700
rect 6210 -30700 6910 -30670
rect 6210 -30730 6220 -30700
rect 4700 -30740 6220 -30730
rect 6900 -30730 6910 -30700
rect 8410 -30700 9110 -30670
rect 8410 -30730 8420 -30700
rect 6900 -30740 8420 -30730
rect 9100 -30730 9110 -30700
rect 10610 -30700 11310 -30670
rect 10610 -30730 10620 -30700
rect 9100 -30740 10620 -30730
rect 11300 -30730 11310 -30700
rect 12810 -30700 13510 -30670
rect 12810 -30730 12820 -30700
rect 11300 -30740 12820 -30730
rect 13500 -30730 13510 -30700
rect 15010 -30700 15710 -30670
rect 15010 -30730 15020 -30700
rect 13500 -30740 15020 -30730
rect 15700 -30730 15710 -30700
rect 17210 -30700 17910 -30670
rect 17210 -30730 17220 -30700
rect 15700 -30740 17220 -30730
rect 17900 -30730 17910 -30700
rect 19410 -30700 20110 -30670
rect 19410 -30730 19420 -30700
rect 20100 -30710 20110 -30700
rect 20290 -30640 20300 -30630
rect 20290 -30700 20320 -30640
rect 20290 -30710 20300 -30700
rect 20100 -30720 20300 -30710
rect 17900 -30740 19420 -30730
rect 28930 -30810 29170 -30800
rect 32950 -30810 33220 -30800
rect 28930 -30880 28940 -30810
rect 29160 -30880 32960 -30810
rect 33210 -30880 33220 -30810
rect 28930 -30890 29170 -30880
rect 32950 -30890 33220 -30880
rect 29060 -30960 29300 -30950
rect 33320 -30960 33590 -30950
rect 29060 -31030 29070 -30960
rect 29290 -31030 33330 -30960
rect 33580 -31030 33590 -30960
rect 29060 -31040 29300 -31030
rect 33320 -31040 33590 -31030
rect 29210 -31110 29450 -31100
rect 35550 -31110 35820 -31100
rect 820 -31150 1020 -31140
rect 20500 -31150 20700 -31140
rect 820 -31160 830 -31150
rect -260 -31220 830 -31160
rect 820 -31230 830 -31220
rect 1010 -31160 1020 -31150
rect 2500 -31160 2700 -31150
rect 3160 -31160 3360 -31150
rect 3820 -31160 4020 -31150
rect 4700 -31160 4900 -31150
rect 5360 -31160 5560 -31150
rect 6020 -31160 6220 -31150
rect 6900 -31160 7100 -31150
rect 7560 -31160 7760 -31150
rect 8220 -31160 8420 -31150
rect 9100 -31160 9300 -31150
rect 9760 -31160 9960 -31150
rect 10420 -31160 10620 -31150
rect 11300 -31160 11500 -31150
rect 11960 -31160 12160 -31150
rect 12620 -31160 12820 -31150
rect 13500 -31160 13700 -31150
rect 14160 -31160 14360 -31150
rect 14820 -31160 15020 -31150
rect 15700 -31160 15900 -31150
rect 16360 -31160 16560 -31150
rect 17020 -31160 17220 -31150
rect 17900 -31160 18100 -31150
rect 18560 -31160 18760 -31150
rect 19220 -31160 19420 -31150
rect 20500 -31160 20510 -31150
rect 1010 -31220 6910 -31160
rect 7090 -31220 7570 -31160
rect 7750 -31220 8230 -31160
rect 8410 -31220 9110 -31160
rect 9290 -31220 9770 -31160
rect 9950 -31220 10430 -31160
rect 10610 -31220 11310 -31160
rect 11490 -31220 11970 -31160
rect 12150 -31220 12630 -31160
rect 12810 -31220 13510 -31160
rect 13690 -31220 14170 -31160
rect 14350 -31220 14830 -31160
rect 15010 -31220 20510 -31160
rect 1010 -31230 1020 -31220
rect 2500 -31230 2700 -31220
rect 3160 -31230 3360 -31220
rect 3820 -31230 4020 -31220
rect 4700 -31230 4900 -31220
rect 5360 -31230 5560 -31220
rect 6020 -31230 6220 -31220
rect 6900 -31230 7100 -31220
rect 7560 -31230 7760 -31220
rect 8220 -31230 8420 -31220
rect 9100 -31230 9300 -31220
rect 9760 -31230 9960 -31220
rect 10420 -31230 10620 -31220
rect 11300 -31230 11500 -31220
rect 11960 -31230 12160 -31220
rect 12620 -31230 12820 -31220
rect 13500 -31230 13700 -31220
rect 14160 -31230 14360 -31220
rect 14820 -31230 15020 -31220
rect 15700 -31230 15900 -31220
rect 16360 -31230 16560 -31220
rect 17020 -31230 17220 -31220
rect 17900 -31230 18100 -31220
rect 18560 -31230 18760 -31220
rect 19220 -31230 19420 -31220
rect 20500 -31230 20510 -31220
rect 20690 -31160 20700 -31150
rect 20690 -31220 22140 -31160
rect 29210 -31180 29220 -31110
rect 29440 -31180 35560 -31110
rect 35810 -31180 35820 -31110
rect 29210 -31190 29450 -31180
rect 35550 -31190 35820 -31180
rect 20690 -31230 20700 -31220
rect 820 -31240 1020 -31230
rect 20500 -31240 20700 -31230
rect 29360 -31260 29600 -31250
rect 37700 -31260 37970 -31250
rect 1220 -31290 1420 -31280
rect 20900 -31290 21100 -31280
rect 1220 -31300 1230 -31290
rect -260 -31360 1230 -31300
rect 1220 -31370 1230 -31360
rect 1410 -31300 1420 -31290
rect 2500 -31300 2700 -31290
rect 3160 -31300 3360 -31290
rect 3820 -31300 4020 -31290
rect 4700 -31300 4900 -31290
rect 5360 -31300 5560 -31290
rect 6020 -31300 6220 -31290
rect 6900 -31300 7100 -31290
rect 7560 -31300 7760 -31290
rect 8220 -31300 8420 -31290
rect 9100 -31300 9300 -31290
rect 9760 -31300 9960 -31290
rect 10420 -31300 10620 -31290
rect 11300 -31300 11500 -31290
rect 11960 -31300 12160 -31290
rect 12620 -31300 12820 -31290
rect 13500 -31300 13700 -31290
rect 14160 -31300 14360 -31290
rect 14820 -31300 15020 -31290
rect 15700 -31300 15900 -31290
rect 16360 -31300 16560 -31290
rect 17020 -31300 17220 -31290
rect 17900 -31300 18100 -31290
rect 18560 -31300 18760 -31290
rect 19220 -31300 19420 -31290
rect 20900 -31300 20910 -31290
rect 1410 -31360 2510 -31300
rect 2690 -31360 3170 -31300
rect 3350 -31360 3830 -31300
rect 4010 -31360 4710 -31300
rect 4890 -31360 5370 -31300
rect 5550 -31360 6030 -31300
rect 6210 -31360 15710 -31300
rect 15890 -31360 16370 -31300
rect 16550 -31360 17030 -31300
rect 17210 -31360 17910 -31300
rect 18090 -31360 18570 -31300
rect 18750 -31360 19230 -31300
rect 19410 -31360 20910 -31300
rect 1410 -31370 1420 -31360
rect 2500 -31370 2700 -31360
rect 3160 -31370 3360 -31360
rect 3820 -31370 4020 -31360
rect 4700 -31370 4900 -31360
rect 5360 -31370 5560 -31360
rect 6020 -31370 6220 -31360
rect 6900 -31370 7100 -31360
rect 7560 -31370 7760 -31360
rect 8220 -31370 8420 -31360
rect 9100 -31370 9300 -31360
rect 9760 -31370 9960 -31360
rect 10420 -31370 10620 -31360
rect 11300 -31370 11500 -31360
rect 11960 -31370 12160 -31360
rect 12620 -31370 12820 -31360
rect 13500 -31370 13700 -31360
rect 14160 -31370 14360 -31360
rect 14820 -31370 15020 -31360
rect 15700 -31370 15900 -31360
rect 16360 -31370 16560 -31360
rect 17020 -31370 17220 -31360
rect 17900 -31370 18100 -31360
rect 18560 -31370 18760 -31360
rect 19220 -31370 19420 -31360
rect 20900 -31370 20910 -31360
rect 21090 -31300 21100 -31290
rect 21090 -31360 22140 -31300
rect 29360 -31330 29370 -31260
rect 29590 -31330 37710 -31260
rect 37960 -31330 37970 -31260
rect 29360 -31340 29600 -31330
rect 37700 -31340 37970 -31330
rect 21090 -31370 21100 -31360
rect 1220 -31380 1420 -31370
rect 20900 -31380 21100 -31370
rect -360 -31450 570 -31440
rect -360 -31830 -350 -31450
rect -170 -31540 570 -31450
rect -170 -31830 -160 -31540
rect 460 -31720 570 -31540
rect 1980 -31710 2120 -31700
rect 1980 -31720 1990 -31710
rect -360 -31840 -160 -31830
rect 80 -31730 280 -31720
rect 80 -32110 90 -31730
rect 270 -32020 280 -31730
rect 460 -31820 1990 -31720
rect 1980 -31830 1990 -31820
rect 2110 -31720 2120 -31710
rect 4180 -31710 4320 -31700
rect 4180 -31720 4190 -31710
rect 2110 -31820 4190 -31720
rect 2110 -31830 2120 -31820
rect 1980 -31840 2120 -31830
rect 4180 -31830 4190 -31820
rect 4310 -31720 4320 -31710
rect 6380 -31710 6520 -31700
rect 6380 -31720 6390 -31710
rect 4310 -31820 6390 -31720
rect 4310 -31830 4320 -31820
rect 4180 -31840 4320 -31830
rect 6380 -31830 6390 -31820
rect 6510 -31720 6520 -31710
rect 8580 -31710 8720 -31700
rect 8580 -31720 8590 -31710
rect 6510 -31820 8590 -31720
rect 6510 -31830 6520 -31820
rect 6380 -31840 6520 -31830
rect 8580 -31830 8590 -31820
rect 8710 -31720 8720 -31710
rect 10780 -31710 10920 -31700
rect 10780 -31720 10790 -31710
rect 8710 -31820 10790 -31720
rect 8710 -31830 8720 -31820
rect 8580 -31840 8720 -31830
rect 10780 -31830 10790 -31820
rect 10910 -31720 10920 -31710
rect 12980 -31710 13120 -31700
rect 12980 -31720 12990 -31710
rect 10910 -31820 12990 -31720
rect 10910 -31830 10920 -31820
rect 10780 -31840 10920 -31830
rect 12980 -31830 12990 -31820
rect 13110 -31720 13120 -31710
rect 15180 -31710 15320 -31700
rect 15180 -31720 15190 -31710
rect 13110 -31820 15190 -31720
rect 13110 -31830 13120 -31820
rect 12980 -31840 13120 -31830
rect 15180 -31830 15190 -31820
rect 15310 -31720 15320 -31710
rect 17380 -31710 17520 -31700
rect 17380 -31720 17390 -31710
rect 15310 -31820 17390 -31720
rect 15310 -31830 15320 -31820
rect 15180 -31840 15320 -31830
rect 17380 -31830 17390 -31820
rect 17510 -31720 17520 -31710
rect 19580 -31710 19720 -31700
rect 19580 -31720 19590 -31710
rect 17510 -31820 19590 -31720
rect 17510 -31830 17520 -31820
rect 17380 -31840 17520 -31830
rect 19580 -31830 19590 -31820
rect 19710 -31720 19720 -31710
rect 19710 -31820 22240 -31720
rect 32530 -31730 33700 -31720
rect 19710 -31830 19720 -31820
rect 19580 -31840 19720 -31830
rect 32530 -31950 32540 -31730
rect 33690 -31950 33700 -31730
rect 32530 -31960 33700 -31950
rect 2200 -32010 2340 -32000
rect 2200 -32020 2210 -32010
rect 270 -32110 2210 -32020
rect 80 -32120 2210 -32110
rect 2200 -32130 2210 -32120
rect 2330 -32020 2340 -32010
rect 4400 -32010 4540 -32000
rect 4400 -32020 4410 -32010
rect 2330 -32120 4410 -32020
rect 2330 -32130 2340 -32120
rect 2200 -32140 2340 -32130
rect 4400 -32130 4410 -32120
rect 4530 -32020 4540 -32010
rect 6600 -32010 6740 -32000
rect 6600 -32020 6610 -32010
rect 4530 -32120 6610 -32020
rect 4530 -32130 4540 -32120
rect 4400 -32140 4540 -32130
rect 6600 -32130 6610 -32120
rect 6730 -32020 6740 -32010
rect 8800 -32010 8940 -32000
rect 8800 -32020 8810 -32010
rect 6730 -32120 8810 -32020
rect 6730 -32130 6740 -32120
rect 6600 -32140 6740 -32130
rect 8800 -32130 8810 -32120
rect 8930 -32020 8940 -32010
rect 11000 -32010 11140 -32000
rect 11000 -32020 11010 -32010
rect 8930 -32120 11010 -32020
rect 8930 -32130 8940 -32120
rect 8800 -32140 8940 -32130
rect 11000 -32130 11010 -32120
rect 11130 -32020 11140 -32010
rect 13200 -32010 13340 -32000
rect 13200 -32020 13210 -32010
rect 11130 -32120 13210 -32020
rect 11130 -32130 11140 -32120
rect 11000 -32140 11140 -32130
rect 13200 -32130 13210 -32120
rect 13330 -32020 13340 -32010
rect 15400 -32010 15540 -32000
rect 15400 -32020 15410 -32010
rect 13330 -32120 15410 -32020
rect 13330 -32130 13340 -32120
rect 13200 -32140 13340 -32130
rect 15400 -32130 15410 -32120
rect 15530 -32020 15540 -32010
rect 17600 -32010 17740 -32000
rect 17600 -32020 17610 -32010
rect 15530 -32120 17610 -32020
rect 15530 -32130 15540 -32120
rect 15400 -32140 15540 -32130
rect 17600 -32130 17610 -32120
rect 17730 -32020 17740 -32010
rect 19800 -32010 19940 -32000
rect 19800 -32020 19810 -32010
rect 17730 -32120 19810 -32020
rect 17730 -32130 17740 -32120
rect 17600 -32140 17740 -32130
rect 19800 -32130 19810 -32120
rect 19930 -32020 19940 -32010
rect 19930 -32120 22240 -32020
rect 19930 -32130 19940 -32120
rect 19800 -32140 19940 -32130
<< via3 >>
rect 36480 11510 36810 11980
rect 830 11170 1010 11250
rect 20510 11170 20690 11250
rect 1230 11030 1410 11110
rect 20910 11030 21090 11110
rect -80 10930 0 10940
rect -80 10870 -70 10930
rect -70 10870 -10 10930
rect -10 10870 0 10930
rect -80 10690 0 10870
rect 2120 10930 2200 10940
rect 2120 10870 2130 10930
rect 2130 10870 2190 10930
rect 2190 10870 2200 10930
rect 2120 10690 2200 10870
rect 4320 10930 4400 10940
rect 4320 10870 4330 10930
rect 4330 10870 4390 10930
rect 4390 10870 4400 10930
rect 4320 10690 4400 10870
rect 6520 10930 6600 10940
rect 6520 10870 6530 10930
rect 6530 10870 6590 10930
rect 6590 10870 6600 10930
rect 6520 10690 6600 10870
rect 8720 10930 8800 10940
rect 8720 10870 8730 10930
rect 8730 10870 8790 10930
rect 8790 10870 8800 10930
rect 8720 10690 8800 10870
rect 10920 10930 11000 10940
rect 10920 10870 10930 10930
rect 10930 10870 10990 10930
rect 10990 10870 11000 10930
rect 10920 10690 11000 10870
rect 13120 10930 13200 10940
rect 13120 10870 13130 10930
rect 13130 10870 13190 10930
rect 13190 10870 13200 10930
rect 13120 10690 13200 10870
rect 15320 10930 15400 10940
rect 15320 10870 15330 10930
rect 15330 10870 15390 10930
rect 15390 10870 15400 10930
rect 15320 10690 15400 10870
rect 17520 10930 17600 10940
rect 17520 10870 17530 10930
rect 17530 10870 17590 10930
rect 17590 10870 17600 10930
rect 17520 10690 17600 10870
rect 19720 10930 19800 10940
rect 19720 10870 19730 10930
rect 19730 10870 19790 10930
rect 19790 10870 19800 10930
rect 19720 10690 19800 10870
rect 21920 10930 22000 10940
rect 21920 10870 21930 10930
rect 21930 10870 21990 10930
rect 21990 10870 22000 10930
rect 21920 10690 22000 10870
rect 1630 10510 1810 10590
rect 20110 10510 20290 10590
rect 830 10370 1010 10450
rect 20510 10370 20690 10450
rect 1230 10230 1410 10310
rect 20910 10230 21090 10310
rect -80 10130 0 10140
rect -80 10070 -70 10130
rect -70 10070 -10 10130
rect -10 10070 0 10130
rect -80 9890 0 10070
rect 2120 10130 2200 10140
rect 2120 10070 2130 10130
rect 2130 10070 2190 10130
rect 2190 10070 2200 10130
rect 2120 9890 2200 10070
rect 4320 10130 4400 10140
rect 4320 10070 4330 10130
rect 4330 10070 4390 10130
rect 4390 10070 4400 10130
rect 4320 9890 4400 10070
rect 6520 10130 6600 10140
rect 6520 10070 6530 10130
rect 6530 10070 6590 10130
rect 6590 10070 6600 10130
rect 6520 9890 6600 10070
rect 8720 10130 8800 10140
rect 8720 10070 8730 10130
rect 8730 10070 8790 10130
rect 8790 10070 8800 10130
rect 8720 9890 8800 10070
rect 10920 10130 11000 10140
rect 10920 10070 10930 10130
rect 10930 10070 10990 10130
rect 10990 10070 11000 10130
rect 10920 9890 11000 10070
rect 13120 10130 13200 10140
rect 13120 10070 13130 10130
rect 13130 10070 13190 10130
rect 13190 10070 13200 10130
rect 13120 9890 13200 10070
rect 15320 10130 15400 10140
rect 15320 10070 15330 10130
rect 15330 10070 15390 10130
rect 15390 10070 15400 10130
rect 15320 9890 15400 10070
rect 17520 10130 17600 10140
rect 17520 10070 17530 10130
rect 17530 10070 17590 10130
rect 17590 10070 17600 10130
rect 17520 9890 17600 10070
rect 19720 10130 19800 10140
rect 19720 10070 19730 10130
rect 19730 10070 19790 10130
rect 19790 10070 19800 10130
rect 19720 9890 19800 10070
rect 21920 10130 22000 10140
rect 21920 10070 21930 10130
rect 21930 10070 21990 10130
rect 21990 10070 22000 10130
rect 21920 9890 22000 10070
rect 1630 9710 1810 9790
rect 20110 9710 20290 9790
rect 830 9570 1010 9650
rect 20510 9570 20690 9650
rect 1230 9430 1410 9510
rect 20910 9430 21090 9510
rect -80 9330 0 9340
rect -80 9270 -70 9330
rect -70 9270 -10 9330
rect -10 9270 0 9330
rect -80 9090 0 9270
rect 2120 9330 2200 9340
rect 2120 9270 2130 9330
rect 2130 9270 2190 9330
rect 2190 9270 2200 9330
rect 2120 9090 2200 9270
rect 4320 9330 4400 9340
rect 4320 9270 4330 9330
rect 4330 9270 4390 9330
rect 4390 9270 4400 9330
rect 4320 9090 4400 9270
rect 6520 9330 6600 9340
rect 6520 9270 6530 9330
rect 6530 9270 6590 9330
rect 6590 9270 6600 9330
rect 6520 9090 6600 9270
rect 8720 9330 8800 9340
rect 8720 9270 8730 9330
rect 8730 9270 8790 9330
rect 8790 9270 8800 9330
rect 8720 9090 8800 9270
rect 10920 9330 11000 9340
rect 10920 9270 10930 9330
rect 10930 9270 10990 9330
rect 10990 9270 11000 9330
rect 10920 9090 11000 9270
rect 13120 9330 13200 9340
rect 13120 9270 13130 9330
rect 13130 9270 13190 9330
rect 13190 9270 13200 9330
rect 13120 9090 13200 9270
rect 15320 9330 15400 9340
rect 15320 9270 15330 9330
rect 15330 9270 15390 9330
rect 15390 9270 15400 9330
rect 15320 9090 15400 9270
rect 17520 9330 17600 9340
rect 17520 9270 17530 9330
rect 17530 9270 17590 9330
rect 17590 9270 17600 9330
rect 17520 9090 17600 9270
rect 19720 9330 19800 9340
rect 19720 9270 19730 9330
rect 19730 9270 19790 9330
rect 19790 9270 19800 9330
rect 19720 9090 19800 9270
rect 21920 9330 22000 9340
rect 21920 9270 21930 9330
rect 21930 9270 21990 9330
rect 21990 9270 22000 9330
rect 21920 9090 22000 9270
rect 37910 9200 38090 9380
rect 430 8910 610 8990
rect 1630 8910 1810 8990
rect 20110 8910 20290 8990
rect 21310 8910 21490 8990
rect 830 8770 1010 8850
rect 20510 8770 20690 8850
rect 1230 8630 1410 8710
rect 20910 8630 21090 8710
rect -80 8530 0 8540
rect -80 8470 -70 8530
rect -70 8470 -10 8530
rect -10 8470 0 8530
rect -80 8290 0 8470
rect 2120 8530 2200 8540
rect 2120 8470 2130 8530
rect 2130 8470 2190 8530
rect 2190 8470 2200 8530
rect 2120 8290 2200 8470
rect 4320 8530 4400 8540
rect 4320 8470 4330 8530
rect 4330 8470 4390 8530
rect 4390 8470 4400 8530
rect 4320 8290 4400 8470
rect 6520 8530 6600 8540
rect 6520 8470 6530 8530
rect 6530 8470 6590 8530
rect 6590 8470 6600 8530
rect 6520 8290 6600 8470
rect 8720 8530 8800 8540
rect 8720 8470 8730 8530
rect 8730 8470 8790 8530
rect 8790 8470 8800 8530
rect 8720 8290 8800 8470
rect 10920 8530 11000 8540
rect 10920 8470 10930 8530
rect 10930 8470 10990 8530
rect 10990 8470 11000 8530
rect 10920 8290 11000 8470
rect 13120 8530 13200 8540
rect 13120 8470 13130 8530
rect 13130 8470 13190 8530
rect 13190 8470 13200 8530
rect 13120 8290 13200 8470
rect 15320 8530 15400 8540
rect 15320 8470 15330 8530
rect 15330 8470 15390 8530
rect 15390 8470 15400 8530
rect 15320 8290 15400 8470
rect 17520 8530 17600 8540
rect 17520 8470 17530 8530
rect 17530 8470 17590 8530
rect 17590 8470 17600 8530
rect 17520 8290 17600 8470
rect 19720 8530 19800 8540
rect 19720 8470 19730 8530
rect 19730 8470 19790 8530
rect 19790 8470 19800 8530
rect 19720 8290 19800 8470
rect 21920 8530 22000 8540
rect 21920 8470 21930 8530
rect 21930 8470 21990 8530
rect 21990 8470 22000 8530
rect 21920 8290 22000 8470
rect 430 8110 610 8190
rect 1630 8110 1810 8190
rect 20110 8110 20290 8190
rect 21310 8110 21490 8190
rect 830 7970 1010 8050
rect 20510 7970 20690 8050
rect 36790 8030 37010 8170
rect 1230 7830 1410 7910
rect 20910 7830 21090 7910
rect 37130 7830 37350 7970
rect -80 7730 0 7740
rect -80 7670 -70 7730
rect -70 7670 -10 7730
rect -10 7670 0 7730
rect -80 7490 0 7670
rect 2120 7730 2200 7740
rect 2120 7670 2130 7730
rect 2130 7670 2190 7730
rect 2190 7670 2200 7730
rect 2120 7490 2200 7670
rect 4320 7730 4400 7740
rect 4320 7670 4330 7730
rect 4330 7670 4390 7730
rect 4390 7670 4400 7730
rect 4320 7490 4400 7670
rect 6520 7730 6600 7740
rect 6520 7670 6530 7730
rect 6530 7670 6590 7730
rect 6590 7670 6600 7730
rect 6520 7490 6600 7670
rect 8720 7730 8800 7740
rect 8720 7670 8730 7730
rect 8730 7670 8790 7730
rect 8790 7670 8800 7730
rect 8720 7490 8800 7670
rect 10920 7730 11000 7740
rect 10920 7670 10930 7730
rect 10930 7670 10990 7730
rect 10990 7670 11000 7730
rect 10920 7490 11000 7670
rect 13120 7730 13200 7740
rect 13120 7670 13130 7730
rect 13130 7670 13190 7730
rect 13190 7670 13200 7730
rect 13120 7490 13200 7670
rect 15320 7730 15400 7740
rect 15320 7670 15330 7730
rect 15330 7670 15390 7730
rect 15390 7670 15400 7730
rect 15320 7490 15400 7670
rect 17520 7730 17600 7740
rect 17520 7670 17530 7730
rect 17530 7670 17590 7730
rect 17590 7670 17600 7730
rect 17520 7490 17600 7670
rect 19720 7730 19800 7740
rect 19720 7670 19730 7730
rect 19730 7670 19790 7730
rect 19790 7670 19800 7730
rect 19720 7490 19800 7670
rect 21920 7730 22000 7740
rect 21920 7670 21930 7730
rect 21930 7670 21990 7730
rect 21990 7670 22000 7730
rect 21920 7490 22000 7670
rect 430 7310 610 7390
rect 1630 7310 1810 7390
rect 20110 7310 20290 7390
rect 21310 7310 21490 7390
rect 830 7170 1010 7250
rect 20510 7170 20690 7250
rect 1230 7030 1410 7110
rect 20910 7030 21090 7110
rect -80 6930 0 6940
rect -80 6870 -70 6930
rect -70 6870 -10 6930
rect -10 6870 0 6930
rect -80 6690 0 6870
rect 2120 6930 2200 6940
rect 2120 6870 2130 6930
rect 2130 6870 2190 6930
rect 2190 6870 2200 6930
rect 2120 6690 2200 6870
rect 4320 6930 4400 6940
rect 4320 6870 4330 6930
rect 4330 6870 4390 6930
rect 4390 6870 4400 6930
rect 4320 6690 4400 6870
rect 6520 6930 6600 6940
rect 6520 6870 6530 6930
rect 6530 6870 6590 6930
rect 6590 6870 6600 6930
rect 6520 6690 6600 6870
rect 8720 6930 8800 6940
rect 8720 6870 8730 6930
rect 8730 6870 8790 6930
rect 8790 6870 8800 6930
rect 8720 6690 8800 6870
rect 10920 6930 11000 6940
rect 10920 6870 10930 6930
rect 10930 6870 10990 6930
rect 10990 6870 11000 6930
rect 10920 6690 11000 6870
rect 13120 6930 13200 6940
rect 13120 6870 13130 6930
rect 13130 6870 13190 6930
rect 13190 6870 13200 6930
rect 13120 6690 13200 6870
rect 15320 6930 15400 6940
rect 15320 6870 15330 6930
rect 15330 6870 15390 6930
rect 15390 6870 15400 6930
rect 15320 6690 15400 6870
rect 17520 6930 17600 6940
rect 17520 6870 17530 6930
rect 17530 6870 17590 6930
rect 17590 6870 17600 6930
rect 17520 6690 17600 6870
rect 19720 6930 19800 6940
rect 19720 6870 19730 6930
rect 19730 6870 19790 6930
rect 19790 6870 19800 6930
rect 19720 6690 19800 6870
rect 21920 6930 22000 6940
rect 21920 6870 21930 6930
rect 21930 6870 21990 6930
rect 21990 6870 22000 6930
rect 21920 6690 22000 6870
rect 430 6510 610 6590
rect 1630 6510 1810 6590
rect 20110 6510 20290 6590
rect 21310 6510 21490 6590
rect 830 6370 1010 6450
rect 20510 6370 20690 6450
rect 1230 6230 1410 6310
rect 20910 6230 21090 6310
rect -80 6130 0 6140
rect -80 6070 -70 6130
rect -70 6070 -10 6130
rect -10 6070 0 6130
rect -80 5890 0 6070
rect 2120 6130 2200 6140
rect 2120 6070 2130 6130
rect 2130 6070 2190 6130
rect 2190 6070 2200 6130
rect 2120 5890 2200 6070
rect 4320 6130 4400 6140
rect 4320 6070 4330 6130
rect 4330 6070 4390 6130
rect 4390 6070 4400 6130
rect 4320 5890 4400 6070
rect 6520 6130 6600 6140
rect 6520 6070 6530 6130
rect 6530 6070 6590 6130
rect 6590 6070 6600 6130
rect 6520 5890 6600 6070
rect 8720 6130 8800 6140
rect 8720 6070 8730 6130
rect 8730 6070 8790 6130
rect 8790 6070 8800 6130
rect 8720 5890 8800 6070
rect 10920 6130 11000 6140
rect 10920 6070 10930 6130
rect 10930 6070 10990 6130
rect 10990 6070 11000 6130
rect 10920 5890 11000 6070
rect 13120 6130 13200 6140
rect 13120 6070 13130 6130
rect 13130 6070 13190 6130
rect 13190 6070 13200 6130
rect 13120 5890 13200 6070
rect 15320 6130 15400 6140
rect 15320 6070 15330 6130
rect 15330 6070 15390 6130
rect 15390 6070 15400 6130
rect 15320 5890 15400 6070
rect 17520 6130 17600 6140
rect 17520 6070 17530 6130
rect 17530 6070 17590 6130
rect 17590 6070 17600 6130
rect 17520 5890 17600 6070
rect 19720 6130 19800 6140
rect 19720 6070 19730 6130
rect 19730 6070 19790 6130
rect 19790 6070 19800 6130
rect 19720 5890 19800 6070
rect 21920 6130 22000 6140
rect 21920 6070 21930 6130
rect 21930 6070 21990 6130
rect 21990 6070 22000 6130
rect 21920 5890 22000 6070
rect 36230 6080 36410 6260
rect 36530 6080 36710 6260
rect 1630 5710 1810 5790
rect 20110 5710 20290 5790
rect 830 5570 1010 5650
rect 20510 5570 20690 5650
rect 1230 5430 1410 5510
rect 20910 5430 21090 5510
rect -80 5330 0 5340
rect -80 5270 -70 5330
rect -70 5270 -10 5330
rect -10 5270 0 5330
rect -80 5090 0 5270
rect 2120 5330 2200 5340
rect 2120 5270 2130 5330
rect 2130 5270 2190 5330
rect 2190 5270 2200 5330
rect 2120 5090 2200 5270
rect 4320 5330 4400 5340
rect 4320 5270 4330 5330
rect 4330 5270 4390 5330
rect 4390 5270 4400 5330
rect 4320 5090 4400 5270
rect 6520 5330 6600 5340
rect 6520 5270 6530 5330
rect 6530 5270 6590 5330
rect 6590 5270 6600 5330
rect 6520 5090 6600 5270
rect 8720 5330 8800 5340
rect 8720 5270 8730 5330
rect 8730 5270 8790 5330
rect 8790 5270 8800 5330
rect 8720 5090 8800 5270
rect 10920 5330 11000 5340
rect 10920 5270 10930 5330
rect 10930 5270 10990 5330
rect 10990 5270 11000 5330
rect 10920 5090 11000 5270
rect 13120 5330 13200 5340
rect 13120 5270 13130 5330
rect 13130 5270 13190 5330
rect 13190 5270 13200 5330
rect 13120 5090 13200 5270
rect 15320 5330 15400 5340
rect 15320 5270 15330 5330
rect 15330 5270 15390 5330
rect 15390 5270 15400 5330
rect 15320 5090 15400 5270
rect 17520 5330 17600 5340
rect 17520 5270 17530 5330
rect 17530 5270 17590 5330
rect 17590 5270 17600 5330
rect 17520 5090 17600 5270
rect 19720 5330 19800 5340
rect 19720 5270 19730 5330
rect 19730 5270 19790 5330
rect 19790 5270 19800 5330
rect 19720 5090 19800 5270
rect 21920 5330 22000 5340
rect 21920 5270 21930 5330
rect 21930 5270 21990 5330
rect 21990 5270 22000 5330
rect 21920 5090 22000 5270
rect 28500 5240 28660 5400
rect 36870 5100 37010 5320
rect 37130 5100 37270 5320
rect 1630 4910 1810 4990
rect 20110 4910 20290 4990
rect 30080 3860 30260 4040
rect 31680 3860 31860 4040
rect 33130 4010 33290 4110
rect 34870 4010 35190 4090
rect 430 3550 610 3730
rect 21310 3550 21490 3730
rect 1630 3150 1810 3330
rect 20110 3150 20290 3330
rect 7810 2810 7930 2930
rect 26210 3240 26370 3400
rect 480 -4780 660 2220
rect 14910 1320 15030 1980
rect 12880 -1260 13240 -1110
rect 2810 -5350 2990 -5170
rect 21280 -5350 21460 -5170
rect 36030 -5350 36210 -5170
rect 1270 -5750 1450 -5570
rect 20510 -5750 20690 -5570
rect 36230 -5750 36410 -5570
rect 31680 -6150 31860 -5970
rect 14910 -6610 15030 -6490
rect 12950 -6990 13110 -6830
rect 30080 -6950 30190 -6770
rect 30190 -6950 30260 -6770
rect 1260 -7350 1440 -7170
rect 20510 -7350 20530 -7170
rect 20530 -7350 20690 -7170
rect 36530 -7350 36710 -7170
rect 2080 -7750 2260 -7570
rect 22070 -7750 22250 -7570
rect 36230 -7750 36410 -7570
rect 7810 -7990 7930 -7870
rect 490 -22380 670 -8090
rect 34910 -16920 35050 -16770
rect 34910 -22610 35050 -22470
rect 1630 -23450 1810 -23270
rect 20110 -23450 20290 -23270
rect 430 -23850 610 -23670
rect 21310 -23850 21490 -23670
rect 28500 -24200 28660 -24040
rect 1630 -25110 1810 -25030
rect 20110 -25110 20290 -25030
rect 36870 -24780 37010 -24640
rect 37130 -24780 37270 -24640
rect 33030 -25000 33290 -24930
rect 33230 -25150 33490 -25080
rect 830 -25630 1010 -25550
rect 20510 -25630 20690 -25550
rect 1230 -25770 1410 -25690
rect 20910 -25770 21090 -25690
rect 1630 -25910 1810 -25830
rect 20110 -25910 20290 -25830
rect 830 -26430 1010 -26350
rect 20510 -26430 20690 -26350
rect 1230 -26570 1410 -26490
rect 20910 -26570 21090 -26490
rect 430 -26710 610 -26630
rect 1630 -26710 1810 -26630
rect 20110 -26710 20290 -26630
rect 21310 -26710 21490 -26630
rect 36030 -27140 36410 -27010
rect 36530 -27140 36910 -27010
rect 830 -27230 1010 -27150
rect 20510 -27230 20690 -27150
rect 1230 -27370 1410 -27290
rect 20910 -27370 21090 -27290
rect 430 -27510 610 -27430
rect 1630 -27510 1810 -27430
rect 20110 -27510 20290 -27430
rect 21310 -27510 21490 -27430
rect 830 -28030 1010 -27950
rect 20510 -28030 20690 -27950
rect 1230 -28170 1410 -28090
rect 20910 -28170 21090 -28090
rect 430 -28310 610 -28230
rect 1630 -28310 1810 -28230
rect 20110 -28310 20290 -28230
rect 21310 -28310 21490 -28230
rect 31820 -28290 33160 -28050
rect 830 -28830 1010 -28750
rect 20510 -28830 20690 -28750
rect 1230 -28970 1410 -28890
rect 20910 -28970 21090 -28890
rect 430 -29110 610 -29030
rect 1630 -29110 1810 -29030
rect 20110 -29110 20290 -29030
rect 21310 -29110 21490 -29030
rect 830 -29630 1010 -29550
rect 20510 -29630 20690 -29550
rect 1230 -29770 1410 -29690
rect 20910 -29770 21090 -29690
rect 1630 -29910 1810 -29830
rect 20110 -29910 20290 -29830
rect 37250 -30110 37690 -29920
rect 830 -30430 1010 -30350
rect 20510 -30430 20690 -30350
rect 1230 -30570 1410 -30490
rect 20910 -30570 21090 -30490
rect 1630 -30710 1810 -30630
rect 20110 -30710 20290 -30630
rect 830 -31230 1010 -31150
rect 20510 -31230 20690 -31150
rect 1230 -31370 1410 -31290
rect 20910 -31370 21090 -31290
rect 32540 -31950 33690 -31730
<< metal4 >>
rect 36470 11980 36820 11990
rect 36470 11900 36480 11980
rect -180 11510 36480 11900
rect 36810 11900 36820 11980
rect 36810 11510 37700 11900
rect -180 11500 37700 11510
rect -180 10940 100 11500
rect -180 10690 -80 10940
rect 0 10690 100 10940
rect -180 10140 100 10690
rect -180 9890 -80 10140
rect 0 9890 100 10140
rect -180 9340 100 9890
rect -180 9090 -80 9340
rect 0 9090 100 9340
rect -180 8540 100 9090
rect -180 8290 -80 8540
rect 0 8290 100 8540
rect -180 7740 100 8290
rect -180 7490 -80 7740
rect 0 7490 100 7740
rect -180 6940 100 7490
rect -180 6690 -80 6940
rect 0 6690 100 6940
rect -180 6140 100 6690
rect -180 5890 -80 6140
rect 0 5890 100 6140
rect -180 5340 100 5890
rect -180 5090 -80 5340
rect 0 5090 100 5340
rect -180 2240 100 5090
rect 420 8990 620 11300
rect 420 8910 430 8990
rect 610 8910 620 8990
rect 420 8190 620 8910
rect 420 8110 430 8190
rect 610 8110 620 8190
rect 420 7390 620 8110
rect 420 7310 430 7390
rect 610 7310 620 7390
rect 420 6590 620 7310
rect 420 6510 430 6590
rect 610 6510 620 6590
rect 420 3730 620 6510
rect 420 3550 430 3730
rect 610 3550 620 3730
rect 420 3540 620 3550
rect 820 11250 1020 11300
rect 820 11170 830 11250
rect 1010 11170 1020 11250
rect 820 10450 1020 11170
rect 820 10370 830 10450
rect 1010 10370 1020 10450
rect 820 9650 1020 10370
rect 820 9570 830 9650
rect 1010 9570 1020 9650
rect 820 8850 1020 9570
rect 820 8770 830 8850
rect 1010 8770 1020 8850
rect 820 8050 1020 8770
rect 820 7970 830 8050
rect 1010 7970 1020 8050
rect 820 7250 1020 7970
rect 820 7170 830 7250
rect 1010 7170 1020 7250
rect 820 6450 1020 7170
rect 820 6370 830 6450
rect 1010 6370 1020 6450
rect 820 5650 1020 6370
rect 820 5570 830 5650
rect 1010 5570 1020 5650
rect -180 2220 670 2240
rect -180 2000 480 2220
rect 470 -4780 480 2000
rect 660 -4780 670 2220
rect 820 2210 1020 5570
rect 1220 11110 1420 11300
rect 1220 11030 1230 11110
rect 1410 11030 1420 11110
rect 1220 10310 1420 11030
rect 1220 10230 1230 10310
rect 1410 10230 1420 10310
rect 1220 9510 1420 10230
rect 1220 9430 1230 9510
rect 1410 9430 1420 9510
rect 1220 8710 1420 9430
rect 1220 8630 1230 8710
rect 1410 8630 1420 8710
rect 1220 7910 1420 8630
rect 1220 7830 1230 7910
rect 1410 7830 1420 7910
rect 1220 7110 1420 7830
rect 1220 7030 1230 7110
rect 1410 7030 1420 7110
rect 1220 6310 1420 7030
rect 1220 6230 1230 6310
rect 1410 6230 1420 6310
rect 1220 5510 1420 6230
rect 1220 5430 1230 5510
rect 1410 5430 1420 5510
rect 1220 2600 1420 5430
rect 1620 10590 1820 11300
rect 1620 10510 1630 10590
rect 1810 10510 1820 10590
rect 1620 9790 1820 10510
rect 1620 9710 1630 9790
rect 1810 9710 1820 9790
rect 1620 8990 1820 9710
rect 1620 8910 1630 8990
rect 1810 8910 1820 8990
rect 1620 8190 1820 8910
rect 1620 8110 1630 8190
rect 1810 8110 1820 8190
rect 1620 7390 1820 8110
rect 1620 7310 1630 7390
rect 1810 7310 1820 7390
rect 1620 6590 1820 7310
rect 1620 6510 1630 6590
rect 1810 6510 1820 6590
rect 1620 5790 1820 6510
rect 1620 5710 1630 5790
rect 1810 5710 1820 5790
rect 1620 4990 1820 5710
rect 1620 4910 1630 4990
rect 1810 4910 1820 4990
rect 1620 3330 1820 4910
rect 2020 10940 2300 11500
rect 2020 10690 2120 10940
rect 2200 10690 2300 10940
rect 2020 10140 2300 10690
rect 2020 9890 2120 10140
rect 2200 9890 2300 10140
rect 2020 9340 2300 9890
rect 2020 9090 2120 9340
rect 2200 9090 2300 9340
rect 2020 8540 2300 9090
rect 2020 8290 2120 8540
rect 2200 8290 2300 8540
rect 2020 7740 2300 8290
rect 2020 7490 2120 7740
rect 2200 7490 2300 7740
rect 2020 6940 2300 7490
rect 2020 6690 2120 6940
rect 2200 6690 2300 6940
rect 2020 6140 2300 6690
rect 2020 5890 2120 6140
rect 2200 5890 2300 6140
rect 2020 5340 2300 5890
rect 2020 5090 2120 5340
rect 2200 5090 2300 5340
rect 2020 3660 2300 5090
rect 4220 10940 4500 11500
rect 4220 10690 4320 10940
rect 4400 10690 4500 10940
rect 4220 10140 4500 10690
rect 4220 9890 4320 10140
rect 4400 9890 4500 10140
rect 4220 9340 4500 9890
rect 4220 9090 4320 9340
rect 4400 9090 4500 9340
rect 4220 8540 4500 9090
rect 4220 8290 4320 8540
rect 4400 8290 4500 8540
rect 4220 7740 4500 8290
rect 4220 7490 4320 7740
rect 4400 7490 4500 7740
rect 4220 6940 4500 7490
rect 4220 6690 4320 6940
rect 4400 6690 4500 6940
rect 4220 6140 4500 6690
rect 4220 5890 4320 6140
rect 4400 5890 4500 6140
rect 4220 5340 4500 5890
rect 4220 5090 4320 5340
rect 4400 5090 4500 5340
rect 4220 3660 4500 5090
rect 6420 10940 6700 11500
rect 6420 10690 6520 10940
rect 6600 10690 6700 10940
rect 6420 10140 6700 10690
rect 6420 9890 6520 10140
rect 6600 9890 6700 10140
rect 6420 9340 6700 9890
rect 6420 9090 6520 9340
rect 6600 9090 6700 9340
rect 6420 8540 6700 9090
rect 6420 8290 6520 8540
rect 6600 8290 6700 8540
rect 6420 7740 6700 8290
rect 6420 7490 6520 7740
rect 6600 7490 6700 7740
rect 6420 6940 6700 7490
rect 6420 6690 6520 6940
rect 6600 6690 6700 6940
rect 6420 6140 6700 6690
rect 6420 5890 6520 6140
rect 6600 5890 6700 6140
rect 6420 5340 6700 5890
rect 6420 5090 6520 5340
rect 6600 5090 6700 5340
rect 6420 3660 6700 5090
rect 8620 10940 8900 11500
rect 8620 10690 8720 10940
rect 8800 10690 8900 10940
rect 8620 10140 8900 10690
rect 8620 9890 8720 10140
rect 8800 9890 8900 10140
rect 8620 9340 8900 9890
rect 8620 9090 8720 9340
rect 8800 9090 8900 9340
rect 8620 8540 8900 9090
rect 8620 8290 8720 8540
rect 8800 8290 8900 8540
rect 8620 7740 8900 8290
rect 8620 7490 8720 7740
rect 8800 7490 8900 7740
rect 8620 6940 8900 7490
rect 8620 6690 8720 6940
rect 8800 6690 8900 6940
rect 8620 6140 8900 6690
rect 8620 5890 8720 6140
rect 8800 5890 8900 6140
rect 8620 5340 8900 5890
rect 8620 5090 8720 5340
rect 8800 5090 8900 5340
rect 8620 3660 8900 5090
rect 10820 10940 11100 11500
rect 10820 10690 10920 10940
rect 11000 10690 11100 10940
rect 10820 10140 11100 10690
rect 10820 9890 10920 10140
rect 11000 9890 11100 10140
rect 10820 9340 11100 9890
rect 10820 9090 10920 9340
rect 11000 9090 11100 9340
rect 10820 8540 11100 9090
rect 10820 8290 10920 8540
rect 11000 8290 11100 8540
rect 10820 7740 11100 8290
rect 10820 7490 10920 7740
rect 11000 7490 11100 7740
rect 10820 6940 11100 7490
rect 10820 6690 10920 6940
rect 11000 6690 11100 6940
rect 10820 6140 11100 6690
rect 10820 5890 10920 6140
rect 11000 5890 11100 6140
rect 10820 5340 11100 5890
rect 10820 5090 10920 5340
rect 11000 5090 11100 5340
rect 10820 3660 11100 5090
rect 13020 10940 13300 11500
rect 13020 10690 13120 10940
rect 13200 10690 13300 10940
rect 13020 10140 13300 10690
rect 13020 9890 13120 10140
rect 13200 9890 13300 10140
rect 13020 9340 13300 9890
rect 13020 9090 13120 9340
rect 13200 9090 13300 9340
rect 13020 8540 13300 9090
rect 13020 8290 13120 8540
rect 13200 8290 13300 8540
rect 13020 7740 13300 8290
rect 13020 7490 13120 7740
rect 13200 7490 13300 7740
rect 13020 6940 13300 7490
rect 13020 6690 13120 6940
rect 13200 6690 13300 6940
rect 13020 6140 13300 6690
rect 13020 5890 13120 6140
rect 13200 5890 13300 6140
rect 13020 5340 13300 5890
rect 13020 5090 13120 5340
rect 13200 5090 13300 5340
rect 13020 3660 13300 5090
rect 15220 10940 15500 11500
rect 15220 10690 15320 10940
rect 15400 10690 15500 10940
rect 15220 10140 15500 10690
rect 15220 9890 15320 10140
rect 15400 9890 15500 10140
rect 15220 9340 15500 9890
rect 15220 9090 15320 9340
rect 15400 9090 15500 9340
rect 15220 8540 15500 9090
rect 15220 8290 15320 8540
rect 15400 8290 15500 8540
rect 15220 7740 15500 8290
rect 15220 7490 15320 7740
rect 15400 7490 15500 7740
rect 15220 6940 15500 7490
rect 15220 6690 15320 6940
rect 15400 6690 15500 6940
rect 15220 6140 15500 6690
rect 15220 5890 15320 6140
rect 15400 5890 15500 6140
rect 15220 5340 15500 5890
rect 15220 5090 15320 5340
rect 15400 5090 15500 5340
rect 15220 3660 15500 5090
rect 17420 10940 17700 11500
rect 17420 10690 17520 10940
rect 17600 10690 17700 10940
rect 17420 10140 17700 10690
rect 17420 9890 17520 10140
rect 17600 9890 17700 10140
rect 17420 9340 17700 9890
rect 17420 9090 17520 9340
rect 17600 9090 17700 9340
rect 17420 8540 17700 9090
rect 17420 8290 17520 8540
rect 17600 8290 17700 8540
rect 17420 7740 17700 8290
rect 17420 7490 17520 7740
rect 17600 7490 17700 7740
rect 17420 6940 17700 7490
rect 17420 6690 17520 6940
rect 17600 6690 17700 6940
rect 17420 6140 17700 6690
rect 17420 5890 17520 6140
rect 17600 5890 17700 6140
rect 17420 5340 17700 5890
rect 17420 5090 17520 5340
rect 17600 5090 17700 5340
rect 17420 3660 17700 5090
rect 19620 10940 19900 11500
rect 19620 10690 19720 10940
rect 19800 10690 19900 10940
rect 19620 10140 19900 10690
rect 19620 9890 19720 10140
rect 19800 9890 19900 10140
rect 19620 9340 19900 9890
rect 19620 9090 19720 9340
rect 19800 9090 19900 9340
rect 19620 8540 19900 9090
rect 19620 8290 19720 8540
rect 19800 8290 19900 8540
rect 19620 7740 19900 8290
rect 19620 7490 19720 7740
rect 19800 7490 19900 7740
rect 19620 6940 19900 7490
rect 19620 6690 19720 6940
rect 19800 6690 19900 6940
rect 19620 6140 19900 6690
rect 19620 5890 19720 6140
rect 19800 5890 19900 6140
rect 19620 5340 19900 5890
rect 19620 5090 19720 5340
rect 19800 5090 19900 5340
rect 19620 3660 19900 5090
rect 20100 10590 20300 11300
rect 20100 10510 20110 10590
rect 20290 10510 20300 10590
rect 20100 9790 20300 10510
rect 20100 9710 20110 9790
rect 20290 9710 20300 9790
rect 20100 8990 20300 9710
rect 20100 8910 20110 8990
rect 20290 8910 20300 8990
rect 20100 8190 20300 8910
rect 20100 8110 20110 8190
rect 20290 8110 20300 8190
rect 20100 7390 20300 8110
rect 20100 7310 20110 7390
rect 20290 7310 20300 7390
rect 20100 6590 20300 7310
rect 20100 6510 20110 6590
rect 20290 6510 20300 6590
rect 20100 5790 20300 6510
rect 20100 5710 20110 5790
rect 20290 5710 20300 5790
rect 20100 4990 20300 5710
rect 20100 4910 20110 4990
rect 20290 4910 20300 4990
rect 1620 3150 1630 3330
rect 1810 3150 1820 3330
rect 1620 3140 1820 3150
rect 20100 3330 20300 4910
rect 20100 3150 20110 3330
rect 20290 3150 20300 3330
rect 20100 3140 20300 3150
rect 20500 11250 20700 11300
rect 20500 11170 20510 11250
rect 20690 11170 20700 11250
rect 20500 10450 20700 11170
rect 20500 10370 20510 10450
rect 20690 10370 20700 10450
rect 20500 9650 20700 10370
rect 20500 9570 20510 9650
rect 20690 9570 20700 9650
rect 20500 8850 20700 9570
rect 20500 8770 20510 8850
rect 20690 8770 20700 8850
rect 20500 8050 20700 8770
rect 20500 7970 20510 8050
rect 20690 7970 20700 8050
rect 20500 7250 20700 7970
rect 20500 7170 20510 7250
rect 20690 7170 20700 7250
rect 20500 6450 20700 7170
rect 20500 6370 20510 6450
rect 20690 6370 20700 6450
rect 20500 5650 20700 6370
rect 20500 5570 20510 5650
rect 20690 5570 20700 5650
rect 7800 2930 7940 2940
rect 7800 2810 7810 2930
rect 7930 2810 7940 2930
rect 1220 2400 2270 2600
rect 820 2010 1460 2210
rect 470 -4800 670 -4780
rect 1260 -5570 1460 2010
rect 1260 -5750 1270 -5570
rect 1450 -5750 1460 -5570
rect 1260 -5760 1460 -5750
rect 1250 -7170 1450 -7160
rect 1250 -7350 1260 -7170
rect 1440 -7350 1450 -7170
rect 480 -8090 680 -8080
rect 480 -22200 490 -8090
rect -260 -22380 490 -22200
rect 670 -22380 680 -8090
rect -260 -22400 680 -22380
rect 1250 -22400 1450 -7350
rect 2070 -7570 2270 2400
rect 2070 -7750 2080 -7570
rect 2260 -7750 2270 -7570
rect 2070 -7760 2270 -7750
rect 2800 -5170 3000 -5160
rect 2800 -5350 2810 -5170
rect 2990 -5350 3000 -5170
rect -260 -31660 -60 -22400
rect 820 -22600 1460 -22400
rect 420 -23670 620 -23660
rect 420 -23850 430 -23670
rect 610 -23850 620 -23670
rect 420 -26630 620 -23850
rect 420 -26710 430 -26630
rect 610 -26710 620 -26630
rect 420 -27430 620 -26710
rect 420 -27510 430 -27430
rect 610 -27510 620 -27430
rect 420 -28230 620 -27510
rect 420 -28310 430 -28230
rect 610 -28310 620 -28230
rect 420 -29030 620 -28310
rect 420 -29110 430 -29030
rect 610 -29110 620 -29030
rect 420 -31420 620 -29110
rect 820 -25550 1020 -22600
rect 2800 -22800 3000 -5350
rect 7800 -7870 7940 2810
rect 14900 1980 15040 1990
rect 14900 1320 14910 1980
rect 15030 1320 15040 1980
rect 12870 -1110 13250 -1100
rect 12870 -1260 12880 -1110
rect 13240 -1260 13250 -1110
rect 12870 -1290 13250 -1260
rect 12980 -6820 13080 -1290
rect 14900 -6490 15040 1320
rect 20500 -5570 20700 5570
rect 20900 11110 21100 11300
rect 20900 11030 20910 11110
rect 21090 11030 21100 11110
rect 20900 10310 21100 11030
rect 20900 10230 20910 10310
rect 21090 10230 21100 10310
rect 20900 9510 21100 10230
rect 20900 9430 20910 9510
rect 21090 9430 21100 9510
rect 20900 8710 21100 9430
rect 20900 8630 20910 8710
rect 21090 8630 21100 8710
rect 20900 7910 21100 8630
rect 20900 7830 20910 7910
rect 21090 7830 21100 7910
rect 20900 7110 21100 7830
rect 20900 7030 20910 7110
rect 21090 7030 21100 7110
rect 20900 6310 21100 7030
rect 20900 6230 20910 6310
rect 21090 6230 21100 6310
rect 20900 5510 21100 6230
rect 20900 5430 20910 5510
rect 21090 5430 21100 5510
rect 20900 3340 21100 5430
rect 21300 8990 21500 11300
rect 21300 8910 21310 8990
rect 21490 8910 21500 8990
rect 21300 8190 21500 8910
rect 21300 8110 21310 8190
rect 21490 8110 21500 8190
rect 21300 7390 21500 8110
rect 21300 7310 21310 7390
rect 21490 7310 21500 7390
rect 21300 6590 21500 7310
rect 21300 6510 21310 6590
rect 21490 6510 21500 6590
rect 21300 3730 21500 6510
rect 21300 3550 21310 3730
rect 21490 3550 21500 3730
rect 21820 10940 22100 11500
rect 21820 10690 21920 10940
rect 22000 10690 22100 10940
rect 21820 10140 22100 10690
rect 21820 9890 21920 10140
rect 22000 9890 22100 10140
rect 21820 9340 22100 9890
rect 21820 9090 21920 9340
rect 22000 9090 22100 9340
rect 21820 8540 22100 9090
rect 21820 8290 21920 8540
rect 22000 8290 22100 8540
rect 21820 7740 22100 8290
rect 36780 8170 37020 8180
rect 36780 8030 36790 8170
rect 37010 8030 37020 8170
rect 36780 8020 37020 8030
rect 21820 7490 21920 7740
rect 22000 7490 22100 7740
rect 21820 6940 22100 7490
rect 21820 6690 21920 6940
rect 22000 6690 22100 6940
rect 21820 6140 22100 6690
rect 21820 5890 21920 6140
rect 22000 5890 22100 6140
rect 36220 6260 36420 6270
rect 36220 6080 36230 6260
rect 36410 6080 36420 6260
rect 36220 6070 36420 6080
rect 21820 5340 22100 5890
rect 21820 5090 21920 5340
rect 22000 5090 22100 5340
rect 28490 5400 28670 5410
rect 28490 5240 28500 5400
rect 28660 5240 28670 5400
rect 28490 5230 28670 5240
rect 21820 3660 22100 5090
rect 21300 3540 21500 3550
rect 26200 3400 26380 3410
rect 20900 3140 22260 3340
rect 26200 3240 26210 3400
rect 26370 3370 26380 3400
rect 28530 3370 28630 5230
rect 33120 4110 33300 4120
rect 26370 3270 28630 3370
rect 26370 3240 26380 3270
rect 26200 3230 26380 3240
rect 20500 -5750 20510 -5570
rect 20690 -5750 20700 -5570
rect 20500 -5760 20700 -5750
rect 21270 -5170 21470 -5160
rect 21270 -5350 21280 -5170
rect 21460 -5350 21470 -5170
rect 14900 -6610 14910 -6490
rect 15030 -6610 15040 -6490
rect 14900 -6620 15040 -6610
rect 12940 -6830 13120 -6820
rect 12940 -6990 12950 -6830
rect 13110 -6990 13120 -6830
rect 12940 -7000 13120 -6990
rect 7800 -7990 7810 -7870
rect 7930 -7990 7940 -7870
rect 7800 -8000 7940 -7990
rect 20500 -7170 20700 -7160
rect 20500 -7350 20510 -7170
rect 20690 -7350 20700 -7170
rect 820 -25630 830 -25550
rect 1010 -25630 1020 -25550
rect 820 -26350 1020 -25630
rect 820 -26430 830 -26350
rect 1010 -26430 1020 -26350
rect 820 -27150 1020 -26430
rect 820 -27230 830 -27150
rect 1010 -27230 1020 -27150
rect 820 -27950 1020 -27230
rect 820 -28030 830 -27950
rect 1010 -28030 1020 -27950
rect 820 -28750 1020 -28030
rect 820 -28830 830 -28750
rect 1010 -28830 1020 -28750
rect 820 -29550 1020 -28830
rect 820 -29630 830 -29550
rect 1010 -29630 1020 -29550
rect 820 -30350 1020 -29630
rect 820 -30430 830 -30350
rect 1010 -30430 1020 -30350
rect 820 -31150 1020 -30430
rect 820 -31230 830 -31150
rect 1010 -31230 1020 -31150
rect 820 -31420 1020 -31230
rect 1220 -23000 3000 -22800
rect 1220 -25690 1420 -23000
rect 1220 -25770 1230 -25690
rect 1410 -25770 1420 -25690
rect 1220 -26490 1420 -25770
rect 1220 -26570 1230 -26490
rect 1410 -26570 1420 -26490
rect 1220 -27290 1420 -26570
rect 1220 -27370 1230 -27290
rect 1410 -27370 1420 -27290
rect 1220 -28090 1420 -27370
rect 1220 -28170 1230 -28090
rect 1410 -28170 1420 -28090
rect 1220 -28890 1420 -28170
rect 1220 -28970 1230 -28890
rect 1410 -28970 1420 -28890
rect 1220 -29690 1420 -28970
rect 1220 -29770 1230 -29690
rect 1410 -29770 1420 -29690
rect 1220 -30490 1420 -29770
rect 1220 -30570 1230 -30490
rect 1410 -30570 1420 -30490
rect 1220 -31290 1420 -30570
rect 1220 -31370 1230 -31290
rect 1410 -31370 1420 -31290
rect 1220 -31420 1420 -31370
rect 1620 -23270 1820 -23260
rect 1620 -23450 1630 -23270
rect 1810 -23450 1820 -23270
rect 1620 -25030 1820 -23450
rect 1620 -25110 1630 -25030
rect 1810 -25110 1820 -25030
rect 1620 -25830 1820 -25110
rect 1620 -25910 1630 -25830
rect 1810 -25910 1820 -25830
rect 1620 -26630 1820 -25910
rect 1620 -26710 1630 -26630
rect 1810 -26710 1820 -26630
rect 1620 -27430 1820 -26710
rect 1620 -27510 1630 -27430
rect 1810 -27510 1820 -27430
rect 1620 -28230 1820 -27510
rect 1620 -28310 1630 -28230
rect 1810 -28310 1820 -28230
rect 1620 -29030 1820 -28310
rect 1620 -29110 1630 -29030
rect 1810 -29110 1820 -29030
rect 1620 -29830 1820 -29110
rect 1620 -29910 1630 -29830
rect 1810 -29910 1820 -29830
rect 1620 -30630 1820 -29910
rect 1620 -30710 1630 -30630
rect 1810 -30710 1820 -30630
rect 1620 -31420 1820 -30710
rect 20100 -23270 20300 -23260
rect 20100 -23450 20110 -23270
rect 20290 -23450 20300 -23270
rect 20100 -25030 20300 -23450
rect 20100 -25110 20110 -25030
rect 20290 -25110 20300 -25030
rect 20100 -25830 20300 -25110
rect 20100 -25910 20110 -25830
rect 20290 -25910 20300 -25830
rect 20100 -26630 20300 -25910
rect 20100 -26710 20110 -26630
rect 20290 -26710 20300 -26630
rect 20100 -27430 20300 -26710
rect 20100 -27510 20110 -27430
rect 20290 -27510 20300 -27430
rect 20100 -28230 20300 -27510
rect 20100 -28310 20110 -28230
rect 20290 -28310 20300 -28230
rect 20100 -29030 20300 -28310
rect 20100 -29110 20110 -29030
rect 20290 -29110 20300 -29030
rect 20100 -29830 20300 -29110
rect 20100 -29910 20110 -29830
rect 20290 -29910 20300 -29830
rect 20100 -30630 20300 -29910
rect 20100 -30710 20110 -30630
rect 20290 -30710 20300 -30630
rect 20100 -31420 20300 -30710
rect 20500 -25550 20700 -7350
rect 21270 -22420 21470 -5350
rect 22060 -7570 22260 3140
rect 22060 -7750 22070 -7570
rect 22250 -7750 22260 -7570
rect 22060 -7760 22260 -7750
rect 20500 -25630 20510 -25550
rect 20690 -25630 20700 -25550
rect 20500 -26350 20700 -25630
rect 20500 -26430 20510 -26350
rect 20690 -26430 20700 -26350
rect 20500 -27150 20700 -26430
rect 20500 -27230 20510 -27150
rect 20690 -27230 20700 -27150
rect 20500 -27950 20700 -27230
rect 20500 -28030 20510 -27950
rect 20690 -28030 20700 -27950
rect 20500 -28750 20700 -28030
rect 20500 -28830 20510 -28750
rect 20690 -28830 20700 -28750
rect 20500 -29550 20700 -28830
rect 20500 -29630 20510 -29550
rect 20690 -29630 20700 -29550
rect 20500 -30350 20700 -29630
rect 20500 -30430 20510 -30350
rect 20690 -30430 20700 -30350
rect 20500 -31150 20700 -30430
rect 20500 -31230 20510 -31150
rect 20690 -31230 20700 -31150
rect 20500 -31420 20700 -31230
rect 20900 -22620 21470 -22420
rect 20900 -25690 21100 -22620
rect 20900 -25770 20910 -25690
rect 21090 -25770 21100 -25690
rect 20900 -26490 21100 -25770
rect 20900 -26570 20910 -26490
rect 21090 -26570 21100 -26490
rect 20900 -27290 21100 -26570
rect 20900 -27370 20910 -27290
rect 21090 -27370 21100 -27290
rect 20900 -28090 21100 -27370
rect 20900 -28170 20910 -28090
rect 21090 -28170 21100 -28090
rect 20900 -28890 21100 -28170
rect 20900 -28970 20910 -28890
rect 21090 -28970 21100 -28890
rect 20900 -29690 21100 -28970
rect 20900 -29770 20910 -29690
rect 21090 -29770 21100 -29690
rect 20900 -30490 21100 -29770
rect 20900 -30570 20910 -30490
rect 21090 -30570 21100 -30490
rect 20900 -31290 21100 -30570
rect 20900 -31370 20910 -31290
rect 21090 -31370 21100 -31290
rect 20900 -31420 21100 -31370
rect 21300 -23670 21500 -23660
rect 21300 -23850 21310 -23670
rect 21490 -23850 21500 -23670
rect 21300 -26630 21500 -23850
rect 28530 -24030 28630 3270
rect 30070 4040 30270 4050
rect 30070 3860 30080 4040
rect 30260 3860 30270 4040
rect 30070 -6770 30270 3860
rect 31670 4040 31870 4050
rect 31670 3860 31680 4040
rect 31860 3860 31870 4040
rect 33120 4010 33130 4110
rect 33290 4010 33300 4110
rect 33120 4000 33300 4010
rect 31670 -5970 31870 3860
rect 31670 -6150 31680 -5970
rect 31860 -6150 31870 -5970
rect 31670 -6160 31870 -6150
rect 30070 -6950 30080 -6770
rect 30260 -6950 30270 -6770
rect 30070 -6960 30270 -6950
rect 28490 -24040 28670 -24030
rect 28490 -24200 28500 -24040
rect 28660 -24200 28670 -24040
rect 28490 -24210 28670 -24200
rect 33200 -24920 33300 4000
rect 33020 -24930 33300 -24920
rect 33020 -25000 33030 -24930
rect 33290 -25000 33300 -24930
rect 33020 -25010 33300 -25000
rect 33400 4090 35200 4100
rect 33400 4010 34870 4090
rect 35190 4010 35200 4090
rect 33400 4000 35200 4010
rect 33400 -25070 33500 4000
rect 36020 -5170 36220 -5160
rect 36020 -5350 36030 -5170
rect 36210 -5350 36220 -5170
rect 36020 -5360 36220 -5350
rect 36020 -7870 36120 -5360
rect 36320 -5560 36420 6070
rect 36220 -5570 36420 -5560
rect 36220 -5750 36230 -5570
rect 36410 -5750 36420 -5570
rect 36220 -5760 36420 -5750
rect 36520 6260 36720 6270
rect 36520 6080 36530 6260
rect 36710 6080 36720 6260
rect 36520 6070 36720 6080
rect 36520 -6900 36620 6070
rect 36920 5330 37020 8020
rect 36860 5320 37020 5330
rect 36860 5100 36870 5320
rect 37010 5100 37020 5320
rect 36860 5090 37020 5100
rect 36320 -7000 36620 -6900
rect 36320 -7560 36420 -7000
rect 36220 -7570 36420 -7560
rect 36220 -7750 36230 -7570
rect 36410 -7750 36420 -7570
rect 36220 -7760 36420 -7750
rect 36520 -7170 36720 -7160
rect 36520 -7350 36530 -7170
rect 36710 -7350 36720 -7170
rect 36520 -7360 36720 -7350
rect 36020 -7970 36420 -7870
rect 34900 -16770 35060 -16740
rect 34900 -16920 34910 -16770
rect 35050 -16920 35060 -16770
rect 34900 -22470 35060 -16920
rect 34900 -22610 34910 -22470
rect 35050 -22610 35060 -22470
rect 34900 -22620 35060 -22610
rect 33220 -25080 33500 -25070
rect 33220 -25150 33230 -25080
rect 33490 -25150 33500 -25080
rect 33220 -25160 33500 -25150
rect 21300 -26710 21310 -26630
rect 21490 -26710 21500 -26630
rect 21300 -27430 21500 -26710
rect 36320 -27000 36420 -7970
rect 36020 -27010 36420 -27000
rect 36020 -27140 36030 -27010
rect 36410 -27140 36420 -27010
rect 36020 -27150 36420 -27140
rect 36520 -27000 36620 -7360
rect 36920 -24630 37020 5090
rect 36860 -24640 37020 -24630
rect 36860 -24780 36870 -24640
rect 37010 -24780 37020 -24640
rect 36860 -24790 37020 -24780
rect 37120 7970 37360 7980
rect 37120 7830 37130 7970
rect 37350 7830 37360 7970
rect 37120 7820 37360 7830
rect 37120 5330 37220 7820
rect 37120 5320 37280 5330
rect 37120 5100 37130 5320
rect 37270 5100 37280 5320
rect 37120 5090 37280 5100
rect 37120 -24630 37220 5090
rect 37120 -24640 37280 -24630
rect 37120 -24780 37130 -24640
rect 37270 -24780 37280 -24640
rect 37120 -24790 37280 -24780
rect 36520 -27010 36920 -27000
rect 36520 -27140 36530 -27010
rect 36910 -27140 36920 -27010
rect 36520 -27150 36920 -27140
rect 21300 -27510 21310 -27430
rect 21490 -27510 21500 -27430
rect 21300 -28230 21500 -27510
rect 21300 -28310 21310 -28230
rect 21490 -28310 21500 -28230
rect 21300 -29030 21500 -28310
rect 21300 -29110 21310 -29030
rect 21490 -29110 21500 -29030
rect 21300 -31420 21500 -29110
rect 31320 -28050 37370 -28020
rect 31320 -28290 31820 -28050
rect 33160 -28290 37370 -28050
rect 31320 -28320 37370 -28290
rect 31320 -31660 31520 -28320
rect 37500 -29910 37700 11500
rect 37240 -29920 37700 -29910
rect 37240 -30110 37250 -29920
rect 37690 -30110 37700 -29920
rect 37240 -30120 37700 -30110
rect 37900 9380 38100 11900
rect 37900 9200 37910 9380
rect 38090 9200 38100 9380
rect 37900 -28020 38100 9200
rect 37900 -28320 38160 -28020
rect 37900 -31660 38100 -28320
rect -260 -31730 38100 -31660
rect -260 -31950 32540 -31730
rect 33690 -31950 38100 -31730
rect -260 -32060 38100 -31950
<< res2p85 >>
rect 22364 4996 22938 11384
rect 23030 4996 23604 11384
rect 23696 4996 24270 11384
rect 24362 4996 24936 11384
rect 25028 4996 25602 11384
rect 25694 4996 26268 11384
rect 26360 4996 26934 11384
rect 22345 -31483 22919 -25095
rect 23011 -31483 23585 -25095
rect 23677 -31483 24251 -25095
rect 24343 -31483 24917 -25095
rect 25009 -31483 25583 -25095
rect 25675 -31483 26249 -25095
rect 26341 -31483 26915 -25095
<< labels >>
flabel metal2 80 -6580 280 -6380 0 FreeSans 320 0 0 0 Vinp
port 0 nsew
flabel metal2 -360 -6580 -160 -6380 0 FreeSans 320 0 0 0 Vinm
port 1 nsew
flabel metal4 35940 11600 36140 11800 0 FreeSans 320 0 0 0 AGND
port 3 nsew
flabel metal3 37980 -27960 38080 -27860 0 FreeSans 320 0 0 0 hyst[1]
port 5 nsew
flabel metal3 37980 -28160 38080 -28060 0 FreeSans 320 0 0 0 hyst[0]
port 6 nsew
flabel metal2 31880 -31880 31980 -31780 0 FreeSans 320 0 0 0 trim[5]
port 7 nsew
flabel metal2 34080 -31880 34180 -31780 0 FreeSans 320 0 0 0 trim[4]
port 8 nsew
flabel metal2 36280 -31880 36380 -31780 0 FreeSans 320 0 0 0 trim[3]
port 9 nsew
flabel metal3 37390 9730 37470 9810 0 FreeSans 320 0 0 0 trim[2]
port 10 nsew
flabel metal3 37390 9910 37470 9990 0 FreeSans 320 0 0 0 trim[1]
port 11 nsew
flabel metal3 37390 10090 37470 10170 0 FreeSans 320 0 0 0 trim[0]
port 12 nsew
flabel metal3 530 2400 680 2530 0 FreeSans 320 0 0 0 ibias
port 15 nsew
flabel metal3 37980 -27760 38080 -27660 0 FreeSans 320 0 0 0 en
port 4 nsew
flabel metal1 36480 7560 36610 7680 0 FreeSans 320 0 0 0 Vout
port 13 nsew
flabel metal3 25908 -6132 26054 -5988 0 FreeSans 160 0 0 0 Vom
flabel metal3 25946 -6922 26060 -6808 0 FreeSans 160 0 0 0 Vop
flabel metal3 34058 -5336 34206 -5190 0 FreeSans 160 0 0 0 Vfold_bot_m
flabel metal3 5232 -23424 5384 -23282 0 FreeSans 160 0 0 0 Vxp
flabel metal3 5272 3160 5424 3302 0 FreeSans 160 0 0 0 Vxm
flabel metal2 11724 -850 11812 -754 0 FreeSans 160 0 0 0 bias_n
flabel metal1 12984 -776 13110 -652 0 FreeSans 160 0 0 0 casc_n
flabel metal1 16736 -8368 16836 -8274 0 FreeSans 160 0 0 0 casc_p
flabel metal1 11734 -10518 11822 -10426 0 FreeSans 160 0 0 0 bias_p
flabel metal1 30102 6544 30204 6644 0 FreeSans 160 0 0 0 Vom_stg2
flabel metal1 31422 6544 31524 6644 0 FreeSans 160 0 0 0 Vop_stg2
flabel metal2 15250 -1268 15372 -1144 0 FreeSans 160 0 0 0 bias_var_n
flabel metal3 31130 -28780 31200 -28710 0 FreeSans 160 0 0 0 enb_hv
flabel metal3 31130 -28930 31200 -28860 0 FreeSans 160 0 0 0 en_hv
flabel metal3 31130 -29080 31200 -29010 0 FreeSans 160 0 0 0 hyst1b_hv
flabel metal3 31130 -29230 31200 -29160 0 FreeSans 160 0 0 0 hyst1_hv
flabel metal3 31130 -29380 31200 -29310 0 FreeSans 160 0 0 0 hyst0b_hv
flabel metal3 31130 -29530 31200 -29460 0 FreeSans 160 0 0 0 hyst0_hv
flabel metal2 26540 -29250 26700 -29080 0 FreeSans 160 0 0 0 res_p_bot
flabel metal2 32090 8740 32180 8820 0 FreeSans 160 0 0 0 bias_stg2
flabel metal1 36460 6800 36620 6930 0 FreeSans 320 0 0 0 DGND
port 16 nsew
flabel metal1 36920 8840 37080 9000 0 FreeSans 320 0 0 0 DVDD
port 14 nsew
flabel metal4 30740 -32020 30870 -31870 0 FreeSans 320 0 0 0 AVDD
port 2 nsew
flabel metal3 30640 -30880 30710 -30810 0 FreeSans 320 0 0 0 trim5_hv
flabel metal3 30640 -31030 30710 -30960 0 FreeSans 320 0 0 0 trim5b_hv
flabel metal3 30640 -31180 30710 -31110 0 FreeSans 320 0 0 0 trim4b_hv
flabel metal3 30640 -31330 30710 -31260 0 FreeSans 320 0 0 0 trim3b_hv
flabel metal1 35770 -28340 35830 -28280 0 FreeSans 320 0 0 0 level_shifter_up_0.VDD_HV
flabel metal1 35830 -29980 35890 -29920 0 FreeSans 320 0 0 0 level_shifter_up_0.GND_HV
flabel metal1 35566 -29280 35650 -29220 0 FreeSans 320 0 0 0 level_shifter_up_0.x_lv
flabel metal2 34190 -29270 34250 -29210 0 FreeSans 320 0 0 0 level_shifter_up_0.xb_hv
flabel metal2 34410 -29270 34470 -29210 0 FreeSans 320 0 0 0 level_shifter_up_0.x_hv
flabel metal1 33992 -31744 34052 -31684 0 FreeSans 320 0 0 0 level_shifter_up_2.VDD_HV
flabel metal1 33932 -30104 33992 -30044 0 FreeSans 320 0 0 0 level_shifter_up_2.GND_HV
flabel metal1 34172 -30804 34256 -30744 0 FreeSans 320 0 0 0 level_shifter_up_2.x_lv
flabel metal2 35572 -30814 35632 -30754 0 FreeSans 320 0 0 0 level_shifter_up_2.xb_hv
flabel metal2 35352 -30814 35412 -30754 0 FreeSans 320 0 0 0 level_shifter_up_2.x_hv
flabel metal1 31792 -31744 31852 -31684 0 FreeSans 320 0 0 0 level_shifter_up_3.VDD_HV
flabel metal1 31732 -30104 31792 -30044 0 FreeSans 320 0 0 0 level_shifter_up_3.GND_HV
flabel metal1 31972 -30804 32056 -30744 0 FreeSans 320 0 0 0 level_shifter_up_3.x_lv
flabel metal2 33372 -30814 33432 -30754 0 FreeSans 320 0 0 0 level_shifter_up_3.xb_hv
flabel metal2 33152 -30814 33212 -30754 0 FreeSans 320 0 0 0 level_shifter_up_3.x_hv
flabel metal1 33570 -28340 33630 -28280 0 FreeSans 320 0 0 0 level_shifter_up_4.VDD_HV
flabel metal1 33630 -29980 33690 -29920 0 FreeSans 320 0 0 0 level_shifter_up_4.GND_HV
flabel metal1 33366 -29280 33450 -29220 0 FreeSans 320 0 0 0 level_shifter_up_4.x_lv
flabel metal2 31990 -29270 32050 -29210 0 FreeSans 320 0 0 0 level_shifter_up_4.xb_hv
flabel metal2 32210 -29270 32270 -29210 0 FreeSans 320 0 0 0 level_shifter_up_4.x_hv
flabel metal1 36192 -31744 36252 -31684 0 FreeSans 320 0 0 0 level_shifter_up_1.VDD_HV
flabel metal1 36132 -30104 36192 -30044 0 FreeSans 320 0 0 0 level_shifter_up_1.GND_HV
flabel metal1 36372 -30804 36456 -30744 0 FreeSans 320 0 0 0 level_shifter_up_1.x_lv
flabel metal2 37772 -30814 37832 -30754 0 FreeSans 320 0 0 0 level_shifter_up_1.xb_hv
flabel metal2 37552 -30814 37612 -30754 0 FreeSans 320 0 0 0 level_shifter_up_1.x_hv
flabel metal1 37970 -28340 38030 -28280 0 FreeSans 320 0 0 0 level_shifter_up_5.VDD_HV
flabel metal1 38030 -29980 38090 -29920 0 FreeSans 320 0 0 0 level_shifter_up_5.GND_HV
flabel metal1 37766 -29280 37850 -29220 0 FreeSans 320 0 0 0 level_shifter_up_5.x_lv
flabel metal2 36390 -29270 36450 -29210 0 FreeSans 320 0 0 0 level_shifter_up_5.xb_hv
flabel metal2 36610 -29270 36670 -29210 0 FreeSans 320 0 0 0 level_shifter_up_5.x_hv
flabel metal1 32312 10266 32372 10326 0 FreeSans 320 0 0 0 level_shifter_up_7.VDD_HV
flabel metal1 32252 11906 32312 11966 0 FreeSans 320 0 0 0 level_shifter_up_7.GND_HV
flabel metal1 32492 11206 32576 11266 0 FreeSans 320 0 0 0 level_shifter_up_7.x_lv
flabel metal2 33892 11196 33952 11256 0 FreeSans 320 0 0 0 level_shifter_up_7.xb_hv
flabel metal2 33672 11196 33732 11256 0 FreeSans 320 0 0 0 level_shifter_up_7.x_hv
flabel metal1 30112 10266 30172 10326 0 FreeSans 320 0 0 0 level_shifter_up_6.VDD_HV
flabel metal1 30052 11906 30112 11966 0 FreeSans 320 0 0 0 level_shifter_up_6.GND_HV
flabel metal1 30292 11206 30376 11266 0 FreeSans 320 0 0 0 level_shifter_up_6.x_lv
flabel metal2 31692 11196 31752 11256 0 FreeSans 320 0 0 0 level_shifter_up_6.xb_hv
flabel metal2 31472 11196 31532 11256 0 FreeSans 320 0 0 0 level_shifter_up_6.x_hv
flabel metal1 34512 10266 34572 10326 0 FreeSans 320 0 0 0 level_shifter_up_8.VDD_HV
flabel metal1 34452 11906 34512 11966 0 FreeSans 320 0 0 0 level_shifter_up_8.GND_HV
flabel metal1 34692 11206 34776 11266 0 FreeSans 320 0 0 0 level_shifter_up_8.x_lv
flabel metal2 36092 11196 36152 11256 0 FreeSans 320 0 0 0 level_shifter_up_8.xb_hv
flabel metal2 35872 11196 35932 11256 0 FreeSans 320 0 0 0 level_shifter_up_8.x_hv
<< end >>
