magic
tech sky130A
magscale 1 2
timestamp 1713585847
<< error_p >>
rect -108 272 -50 278
rect 50 272 108 278
rect -108 238 -96 272
rect 50 238 62 272
rect -108 232 -50 238
rect 50 232 108 238
rect -108 -238 -50 -232
rect 50 -238 108 -232
rect -108 -272 -96 -238
rect 50 -272 62 -238
rect -108 -278 -50 -272
rect 50 -278 108 -272
<< pwell >>
rect -357 -458 357 458
<< mvnmos >>
rect -129 -200 -29 200
rect 29 -200 129 200
<< mvndiff >>
rect -187 188 -129 200
rect -187 -188 -175 188
rect -141 -188 -129 188
rect -187 -200 -129 -188
rect -29 188 29 200
rect -29 -188 -17 188
rect 17 -188 29 188
rect -29 -200 29 -188
rect 129 188 187 200
rect 129 -188 141 188
rect 175 -188 187 188
rect 129 -200 187 -188
<< mvndiffc >>
rect -175 -188 -141 188
rect -17 -188 17 188
rect 141 -188 175 188
<< mvpsubdiff >>
rect -321 410 321 422
rect -321 376 -213 410
rect 213 376 321 410
rect -321 364 321 376
rect -321 314 -263 364
rect -321 -314 -309 314
rect -275 -314 -263 314
rect 263 314 321 364
rect -321 -364 -263 -314
rect 263 -314 275 314
rect 309 -314 321 314
rect 263 -364 321 -314
rect -321 -376 321 -364
rect -321 -410 -213 -376
rect 213 -410 321 -376
rect -321 -422 321 -410
<< mvpsubdiffcont >>
rect -213 376 213 410
rect -309 -314 -275 314
rect 275 -314 309 314
rect -213 -410 213 -376
<< poly >>
rect -129 272 -29 288
rect -129 238 -113 272
rect -45 238 -29 272
rect -129 200 -29 238
rect 29 272 129 288
rect 29 238 45 272
rect 113 238 129 272
rect 29 200 129 238
rect -129 -238 -29 -200
rect -129 -272 -113 -238
rect -45 -272 -29 -238
rect -129 -288 -29 -272
rect 29 -238 129 -200
rect 29 -272 45 -238
rect 113 -272 129 -238
rect 29 -288 129 -272
<< polycont >>
rect -113 238 -45 272
rect 45 238 113 272
rect -113 -272 -45 -238
rect 45 -272 113 -238
<< locali >>
rect -309 376 -220 410
rect 220 376 309 410
rect -309 314 -275 376
rect 275 314 309 376
rect -129 238 -113 272
rect -45 238 -29 272
rect 29 238 45 272
rect 113 238 129 272
rect -175 188 -141 204
rect -175 -204 -141 -188
rect -17 188 17 204
rect -17 -204 17 -188
rect 141 188 175 204
rect 141 -204 175 -188
rect -129 -272 -113 -238
rect -45 -272 -29 -238
rect 29 -272 45 -238
rect 113 -272 129 -238
rect -309 -376 -275 -314
rect 275 -376 309 -314
rect -309 -410 -213 -376
rect 213 -410 309 -376
<< viali >>
rect -220 376 -213 410
rect -213 376 213 410
rect 213 376 220 410
rect -309 -301 -275 301
rect -96 238 -62 272
rect 62 238 96 272
rect -175 -188 -141 188
rect -17 -188 17 188
rect 141 -188 175 188
rect -96 -272 -62 -238
rect 62 -272 96 -238
rect 275 -301 309 301
<< metal1 >>
rect -232 410 232 416
rect -232 376 -220 410
rect 220 376 232 410
rect -232 370 232 376
rect -315 301 -269 313
rect -315 -301 -309 301
rect -275 -301 -269 301
rect 269 301 315 313
rect -108 272 -50 278
rect -108 238 -96 272
rect -62 238 -50 272
rect -108 232 -50 238
rect 50 272 108 278
rect 50 238 62 272
rect 96 238 108 272
rect 50 232 108 238
rect -181 188 -135 200
rect -181 -188 -175 188
rect -141 -188 -135 188
rect -181 -200 -135 -188
rect -23 188 23 200
rect -23 -188 -17 188
rect 17 -188 23 188
rect -23 -200 23 -188
rect 135 188 181 200
rect 135 -188 141 188
rect 175 -188 181 188
rect 135 -200 181 -188
rect -108 -238 -50 -232
rect -108 -272 -96 -238
rect -62 -272 -50 -238
rect -108 -278 -50 -272
rect 50 -238 108 -232
rect 50 -272 62 -238
rect 96 -272 108 -238
rect 50 -278 108 -272
rect -315 -313 -269 -301
rect 269 -301 275 301
rect 309 -301 315 301
rect 269 -313 315 -301
<< properties >>
string FIXED_BBOX -292 -393 292 393
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 2 l 0.50 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 80 viagl 80 viagt 80
<< end >>
