magic
tech sky130A
magscale 1 2
timestamp 1713594949
<< pwell >>
rect -533 -1182 533 1182
<< psubdiff >>
rect -497 1112 -401 1146
rect 401 1112 497 1146
rect -497 1050 -463 1112
rect 463 1050 497 1112
rect -497 -1112 -463 -1050
rect 463 -1112 497 -1050
rect -497 -1146 -401 -1112
rect 401 -1146 497 -1112
<< psubdiffcont >>
rect -401 1112 401 1146
rect -497 -1050 -463 1050
rect 463 -1050 497 1050
rect -401 -1146 401 -1112
<< xpolycontact >>
rect -367 584 -297 1016
rect -367 52 -297 484
rect -201 584 -131 1016
rect -201 52 -131 484
rect -35 584 35 1016
rect -35 52 35 484
rect 131 584 201 1016
rect 131 52 201 484
rect 297 584 367 1016
rect 297 52 367 484
rect -367 -484 -297 -52
rect -367 -1016 -297 -584
rect -201 -484 -131 -52
rect -201 -1016 -131 -584
rect -35 -484 35 -52
rect -35 -1016 35 -584
rect 131 -484 201 -52
rect 131 -1016 201 -584
rect 297 -484 367 -52
rect 297 -1016 367 -584
<< xpolyres >>
rect -367 484 -297 584
rect -201 484 -131 584
rect -35 484 35 584
rect 131 484 201 584
rect 297 484 367 584
rect -367 -584 -297 -484
rect -201 -584 -131 -484
rect -35 -584 35 -484
rect 131 -584 201 -484
rect 297 -584 367 -484
<< locali >>
rect -497 1112 -401 1146
rect 401 1112 497 1146
rect -497 1050 -463 1112
rect 463 1050 497 1112
rect -497 -1112 -463 -1050
rect 463 -1112 497 -1050
rect -497 -1146 -401 -1112
rect 401 -1146 497 -1112
<< viali >>
rect -351 601 -313 998
rect -185 601 -147 998
rect -19 601 19 998
rect 147 601 185 998
rect 313 601 351 998
rect -351 70 -313 467
rect -185 70 -147 467
rect -19 70 19 467
rect 147 70 185 467
rect 313 70 351 467
rect -351 -467 -313 -70
rect -185 -467 -147 -70
rect -19 -467 19 -70
rect 147 -467 185 -70
rect 313 -467 351 -70
rect -351 -998 -313 -601
rect -185 -998 -147 -601
rect -19 -998 19 -601
rect 147 -998 185 -601
rect 313 -998 351 -601
<< metal1 >>
rect -357 998 -307 1010
rect -357 601 -351 998
rect -313 601 -307 998
rect -357 589 -307 601
rect -191 998 -141 1010
rect -191 601 -185 998
rect -147 601 -141 998
rect -191 589 -141 601
rect -25 998 25 1010
rect -25 601 -19 998
rect 19 601 25 998
rect -25 589 25 601
rect 141 998 191 1010
rect 141 601 147 998
rect 185 601 191 998
rect 141 589 191 601
rect 307 998 357 1010
rect 307 601 313 998
rect 351 601 357 998
rect 307 589 357 601
rect -357 467 -307 479
rect -357 70 -351 467
rect -313 70 -307 467
rect -357 58 -307 70
rect -191 467 -141 479
rect -191 70 -185 467
rect -147 70 -141 467
rect -191 58 -141 70
rect -25 467 25 479
rect -25 70 -19 467
rect 19 70 25 467
rect -25 58 25 70
rect 141 467 191 479
rect 141 70 147 467
rect 185 70 191 467
rect 141 58 191 70
rect 307 467 357 479
rect 307 70 313 467
rect 351 70 357 467
rect 307 58 357 70
rect -357 -70 -307 -58
rect -357 -467 -351 -70
rect -313 -467 -307 -70
rect -357 -479 -307 -467
rect -191 -70 -141 -58
rect -191 -467 -185 -70
rect -147 -467 -141 -70
rect -191 -479 -141 -467
rect -25 -70 25 -58
rect -25 -467 -19 -70
rect 19 -467 25 -70
rect -25 -479 25 -467
rect 141 -70 191 -58
rect 141 -467 147 -70
rect 185 -467 191 -70
rect 141 -479 191 -467
rect 307 -70 357 -58
rect 307 -467 313 -70
rect 351 -467 357 -70
rect 307 -479 357 -467
rect -357 -601 -307 -589
rect -357 -998 -351 -601
rect -313 -998 -307 -601
rect -357 -1010 -307 -998
rect -191 -601 -141 -589
rect -191 -998 -185 -601
rect -147 -998 -141 -601
rect -191 -1010 -141 -998
rect -25 -601 25 -589
rect -25 -998 -19 -601
rect 19 -998 25 -601
rect -25 -1010 25 -998
rect 141 -601 191 -589
rect 141 -998 147 -601
rect 185 -998 191 -601
rect 141 -1010 191 -998
rect 307 -601 357 -589
rect 307 -998 313 -601
rect 351 -998 357 -601
rect 307 -1010 357 -998
<< res0p35 >>
rect -369 482 -295 586
rect -203 482 -129 586
rect -37 482 37 586
rect 129 482 203 586
rect 295 482 369 586
rect -369 -586 -295 -482
rect -203 -586 -129 -482
rect -37 -586 37 -482
rect 129 -586 203 -482
rect 295 -586 369 -482
<< properties >>
string FIXED_BBOX -480 -1129 480 1129
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 0.50 m 2 nx 5 wmin 0.350 lmin 0.50 rho 2000 val 3.932k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
