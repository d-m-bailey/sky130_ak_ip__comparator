magic
tech sky130A
magscale 1 2
timestamp 1713587824
<< pwell >>
rect -428 -308 428 308
<< mvnmos >>
rect -200 -50 200 50
<< mvndiff >>
rect -258 38 -200 50
rect -258 -38 -246 38
rect -212 -38 -200 38
rect -258 -50 -200 -38
rect 200 38 258 50
rect 200 -38 212 38
rect 246 -38 258 38
rect 200 -50 258 -38
<< mvndiffc >>
rect -246 -38 -212 38
rect 212 -38 246 38
<< mvpsubdiff >>
rect -392 260 392 272
rect -392 226 -284 260
rect 284 226 392 260
rect -392 214 392 226
rect -392 164 -334 214
rect -392 -164 -380 164
rect -346 -164 -334 164
rect 334 164 392 214
rect -392 -214 -334 -164
rect 334 -164 346 164
rect 380 -164 392 164
rect 334 -214 392 -164
rect -392 -226 392 -214
rect -392 -260 -284 -226
rect 284 -260 392 -226
rect -392 -272 392 -260
<< mvpsubdiffcont >>
rect -284 226 284 260
rect -380 -164 -346 164
rect 346 -164 380 164
rect -284 -260 284 -226
<< poly >>
rect -200 122 200 138
rect -200 88 -184 122
rect 184 88 200 122
rect -200 50 200 88
rect -200 -88 200 -50
rect -200 -122 -184 -88
rect 184 -122 200 -88
rect -200 -138 200 -122
<< polycont >>
rect -184 88 184 122
rect -184 -122 184 -88
<< locali >>
rect -380 226 -284 260
rect 284 226 380 260
rect -380 164 -346 226
rect 346 181 380 226
rect -200 88 -184 122
rect 184 88 200 122
rect -246 38 -212 54
rect -246 -54 -212 -38
rect 212 38 246 54
rect 212 -54 246 -38
rect -200 -122 -184 -88
rect 184 -122 200 -88
rect -380 -226 -346 -164
rect 346 -226 380 -181
rect -380 -260 -284 -226
rect 284 -260 380 -226
<< viali >>
rect 346 164 380 181
rect -184 88 184 122
rect -246 -38 -212 38
rect 212 -38 246 38
rect -184 -122 184 -88
rect 346 -164 380 164
rect 346 -181 380 -164
<< metal1 >>
rect 340 181 386 193
rect -196 122 196 128
rect -196 88 -184 122
rect 184 88 196 122
rect -196 82 196 88
rect -252 38 -206 50
rect -252 -38 -246 38
rect -212 -38 -206 38
rect -252 -50 -206 -38
rect 206 38 252 50
rect 206 -38 212 38
rect 246 -38 252 38
rect 206 -50 252 -38
rect -196 -88 196 -82
rect -196 -122 -184 -88
rect 184 -122 196 -88
rect -196 -128 196 -122
rect 340 -181 346 181
rect 380 -181 386 181
rect 340 -193 386 -181
<< properties >>
string FIXED_BBOX -363 -243 363 243
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 0.5 l 2 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 80 viagl 0 viagt 0
<< end >>
