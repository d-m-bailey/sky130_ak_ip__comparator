magic
tech sky130A
magscale 1 2
timestamp 1713598147
<< pwell >>
rect -696 -710 696 710
<< nmos >>
rect -500 -500 500 500
<< ndiff >>
rect -558 488 -500 500
rect -558 -488 -546 488
rect -512 -488 -500 488
rect -558 -500 -500 -488
rect 500 488 558 500
rect 500 -488 512 488
rect 546 -488 558 488
rect 500 -500 558 -488
<< ndiffc >>
rect -546 -488 -512 488
rect 512 -488 546 488
<< psubdiff >>
rect -660 640 -564 674
rect 564 640 660 674
rect -660 578 -626 640
rect 626 578 660 640
rect -660 -640 -626 -578
rect 626 -640 660 -578
rect -660 -674 -564 -640
rect 564 -674 660 -640
<< psubdiffcont >>
rect -564 640 564 674
rect -660 -578 -626 578
rect 626 -578 660 578
rect -564 -674 564 -640
<< poly >>
rect -500 572 500 588
rect -500 538 -484 572
rect 484 538 500 572
rect -500 500 500 538
rect -500 -538 500 -500
rect -500 -572 -484 -538
rect 484 -572 500 -538
rect -500 -588 500 -572
<< polycont >>
rect -484 538 484 572
rect -484 -572 484 -538
<< locali >>
rect -660 640 -564 674
rect 564 640 660 674
rect -660 578 -626 640
rect 626 578 660 640
rect -500 538 -484 572
rect 484 538 500 572
rect -546 488 -512 504
rect -546 -504 -512 -488
rect 512 488 546 504
rect 512 -504 546 -488
rect -500 -572 -484 -538
rect 484 -572 500 -538
rect -660 -640 -626 -578
rect 626 -640 660 -578
rect -660 -674 -564 -640
rect 564 -674 660 -640
<< viali >>
rect -501 640 501 674
rect -484 538 484 572
rect -660 -512 -626 512
rect -546 -488 -512 488
rect 512 -488 546 488
rect 626 -512 660 512
rect -484 -572 484 -538
rect -501 -674 501 -640
<< metal1 >>
rect -513 674 513 680
rect -513 640 -501 674
rect 501 640 513 674
rect -513 634 513 640
rect -496 572 496 578
rect -496 538 -484 572
rect 484 538 496 572
rect -496 532 496 538
rect -666 512 -620 524
rect -666 -512 -660 512
rect -626 -512 -620 512
rect 620 512 666 524
rect -552 488 -506 500
rect -552 -488 -546 488
rect -512 -488 -506 488
rect -552 -500 -506 -488
rect 506 488 552 500
rect 506 -488 512 488
rect 546 -488 552 488
rect 506 -500 552 -488
rect -666 -524 -620 -512
rect 620 -512 626 512
rect 660 -512 666 512
rect 620 -524 666 -512
rect -496 -538 496 -532
rect -496 -572 -484 -538
rect 484 -572 496 -538
rect -496 -578 496 -572
rect -513 -640 513 -634
rect -513 -674 -501 -640
rect 501 -674 513 -640
rect -513 -680 513 -674
<< properties >>
string FIXED_BBOX -643 -657 643 657
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 5 l 5 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 80 viagr 80 viagl 80 viagt 80
<< end >>
