magic
tech sky130A
magscale 1 2
timestamp 1713215442
<< error_p >>
rect -111 172 -47 178
rect 47 172 111 178
rect -111 138 -99 172
rect 47 138 59 172
rect -111 132 -47 138
rect 47 132 111 138
rect -111 -138 -47 -132
rect 47 -138 111 -132
rect -111 -172 -99 -138
rect 47 -172 59 -138
rect -111 -178 -47 -172
rect 47 -178 111 -172
<< pwell >>
rect -357 -358 357 358
<< mvnmos >>
rect -129 -100 -29 100
rect 29 -100 129 100
<< mvndiff >>
rect -187 88 -129 100
rect -187 -88 -175 88
rect -141 -88 -129 88
rect -187 -100 -129 -88
rect -29 88 29 100
rect -29 -88 -17 88
rect 17 -88 29 88
rect -29 -100 29 -88
rect 129 88 187 100
rect 129 -88 141 88
rect 175 -88 187 88
rect 129 -100 187 -88
<< mvndiffc >>
rect -175 -88 -141 88
rect -17 -88 17 88
rect 141 -88 175 88
<< mvpsubdiff >>
rect -321 310 321 322
rect -321 276 -213 310
rect 213 276 321 310
rect -321 264 321 276
rect -321 214 -263 264
rect -321 -214 -309 214
rect -275 -214 -263 214
rect 263 214 321 264
rect -321 -264 -263 -214
rect 263 -214 275 214
rect 309 -214 321 214
rect 263 -264 321 -214
rect -321 -276 321 -264
rect -321 -310 -213 -276
rect 213 -310 321 -276
rect -321 -322 321 -310
<< mvpsubdiffcont >>
rect -213 276 213 310
rect -309 -214 -275 214
rect 275 -214 309 214
rect -213 -310 213 -276
<< poly >>
rect -129 172 -29 188
rect -129 138 -113 172
rect -45 138 -29 172
rect -129 100 -29 138
rect 29 172 129 188
rect 29 138 45 172
rect 113 138 129 172
rect 29 100 129 138
rect -129 -138 -29 -100
rect -129 -172 -113 -138
rect -45 -172 -29 -138
rect -129 -188 -29 -172
rect 29 -138 129 -100
rect 29 -172 45 -138
rect 113 -172 129 -138
rect 29 -188 129 -172
<< polycont >>
rect -113 138 -45 172
rect 45 138 113 172
rect -113 -172 -45 -138
rect 45 -172 113 -138
<< locali >>
rect -309 276 -213 310
rect 213 276 309 310
rect -309 221 -275 276
rect 275 214 309 276
rect -129 138 -113 172
rect -45 138 -29 172
rect 29 138 45 172
rect 113 138 129 172
rect -175 88 -141 104
rect -175 -104 -141 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 141 88 175 104
rect 141 -104 175 -88
rect -129 -172 -113 -138
rect -45 -172 -29 -138
rect 29 -172 45 -138
rect 113 -172 129 -138
rect -309 -276 -275 -221
rect 275 -276 309 -214
rect -309 -310 -220 -276
rect 220 -310 309 -276
<< viali >>
rect -309 214 -275 221
rect -309 -214 -275 214
rect -99 138 -59 172
rect 59 138 99 172
rect -175 -88 -141 88
rect -17 -88 17 88
rect 141 -88 175 88
rect -99 -172 -59 -138
rect 59 -172 99 -138
rect -309 -221 -275 -214
rect -220 -310 -213 -276
rect -213 -310 213 -276
rect 213 -310 220 -276
<< metal1 >>
rect -315 221 -269 233
rect -315 -221 -309 221
rect -275 -221 -269 221
rect -111 172 -47 178
rect -111 138 -99 172
rect -59 138 -47 172
rect -111 132 -47 138
rect 47 172 111 178
rect 47 138 59 172
rect 99 138 111 172
rect 47 132 111 138
rect -181 88 -135 100
rect -181 -88 -175 88
rect -141 -88 -135 88
rect -181 -100 -135 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 135 88 181 100
rect 135 -88 141 88
rect 175 -88 181 88
rect 135 -100 181 -88
rect -111 -138 -47 -132
rect -111 -172 -99 -138
rect -59 -172 -47 -138
rect -111 -178 -47 -172
rect 47 -138 111 -132
rect 47 -172 59 -138
rect 99 -172 111 -138
rect 47 -178 111 -172
rect -315 -233 -269 -221
rect -232 -276 232 -270
rect -232 -310 -220 -276
rect 220 -310 232 -276
rect -232 -316 232 -310
<< properties >>
string FIXED_BBOX -292 -293 292 293
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 1 l 0.5 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 60 viagb 80 viagr 0 viagl 80 viagt 0
<< end >>
