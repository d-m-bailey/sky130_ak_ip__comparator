magic
tech sky130A
magscale 1 2
timestamp 1726751280
<< pwell >>
rect -2503 -3844 2503 3844
<< mvpsubdiff >>
rect -2437 3766 2437 3778
rect -2437 3732 -2329 3766
rect 2329 3732 2437 3766
rect -2437 3720 2437 3732
rect -2437 3670 -2379 3720
rect -2437 -3670 -2425 3670
rect -2391 -3670 -2379 3670
rect 2379 3670 2437 3720
rect -2437 -3720 -2379 -3670
rect 2379 -3670 2391 3670
rect 2425 -3670 2437 3670
rect 2379 -3720 2437 -3670
rect -2437 -3732 2437 -3720
rect -2437 -3766 -2329 -3732
rect 2329 -3766 2437 -3732
rect -2437 -3778 2437 -3766
<< mvpsubdiffcont >>
rect -2329 3732 2329 3766
rect -2425 -3670 -2391 3670
rect 2391 -3670 2425 3670
rect -2329 -3766 2329 -3732
<< xpolycontact >>
rect -2283 3192 -1713 3624
rect -2283 -3624 -1713 -3192
rect -1617 3192 -1047 3624
rect -1617 -3624 -1047 -3192
rect -951 3192 -381 3624
rect -951 -3624 -381 -3192
rect -285 3192 285 3624
rect -285 -3624 285 -3192
rect 381 3192 951 3624
rect 381 -3624 951 -3192
rect 1047 3192 1617 3624
rect 1047 -3624 1617 -3192
rect 1713 3192 2283 3624
rect 1713 -3624 2283 -3192
<< ppolyres >>
rect -2283 -3192 -1713 3192
rect -1617 -3192 -1047 3192
rect -951 -3192 -381 3192
rect -285 -3192 285 3192
rect 381 -3192 951 3192
rect 1047 -3192 1617 3192
rect 1713 -3192 2283 3192
<< locali >>
rect -2425 3732 -2329 3766
rect 2329 3732 2425 3766
rect -2425 3670 -2391 3732
rect 2391 3670 2425 3732
rect -2425 -3732 -2391 -3670
rect 2391 -3732 2425 -3670
rect -2425 -3766 -2329 -3732
rect 2329 -3766 2425 -3732
<< viali >>
rect -2152 3732 2152 3766
rect -2425 -3359 -2391 3359
rect -2267 3209 -1729 3606
rect -1601 3209 -1063 3606
rect -935 3209 -397 3606
rect -269 3209 269 3606
rect 397 3209 935 3606
rect 1063 3209 1601 3606
rect 1729 3209 2267 3606
rect -2267 -3606 -1729 -3209
rect -1601 -3606 -1063 -3209
rect -935 -3606 -397 -3209
rect -269 -3606 269 -3209
rect 397 -3606 935 -3209
rect 1063 -3606 1601 -3209
rect 1729 -3606 2267 -3209
rect 2391 -3359 2425 3359
rect -2152 -3766 2152 -3732
<< metal1 >>
rect -2164 3766 2164 3772
rect -2164 3732 -2152 3766
rect 2152 3732 2164 3766
rect -2164 3726 2164 3732
rect -2279 3606 -1717 3612
rect -2431 3359 -2385 3371
rect -2431 -3359 -2425 3359
rect -2391 -3359 -2385 3359
rect -2279 3209 -2267 3606
rect -1729 3209 -1717 3606
rect -2279 3203 -1717 3209
rect -1613 3606 -1051 3612
rect -1613 3209 -1601 3606
rect -1063 3209 -1051 3606
rect -1613 3203 -1051 3209
rect -947 3606 -385 3612
rect -947 3209 -935 3606
rect -397 3209 -385 3606
rect -947 3203 -385 3209
rect -281 3606 281 3612
rect -281 3209 -269 3606
rect 269 3209 281 3606
rect -281 3203 281 3209
rect 385 3606 947 3612
rect 385 3209 397 3606
rect 935 3209 947 3606
rect 385 3203 947 3209
rect 1051 3606 1613 3612
rect 1051 3209 1063 3606
rect 1601 3209 1613 3606
rect 1051 3203 1613 3209
rect 1717 3606 2279 3612
rect 1717 3209 1729 3606
rect 2267 3209 2279 3606
rect 1717 3203 2279 3209
rect 2385 3359 2431 3371
rect -2431 -3371 -2385 -3359
rect -2279 -3209 -1717 -3203
rect -2279 -3606 -2267 -3209
rect -1729 -3606 -1717 -3209
rect -2279 -3612 -1717 -3606
rect -1613 -3209 -1051 -3203
rect -1613 -3606 -1601 -3209
rect -1063 -3606 -1051 -3209
rect -1613 -3612 -1051 -3606
rect -947 -3209 -385 -3203
rect -947 -3606 -935 -3209
rect -397 -3606 -385 -3209
rect -947 -3612 -385 -3606
rect -281 -3209 281 -3203
rect -281 -3606 -269 -3209
rect 269 -3606 281 -3209
rect -281 -3612 281 -3606
rect 385 -3209 947 -3203
rect 385 -3606 397 -3209
rect 935 -3606 947 -3209
rect 385 -3612 947 -3606
rect 1051 -3209 1613 -3203
rect 1051 -3606 1063 -3209
rect 1601 -3606 1613 -3209
rect 1051 -3612 1613 -3606
rect 1717 -3209 2279 -3203
rect 1717 -3606 1729 -3209
rect 2267 -3606 2279 -3209
rect 2385 -3359 2391 3359
rect 2425 -3359 2431 3359
rect 2385 -3371 2431 -3359
rect 1717 -3612 2279 -3606
rect -2164 -3732 2164 -3726
rect -2164 -3766 -2152 -3732
rect 2152 -3766 2164 -3732
rect -2164 -3772 2164 -3766
<< properties >>
string FIXED_BBOX -2408 -3749 2408 3749
string gencell sky130_fd_pr__res_high_po_2p85
string library sky130
string MASKHINTS_HVI -2562 -3833 2492 -3665 -2562 3664 2492 3832
string parameters w 2.85 l 31.92 m 1 nx 7 wmin 2.850 lmin 0.50 rho 319.8 val 3.718k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 2.850 n_guard 0 hv_guard 1 vias 1 viagb 90 viagt 90 viagl 90 viagr 90
<< end >>
