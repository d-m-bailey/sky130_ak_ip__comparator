magic
tech sky130A
magscale 1 2
timestamp 1726591983
<< dnwell >>
rect -1360 11270 30240 13200
rect -1360 9062 34264 11270
rect -1360 -31160 39240 9062
rect -1360 -33200 31650 -31160
<< nwell >>
rect -1440 12994 30320 13280
rect -1440 -32994 -1154 12994
rect 27680 8060 29480 11700
rect 30034 11350 30320 12994
rect 31240 12170 33620 12900
rect 30034 11064 34347 11350
rect 35540 11200 35670 11250
rect 36420 11090 36690 11150
rect 30730 9350 33510 10050
rect 34044 9145 34347 11064
rect 34044 8820 39320 9145
rect 27680 4060 32020 8060
rect -600 -23770 38400 -7600
rect -600 -23800 22060 -23770
rect 27290 -23800 38400 -23770
rect -400 -32400 22060 -23800
rect 31600 -27526 38400 -23800
rect 32796 -29221 38390 -29220
rect 32600 -29960 38390 -29221
rect 39034 -30954 39320 8820
rect 31441 -31240 39320 -30954
rect 31441 -32994 31740 -31240
rect 32638 -32800 38380 -32070
rect -1440 -33280 31740 -32994
<< pwell >>
rect -200 -4910 27100 11990
rect 36920 10710 37020 10880
rect 35530 9720 35660 9780
rect 35554 7670 35850 7750
<< psubdiff >>
rect -1800 13566 -1704 13600
rect 39504 13566 39600 13600
rect -1800 13504 -1766 13566
rect 39566 13504 39600 13566
rect -1800 -33566 -1766 -33504
rect 39566 -33566 39600 -33504
rect -1800 -33600 -1704 -33566
rect 39504 -33600 39600 -33566
<< nsubdiff >>
rect -1403 13223 30283 13243
rect -1403 13189 -1323 13223
rect 30203 13189 30283 13223
rect -1403 13169 30283 13189
rect -1403 13163 -1329 13169
rect -1403 -33163 -1383 13163
rect -1349 -33163 -1329 13163
rect 30209 13163 30283 13169
rect 30209 11319 30229 13163
rect 30263 11319 30283 13163
rect 30209 11313 30283 11319
rect 30209 11293 34310 11313
rect 30209 11259 30289 11293
rect 34230 11259 34310 11293
rect 30209 11239 34310 11259
rect 34236 11233 34310 11239
rect 34236 9084 34256 11233
rect 34290 9084 34310 11233
rect 34236 9078 34310 9084
rect 34236 9058 39283 9078
rect 34236 9024 34316 9058
rect 39203 9024 39283 9058
rect 34236 9004 39283 9024
rect 39209 8998 39283 9004
rect 39209 -31123 39229 8998
rect 39263 -31123 39283 8998
rect 39209 -31129 39283 -31123
rect -1403 -33169 -1329 -33163
rect 31616 -31149 39283 -31129
rect 31616 -31183 31696 -31149
rect 39203 -31183 39283 -31149
rect 31616 -31203 39283 -31183
rect 31616 -31209 31690 -31203
rect 31616 -33163 31636 -31209
rect 31670 -33163 31690 -31209
rect 31616 -33169 31690 -33163
rect -1403 -33189 31690 -33169
rect -1403 -33223 -1323 -33189
rect 31610 -33223 31690 -33189
rect -1403 -33243 31690 -33223
<< psubdiffcont >>
rect -1704 13566 39504 13600
rect -1800 -33504 -1766 13504
rect 39566 -33504 39600 13504
rect -1704 -33600 39504 -33566
<< nsubdiffcont >>
rect -1323 13189 30203 13223
rect -1383 -33163 -1349 13163
rect 30229 11319 30263 13163
rect 30289 11259 34230 11293
rect 34256 9084 34290 11233
rect 34316 9024 39203 9058
rect 39229 -31123 39263 8998
rect 31696 -31183 39203 -31149
rect 31636 -33163 31670 -31209
rect -1323 -33223 31610 -33189
<< locali >>
rect -1900 13600 39700 13700
rect -1900 13566 -1704 13600
rect 39504 13566 39700 13600
rect -1900 13504 39700 13566
rect -1900 -33504 -1800 13504
rect -1766 13500 39566 13504
rect -1766 -33500 -1700 13500
rect -1500 13223 30300 13300
rect -1500 13189 -1323 13223
rect 30203 13189 30300 13223
rect -1500 13163 30300 13189
rect -1500 -33163 -1383 13163
rect -1349 13100 30229 13163
rect -1349 -7400 -1300 13100
rect -300 11920 27280 12100
rect -300 11900 22920 11920
rect -300 11620 60 11900
rect 300 11760 500 11900
rect 960 11760 1160 11900
rect 1620 11760 1820 11900
rect 2060 11620 2260 11900
rect 2500 11760 2700 11900
rect 3160 11760 3360 11900
rect 3820 11760 4020 11900
rect 4260 11620 4460 11900
rect 4700 11760 4900 11900
rect 5360 11760 5560 11900
rect 6020 11760 6220 11900
rect 6460 11620 6660 11900
rect 6900 11760 7100 11900
rect 7560 11760 7760 11900
rect 8220 11760 8420 11900
rect 8660 11620 8860 11900
rect 9100 11760 9300 11900
rect 9760 11760 9960 11900
rect 10420 11760 10620 11900
rect 10860 11620 11060 11900
rect 11300 11760 11500 11900
rect 11960 11760 12160 11900
rect 12620 11760 12820 11900
rect 13060 11620 13260 11900
rect 13500 11760 13700 11900
rect 14160 11760 14360 11900
rect 14820 11760 15020 11900
rect 15260 11620 15460 11900
rect 15700 11760 15900 11900
rect 16360 11760 16560 11900
rect 17020 11760 17220 11900
rect 17460 11620 17660 11900
rect 17900 11760 18100 11900
rect 18560 11760 18760 11900
rect 19220 11760 19420 11900
rect 19660 11620 19860 11900
rect 20100 11760 20300 11900
rect 20760 11760 20960 11900
rect 21420 11760 21620 11900
rect 21860 11620 22920 11900
rect -300 11520 200 11620
rect 1920 11520 2400 11620
rect 4120 11520 4600 11620
rect 6320 11520 6800 11620
rect 8520 11520 9000 11620
rect 10720 11520 11200 11620
rect 12920 11520 13400 11620
rect 15120 11520 15600 11620
rect 17320 11520 17800 11620
rect 19520 11520 20000 11620
rect 21720 11520 22920 11620
rect -300 11260 60 11520
rect 280 11260 480 11400
rect 960 11260 1160 11400
rect 1620 11260 1820 11400
rect 2060 11260 2260 11520
rect 2480 11260 2680 11400
rect 3160 11260 3360 11400
rect 3820 11260 4020 11400
rect 4260 11260 4460 11520
rect 4680 11260 4880 11400
rect 5360 11260 5560 11400
rect 6020 11260 6220 11400
rect 6460 11260 6660 11520
rect 6880 11260 7080 11400
rect 7560 11260 7760 11400
rect 8220 11260 8420 11400
rect 8660 11260 8860 11520
rect 9080 11260 9280 11400
rect 9760 11260 9960 11400
rect 10420 11260 10620 11400
rect 10860 11260 11060 11520
rect 11280 11260 11480 11400
rect 11960 11260 12160 11400
rect 12620 11260 12820 11400
rect 13060 11260 13260 11520
rect 13480 11260 13680 11400
rect 14160 11260 14360 11400
rect 14820 11260 15020 11400
rect 15260 11260 15460 11520
rect 15680 11260 15880 11400
rect 16360 11260 16560 11400
rect 17020 11260 17220 11400
rect 17460 11260 17660 11520
rect 17880 11260 18080 11400
rect 18560 11260 18760 11400
rect 19220 11260 19420 11400
rect 19660 11260 19860 11520
rect 21860 11400 22920 11520
rect 26380 11400 27280 11920
rect 20080 11260 20280 11400
rect 20760 11260 20960 11400
rect 21420 11260 21620 11400
rect 21860 11260 22260 11400
rect -300 11100 22260 11260
rect -300 10930 60 11100
rect 300 10960 500 11100
rect 960 10960 1160 11100
rect 1620 10960 1820 11100
rect -300 10870 -70 10930
rect -10 10870 60 10930
rect -300 10820 60 10870
rect 2060 10930 2260 11100
rect 2060 10870 2130 10930
rect 2190 10870 2260 10930
rect 2060 10820 2260 10870
rect -300 10720 200 10820
rect 1920 10720 2260 10820
rect -300 10460 60 10720
rect 280 10460 480 10600
rect 960 10460 1160 10600
rect 1620 10460 1820 10600
rect 2060 10460 2260 10720
rect 4260 10930 4460 11100
rect 4260 10870 4330 10930
rect 4390 10870 4460 10930
rect 4260 10460 4460 10870
rect 6460 10930 6660 11100
rect 6460 10870 6530 10930
rect 6590 10870 6660 10930
rect 6460 10460 6660 10870
rect 8660 10930 8860 11100
rect 8660 10870 8730 10930
rect 8790 10870 8860 10930
rect 8660 10460 8860 10870
rect 10860 10930 11060 11100
rect 10860 10870 10930 10930
rect 10990 10870 11060 10930
rect 10860 10460 11060 10870
rect 13060 10930 13260 11100
rect 13060 10870 13130 10930
rect 13190 10870 13260 10930
rect 13060 10460 13260 10870
rect 15260 10930 15460 11100
rect 15260 10870 15330 10930
rect 15390 10870 15460 10930
rect 15260 10460 15460 10870
rect 17460 10930 17660 11100
rect 17460 10870 17530 10930
rect 17590 10870 17660 10930
rect 17460 10460 17660 10870
rect 19660 10930 19860 11100
rect 20100 10960 20300 11100
rect 20760 10960 20960 11100
rect 21420 10960 21620 11100
rect 19660 10870 19730 10930
rect 19790 10870 19860 10930
rect 19660 10820 19860 10870
rect 21860 10930 22260 11100
rect 21860 10870 21930 10930
rect 21990 10870 22260 10930
rect 21860 10820 22260 10870
rect 19660 10720 20000 10820
rect 21720 10720 22260 10820
rect 19660 10460 19860 10720
rect 20080 10460 20280 10600
rect 20760 10460 20960 10600
rect 21420 10460 21620 10600
rect 21860 10460 22260 10720
rect -300 10300 22260 10460
rect -300 10130 60 10300
rect 300 10160 500 10300
rect 960 10160 1160 10300
rect 1620 10160 1820 10300
rect -300 10070 -70 10130
rect -10 10070 60 10130
rect -300 10020 60 10070
rect 2060 10130 2260 10300
rect 2060 10070 2130 10130
rect 2190 10070 2260 10130
rect 2060 10020 2260 10070
rect -300 9920 200 10020
rect 1920 9920 2260 10020
rect -300 9660 60 9920
rect 280 9660 480 9800
rect 960 9660 1160 9800
rect 1620 9660 1820 9800
rect 2060 9660 2260 9920
rect 4260 10130 4460 10300
rect 4260 10070 4330 10130
rect 4390 10070 4460 10130
rect 4260 9660 4460 10070
rect 6460 10130 6660 10300
rect 6460 10070 6530 10130
rect 6590 10070 6660 10130
rect 6460 9660 6660 10070
rect 8660 10130 8860 10300
rect 8660 10070 8730 10130
rect 8790 10070 8860 10130
rect 8660 9660 8860 10070
rect 10860 10130 11060 10300
rect 10860 10070 10930 10130
rect 10990 10070 11060 10130
rect 10860 9660 11060 10070
rect 13060 10130 13260 10300
rect 13060 10070 13130 10130
rect 13190 10070 13260 10130
rect 13060 9660 13260 10070
rect 15260 10130 15460 10300
rect 15260 10070 15330 10130
rect 15390 10070 15460 10130
rect 15260 9660 15460 10070
rect 17460 10130 17660 10300
rect 17460 10070 17530 10130
rect 17590 10070 17660 10130
rect 17460 9660 17660 10070
rect 19660 10130 19860 10300
rect 20100 10160 20300 10300
rect 20760 10160 20960 10300
rect 21420 10160 21620 10300
rect 19660 10070 19730 10130
rect 19790 10070 19860 10130
rect 19660 10020 19860 10070
rect 21860 10130 22260 10300
rect 21860 10070 21930 10130
rect 21990 10070 22260 10130
rect 21860 10020 22260 10070
rect 19660 9920 20000 10020
rect 21720 9920 22260 10020
rect 19660 9660 19860 9920
rect 20080 9660 20280 9800
rect 20760 9660 20960 9800
rect 21420 9660 21620 9800
rect 21860 9660 22260 9920
rect -300 9500 22260 9660
rect -300 9330 60 9500
rect 300 9360 500 9500
rect 960 9360 1160 9500
rect 1620 9360 1820 9500
rect -300 9270 -70 9330
rect -10 9270 60 9330
rect -300 9220 60 9270
rect 2060 9330 2260 9500
rect 2060 9270 2130 9330
rect 2190 9270 2260 9330
rect 2060 9220 2260 9270
rect -300 9120 200 9220
rect 1920 9120 2260 9220
rect -300 8860 60 9120
rect 280 8860 480 9000
rect 960 8860 1160 9000
rect 1620 8860 1820 9000
rect 2060 8860 2260 9120
rect 4260 9330 4460 9500
rect 4260 9270 4330 9330
rect 4390 9270 4460 9330
rect 4260 8860 4460 9270
rect 6460 9330 6660 9500
rect 6460 9270 6530 9330
rect 6590 9270 6660 9330
rect 6460 8860 6660 9270
rect 8660 9330 8860 9500
rect 8660 9270 8730 9330
rect 8790 9270 8860 9330
rect 8660 8860 8860 9270
rect 10860 9330 11060 9500
rect 10860 9270 10930 9330
rect 10990 9270 11060 9330
rect 10860 8860 11060 9270
rect 13060 9330 13260 9500
rect 13060 9270 13130 9330
rect 13190 9270 13260 9330
rect 13060 8860 13260 9270
rect 15260 9330 15460 9500
rect 15260 9270 15330 9330
rect 15390 9270 15460 9330
rect 15260 8860 15460 9270
rect 17460 9330 17660 9500
rect 17460 9270 17530 9330
rect 17590 9270 17660 9330
rect 17460 8860 17660 9270
rect 19660 9330 19860 9500
rect 20100 9360 20300 9500
rect 20760 9360 20960 9500
rect 21420 9360 21620 9500
rect 19660 9270 19730 9330
rect 19790 9270 19860 9330
rect 19660 9220 19860 9270
rect 21860 9330 22260 9500
rect 21860 9270 21930 9330
rect 21990 9270 22260 9330
rect 21860 9220 22260 9270
rect 19660 9120 20000 9220
rect 21720 9120 22260 9220
rect 19660 8860 19860 9120
rect 20080 8860 20280 9000
rect 20760 8860 20960 9000
rect 21420 8860 21620 9000
rect 21860 8860 22260 9120
rect -300 8700 22260 8860
rect -300 8530 60 8700
rect 300 8560 500 8700
rect 960 8560 1160 8700
rect 1620 8560 1820 8700
rect -300 8470 -70 8530
rect -10 8470 60 8530
rect -300 8420 60 8470
rect 2060 8530 2260 8700
rect 2060 8470 2130 8530
rect 2190 8470 2260 8530
rect 2060 8420 2260 8470
rect -300 8320 200 8420
rect 1920 8320 2260 8420
rect -300 8060 60 8320
rect 280 8060 480 8200
rect 960 8060 1160 8200
rect 1620 8060 1820 8200
rect 2060 8060 2260 8320
rect 4260 8530 4460 8700
rect 4260 8470 4330 8530
rect 4390 8470 4460 8530
rect 4260 8060 4460 8470
rect 6460 8530 6660 8700
rect 6460 8470 6530 8530
rect 6590 8470 6660 8530
rect 6460 8060 6660 8470
rect 8660 8530 8860 8700
rect 8660 8470 8730 8530
rect 8790 8470 8860 8530
rect 8660 8060 8860 8470
rect 10860 8530 11060 8700
rect 10860 8470 10930 8530
rect 10990 8470 11060 8530
rect 10860 8060 11060 8470
rect 13060 8530 13260 8700
rect 13060 8470 13130 8530
rect 13190 8470 13260 8530
rect 13060 8060 13260 8470
rect 15260 8530 15460 8700
rect 15260 8470 15330 8530
rect 15390 8470 15460 8530
rect 15260 8060 15460 8470
rect 17460 8530 17660 8700
rect 17460 8470 17530 8530
rect 17590 8470 17660 8530
rect 17460 8060 17660 8470
rect 19660 8530 19860 8700
rect 20100 8560 20300 8700
rect 20760 8560 20960 8700
rect 21420 8560 21620 8700
rect 19660 8470 19730 8530
rect 19790 8470 19860 8530
rect 19660 8420 19860 8470
rect 21860 8530 22260 8700
rect 21860 8470 21930 8530
rect 21990 8470 22260 8530
rect 21860 8420 22260 8470
rect 19660 8320 20000 8420
rect 21720 8320 22260 8420
rect 19660 8060 19860 8320
rect 20080 8060 20280 8200
rect 20760 8060 20960 8200
rect 21420 8060 21620 8200
rect 21860 8060 22260 8320
rect -300 7900 22260 8060
rect -300 7730 60 7900
rect 300 7760 500 7900
rect 960 7760 1160 7900
rect 1620 7760 1820 7900
rect -300 7670 -70 7730
rect -10 7670 60 7730
rect -300 7620 60 7670
rect 2060 7730 2260 7900
rect 2060 7670 2130 7730
rect 2190 7670 2260 7730
rect 2060 7620 2260 7670
rect -300 7520 200 7620
rect 1920 7520 2260 7620
rect -300 7260 60 7520
rect 280 7260 480 7400
rect 960 7260 1160 7400
rect 1620 7260 1820 7400
rect 2060 7260 2260 7520
rect 4260 7730 4460 7900
rect 4260 7670 4330 7730
rect 4390 7670 4460 7730
rect 4260 7260 4460 7670
rect 6460 7730 6660 7900
rect 6460 7670 6530 7730
rect 6590 7670 6660 7730
rect 6460 7260 6660 7670
rect 8660 7730 8860 7900
rect 8660 7670 8730 7730
rect 8790 7670 8860 7730
rect 8660 7260 8860 7670
rect 10860 7730 11060 7900
rect 10860 7670 10930 7730
rect 10990 7670 11060 7730
rect 10860 7260 11060 7670
rect 13060 7730 13260 7900
rect 13060 7670 13130 7730
rect 13190 7670 13260 7730
rect 13060 7260 13260 7670
rect 15260 7730 15460 7900
rect 15260 7670 15330 7730
rect 15390 7670 15460 7730
rect 15260 7260 15460 7670
rect 17460 7730 17660 7900
rect 17460 7670 17530 7730
rect 17590 7670 17660 7730
rect 17460 7260 17660 7670
rect 19660 7730 19860 7900
rect 20100 7760 20300 7900
rect 20760 7760 20960 7900
rect 21420 7760 21620 7900
rect 19660 7670 19730 7730
rect 19790 7670 19860 7730
rect 19660 7620 19860 7670
rect 21860 7730 22260 7900
rect 21860 7670 21930 7730
rect 21990 7670 22260 7730
rect 21860 7620 22260 7670
rect 19660 7520 20000 7620
rect 21720 7520 22260 7620
rect 19660 7260 19860 7520
rect 20080 7260 20280 7400
rect 20760 7260 20960 7400
rect 21420 7260 21620 7400
rect 21860 7260 22260 7520
rect -300 7100 22260 7260
rect -300 6930 60 7100
rect 300 6960 500 7100
rect 960 6960 1160 7100
rect 1620 6960 1820 7100
rect -300 6870 -70 6930
rect -10 6870 60 6930
rect -300 6820 60 6870
rect 2060 6930 2260 7100
rect 2060 6870 2130 6930
rect 2190 6870 2260 6930
rect 2060 6820 2260 6870
rect -300 6720 200 6820
rect 1920 6720 2260 6820
rect -300 6460 60 6720
rect 280 6460 480 6600
rect 960 6460 1160 6600
rect 1620 6460 1820 6600
rect 2060 6460 2260 6720
rect 4260 6930 4460 7100
rect 4260 6870 4330 6930
rect 4390 6870 4460 6930
rect 4260 6460 4460 6870
rect 6460 6930 6660 7100
rect 6460 6870 6530 6930
rect 6590 6870 6660 6930
rect 6460 6460 6660 6870
rect 8660 6930 8860 7100
rect 8660 6870 8730 6930
rect 8790 6870 8860 6930
rect 8660 6460 8860 6870
rect 10860 6930 11060 7100
rect 10860 6870 10930 6930
rect 10990 6870 11060 6930
rect 10860 6460 11060 6870
rect 13060 6930 13260 7100
rect 13060 6870 13130 6930
rect 13190 6870 13260 6930
rect 13060 6460 13260 6870
rect 15260 6930 15460 7100
rect 15260 6870 15330 6930
rect 15390 6870 15460 6930
rect 15260 6460 15460 6870
rect 17460 6930 17660 7100
rect 17460 6870 17530 6930
rect 17590 6870 17660 6930
rect 17460 6460 17660 6870
rect 19660 6930 19860 7100
rect 20100 6960 20300 7100
rect 20760 6960 20960 7100
rect 21420 6960 21620 7100
rect 19660 6870 19730 6930
rect 19790 6870 19860 6930
rect 19660 6820 19860 6870
rect 21860 6930 22260 7100
rect 21860 6870 21930 6930
rect 21990 6870 22260 6930
rect 21860 6820 22260 6870
rect 19660 6720 20000 6820
rect 21720 6720 22260 6820
rect 19660 6460 19860 6720
rect 20080 6460 20280 6600
rect 20760 6460 20960 6600
rect 21420 6460 21620 6600
rect 21860 6460 22260 6720
rect -300 6300 22260 6460
rect -300 6130 60 6300
rect 300 6160 500 6300
rect 960 6160 1160 6300
rect 1620 6160 1820 6300
rect -300 6070 -70 6130
rect -10 6070 60 6130
rect -300 6020 60 6070
rect 2060 6130 2260 6300
rect 2060 6070 2130 6130
rect 2190 6070 2260 6130
rect 2060 6020 2260 6070
rect -300 5920 200 6020
rect 1920 5920 2260 6020
rect -300 5660 60 5920
rect 280 5660 480 5800
rect 960 5660 1160 5800
rect 1620 5660 1820 5800
rect 2060 5660 2260 5920
rect 4260 6130 4460 6300
rect 4260 6070 4330 6130
rect 4390 6070 4460 6130
rect 4260 5660 4460 6070
rect 6460 6130 6660 6300
rect 6460 6070 6530 6130
rect 6590 6070 6660 6130
rect 6460 5660 6660 6070
rect 8660 6130 8860 6300
rect 8660 6070 8730 6130
rect 8790 6070 8860 6130
rect 8660 5660 8860 6070
rect 10860 6130 11060 6300
rect 10860 6070 10930 6130
rect 10990 6070 11060 6130
rect 10860 5660 11060 6070
rect 13060 6130 13260 6300
rect 13060 6070 13130 6130
rect 13190 6070 13260 6130
rect 13060 5660 13260 6070
rect 15260 6130 15460 6300
rect 15260 6070 15330 6130
rect 15390 6070 15460 6130
rect 15260 5660 15460 6070
rect 17460 6130 17660 6300
rect 17460 6070 17530 6130
rect 17590 6070 17660 6130
rect 17460 5660 17660 6070
rect 19660 6130 19860 6300
rect 20100 6160 20300 6300
rect 20760 6160 20960 6300
rect 21420 6160 21620 6300
rect 19660 6070 19730 6130
rect 19790 6070 19860 6130
rect 19660 6020 19860 6070
rect 21860 6130 22260 6300
rect 21860 6070 21930 6130
rect 21990 6070 22260 6130
rect 21860 6020 22260 6070
rect 19660 5920 20000 6020
rect 21720 5920 22260 6020
rect 19660 5660 19860 5920
rect 20080 5660 20280 5800
rect 20760 5660 20960 5800
rect 21420 5660 21620 5800
rect 21860 5660 22260 5920
rect -300 5500 22260 5660
rect -300 5330 60 5500
rect 300 5360 500 5500
rect 960 5360 1160 5500
rect 1620 5360 1820 5500
rect -300 5270 -70 5330
rect -10 5270 60 5330
rect -300 5220 60 5270
rect 2060 5330 2260 5500
rect 2060 5270 2130 5330
rect 2190 5270 2260 5330
rect 2060 5220 2260 5270
rect -300 5120 200 5220
rect 1920 5120 2260 5220
rect -300 4860 60 5120
rect 280 4860 480 5000
rect 960 4860 1160 5000
rect 1620 4860 1820 5000
rect 2060 4860 2260 5120
rect 4260 5330 4460 5500
rect 4260 5270 4330 5330
rect 4390 5270 4460 5330
rect 4260 4860 4460 5270
rect 6460 5330 6660 5500
rect 6460 5270 6530 5330
rect 6590 5270 6660 5330
rect 6460 4860 6660 5270
rect 8660 5330 8860 5500
rect 8660 5270 8730 5330
rect 8790 5270 8860 5330
rect 8660 4860 8860 5270
rect 10860 5330 11060 5500
rect 10860 5270 10930 5330
rect 10990 5270 11060 5330
rect 10860 4970 11060 5270
rect 13060 5330 13260 5500
rect 13060 5270 13130 5330
rect 13190 5270 13260 5330
rect 10850 4860 11070 4970
rect 13060 4860 13260 5270
rect 15260 5330 15460 5500
rect 15260 5270 15330 5330
rect 15390 5270 15460 5330
rect 15260 4860 15460 5270
rect 17460 5330 17660 5500
rect 17460 5270 17530 5330
rect 17590 5270 17660 5330
rect 17460 4860 17660 5270
rect 19660 5330 19860 5500
rect 20100 5360 20300 5500
rect 20760 5360 20960 5500
rect 21420 5360 21620 5500
rect 19660 5270 19730 5330
rect 19790 5270 19860 5330
rect 19660 5220 19860 5270
rect 21860 5330 22260 5500
rect 21860 5270 21930 5330
rect 21990 5270 22260 5330
rect 21860 5220 22260 5270
rect 19660 5120 20000 5220
rect 21720 5120 22260 5220
rect 19660 4860 19860 5120
rect 20080 4860 20280 5000
rect 20760 4860 20960 5000
rect 21420 4860 21620 5000
rect 21860 4980 22260 5120
rect 27040 4980 27280 11400
rect 21860 4860 22920 4980
rect -300 4700 22920 4860
rect -300 4420 60 4700
rect 300 4560 500 4700
rect 960 4560 1160 4700
rect 1620 4560 1820 4700
rect 2060 4420 2260 4700
rect 2500 4560 2700 4700
rect 3160 4560 3360 4700
rect 3820 4560 4020 4700
rect 4260 4420 4460 4700
rect 4700 4560 4900 4700
rect 5360 4560 5560 4700
rect 6020 4560 6220 4700
rect 6460 4420 6660 4700
rect 6900 4560 7100 4700
rect 7560 4560 7760 4700
rect 8220 4560 8420 4700
rect 8660 4420 8860 4700
rect -300 4320 200 4420
rect 1920 4320 2400 4420
rect 4120 4320 4600 4420
rect 6320 4320 6800 4420
rect 8520 4320 8860 4420
rect -300 4060 60 4320
rect 280 4060 480 4200
rect 960 4060 1160 4200
rect 1620 4060 1820 4200
rect 2060 4060 2260 4320
rect 2480 4060 2680 4200
rect 3160 4060 3360 4200
rect 3820 4060 4020 4200
rect 4260 4060 4460 4320
rect 4680 4060 4880 4200
rect 5360 4060 5560 4200
rect 6020 4060 6220 4200
rect 6460 4060 6660 4320
rect 6880 4060 7080 4200
rect 7560 4060 7760 4200
rect 8220 4060 8420 4200
rect 8660 4060 8860 4320
rect 10850 4060 11070 4700
rect 13060 4420 13260 4700
rect 13500 4560 13700 4700
rect 14160 4560 14360 4700
rect 14820 4560 15020 4700
rect 15260 4420 15460 4700
rect 15700 4560 15900 4700
rect 16360 4560 16560 4700
rect 17020 4560 17220 4700
rect 17460 4420 17660 4700
rect 17900 4560 18100 4700
rect 18560 4560 18760 4700
rect 19220 4560 19420 4700
rect 19660 4420 19860 4700
rect 20100 4560 20300 4700
rect 20760 4560 20960 4700
rect 21420 4560 21620 4700
rect 21860 4460 22920 4700
rect 26380 4460 27280 4980
rect 21860 4420 27280 4460
rect 13060 4320 13400 4420
rect 15120 4320 15600 4420
rect 17320 4320 17800 4420
rect 19520 4320 20000 4420
rect 21720 4320 27280 4420
rect 13060 4060 13260 4320
rect 13480 4060 13680 4200
rect 14160 4060 14360 4200
rect 14820 4060 15020 4200
rect 15260 4060 15460 4320
rect 15680 4060 15880 4200
rect 16360 4060 16560 4200
rect 17020 4060 17220 4200
rect 17460 4060 17660 4320
rect 17880 4060 18080 4200
rect 18560 4060 18760 4200
rect 19220 4060 19420 4200
rect 19660 4060 19860 4320
rect 20080 4060 20280 4200
rect 20760 4060 20960 4200
rect 21420 4060 21620 4200
rect 21860 4060 27280 4320
rect 28910 11120 29150 11570
rect 30100 11319 30229 13100
rect 30263 11370 30300 13163
rect 30263 11319 34327 11370
rect 30100 11308 34327 11319
rect 30100 11293 30330 11308
rect 34142 11293 34327 11308
rect 30100 11259 30289 11293
rect 34230 11259 34327 11293
rect 30100 11256 30330 11259
rect 34142 11256 34327 11259
rect 30100 11233 34327 11256
rect 30100 11170 34256 11233
rect 30100 11169 30420 11170
rect 28910 7220 29460 11120
rect 34127 9200 34256 11170
rect 34126 9084 34256 9200
rect 34290 9135 34327 11233
rect 36426 9326 36546 9986
rect 34290 9084 39300 9135
rect 34126 9058 39300 9084
rect 34126 9024 34316 9058
rect 39203 9024 39300 9058
rect 34126 8998 39300 9024
rect 34126 8935 39229 8998
rect 36426 8092 36546 8628
rect 35238 7958 37732 8092
rect 35380 7470 35706 7958
rect 36426 7470 36566 7958
rect 37288 7470 37600 7958
rect 28910 4110 29150 7220
rect 35380 7176 37600 7470
rect 35380 6982 36128 7176
rect 36810 6982 37600 7176
rect 35380 6440 37600 6982
rect 35380 6120 38400 6440
rect 35380 4330 36240 6120
rect 35340 4310 36240 4330
rect 32040 4160 36240 4310
rect 32040 4152 32600 4160
rect -300 3640 27280 4060
rect 32040 3640 32606 4152
rect -300 3500 32606 3640
rect -300 2430 16970 3500
rect 17880 3358 32606 3500
rect 32846 3364 33184 3374
rect 34138 3364 34796 4160
rect 35540 4120 36240 4160
rect 35544 3780 36240 4120
rect 37840 3780 38400 6120
rect 35544 3366 38400 3780
rect 35434 3364 38400 3366
rect 32846 3358 33878 3364
rect 17880 3352 33878 3358
rect 34138 3352 38400 3364
rect 17880 3220 38400 3352
rect 17880 3210 33878 3220
rect 17880 2446 32284 3210
rect 32846 2446 33878 3210
rect 17880 2434 33878 2446
rect 34426 2440 35464 3220
rect 36060 2440 38400 3220
rect 34426 2434 38400 2440
rect 17880 2430 38400 2434
rect -300 2220 38400 2430
rect -300 2210 36660 2220
rect -300 2200 1470 2210
rect -300 1120 0 2200
rect 180 2080 340 2200
rect 180 1120 340 1220
rect 520 1120 620 2200
rect 800 2080 960 2200
rect 800 1120 960 1220
rect 1140 1120 1470 2200
rect -300 1020 1470 1120
rect -300 540 0 1020
rect 180 940 340 1020
rect 180 540 340 680
rect 520 540 620 1020
rect 800 940 960 1020
rect 1140 920 1470 1020
rect 1140 900 1460 920
rect 800 540 960 680
rect 1140 550 1470 900
rect 2860 550 3070 2210
rect 4460 550 4670 2210
rect 6060 550 6270 2210
rect 7660 550 7870 2210
rect 9260 550 9470 2210
rect 10860 550 11070 2210
rect 12460 550 12670 2210
rect 14060 550 14270 2210
rect 15660 550 15870 2210
rect 17260 550 17470 2210
rect 18860 550 19070 2210
rect 20460 550 20670 2210
rect 22060 550 22270 2210
rect 23660 550 23870 2210
rect 25260 550 25470 2210
rect 26860 550 27070 2210
rect 28460 550 28670 2210
rect 30060 550 30270 2210
rect 31660 550 31870 2210
rect 33260 550 33470 2210
rect 34860 550 35070 2210
rect 36460 550 36660 2210
rect 1140 540 36660 550
rect 38060 540 38400 2220
rect -300 420 38400 540
rect -300 -680 0 420
rect 180 280 340 420
rect 180 -680 340 -580
rect 520 -680 620 420
rect 800 280 960 420
rect 1140 410 36800 420
rect 800 -680 960 -580
rect 1140 -680 1470 410
rect -300 -780 1470 -680
rect -300 -1260 0 -780
rect 180 -860 340 -780
rect 180 -1260 340 -1120
rect 520 -1260 620 -780
rect 800 -860 960 -780
rect 1140 -880 1470 -780
rect 1140 -900 1460 -880
rect 800 -1260 960 -1120
rect 1140 -1250 1470 -900
rect 2860 -1250 3070 410
rect 4460 -1250 4670 410
rect 6060 -1250 6270 410
rect 7660 -1250 7870 410
rect 9260 -1250 9470 410
rect 10860 -1250 11070 410
rect 12460 -1250 12670 410
rect 14060 -1250 14270 410
rect 15660 -1250 15870 410
rect 17260 -1250 17470 410
rect 18860 -1250 19070 410
rect 20460 -1250 20670 410
rect 22060 -1250 22270 410
rect 23660 -1250 23870 410
rect 25260 -1250 25470 410
rect 26860 -1250 27070 410
rect 28460 -1250 28670 410
rect 30060 -1250 30270 410
rect 31660 -1250 31870 410
rect 33260 -1250 33470 410
rect 34860 -1250 35070 410
rect 36460 249 36800 410
rect 36855 261 36871 295
rect 36980 280 37140 420
rect 37247 261 37263 295
rect 37320 249 37420 420
rect 37473 261 37489 295
rect 37600 280 37760 420
rect 37865 261 37881 295
rect 37940 249 38400 420
rect 36460 233 36821 249
rect 37297 233 37439 249
rect 37915 233 38400 249
rect 36460 -535 36800 233
rect 37320 -535 37420 233
rect 37940 -535 38400 233
rect 36460 -551 36821 -535
rect 37297 -551 37439 -535
rect 37915 -551 38400 -535
rect 36460 -680 36800 -551
rect 36855 -597 36871 -563
rect 36980 -680 37140 -580
rect 37247 -597 37263 -563
rect 37320 -680 37420 -551
rect 37473 -597 37489 -563
rect 37600 -680 37760 -580
rect 37865 -597 37881 -563
rect 37940 -680 38400 -551
rect 36460 -780 38400 -680
rect 36460 -897 36800 -780
rect 36855 -885 36871 -851
rect 36980 -860 37140 -780
rect 37247 -885 37263 -851
rect 37320 -897 37420 -780
rect 37473 -885 37489 -851
rect 37600 -860 37760 -780
rect 37865 -885 37881 -851
rect 37940 -897 38400 -780
rect 36460 -913 36821 -897
rect 37297 -913 37439 -897
rect 37915 -913 38400 -897
rect 36460 -1081 36800 -913
rect 37320 -1081 37420 -913
rect 37940 -1081 38400 -913
rect 36460 -1097 36821 -1081
rect 37297 -1097 37439 -1081
rect 37915 -1097 38400 -1081
rect 36460 -1243 36800 -1097
rect 36855 -1143 36871 -1109
rect 36980 -1243 37140 -1120
rect 37247 -1143 37263 -1109
rect 37320 -1243 37420 -1097
rect 37473 -1143 37489 -1109
rect 37600 -1243 37760 -1120
rect 37865 -1143 37881 -1109
rect 37940 -1243 38400 -1097
rect 36460 -1250 38400 -1243
rect 1140 -1260 38400 -1250
rect -300 -1380 38400 -1260
rect -300 -2480 0 -1380
rect 180 -1520 340 -1380
rect 180 -2480 340 -2380
rect 520 -2480 620 -1380
rect 800 -1520 960 -1380
rect 1140 -1390 36800 -1380
rect 800 -2480 960 -2380
rect 1140 -2480 1470 -1390
rect -300 -2580 1470 -2480
rect -300 -3060 0 -2580
rect 180 -2660 340 -2580
rect 180 -3060 340 -2920
rect 520 -3060 620 -2580
rect 800 -2660 960 -2580
rect 1140 -2680 1470 -2580
rect 1140 -2700 1460 -2680
rect 800 -3060 960 -2920
rect 1140 -3050 1470 -2700
rect 2860 -3050 3070 -1390
rect 4460 -3050 4670 -1390
rect 6060 -3050 6270 -1390
rect 7660 -3050 7870 -1390
rect 9260 -3050 9470 -1390
rect 10860 -3050 11070 -1390
rect 12460 -3050 12670 -1390
rect 14060 -3050 14270 -1390
rect 15660 -3050 15870 -1390
rect 17260 -3050 17470 -1390
rect 18860 -3050 19070 -1390
rect 20460 -3050 20670 -1390
rect 22060 -3050 22270 -1390
rect 23660 -3050 23870 -1390
rect 25260 -3050 25470 -1390
rect 26860 -3050 27070 -1390
rect 28460 -3050 28670 -1390
rect 30060 -3050 30270 -1390
rect 31660 -3050 31870 -1390
rect 33260 -3050 33470 -1390
rect 34860 -3050 35070 -1390
rect 36460 -1551 36800 -1390
rect 36855 -1539 36871 -1505
rect 36980 -1520 37140 -1380
rect 37247 -1539 37263 -1505
rect 37320 -1551 37420 -1380
rect 37473 -1539 37489 -1505
rect 37600 -1520 37760 -1380
rect 37865 -1539 37881 -1505
rect 37940 -1551 38400 -1380
rect 36460 -1567 36821 -1551
rect 37297 -1567 37439 -1551
rect 37915 -1567 38400 -1551
rect 36460 -2335 36800 -1567
rect 37320 -2335 37420 -1567
rect 37940 -2335 38400 -1567
rect 36460 -2351 36821 -2335
rect 37297 -2351 37439 -2335
rect 37915 -2351 38400 -2335
rect 36460 -2480 36800 -2351
rect 36855 -2397 36871 -2363
rect 36980 -2480 37140 -2380
rect 37247 -2397 37263 -2363
rect 37320 -2480 37420 -2351
rect 37473 -2397 37489 -2363
rect 37600 -2480 37760 -2380
rect 37865 -2397 37881 -2363
rect 37940 -2480 38400 -2351
rect 36460 -2580 38400 -2480
rect 36460 -2697 36800 -2580
rect 36855 -2685 36871 -2651
rect 36980 -2660 37140 -2580
rect 37247 -2685 37263 -2651
rect 37320 -2697 37420 -2580
rect 37473 -2685 37489 -2651
rect 37600 -2660 37760 -2580
rect 37865 -2685 37881 -2651
rect 37940 -2697 38400 -2580
rect 36460 -2713 36821 -2697
rect 37297 -2713 37439 -2697
rect 37915 -2713 38400 -2697
rect 36460 -2881 36800 -2713
rect 37320 -2881 37420 -2713
rect 37940 -2881 38400 -2713
rect 36460 -2897 36821 -2881
rect 37297 -2897 37439 -2881
rect 37915 -2897 38400 -2881
rect 36460 -3043 36800 -2897
rect 36855 -2943 36871 -2909
rect 36980 -3043 37140 -2920
rect 37247 -2943 37263 -2909
rect 37320 -3043 37420 -2897
rect 37473 -2943 37489 -2909
rect 37600 -3043 37760 -2920
rect 37865 -2943 37881 -2909
rect 37940 -3043 38400 -2897
rect 36460 -3050 38400 -3043
rect 1140 -3060 38400 -3050
rect -300 -3180 38400 -3060
rect -300 -4280 0 -3180
rect 180 -3320 340 -3180
rect 180 -4280 340 -4180
rect 520 -4280 620 -3180
rect 800 -3320 960 -3180
rect 1140 -3190 36800 -3180
rect 800 -4280 960 -4180
rect 1140 -4280 1470 -3190
rect -300 -4380 1470 -4280
rect -300 -4860 0 -4380
rect 180 -4460 340 -4380
rect 180 -4860 340 -4720
rect 520 -4860 620 -4380
rect 800 -4460 960 -4380
rect 1140 -4460 1470 -4380
rect 1140 -4480 1460 -4460
rect 800 -4860 960 -4720
rect 1140 -4850 1470 -4480
rect 2860 -4850 3070 -3190
rect 4460 -4850 4670 -3190
rect 6060 -4850 6270 -3190
rect 7660 -4850 7870 -3190
rect 9260 -4850 9470 -3190
rect 10860 -4850 11070 -3190
rect 12460 -4850 12670 -3190
rect 14060 -4850 14270 -3190
rect 15660 -4850 15870 -3190
rect 17260 -4850 17470 -3190
rect 18860 -4850 19070 -3190
rect 20460 -4850 20670 -3190
rect 22060 -4850 22270 -3190
rect 23660 -4850 23870 -3190
rect 25260 -4850 25470 -3190
rect 26860 -4850 27070 -3190
rect 28460 -4850 28670 -3190
rect 30060 -4850 30270 -3190
rect 31660 -4850 31870 -3190
rect 33260 -4850 33470 -3190
rect 34860 -4850 35070 -3190
rect 36460 -3351 36800 -3190
rect 36855 -3339 36871 -3305
rect 36980 -3320 37140 -3180
rect 37247 -3339 37263 -3305
rect 37320 -3351 37420 -3180
rect 37473 -3339 37489 -3305
rect 37600 -3320 37760 -3180
rect 37865 -3339 37881 -3305
rect 37940 -3351 38400 -3180
rect 36460 -3367 36821 -3351
rect 37297 -3367 37439 -3351
rect 37915 -3367 38400 -3351
rect 36460 -4135 36800 -3367
rect 37320 -4135 37420 -3367
rect 37940 -4135 38400 -3367
rect 36460 -4151 36821 -4135
rect 37297 -4151 37439 -4135
rect 37915 -4151 38400 -4135
rect 36460 -4280 36800 -4151
rect 36855 -4197 36871 -4163
rect 36980 -4280 37140 -4180
rect 37247 -4197 37263 -4163
rect 37320 -4280 37420 -4151
rect 37473 -4197 37489 -4163
rect 37600 -4280 37760 -4180
rect 37865 -4197 37881 -4163
rect 37940 -4280 38400 -4151
rect 36460 -4380 38400 -4280
rect 36460 -4497 36800 -4380
rect 36855 -4485 36871 -4451
rect 36980 -4460 37140 -4380
rect 37247 -4485 37263 -4451
rect 37320 -4497 37420 -4380
rect 37473 -4485 37489 -4451
rect 37600 -4460 37760 -4380
rect 37865 -4485 37881 -4451
rect 37940 -4497 38400 -4380
rect 36460 -4513 36821 -4497
rect 37297 -4513 37439 -4497
rect 37915 -4513 38400 -4497
rect 36460 -4681 36800 -4513
rect 37320 -4681 37420 -4513
rect 37940 -4681 38400 -4513
rect 36460 -4697 36821 -4681
rect 37297 -4697 37439 -4681
rect 37915 -4697 38400 -4681
rect 36460 -4843 36800 -4697
rect 36855 -4743 36871 -4709
rect 36980 -4843 37140 -4720
rect 37247 -4743 37263 -4709
rect 37320 -4843 37420 -4697
rect 37473 -4743 37489 -4709
rect 37600 -4843 37760 -4720
rect 37865 -4743 37881 -4709
rect 37940 -4843 38400 -4697
rect 36460 -4850 38400 -4843
rect 1140 -4860 38400 -4850
rect -300 -5600 38400 -4860
rect 39100 -7400 39229 8935
rect -1349 -8060 39229 -7400
rect -1349 -9700 1460 -8060
rect 2900 -9700 3060 -8060
rect 4500 -9700 4660 -8060
rect 6100 -9700 6260 -8060
rect 7700 -9700 7860 -8060
rect 9300 -9700 9460 -8060
rect 10900 -9700 11060 -8060
rect 12500 -9700 12660 -8060
rect 14100 -9700 14260 -8060
rect 15700 -9700 15860 -8060
rect 17300 -9700 17460 -8060
rect 18900 -9700 19060 -8060
rect 20500 -9700 20660 -8060
rect 22100 -9700 22260 -8060
rect 23700 -9700 23860 -8060
rect 25300 -9700 25460 -8060
rect 26900 -9700 27060 -8060
rect 28500 -9700 28660 -8060
rect 30100 -9700 30260 -8060
rect 31700 -9700 31860 -8060
rect 33300 -9700 33460 -8060
rect 34900 -9700 35060 -8060
rect 36500 -9700 39229 -8060
rect -1349 -9860 39229 -9700
rect -1349 -11500 1460 -9860
rect 2900 -11500 3060 -9860
rect 4500 -11500 4660 -9860
rect 6100 -11500 6260 -9860
rect 7700 -11500 7860 -9860
rect 9300 -11500 9460 -9860
rect 10900 -11500 11060 -9860
rect 12500 -11500 12660 -9860
rect 14100 -11500 14260 -9860
rect 15700 -11500 15860 -9860
rect 17300 -11500 17460 -9860
rect 18900 -11500 19060 -9860
rect 20500 -11500 20660 -9860
rect 22100 -11500 22260 -9860
rect 23700 -11500 23860 -9860
rect 25300 -11500 25460 -9860
rect 26900 -11500 27060 -9860
rect 28500 -11500 28660 -9860
rect 30100 -11500 30260 -9860
rect 31700 -11500 31860 -9860
rect 33300 -11500 33460 -9860
rect 34900 -11500 35060 -9860
rect 36500 -11500 39229 -9860
rect -1349 -11660 39229 -11500
rect -1349 -13300 1460 -11660
rect 2900 -13300 3060 -11660
rect 4500 -13300 4660 -11660
rect 6100 -13300 6260 -11660
rect 7700 -13300 7860 -11660
rect 9300 -13300 9460 -11660
rect 10900 -13300 11060 -11660
rect 12500 -13300 12660 -11660
rect 14100 -13300 14260 -11660
rect 15700 -13300 15860 -11660
rect 17300 -13300 17460 -11660
rect 18900 -13300 19060 -11660
rect 20500 -13300 20660 -11660
rect 22100 -13300 22260 -11660
rect 23700 -13300 23860 -11660
rect 25300 -13300 25460 -11660
rect 26900 -13300 27060 -11660
rect 28500 -13300 28660 -11660
rect 30100 -13300 30260 -11660
rect 31700 -13300 31860 -11660
rect 33300 -13300 33460 -11660
rect 34900 -13300 35060 -11660
rect 36500 -13300 39229 -11660
rect -1349 -13460 39229 -13300
rect -1349 -15100 1460 -13460
rect 2900 -15100 3060 -13460
rect 4500 -15100 4660 -13460
rect 6100 -15100 6260 -13460
rect 7700 -15100 7860 -13460
rect 9300 -15100 9460 -13460
rect 10900 -15100 11060 -13460
rect 12500 -15100 12660 -13460
rect 14100 -15100 14260 -13460
rect 15700 -15100 15860 -13460
rect 17300 -15100 17460 -13460
rect 18900 -15100 19060 -13460
rect 20500 -15100 20660 -13460
rect 22100 -15100 22260 -13460
rect 23700 -15100 23860 -13460
rect 25300 -15100 25460 -13460
rect 26900 -15100 27060 -13460
rect 28500 -15100 28660 -13460
rect 30100 -15100 30260 -13460
rect 31700 -15100 31860 -13460
rect 33300 -15100 33460 -13460
rect 34900 -15100 35060 -13460
rect 36500 -15100 39229 -13460
rect -1349 -15260 39229 -15100
rect -1349 -16900 1460 -15260
rect 2900 -16900 3060 -15260
rect 4500 -16900 4660 -15260
rect 6100 -16900 6260 -15260
rect 7700 -16900 7860 -15260
rect 9300 -16900 9460 -15260
rect 10900 -16900 11060 -15260
rect 12500 -16900 12660 -15260
rect 14100 -16900 14260 -15260
rect 15700 -16900 15860 -15260
rect 17300 -16900 17460 -15260
rect 18900 -16900 19060 -15260
rect 20500 -16900 20660 -15260
rect 22100 -16900 22260 -15260
rect 23700 -16900 23860 -15260
rect 25300 -16900 25460 -15260
rect 26900 -16900 27060 -15260
rect 28500 -16900 28660 -15260
rect 30100 -16900 30260 -15260
rect 31700 -16900 31860 -15260
rect 33300 -16900 33460 -15260
rect 34900 -16900 35060 -15260
rect 36500 -16900 39229 -15260
rect -1349 -17060 39229 -16900
rect -1349 -18700 1460 -17060
rect 2900 -18700 3060 -17060
rect 4500 -18700 4660 -17060
rect 6100 -18700 6260 -17060
rect 7700 -18700 7860 -17060
rect 9300 -18700 9460 -17060
rect 10900 -18700 11060 -17060
rect 12500 -18700 12660 -17060
rect 14100 -18700 14260 -17060
rect 15700 -18700 15860 -17060
rect 17300 -18700 17460 -17060
rect 18900 -18700 19060 -17060
rect 20500 -18700 20660 -17060
rect 22100 -18700 22260 -17060
rect 23700 -18700 23860 -17060
rect 25300 -18700 25460 -17060
rect 26900 -18700 27060 -17060
rect 28500 -18700 28660 -17060
rect 30100 -18700 30260 -17060
rect 31700 -18700 31860 -17060
rect 33300 -18700 33460 -17060
rect 34900 -18700 35060 -17060
rect 36500 -18700 39229 -17060
rect -1349 -18860 39229 -18700
rect -1349 -20500 1460 -18860
rect 2900 -20500 3060 -18860
rect 4500 -20500 4660 -18860
rect 6100 -20500 6260 -18860
rect 7700 -20500 7860 -18860
rect 9300 -20500 9460 -18860
rect 10900 -20500 11060 -18860
rect 12500 -20500 12660 -18860
rect 14100 -20500 14260 -18860
rect 15700 -20500 15860 -18860
rect 17300 -20500 17460 -18860
rect 18900 -20500 19060 -18860
rect 20500 -20500 20660 -18860
rect 22100 -20500 22260 -18860
rect 23700 -20500 23860 -18860
rect 25300 -20500 25460 -18860
rect 26900 -20500 27060 -18860
rect 28500 -20500 28660 -18860
rect 30100 -20500 30260 -18860
rect 31700 -20500 31860 -18860
rect 33300 -20500 33460 -18860
rect 34900 -20500 35060 -18860
rect 36500 -20500 39229 -18860
rect -1349 -20660 39229 -20500
rect -1349 -22300 1460 -20660
rect 2900 -22300 3060 -20660
rect 4500 -22280 4660 -20660
rect 6100 -22280 6260 -20660
rect 7700 -22280 7860 -20660
rect 9300 -22280 9460 -20660
rect 10900 -22280 11060 -20660
rect 12500 -22280 12660 -20660
rect 14100 -22280 14260 -20660
rect 15700 -22280 15860 -20660
rect 17300 -22280 17460 -20660
rect 18900 -22280 19060 -20660
rect 20500 -22280 20660 -20660
rect 22100 -22280 22260 -20660
rect 3300 -22300 22260 -22280
rect 23700 -22300 23860 -20660
rect 25300 -22300 25460 -20660
rect 26900 -22300 27060 -20660
rect 28500 -22300 28660 -20660
rect 30100 -22300 30260 -20660
rect 31700 -22300 31860 -20660
rect 33300 -22300 33460 -20660
rect 34900 -22300 35060 -20660
rect 36500 -22300 39229 -20660
rect -1349 -22430 39229 -22300
rect -1349 -22540 32520 -22430
rect -1349 -23660 28240 -22540
rect 29140 -23240 32520 -22540
rect 33410 -23240 33880 -22430
rect 34040 -22440 39229 -22430
rect 34480 -23240 39229 -22440
rect 29140 -23560 39229 -23240
rect 29140 -23660 33060 -23560
rect -1349 -23890 33060 -23660
rect -1349 -24980 21950 -23890
rect 27460 -23900 33060 -23890
rect -1349 -25620 2260 -24980
rect 4240 -25620 4460 -24980
rect 6440 -25620 6660 -24980
rect 8640 -25620 8860 -24980
rect 10840 -25620 11060 -24980
rect 13040 -25620 13260 -24980
rect 15240 -25620 15460 -24980
rect 17440 -25620 17660 -24980
rect 19640 -25620 21950 -24980
rect -1349 -25780 21950 -25620
rect -1349 -26420 2260 -25780
rect 4240 -26420 4460 -25780
rect 6440 -26420 6660 -25780
rect 8640 -26420 8860 -25780
rect 10840 -26420 11060 -25780
rect 13040 -26420 13260 -25780
rect 15240 -26420 15460 -25780
rect 17440 -26420 17660 -25780
rect 19640 -26420 21950 -25780
rect -1349 -26580 21950 -26420
rect -1349 -27220 2260 -26580
rect 4240 -27220 4460 -26580
rect 6440 -27220 6660 -26580
rect 8640 -27220 8860 -26580
rect 10840 -27220 11060 -26580
rect 13040 -27220 13260 -26580
rect 15240 -27220 15460 -26580
rect 17440 -27220 17660 -26580
rect 19640 -27220 21950 -26580
rect -1349 -27380 21950 -27220
rect -1349 -28020 2260 -27380
rect 4240 -28020 4460 -27380
rect 6440 -28020 6660 -27380
rect 8640 -28020 8860 -27380
rect 10840 -28020 11060 -27380
rect 13040 -28020 13260 -27380
rect 15240 -28020 15460 -27380
rect 17440 -28020 17660 -27380
rect 19640 -28020 21950 -27380
rect -1349 -28180 21950 -28020
rect -1349 -28820 2260 -28180
rect 4240 -28820 4460 -28180
rect 6440 -28820 6660 -28180
rect 8640 -28820 8860 -28180
rect 10840 -28820 11060 -28180
rect 13040 -28820 13260 -28180
rect 15240 -28820 15460 -28180
rect 17440 -28820 17660 -28180
rect 19640 -28820 21950 -28180
rect -1349 -28980 21950 -28820
rect -1349 -29620 2260 -28980
rect 4240 -29620 4460 -28980
rect 6440 -29620 6660 -28980
rect 8640 -29620 8860 -28980
rect 10840 -29620 11060 -28980
rect 13040 -29620 13260 -28980
rect 15240 -29620 15460 -28980
rect 17440 -29620 17660 -28980
rect 19640 -29620 21950 -28980
rect -1349 -29780 21950 -29620
rect -1349 -30420 2260 -29780
rect 4240 -30420 4460 -29780
rect 6440 -30420 6660 -29780
rect 8640 -30420 8860 -29780
rect 10840 -30420 11060 -29780
rect 13040 -30420 13260 -29780
rect 15240 -30420 15460 -29780
rect 17440 -30420 17660 -29780
rect 19640 -30420 21950 -29780
rect -1349 -30580 21950 -30420
rect -1349 -31220 2260 -30580
rect 4240 -31220 4460 -30580
rect 6440 -31220 6660 -30580
rect 8640 -31220 8860 -30580
rect 10840 -31220 11060 -30580
rect 13040 -31220 13260 -30580
rect 15240 -31220 15460 -30580
rect 17440 -31220 17660 -30580
rect 19640 -31220 21950 -30580
rect -1349 -32410 21950 -31220
rect 22110 -24300 27700 -24130
rect 22110 -24520 29820 -24300
rect 22110 -24600 27800 -24520
rect 22110 -25060 22900 -24600
rect 22110 -31500 22220 -25060
rect 26360 -25080 27800 -24600
rect 27020 -25300 27800 -25080
rect 28920 -25300 29820 -24520
rect 27020 -25420 29820 -25300
rect 27020 -26340 27800 -25420
rect 28774 -25604 28808 -25588
rect 28774 -25688 28808 -25672
rect 28774 -25762 28808 -25746
rect 28774 -25846 28808 -25830
rect 28774 -25920 28808 -25904
rect 28774 -26004 28808 -25988
rect 28774 -26078 28808 -26062
rect 28774 -26162 28808 -26146
rect 28920 -26340 29820 -25420
rect 27020 -26460 29820 -26340
rect 27020 -27360 27800 -26460
rect 28920 -27360 29820 -26460
rect 27020 -27500 29820 -27360
rect 27020 -28400 27800 -27500
rect 28920 -28400 29820 -27500
rect 31500 -24360 33060 -23900
rect 31500 -24380 33040 -24360
rect 34260 -24380 34440 -23560
rect 37220 -24340 39229 -23560
rect 34720 -24380 39229 -24340
rect 31500 -24700 39229 -24380
rect 31500 -24900 34780 -24700
rect 31500 -27060 34760 -24900
rect 35980 -27060 36120 -24700
rect 37320 -27060 39229 -24700
rect 31500 -27526 39229 -27060
rect 27020 -28540 29820 -28400
rect 27020 -29440 27800 -28540
rect 28920 -29440 29820 -28540
rect 27020 -29580 29820 -29440
rect 27020 -30480 27800 -29580
rect 28920 -30480 29820 -29580
rect 27020 -30620 29820 -30480
rect 27020 -31500 27800 -30620
rect 22110 -32000 22900 -31500
rect 26360 -31520 27800 -31500
rect 28920 -31520 29820 -30620
rect 39140 -31060 39229 -27526
rect 26360 -31660 29820 -31520
rect 31560 -31123 39229 -31060
rect 39263 -31123 39300 8998
rect 31560 -31142 39300 -31123
rect 31560 -31149 31742 -31142
rect 39152 -31149 39300 -31142
rect 31560 -31183 31696 -31149
rect 39203 -31183 39300 -31149
rect 31560 -31206 31742 -31183
rect 39152 -31206 39300 -31183
rect 31560 -31209 39300 -31206
rect 26360 -32000 27700 -31660
rect 22110 -32260 27700 -32000
rect -1349 -32500 22030 -32410
rect -1349 -33100 27100 -32500
rect 31560 -33100 31636 -31209
rect -1349 -33163 31636 -33100
rect 31670 -31260 39300 -31209
rect 31670 -33163 31760 -31260
rect -1500 -33189 31760 -33163
rect -1500 -33223 -1323 -33189
rect 31610 -33223 31760 -33189
rect -1500 -33300 31760 -33223
rect 39500 -33500 39566 13500
rect -1766 -33504 39566 -33500
rect 39600 -33504 39700 13504
rect -1900 -33566 39700 -33504
rect -1900 -33600 -1704 -33566
rect 39504 -33600 39700 -33566
rect -1900 -33700 39700 -33600
<< viali >>
rect -1704 13566 39504 13600
rect -1800 -33504 -1766 13504
rect -1283 13189 30163 13223
rect -1383 -33123 -1349 13123
rect -70 10870 -10 10930
rect 2130 10870 2190 10930
rect 4330 10870 4390 10930
rect 6530 10870 6590 10930
rect 8730 10870 8790 10930
rect 10930 10870 10990 10930
rect 13130 10870 13190 10930
rect 15330 10870 15390 10930
rect 17530 10870 17590 10930
rect 19730 10870 19790 10930
rect 21930 10870 21990 10930
rect -70 10070 -10 10130
rect 2130 10070 2190 10130
rect 4330 10070 4390 10130
rect 6530 10070 6590 10130
rect 8730 10070 8790 10130
rect 10930 10070 10990 10130
rect 13130 10070 13190 10130
rect 15330 10070 15390 10130
rect 17530 10070 17590 10130
rect 19730 10070 19790 10130
rect 21930 10070 21990 10130
rect -70 9270 -10 9330
rect 2130 9270 2190 9330
rect 4330 9270 4390 9330
rect 6530 9270 6590 9330
rect 8730 9270 8790 9330
rect 10930 9270 10990 9330
rect 13130 9270 13190 9330
rect 15330 9270 15390 9330
rect 17530 9270 17590 9330
rect 19730 9270 19790 9330
rect 21930 9270 21990 9330
rect -70 8470 -10 8530
rect 2130 8470 2190 8530
rect 4330 8470 4390 8530
rect 6530 8470 6590 8530
rect 8730 8470 8790 8530
rect 10930 8470 10990 8530
rect 13130 8470 13190 8530
rect 15330 8470 15390 8530
rect 17530 8470 17590 8530
rect 19730 8470 19790 8530
rect 21930 8470 21990 8530
rect -70 7670 -10 7730
rect 2130 7670 2190 7730
rect 4330 7670 4390 7730
rect 6530 7670 6590 7730
rect 8730 7670 8790 7730
rect 10930 7670 10990 7730
rect 13130 7670 13190 7730
rect 15330 7670 15390 7730
rect 17530 7670 17590 7730
rect 19730 7670 19790 7730
rect 21930 7670 21990 7730
rect -70 6870 -10 6930
rect 2130 6870 2190 6930
rect 4330 6870 4390 6930
rect 6530 6870 6590 6930
rect 8730 6870 8790 6930
rect 10930 6870 10990 6930
rect 13130 6870 13190 6930
rect 15330 6870 15390 6930
rect 17530 6870 17590 6930
rect 19730 6870 19790 6930
rect 21930 6870 21990 6930
rect -70 6070 -10 6130
rect 2130 6070 2190 6130
rect 4330 6070 4390 6130
rect 6530 6070 6590 6130
rect 8730 6070 8790 6130
rect 10930 6070 10990 6130
rect 13130 6070 13190 6130
rect 15330 6070 15390 6130
rect 17530 6070 17590 6130
rect 19730 6070 19790 6130
rect 21930 6070 21990 6130
rect -70 5270 -10 5330
rect 2130 5270 2190 5330
rect 4330 5270 4390 5330
rect 6530 5270 6590 5330
rect 8730 5270 8790 5330
rect 10930 5270 10990 5330
rect 13130 5270 13190 5330
rect 15330 5270 15390 5330
rect 17530 5270 17590 5330
rect 19730 5270 19790 5330
rect 21930 5270 21990 5330
rect 30229 11359 30263 13123
rect 30330 11293 34142 11308
rect 30330 11259 34142 11293
rect 30330 11256 34142 11259
rect 34256 9124 34290 11193
rect 34352 9024 39163 9058
rect 36128 6982 36810 7176
rect 39229 -31083 39263 8958
rect 31742 -31149 39152 -31142
rect 31742 -31183 39152 -31149
rect 31742 -31206 39152 -31183
rect 31636 -33123 31670 -31249
rect -1283 -33223 31570 -33189
rect 39566 -33504 39600 13504
rect -1704 -33600 39504 -33566
<< metal1 >>
rect -1900 13600 39700 13700
rect -1900 13566 -1704 13600
rect 39504 13566 39700 13600
rect -1900 13504 39700 13566
rect -1900 -33504 -1800 13504
rect -1766 13500 39566 13504
rect -1766 -33500 -1700 13500
rect -1500 13223 30300 13300
rect -1500 13189 -1283 13223
rect 30163 13189 30300 13223
rect -1500 13123 30300 13189
rect -1500 -33123 -1383 13123
rect -1349 13100 30229 13123
rect -1349 -9600 -1300 13100
rect 23050 11400 24240 11790
rect 24380 11400 25590 11790
rect 25710 11780 26250 11790
rect 25710 11410 25720 11780
rect 26240 11410 26250 11780
rect 29280 11660 29500 13100
rect 27920 11560 29500 11660
rect 25710 11400 26250 11410
rect 27250 11490 27330 11500
rect 27250 11400 27260 11490
rect 27320 11464 27330 11490
rect 27320 11418 27950 11464
rect 27320 11400 27330 11418
rect 27250 11390 27330 11400
rect 27730 11330 27810 11340
rect 27730 11306 27740 11330
rect 27260 11260 27740 11306
rect 27730 11240 27740 11260
rect 27800 11306 27810 11330
rect 27800 11260 27950 11306
rect 27800 11240 27810 11260
rect 2500 11180 2510 11240
rect 2690 11180 2700 11240
rect 2500 10940 2700 11180
rect 3160 11180 3170 11240
rect 3350 11180 3360 11240
rect 3160 10940 3360 11180
rect 3820 11180 3830 11240
rect 4010 11180 4020 11240
rect 3820 10940 4020 11180
rect 4700 11180 4710 11240
rect 4890 11180 4900 11240
rect 4700 10940 4900 11180
rect 5360 11180 5370 11240
rect 5550 11180 5560 11240
rect 5360 10940 5560 11180
rect 6020 11180 6030 11240
rect 6210 11180 6220 11240
rect 6020 10940 6220 11180
rect 6900 11100 7100 11240
rect 6900 11040 6910 11100
rect 7090 11040 7100 11100
rect 6900 10940 7100 11040
rect 7560 11100 7760 11240
rect 7560 11040 7570 11100
rect 7750 11040 7760 11100
rect 7560 10940 7760 11040
rect 8220 11100 8420 11240
rect 8220 11040 8230 11100
rect 8410 11040 8420 11100
rect 8220 10940 8420 11040
rect 9100 11100 9300 11240
rect 9100 11040 9110 11100
rect 9290 11040 9300 11100
rect 9100 10940 9300 11040
rect 9760 11100 9960 11240
rect 9760 11040 9770 11100
rect 9950 11040 9960 11100
rect 9760 10940 9960 11040
rect 10420 11100 10620 11240
rect 10420 11040 10430 11100
rect 10610 11040 10620 11100
rect 10420 10940 10620 11040
rect 11300 11100 11500 11240
rect 11300 11040 11310 11100
rect 11490 11040 11500 11100
rect 11300 10940 11500 11040
rect 11960 11100 12160 11240
rect 11960 11040 11970 11100
rect 12150 11040 12160 11100
rect 11960 10940 12160 11040
rect 12620 11100 12820 11240
rect 12620 11040 12630 11100
rect 12810 11040 12820 11100
rect 12620 10940 12820 11040
rect 13500 11100 13700 11240
rect 13500 11040 13510 11100
rect 13690 11040 13700 11100
rect 13500 10940 13700 11040
rect 14160 11100 14360 11240
rect 14160 11040 14170 11100
rect 14350 11040 14360 11100
rect 14160 10940 14360 11040
rect 14820 11100 15020 11240
rect 14820 11040 14830 11100
rect 15010 11040 15020 11100
rect 14820 10940 15020 11040
rect 15700 11180 15710 11240
rect 15890 11180 15900 11240
rect 15700 10940 15900 11180
rect 16360 11180 16370 11240
rect 16550 11180 16560 11240
rect 16360 10940 16560 11180
rect 17020 11180 17030 11240
rect 17210 11180 17220 11240
rect 17020 10940 17220 11180
rect 17900 11180 17910 11240
rect 18090 11180 18100 11240
rect 17900 10940 18100 11180
rect 18560 11180 18570 11240
rect 18750 11180 18760 11240
rect 18560 10940 18760 11180
rect 19220 11180 19230 11240
rect 19410 11180 19420 11240
rect 27730 11230 27810 11240
rect 28770 11180 28820 11400
rect 29260 11280 29340 11290
rect 29260 11180 29270 11280
rect 19220 10940 19420 11180
rect 27250 11170 27330 11180
rect 27250 11080 27260 11170
rect 27320 11148 27330 11170
rect 27320 11102 27950 11148
rect 27320 11080 27330 11102
rect 27250 11070 27330 11080
rect 28770 11100 29270 11180
rect 27730 11015 27810 11025
rect 27730 10990 27740 11015
rect 27260 10944 27740 10990
rect -90 10930 10 10940
rect -90 10870 -70 10930
rect -10 10870 10 10930
rect -90 10860 10 10870
rect 2110 10930 2210 10940
rect 2110 10870 2130 10930
rect 2190 10870 2210 10930
rect 2110 10860 2210 10870
rect 4310 10930 4410 10940
rect 4310 10870 4330 10930
rect 4390 10870 4410 10930
rect 4310 10860 4410 10870
rect 6510 10930 6610 10940
rect 6510 10870 6530 10930
rect 6590 10870 6610 10930
rect 6510 10860 6610 10870
rect 8710 10930 8810 10940
rect 8710 10870 8730 10930
rect 8790 10870 8810 10930
rect 8710 10860 8810 10870
rect 10910 10930 11010 10940
rect 10910 10870 10930 10930
rect 10990 10870 11010 10930
rect 10910 10860 11010 10870
rect 13110 10930 13210 10940
rect 13110 10870 13130 10930
rect 13190 10870 13210 10930
rect 13110 10860 13210 10870
rect 15310 10930 15410 10940
rect 15310 10870 15330 10930
rect 15390 10870 15410 10930
rect 15310 10860 15410 10870
rect 17510 10930 17610 10940
rect 17510 10870 17530 10930
rect 17590 10870 17610 10930
rect 17510 10860 17610 10870
rect 19710 10930 19810 10940
rect 19710 10870 19730 10930
rect 19790 10870 19810 10930
rect 19710 10860 19810 10870
rect 21910 10930 22010 10940
rect 21910 10870 21930 10930
rect 21990 10870 22010 10930
rect 27730 10925 27740 10944
rect 27800 10990 27810 11015
rect 27800 10944 27950 10990
rect 27800 10925 27810 10944
rect 27730 10915 27810 10925
rect 21910 10860 22010 10870
rect 27250 10855 27330 10865
rect 4100 10760 4220 10820
rect 4280 10760 4510 10820
rect 6300 10760 6420 10820
rect 6480 10760 6710 10820
rect 8500 10760 8840 10820
rect 8900 10760 8910 10820
rect 10700 10760 11040 10820
rect 11100 10760 11110 10820
rect 12900 10760 13240 10820
rect 13300 10760 13310 10820
rect 15100 10760 15440 10820
rect 15500 10760 15510 10820
rect 17300 10760 17420 10820
rect 17480 10760 17710 10820
rect 19500 10740 19620 10800
rect 19680 10740 19910 10800
rect 27250 10765 27260 10855
rect 27320 10832 27330 10855
rect 28770 10850 28820 11100
rect 29260 11060 29270 11100
rect 29330 11060 29340 11280
rect 29260 11050 29340 11060
rect 27320 10786 27950 10832
rect 27320 10765 27330 10786
rect 27250 10755 27330 10765
rect 2010 10650 2020 10710
rect 2080 10650 2420 10710
rect 4210 10650 4220 10710
rect 4280 10650 4620 10710
rect 6410 10650 6640 10710
rect 6700 10650 6820 10710
rect 8610 10650 8840 10710
rect 8900 10650 9020 10710
rect 10810 10650 11040 10710
rect 11100 10650 11220 10710
rect 13010 10650 13240 10710
rect 13300 10650 13420 10710
rect 15210 10650 15220 10710
rect 15280 10650 15620 10710
rect 17410 10650 17420 10710
rect 17480 10650 17820 10710
rect 29400 10680 29500 11560
rect 2500 10610 4020 10620
rect 2500 10550 2510 10610
rect 4010 10550 4020 10610
rect 2500 10540 4020 10550
rect 4700 10610 6220 10622
rect 4700 10550 4710 10610
rect 6210 10550 6220 10610
rect 4700 10540 6220 10550
rect 6900 10610 8420 10622
rect 6900 10550 6910 10610
rect 8410 10550 8420 10610
rect 6900 10540 8420 10550
rect 9100 10610 10620 10622
rect 9100 10550 9110 10610
rect 10610 10550 10620 10610
rect 9100 10540 10620 10550
rect 11300 10610 12820 10622
rect 11300 10550 11310 10610
rect 12810 10550 12820 10610
rect 11300 10540 12820 10550
rect 13500 10610 15020 10622
rect 13500 10550 13510 10610
rect 15010 10550 15020 10610
rect 13500 10540 15020 10550
rect 15700 10610 17220 10622
rect 15700 10550 15710 10610
rect 17210 10550 17220 10610
rect 15700 10540 17220 10550
rect 17900 10610 19420 10622
rect 17900 10550 17910 10610
rect 19410 10550 19420 10610
rect 17900 10540 19420 10550
rect 27920 10520 29500 10680
rect 27730 10450 27810 10460
rect 2500 10300 2700 10440
rect 2500 10240 2510 10300
rect 2690 10240 2700 10300
rect 2500 10140 2700 10240
rect 3160 10300 3360 10440
rect 3160 10240 3170 10300
rect 3350 10240 3360 10300
rect 3160 10140 3360 10240
rect 3820 10300 4020 10440
rect 3820 10240 3830 10300
rect 4010 10240 4020 10300
rect 3820 10140 4020 10240
rect 4700 10300 4900 10440
rect 4700 10240 4710 10300
rect 4890 10240 4900 10300
rect 4700 10140 4900 10240
rect 5360 10300 5560 10440
rect 5360 10240 5370 10300
rect 5550 10240 5560 10300
rect 5360 10140 5560 10240
rect 6020 10300 6220 10440
rect 6020 10240 6030 10300
rect 6210 10240 6220 10300
rect 6020 10140 6220 10240
rect 6900 10380 6910 10440
rect 7090 10380 7100 10440
rect 6900 10140 7100 10380
rect 7560 10380 7570 10440
rect 7750 10380 7760 10440
rect 7560 10140 7760 10380
rect 8220 10380 8230 10440
rect 8410 10380 8420 10440
rect 8220 10140 8420 10380
rect 9100 10380 9110 10440
rect 9290 10380 9300 10440
rect 9100 10140 9300 10380
rect 9760 10380 9770 10440
rect 9950 10380 9960 10440
rect 9760 10140 9960 10380
rect 10420 10380 10430 10440
rect 10610 10380 10620 10440
rect 10420 10140 10620 10380
rect 11300 10380 11310 10440
rect 11490 10380 11500 10440
rect 11300 10140 11500 10380
rect 11960 10380 11970 10440
rect 12150 10380 12160 10440
rect 11960 10140 12160 10380
rect 12620 10380 12630 10440
rect 12810 10380 12820 10440
rect 12620 10140 12820 10380
rect 13500 10380 13510 10440
rect 13690 10380 13700 10440
rect 13500 10140 13700 10380
rect 14160 10380 14170 10440
rect 14350 10380 14360 10440
rect 14160 10140 14360 10380
rect 14820 10380 14830 10440
rect 15010 10380 15020 10440
rect 14820 10140 15020 10380
rect 15700 10300 15900 10440
rect 15700 10240 15710 10300
rect 15890 10240 15900 10300
rect 15700 10140 15900 10240
rect 16360 10300 16560 10440
rect 16360 10240 16370 10300
rect 16550 10240 16560 10300
rect 16360 10140 16560 10240
rect 17020 10300 17220 10440
rect 17020 10240 17030 10300
rect 17210 10240 17220 10300
rect 17020 10140 17220 10240
rect 17900 10300 18100 10440
rect 17900 10240 17910 10300
rect 18090 10240 18100 10300
rect 17900 10140 18100 10240
rect 18560 10300 18760 10440
rect 18560 10240 18570 10300
rect 18750 10240 18760 10300
rect 18560 10140 18760 10240
rect 19220 10300 19420 10440
rect 27730 10424 27740 10450
rect 27260 10378 27740 10424
rect 27730 10360 27740 10378
rect 27800 10424 27810 10450
rect 27800 10378 27950 10424
rect 27800 10360 27810 10378
rect 27730 10350 27810 10360
rect 19220 10240 19230 10300
rect 19410 10240 19420 10300
rect 27370 10290 27450 10300
rect 27370 10266 27380 10290
rect 19220 10140 19420 10240
rect 27260 10220 27380 10266
rect 27370 10200 27380 10220
rect 27440 10266 27450 10290
rect 27440 10220 27950 10266
rect 27440 10200 27450 10220
rect 27370 10190 27450 10200
rect -90 10130 10 10140
rect -90 10070 -70 10130
rect -10 10070 10 10130
rect -90 10060 10 10070
rect 2110 10130 2210 10140
rect 2110 10070 2130 10130
rect 2190 10070 2210 10130
rect 2110 10060 2210 10070
rect 4310 10130 4410 10140
rect 4310 10070 4330 10130
rect 4390 10070 4410 10130
rect 4310 10060 4410 10070
rect 6510 10130 6610 10140
rect 6510 10070 6530 10130
rect 6590 10070 6610 10130
rect 6510 10060 6610 10070
rect 8710 10130 8810 10140
rect 8710 10070 8730 10130
rect 8790 10070 8810 10130
rect 8710 10060 8810 10070
rect 10910 10130 11010 10140
rect 10910 10070 10930 10130
rect 10990 10070 11010 10130
rect 10910 10060 11010 10070
rect 13110 10130 13210 10140
rect 13110 10070 13130 10130
rect 13190 10070 13210 10130
rect 13110 10060 13210 10070
rect 15310 10130 15410 10140
rect 15310 10070 15330 10130
rect 15390 10070 15410 10130
rect 15310 10060 15410 10070
rect 17510 10130 17610 10140
rect 17510 10070 17530 10130
rect 17590 10070 17610 10130
rect 17510 10060 17610 10070
rect 19710 10130 19810 10140
rect 19710 10070 19730 10130
rect 19790 10070 19810 10130
rect 19710 10060 19810 10070
rect 21910 10130 22010 10140
rect 21910 10070 21930 10130
rect 21990 10070 22010 10130
rect 27730 10130 27810 10140
rect 27730 10108 27740 10130
rect 21910 10060 22010 10070
rect 27260 10062 27740 10108
rect 27730 10040 27740 10062
rect 27800 10108 27810 10130
rect 28770 10120 28820 10360
rect 29130 10190 29210 10200
rect 29130 10120 29140 10190
rect 27800 10062 27950 10108
rect 27800 10040 27810 10062
rect 27730 10030 27810 10040
rect 28770 10040 29140 10120
rect 4100 9960 4440 10020
rect 4500 9960 4510 10020
rect 6300 9960 6640 10020
rect 6700 9960 6710 10020
rect 8500 9960 8620 10020
rect 8680 9960 8910 10020
rect 10700 9960 10820 10020
rect 10880 9960 11110 10020
rect 12900 9960 13020 10020
rect 13080 9960 13310 10020
rect 15100 9960 15220 10020
rect 15280 9960 15510 10020
rect 17300 9960 17640 10020
rect 17700 9960 17710 10020
rect 19500 9940 19840 10000
rect 19900 9940 19910 10000
rect 27370 9975 27450 9985
rect 27370 9950 27380 9975
rect 2010 9850 2240 9910
rect 2300 9850 2420 9910
rect 4210 9850 4440 9910
rect 4500 9850 4620 9910
rect 6410 9850 6420 9910
rect 6480 9850 6820 9910
rect 8610 9850 8620 9910
rect 8680 9850 9020 9910
rect 10810 9850 10820 9910
rect 10880 9850 11220 9910
rect 13010 9850 13020 9910
rect 13080 9850 13420 9910
rect 15210 9850 15440 9910
rect 15500 9850 15620 9910
rect 17410 9850 17640 9910
rect 17700 9850 17820 9910
rect 27260 9904 27380 9950
rect 27370 9885 27380 9904
rect 27440 9950 27450 9975
rect 27440 9904 27950 9950
rect 27440 9885 27450 9904
rect 27370 9875 27450 9885
rect 2500 9810 4020 9822
rect 2500 9750 2510 9810
rect 4010 9750 4020 9810
rect 2500 9740 4020 9750
rect 4700 9810 6220 9822
rect 4700 9750 4710 9810
rect 6210 9750 6220 9810
rect 4700 9740 6220 9750
rect 6900 9810 8420 9822
rect 6900 9750 6910 9810
rect 8410 9750 8420 9810
rect 6900 9740 8420 9750
rect 9100 9810 10620 9822
rect 9100 9750 9110 9810
rect 10610 9750 10620 9810
rect 9100 9740 10620 9750
rect 11300 9810 12820 9822
rect 11300 9750 11310 9810
rect 12810 9750 12820 9810
rect 11300 9740 12820 9750
rect 13500 9810 15020 9822
rect 13500 9750 13510 9810
rect 15010 9750 15020 9810
rect 13500 9740 15020 9750
rect 15700 9810 17220 9822
rect 15700 9750 15710 9810
rect 17210 9750 17220 9810
rect 15700 9740 17220 9750
rect 17900 9810 19420 9822
rect 17900 9750 17910 9810
rect 19410 9750 19420 9810
rect 27730 9815 27810 9825
rect 27730 9792 27740 9815
rect 17900 9740 19420 9750
rect 27260 9746 27740 9792
rect 27730 9725 27740 9746
rect 27800 9792 27810 9815
rect 28770 9810 28820 10040
rect 29130 9970 29140 10040
rect 29200 9970 29210 10190
rect 29130 9960 29210 9970
rect 27800 9746 27950 9792
rect 27800 9725 27810 9746
rect 27730 9715 27810 9725
rect 29320 9640 29500 10520
rect 30100 11359 30229 13100
rect 30263 11380 30300 13123
rect 31260 12780 33820 12980
rect 31260 12260 31340 12780
rect 31920 12260 32140 12780
rect 32690 12280 32940 12780
rect 33520 12560 33820 12780
rect 33520 12540 38300 12560
rect 33520 12280 36920 12540
rect 38280 12280 38300 12540
rect 33520 12260 38300 12280
rect 35220 12230 38100 12260
rect 31220 11682 31340 11980
rect 31900 11682 32140 12000
rect 32690 11682 32950 12000
rect 33520 11900 33640 11980
rect 33520 11682 34874 11900
rect 31220 11660 31362 11682
rect 31532 11660 31712 11682
rect 31892 11660 32162 11682
rect 32332 11660 32512 11682
rect 32690 11660 32962 11682
rect 33132 11660 33312 11682
rect 33492 11660 34874 11682
rect 31220 11644 32680 11660
rect 32690 11644 34874 11660
rect 31220 11574 34874 11644
rect 31230 11500 34874 11574
rect 30263 11359 34324 11380
rect 30100 11308 34324 11359
rect 30100 11256 30330 11308
rect 34142 11256 34324 11308
rect 30100 11193 34324 11256
rect 30100 11172 34256 11193
rect 30100 9900 30300 11172
rect 30802 10876 33752 10896
rect 30802 10346 30826 10876
rect 31190 10826 33752 10876
rect 31190 10800 32680 10826
rect 32690 10800 33752 10826
rect 31190 10374 31340 10800
rect 31190 10346 31318 10374
rect 30802 10320 31318 10346
rect 31900 10320 32140 10800
rect 32690 10660 32950 10800
rect 32690 10322 32940 10660
rect 33520 10500 33752 10800
rect 32730 10320 32940 10322
rect 33530 10320 33752 10500
rect 31414 10262 31502 10280
rect 31414 10082 31422 10262
rect 31494 10082 31502 10262
rect 31414 10076 31502 10082
rect 31748 10262 31836 10280
rect 31748 10082 31756 10262
rect 31828 10082 31836 10262
rect 31748 10076 31836 10082
rect 32548 10262 32636 10280
rect 32548 10082 32556 10262
rect 32628 10082 32636 10262
rect 32548 10076 32636 10082
rect 33348 10262 33436 10280
rect 33348 10082 33356 10262
rect 33428 10082 33436 10262
rect 33348 10076 33436 10082
rect 34124 9900 34256 11172
rect 30100 9640 31340 9900
rect 2500 9580 2510 9640
rect 2690 9580 2700 9640
rect 2500 9340 2700 9580
rect 3160 9580 3170 9640
rect 3350 9580 3360 9640
rect 3160 9340 3360 9580
rect 3820 9580 3830 9640
rect 4010 9580 4020 9640
rect 3820 9340 4020 9580
rect 4700 9580 4710 9640
rect 4890 9580 4900 9640
rect 4700 9340 4900 9580
rect 5360 9580 5370 9640
rect 5550 9580 5560 9640
rect 5360 9340 5560 9580
rect 6020 9580 6030 9640
rect 6210 9580 6220 9640
rect 6020 9340 6220 9580
rect 6900 9500 7100 9640
rect 6900 9440 6910 9500
rect 7090 9440 7100 9500
rect 6900 9340 7100 9440
rect 7560 9500 7760 9640
rect 7560 9440 7570 9500
rect 7750 9440 7760 9500
rect 7560 9340 7760 9440
rect 8220 9500 8420 9640
rect 8220 9440 8230 9500
rect 8410 9440 8420 9500
rect 8220 9340 8420 9440
rect 9100 9500 9300 9640
rect 9100 9440 9110 9500
rect 9290 9440 9300 9500
rect 9100 9340 9300 9440
rect 9760 9500 9960 9640
rect 9760 9440 9770 9500
rect 9950 9440 9960 9500
rect 9760 9340 9960 9440
rect 10420 9500 10620 9640
rect 10420 9440 10430 9500
rect 10610 9440 10620 9500
rect 10420 9340 10620 9440
rect 11300 9500 11500 9640
rect 11300 9440 11310 9500
rect 11490 9440 11500 9500
rect 11300 9340 11500 9440
rect 11960 9500 12160 9640
rect 11960 9440 11970 9500
rect 12150 9440 12160 9500
rect 11960 9340 12160 9440
rect 12620 9500 12820 9640
rect 12620 9440 12630 9500
rect 12810 9440 12820 9500
rect 12620 9340 12820 9440
rect 13500 9500 13700 9640
rect 13500 9440 13510 9500
rect 13690 9440 13700 9500
rect 13500 9340 13700 9440
rect 14160 9500 14360 9640
rect 14160 9440 14170 9500
rect 14350 9440 14360 9500
rect 14160 9340 14360 9440
rect 14820 9500 15020 9640
rect 14820 9440 14830 9500
rect 15010 9440 15020 9500
rect 14820 9340 15020 9440
rect 15700 9580 15710 9640
rect 15890 9580 15900 9640
rect 15700 9340 15900 9580
rect 16360 9580 16370 9640
rect 16550 9580 16560 9640
rect 16360 9340 16560 9580
rect 17020 9580 17030 9640
rect 17210 9580 17220 9640
rect 17020 9340 17220 9580
rect 17900 9580 17910 9640
rect 18090 9580 18100 9640
rect 17900 9340 18100 9580
rect 18560 9580 18570 9640
rect 18750 9580 18760 9640
rect 18560 9340 18760 9580
rect 19220 9580 19230 9640
rect 19410 9580 19420 9640
rect 19220 9340 19420 9580
rect 27920 9480 31340 9640
rect 31900 9480 32140 9900
rect 32690 9480 32940 9900
rect 33500 9480 34256 9900
rect 27250 9405 27330 9415
rect -90 9330 10 9340
rect -90 9270 -70 9330
rect -10 9270 10 9330
rect -90 9260 10 9270
rect 2110 9330 2210 9340
rect 2110 9270 2130 9330
rect 2190 9270 2210 9330
rect 2110 9260 2210 9270
rect 4310 9330 4410 9340
rect 4310 9270 4330 9330
rect 4390 9270 4410 9330
rect 4310 9260 4410 9270
rect 6510 9330 6610 9340
rect 6510 9270 6530 9330
rect 6590 9270 6610 9330
rect 6510 9260 6610 9270
rect 8710 9330 8810 9340
rect 8710 9270 8730 9330
rect 8790 9270 8810 9330
rect 8710 9260 8810 9270
rect 10910 9330 11010 9340
rect 10910 9270 10930 9330
rect 10990 9270 11010 9330
rect 10910 9260 11010 9270
rect 13110 9330 13210 9340
rect 13110 9270 13130 9330
rect 13190 9270 13210 9330
rect 13110 9260 13210 9270
rect 15310 9330 15410 9340
rect 15310 9270 15330 9330
rect 15390 9270 15410 9330
rect 15310 9260 15410 9270
rect 17510 9330 17610 9340
rect 17510 9270 17530 9330
rect 17590 9270 17610 9330
rect 17510 9260 17610 9270
rect 19710 9330 19810 9340
rect 19710 9270 19730 9330
rect 19790 9270 19810 9330
rect 21910 9330 22010 9340
rect 19710 9260 19810 9270
rect 20230 9300 20310 9310
rect 1410 9210 1490 9220
rect 1410 9060 1420 9210
rect 1480 9110 1490 9210
rect 4100 9160 4510 9220
rect 6300 9160 6420 9220
rect 6480 9160 6710 9220
rect 8500 9160 8840 9220
rect 8900 9160 8910 9220
rect 10700 9160 11040 9220
rect 11100 9160 11110 9220
rect 12900 9160 13240 9220
rect 13300 9160 13310 9220
rect 15100 9160 15440 9220
rect 15500 9160 15510 9220
rect 17300 9160 17420 9220
rect 17480 9160 17710 9220
rect 20230 9200 20240 9300
rect 19500 9150 20240 9200
rect 20300 9150 20310 9300
rect 21910 9270 21930 9330
rect 21990 9270 22010 9330
rect 27250 9315 27260 9405
rect 27320 9384 27330 9405
rect 27320 9338 27950 9384
rect 27320 9315 27330 9338
rect 30100 9320 34256 9480
rect 27250 9305 27330 9315
rect 21910 9260 22010 9270
rect 27490 9250 27570 9260
rect 27490 9226 27500 9250
rect 27260 9180 27500 9226
rect 27490 9160 27500 9180
rect 27560 9226 27570 9250
rect 27560 9180 27950 9226
rect 27560 9160 27570 9180
rect 27490 9150 27570 9160
rect 19500 9140 20310 9150
rect 1480 9060 2420 9110
rect 1410 9050 2420 9060
rect 4210 9050 4220 9110
rect 4280 9050 4620 9110
rect 6410 9050 6640 9110
rect 6700 9050 6820 9110
rect 8610 9050 8840 9110
rect 8900 9050 9020 9110
rect 10810 9050 11040 9110
rect 11100 9050 11220 9110
rect 13010 9050 13240 9110
rect 13300 9050 13420 9110
rect 15210 9050 15220 9110
rect 15280 9050 15620 9110
rect 17410 9050 17820 9110
rect 28770 9100 28810 9320
rect 28870 9160 28950 9170
rect 28870 9100 28880 9160
rect 27250 9090 27330 9100
rect 4700 9010 6220 9022
rect 420 8990 620 9000
rect 420 8910 430 8990
rect 610 8980 620 8990
rect 610 8920 4040 8980
rect 4700 8950 4710 9010
rect 6210 8950 6220 9010
rect 4700 8940 6220 8950
rect 6900 9010 8420 9022
rect 6900 8950 6910 9010
rect 8410 8950 8420 9010
rect 6900 8940 8420 8950
rect 9100 9010 10620 9022
rect 9100 8950 9110 9010
rect 10610 8950 10620 9010
rect 9100 8940 10620 8950
rect 11300 9010 12820 9022
rect 11300 8950 11310 9010
rect 12810 8950 12820 9010
rect 11300 8940 12820 8950
rect 13500 9010 15020 9022
rect 13500 8950 13510 9010
rect 15010 8950 15020 9010
rect 13500 8940 15020 8950
rect 15700 9010 17220 9022
rect 15700 8950 15710 9010
rect 17210 8950 17220 9010
rect 27250 9000 27260 9090
rect 27320 9068 27330 9090
rect 27320 9022 27950 9068
rect 27320 9000 27330 9022
rect 21300 8990 21500 9000
rect 27250 8990 27330 9000
rect 28770 9000 28880 9100
rect 21300 8980 21310 8990
rect 15700 8940 17220 8950
rect 17880 8920 21310 8980
rect 610 8910 620 8920
rect 420 8900 620 8910
rect 21300 8910 21310 8920
rect 21490 8910 21500 8990
rect 27490 8935 27570 8945
rect 27490 8910 27500 8935
rect 21300 8900 21500 8910
rect 27260 8864 27500 8910
rect 27490 8845 27500 8864
rect 27560 8910 27570 8935
rect 27560 8864 27950 8910
rect 27560 8845 27570 8864
rect 2500 8700 2700 8840
rect 2500 8640 2510 8700
rect 2690 8640 2700 8700
rect 2500 8540 2700 8640
rect 3160 8700 3360 8840
rect 3160 8640 3170 8700
rect 3350 8640 3360 8700
rect 3160 8540 3360 8640
rect 3820 8700 4020 8840
rect 3820 8640 3830 8700
rect 4010 8640 4020 8700
rect 3820 8540 4020 8640
rect 4700 8700 4900 8840
rect 4700 8640 4710 8700
rect 4890 8640 4900 8700
rect 4700 8540 4900 8640
rect 5360 8700 5560 8840
rect 5360 8640 5370 8700
rect 5550 8640 5560 8700
rect 5360 8540 5560 8640
rect 6020 8700 6220 8840
rect 6020 8640 6030 8700
rect 6210 8640 6220 8700
rect 6020 8540 6220 8640
rect 6900 8780 6910 8840
rect 7090 8780 7100 8840
rect 6900 8540 7100 8780
rect 7560 8780 7570 8840
rect 7750 8780 7760 8840
rect 7560 8540 7760 8780
rect 8220 8780 8230 8840
rect 8410 8780 8420 8840
rect 8220 8540 8420 8780
rect 9100 8780 9110 8840
rect 9290 8780 9300 8840
rect 9100 8540 9300 8780
rect 9760 8780 9770 8840
rect 9950 8780 9960 8840
rect 9760 8540 9960 8780
rect 10420 8780 10430 8840
rect 10610 8780 10620 8840
rect 10420 8540 10620 8780
rect 11300 8780 11310 8840
rect 11490 8780 11500 8840
rect 11300 8540 11500 8780
rect 11960 8780 11970 8840
rect 12150 8780 12160 8840
rect 11960 8540 12160 8780
rect 12620 8780 12630 8840
rect 12810 8780 12820 8840
rect 12620 8540 12820 8780
rect 13500 8780 13510 8840
rect 13690 8780 13700 8840
rect 13500 8540 13700 8780
rect 14160 8780 14170 8840
rect 14350 8780 14360 8840
rect 14160 8540 14360 8780
rect 14820 8780 14830 8840
rect 15010 8780 15020 8840
rect 14820 8540 15020 8780
rect 15700 8700 15900 8840
rect 15700 8640 15710 8700
rect 15890 8640 15900 8700
rect 15700 8540 15900 8640
rect 16360 8700 16560 8840
rect 16360 8640 16370 8700
rect 16550 8640 16560 8700
rect 16360 8540 16560 8640
rect 17020 8700 17220 8840
rect 17020 8640 17030 8700
rect 17210 8640 17220 8700
rect 17020 8540 17220 8640
rect 17900 8700 18100 8840
rect 17900 8640 17910 8700
rect 18090 8640 18100 8700
rect 17900 8540 18100 8640
rect 18560 8700 18760 8840
rect 18560 8640 18570 8700
rect 18750 8640 18760 8700
rect 18560 8540 18760 8640
rect 19220 8700 19420 8840
rect 27490 8835 27570 8845
rect 19220 8640 19230 8700
rect 19410 8640 19420 8700
rect 27250 8775 27330 8785
rect 27250 8685 27260 8775
rect 27320 8752 27330 8775
rect 28770 8770 28810 9000
rect 28870 8940 28880 9000
rect 28940 8940 28950 9160
rect 28870 8930 28950 8940
rect 31180 9160 34256 9320
rect 27320 8706 27950 8752
rect 27320 8685 27330 8706
rect 27250 8675 27330 8685
rect 19220 8540 19420 8640
rect 31180 8620 32020 9160
rect 34124 9124 34256 9160
rect 34290 9140 34324 11193
rect 34474 11022 34874 11500
rect 35220 11290 35350 12230
rect 35400 12130 35800 12180
rect 35430 11250 35510 12130
rect 35570 11250 35620 12090
rect 35690 11250 35770 12130
rect 35990 12090 36050 12230
rect 36240 12130 36640 12180
rect 35840 11290 36200 12090
rect 36280 11250 36360 12130
rect 35390 11200 36370 11250
rect 34474 10846 34490 11022
rect 34848 10846 34874 11022
rect 34474 10820 34874 10846
rect 35450 9780 35520 11200
rect 36420 11150 36470 11420
rect 36530 11210 36610 12130
rect 36700 12030 38100 12230
rect 36700 11850 36940 12030
rect 37070 11850 37360 12030
rect 37490 11850 37780 12030
rect 37910 11850 38100 12030
rect 36700 11840 38100 11850
rect 36700 11290 36820 11840
rect 36870 11730 37110 11772
rect 37150 11740 37530 11770
rect 37570 11740 37950 11770
rect 36870 11150 36900 11730
rect 37150 11690 37190 11740
rect 37570 11690 37610 11740
rect 36980 11680 37060 11690
rect 36980 11300 36990 11680
rect 37050 11300 37060 11680
rect 36980 11290 37060 11300
rect 36420 11110 36900 11150
rect 36420 11050 36730 11110
rect 36640 10780 36730 11050
rect 37060 10780 37100 11240
rect 35900 10730 37100 10780
rect 35600 10570 35650 10690
rect 35600 10190 35780 10570
rect 35600 10010 35650 10190
rect 35810 10150 35860 10650
rect 35900 10510 35930 10730
rect 35970 10150 36020 10650
rect 35810 10140 36020 10150
rect 35810 10070 35820 10140
rect 36010 10070 36020 10140
rect 35810 10060 36020 10070
rect 36060 10010 36090 10310
rect 36130 10150 36180 10650
rect 36220 10500 36250 10730
rect 36290 10150 36340 10650
rect 36490 10570 36540 10690
rect 36380 10190 36540 10570
rect 36130 10140 36340 10150
rect 36130 10070 36140 10140
rect 36330 10070 36340 10140
rect 36130 10060 36340 10070
rect 36490 10012 36540 10190
rect 36640 10270 36730 10730
rect 37060 10550 37100 10730
rect 37140 11020 37190 11690
rect 37400 11680 37480 11690
rect 37400 11300 37410 11680
rect 37470 11300 37480 11680
rect 37400 11290 37480 11300
rect 37140 11010 37350 11020
rect 37140 10860 37190 11010
rect 37340 10860 37350 11010
rect 37140 10850 37350 10860
rect 37140 10780 37190 10850
rect 37480 10780 37520 11240
rect 37140 10730 37520 10780
rect 36980 10500 37060 10510
rect 36980 10320 36990 10500
rect 37050 10320 37060 10500
rect 36980 10310 37060 10320
rect 37140 10310 37190 10730
rect 37480 10550 37520 10730
rect 37560 10780 37610 11690
rect 37820 11680 37900 11690
rect 37820 11300 37830 11680
rect 37890 11300 37900 11680
rect 37820 11290 37900 11300
rect 37900 10780 37940 11240
rect 37560 10750 37940 10780
rect 37560 10600 37610 10750
rect 37760 10730 37940 10750
rect 37760 10600 37770 10730
rect 37560 10590 37770 10600
rect 37400 10500 37480 10510
rect 37400 10320 37410 10500
rect 37470 10320 37480 10500
rect 37400 10310 37480 10320
rect 37560 10310 37610 10590
rect 37900 10550 37940 10730
rect 37980 10970 38030 11690
rect 37980 10960 38130 10970
rect 37980 10780 37990 10960
rect 38120 10780 38130 10960
rect 37980 10770 38130 10780
rect 37820 10500 37900 10510
rect 37820 10320 37830 10500
rect 37890 10320 37900 10500
rect 37820 10310 37900 10320
rect 37980 10310 38030 10770
rect 39500 10434 39566 13500
rect 38268 10406 39566 10434
rect 37150 10270 37190 10310
rect 37570 10270 37610 10310
rect 36640 10240 37110 10270
rect 37150 10240 37520 10270
rect 37570 10240 37950 10270
rect 36640 10040 36730 10240
rect 36930 10160 38070 10170
rect 38268 10160 38298 10406
rect 36410 10010 36560 10012
rect 35600 9960 36560 10010
rect 36410 9924 36560 9960
rect 36640 9940 36840 10040
rect 36930 9980 36950 10160
rect 37080 9980 37370 10160
rect 37500 9980 37790 10160
rect 37920 9980 38298 10160
rect 36930 9970 38298 9980
rect 35450 9720 36220 9780
rect 35250 9664 35394 9676
rect 35250 9542 35266 9664
rect 35384 9660 35394 9664
rect 35384 9560 36300 9660
rect 35384 9542 35400 9560
rect 35250 9526 35400 9542
rect 35360 9520 35400 9526
rect 35440 9496 36240 9500
rect 36410 9496 36430 9924
rect 35438 9434 36430 9496
rect 36542 9496 36560 9924
rect 36750 9780 36840 9940
rect 38266 9848 38298 9970
rect 39274 9848 39566 10406
rect 38266 9820 39566 9848
rect 36750 9720 37520 9780
rect 37572 9664 37716 9680
rect 37572 9660 37584 9664
rect 36680 9560 37584 9660
rect 37572 9542 37584 9560
rect 37702 9542 37716 9664
rect 37572 9530 37716 9542
rect 36750 9496 37520 9500
rect 36542 9434 37534 9496
rect 35438 9384 37534 9434
rect 34290 9124 39350 9140
rect 34124 9058 39350 9124
rect 34124 9024 34352 9058
rect 39163 9024 39350 9058
rect 34124 8958 39350 9024
rect 34124 8940 39229 8958
rect -90 8530 10 8540
rect -90 8470 -70 8530
rect -10 8470 10 8530
rect -90 8460 10 8470
rect 2110 8530 2210 8540
rect 2110 8470 2130 8530
rect 2190 8470 2210 8530
rect 2110 8460 2210 8470
rect 4310 8530 4410 8540
rect 4310 8470 4330 8530
rect 4390 8470 4410 8530
rect 4310 8460 4410 8470
rect 6510 8530 6610 8540
rect 6510 8470 6530 8530
rect 6590 8470 6610 8530
rect 6510 8460 6610 8470
rect 8710 8530 8810 8540
rect 8710 8470 8730 8530
rect 8790 8470 8810 8530
rect 8710 8460 8810 8470
rect 10910 8530 11010 8540
rect 10910 8470 10930 8530
rect 10990 8470 11010 8530
rect 10910 8460 11010 8470
rect 13110 8530 13210 8540
rect 13110 8470 13130 8530
rect 13190 8470 13210 8530
rect 13110 8460 13210 8470
rect 15310 8530 15410 8540
rect 15310 8470 15330 8530
rect 15390 8470 15410 8530
rect 15310 8460 15410 8470
rect 17510 8530 17610 8540
rect 17510 8470 17530 8530
rect 17590 8470 17610 8530
rect 17510 8460 17610 8470
rect 19710 8530 19810 8540
rect 19710 8470 19730 8530
rect 19790 8470 19810 8530
rect 21910 8530 22010 8540
rect 19710 8460 19810 8470
rect 20430 8500 20510 8510
rect 1610 8410 1690 8420
rect 1610 8260 1620 8410
rect 1680 8310 1690 8410
rect 4100 8360 4510 8420
rect 6300 8360 6640 8420
rect 6700 8360 6710 8420
rect 8500 8360 8620 8420
rect 8680 8360 8910 8420
rect 10700 8360 10820 8420
rect 10880 8360 11110 8420
rect 12900 8360 13020 8420
rect 13080 8360 13310 8420
rect 15100 8360 15220 8420
rect 15280 8360 15510 8420
rect 17300 8360 17640 8420
rect 17700 8360 17710 8420
rect 20430 8400 20440 8500
rect 19500 8350 20440 8400
rect 20500 8350 20510 8500
rect 21910 8470 21930 8530
rect 21990 8470 22010 8530
rect 21910 8460 22010 8470
rect 27920 8460 32020 8620
rect 35444 8558 37528 8670
rect 35442 8482 37530 8558
rect 19500 8340 20510 8350
rect 27250 8370 27330 8380
rect 1680 8260 2420 8310
rect 1610 8250 2420 8260
rect 4210 8250 4440 8310
rect 4500 8250 4620 8310
rect 6410 8250 6420 8310
rect 6480 8250 6820 8310
rect 8610 8250 8620 8310
rect 8680 8250 9020 8310
rect 10810 8250 10820 8310
rect 10880 8250 11220 8310
rect 13010 8250 13020 8310
rect 13080 8250 13420 8310
rect 15210 8250 15440 8310
rect 15500 8250 15620 8310
rect 17410 8250 17820 8310
rect 27250 8280 27260 8370
rect 27320 8344 27330 8370
rect 27320 8298 27950 8344
rect 27320 8280 27330 8298
rect 27250 8270 27330 8280
rect 4700 8210 6220 8222
rect 420 8190 620 8200
rect 420 8110 430 8190
rect 610 8180 620 8190
rect 610 8120 4040 8180
rect 4700 8150 4710 8210
rect 6210 8150 6220 8210
rect 4700 8140 6220 8150
rect 6900 8210 8420 8222
rect 6900 8150 6910 8210
rect 8410 8150 8420 8210
rect 6900 8140 8420 8150
rect 9100 8210 10620 8222
rect 9100 8150 9110 8210
rect 10610 8150 10620 8210
rect 9100 8140 10620 8150
rect 11300 8210 12820 8222
rect 11300 8150 11310 8210
rect 12810 8150 12820 8210
rect 11300 8140 12820 8150
rect 13500 8210 15020 8222
rect 13500 8150 13510 8210
rect 15010 8150 15020 8210
rect 13500 8140 15020 8150
rect 15700 8210 17220 8222
rect 15700 8150 15710 8210
rect 17210 8150 17220 8210
rect 27610 8210 27690 8220
rect 21300 8190 21500 8200
rect 21300 8180 21310 8190
rect 15700 8140 17220 8150
rect 17880 8120 21310 8180
rect 610 8110 620 8120
rect 420 8100 620 8110
rect 21300 8110 21310 8120
rect 21490 8110 21500 8190
rect 27610 8186 27620 8210
rect 27260 8140 27620 8186
rect 27610 8120 27620 8140
rect 27680 8186 27690 8210
rect 27680 8140 27950 8186
rect 27680 8120 27690 8140
rect 27610 8110 27690 8120
rect 21300 8100 21500 8110
rect 27250 8050 27330 8060
rect 2500 7900 2700 8040
rect 2500 7840 2510 7900
rect 2690 7840 2700 7900
rect 2500 7740 2700 7840
rect 3160 7900 3360 8040
rect 3160 7840 3170 7900
rect 3350 7840 3360 7900
rect 3160 7740 3360 7840
rect 3820 7900 4020 8040
rect 3820 7840 3830 7900
rect 4010 7840 4020 7900
rect 3820 7740 4020 7840
rect 4700 7900 4900 8040
rect 4700 7840 4710 7900
rect 4890 7840 4900 7900
rect 4700 7740 4900 7840
rect 5360 7900 5560 8040
rect 5360 7840 5370 7900
rect 5550 7840 5560 7900
rect 5360 7740 5560 7840
rect 6020 7900 6220 8040
rect 6020 7840 6030 7900
rect 6210 7840 6220 7900
rect 6020 7740 6220 7840
rect 6900 7980 6910 8040
rect 7090 7980 7100 8040
rect 6900 7740 7100 7980
rect 7560 7980 7570 8040
rect 7750 7980 7760 8040
rect 7560 7740 7760 7980
rect 8220 7980 8230 8040
rect 8410 7980 8420 8040
rect 8220 7740 8420 7980
rect 9100 7980 9110 8040
rect 9290 7980 9300 8040
rect 9100 7740 9300 7980
rect 9760 7980 9770 8040
rect 9950 7980 9960 8040
rect 9760 7740 9960 7980
rect 10420 7980 10430 8040
rect 10610 7980 10620 8040
rect 10420 7740 10620 7980
rect 11300 7980 11310 8040
rect 11490 7980 11500 8040
rect 11300 7740 11500 7980
rect 11960 7980 11970 8040
rect 12150 7980 12160 8040
rect 11960 7740 12160 7980
rect 12620 7980 12630 8040
rect 12810 7980 12820 8040
rect 12620 7740 12820 7980
rect 13500 7980 13510 8040
rect 13690 7980 13700 8040
rect 13500 7740 13700 7980
rect 14160 7980 14170 8040
rect 14350 7980 14360 8040
rect 14160 7740 14360 7980
rect 14820 7980 14830 8040
rect 15010 7980 15020 8040
rect 14820 7740 15020 7980
rect 15700 7900 15900 8040
rect 15700 7840 15710 7900
rect 15890 7840 15900 7900
rect 15700 7740 15900 7840
rect 16360 7900 16560 8040
rect 16360 7840 16370 7900
rect 16550 7840 16560 7900
rect 16360 7740 16560 7840
rect 17020 7900 17220 8040
rect 17020 7840 17030 7900
rect 17210 7840 17220 7900
rect 17020 7740 17220 7840
rect 17900 7900 18100 8040
rect 17900 7840 17910 7900
rect 18090 7840 18100 7900
rect 17900 7740 18100 7840
rect 18560 7900 18760 8040
rect 18560 7840 18570 7900
rect 18750 7840 18760 7900
rect 18560 7740 18760 7840
rect 19220 7900 19420 8040
rect 27250 7960 27260 8050
rect 27320 8028 27330 8050
rect 28770 8050 28810 8280
rect 29000 8110 29080 8120
rect 29000 8050 29010 8110
rect 27320 7982 27950 8028
rect 27320 7960 27330 7982
rect 27250 7950 27330 7960
rect 28770 7960 29010 8050
rect 19220 7840 19230 7900
rect 19410 7840 19420 7900
rect 27610 7890 27690 7900
rect 27610 7870 27620 7890
rect 19220 7740 19420 7840
rect 27260 7824 27620 7870
rect 27610 7800 27620 7824
rect 27680 7870 27690 7890
rect 27680 7824 27950 7870
rect 27680 7800 27690 7824
rect 27610 7790 27690 7800
rect 27250 7740 27330 7750
rect -90 7730 10 7740
rect -90 7670 -70 7730
rect -10 7670 10 7730
rect -90 7660 10 7670
rect 2110 7730 2210 7740
rect 2110 7670 2130 7730
rect 2190 7670 2210 7730
rect 2110 7660 2210 7670
rect 4310 7730 4410 7740
rect 4310 7670 4330 7730
rect 4390 7670 4410 7730
rect 4310 7660 4410 7670
rect 6510 7730 6610 7740
rect 6510 7670 6530 7730
rect 6590 7670 6610 7730
rect 6510 7660 6610 7670
rect 8710 7730 8810 7740
rect 8710 7670 8730 7730
rect 8790 7670 8810 7730
rect 8710 7660 8810 7670
rect 10910 7730 11010 7740
rect 10910 7670 10930 7730
rect 10990 7670 11010 7730
rect 10910 7660 11010 7670
rect 13110 7730 13210 7740
rect 13110 7670 13130 7730
rect 13190 7670 13210 7730
rect 13110 7660 13210 7670
rect 15310 7730 15410 7740
rect 15310 7670 15330 7730
rect 15390 7670 15410 7730
rect 15310 7660 15410 7670
rect 17510 7730 17610 7740
rect 17510 7670 17530 7730
rect 17590 7670 17610 7730
rect 17510 7660 17610 7670
rect 19710 7730 19810 7740
rect 19710 7670 19730 7730
rect 19790 7670 19810 7730
rect 21910 7730 22010 7740
rect 19710 7660 19810 7670
rect 20430 7700 20510 7710
rect 1610 7610 1690 7620
rect 1610 7460 1620 7610
rect 1680 7510 1690 7610
rect 4100 7560 4510 7620
rect 6300 7560 6640 7620
rect 6700 7560 6710 7620
rect 8500 7560 8620 7620
rect 8680 7560 8910 7620
rect 10700 7560 10820 7620
rect 10880 7560 11110 7620
rect 12900 7560 13020 7620
rect 13080 7560 13310 7620
rect 15100 7560 15220 7620
rect 15280 7560 15510 7620
rect 17300 7560 17640 7620
rect 17700 7560 17710 7620
rect 20430 7600 20440 7700
rect 19500 7550 20440 7600
rect 20500 7550 20510 7700
rect 21910 7670 21930 7730
rect 21990 7670 22010 7730
rect 21910 7660 22010 7670
rect 27250 7650 27260 7740
rect 27320 7712 27330 7740
rect 28770 7730 28810 7960
rect 29000 7890 29010 7960
rect 29070 7890 29080 8110
rect 31180 7980 32020 8460
rect 35360 8426 35400 8428
rect 35238 8414 35400 8426
rect 35238 8292 35254 8414
rect 35372 8400 35400 8414
rect 36270 8400 36320 8448
rect 35372 8300 36320 8400
rect 35372 8292 35400 8300
rect 35238 8280 35400 8292
rect 29000 7880 29080 7890
rect 29540 7860 32020 7980
rect 27320 7666 27950 7712
rect 27320 7650 27330 7666
rect 27250 7640 27330 7650
rect 29540 7660 29900 7860
rect 29540 7560 29920 7660
rect 19500 7540 20510 7550
rect 1680 7460 2420 7510
rect 1610 7450 2420 7460
rect 4210 7450 4440 7510
rect 4500 7450 4620 7510
rect 6410 7450 6420 7510
rect 6480 7450 6820 7510
rect 8610 7450 8620 7510
rect 8680 7450 9020 7510
rect 10810 7450 10820 7510
rect 10880 7450 11220 7510
rect 13010 7450 13020 7510
rect 13080 7450 13420 7510
rect 15210 7450 15440 7510
rect 15500 7450 15620 7510
rect 17410 7450 17820 7510
rect 4700 7410 6220 7422
rect 420 7390 620 7400
rect 420 7310 430 7390
rect 610 7380 620 7390
rect 610 7320 4040 7380
rect 4700 7350 4710 7410
rect 6210 7350 6220 7410
rect 4700 7340 6220 7350
rect 6900 7410 8420 7422
rect 6900 7350 6910 7410
rect 8410 7350 8420 7410
rect 6900 7340 8420 7350
rect 9100 7410 10620 7422
rect 9100 7350 9110 7410
rect 10610 7350 10620 7410
rect 9100 7340 10620 7350
rect 11300 7410 12820 7422
rect 11300 7350 11310 7410
rect 12810 7350 12820 7410
rect 11300 7340 12820 7350
rect 13500 7410 15020 7422
rect 13500 7350 13510 7410
rect 15010 7350 15020 7410
rect 13500 7340 15020 7350
rect 15700 7410 17220 7422
rect 15700 7350 15710 7410
rect 17210 7350 17220 7410
rect 27920 7400 29920 7560
rect 21300 7390 21500 7400
rect 21300 7380 21310 7390
rect 15700 7340 17220 7350
rect 17880 7320 21310 7380
rect 610 7310 620 7320
rect 420 7300 620 7310
rect 21300 7310 21310 7320
rect 21490 7310 21500 7390
rect 21300 7300 21500 7310
rect 27370 7330 27450 7340
rect 27370 7304 27380 7330
rect 27260 7258 27380 7304
rect 27370 7240 27380 7258
rect 27440 7304 27450 7330
rect 27440 7258 27950 7304
rect 29540 7300 29920 7400
rect 29540 7260 29900 7300
rect 27440 7240 27450 7258
rect 2500 7180 2510 7240
rect 2690 7180 2700 7240
rect 2500 6940 2700 7180
rect 3160 7180 3170 7240
rect 3350 7180 3360 7240
rect 3160 6940 3360 7180
rect 3820 7180 3830 7240
rect 4010 7180 4020 7240
rect 3820 6940 4020 7180
rect 4700 7180 4710 7240
rect 4890 7180 4900 7240
rect 4700 6940 4900 7180
rect 5360 7180 5370 7240
rect 5550 7180 5560 7240
rect 5360 6940 5560 7180
rect 6020 7180 6030 7240
rect 6210 7180 6220 7240
rect 6020 6940 6220 7180
rect 6900 7100 7100 7240
rect 6900 7040 6910 7100
rect 7090 7040 7100 7100
rect 6900 6940 7100 7040
rect 7560 7100 7760 7240
rect 7560 7040 7570 7100
rect 7750 7040 7760 7100
rect 7560 6940 7760 7040
rect 8220 7100 8420 7240
rect 8220 7040 8230 7100
rect 8410 7040 8420 7100
rect 8220 6940 8420 7040
rect 9100 7100 9300 7240
rect 9100 7040 9110 7100
rect 9290 7040 9300 7100
rect 9100 6940 9300 7040
rect 9760 7100 9960 7240
rect 9760 7040 9770 7100
rect 9950 7040 9960 7100
rect 9760 6940 9960 7040
rect 10420 7100 10620 7240
rect 10420 7040 10430 7100
rect 10610 7040 10620 7100
rect 10420 6940 10620 7040
rect 11300 7100 11500 7240
rect 11300 7040 11310 7100
rect 11490 7040 11500 7100
rect 11300 6940 11500 7040
rect 11960 7100 12160 7240
rect 11960 7040 11970 7100
rect 12150 7040 12160 7100
rect 11960 6940 12160 7040
rect 12620 7100 12820 7240
rect 12620 7040 12630 7100
rect 12810 7040 12820 7100
rect 12620 6940 12820 7040
rect 13500 7100 13700 7240
rect 13500 7040 13510 7100
rect 13690 7040 13700 7100
rect 13500 6940 13700 7040
rect 14160 7100 14360 7240
rect 14160 7040 14170 7100
rect 14350 7040 14360 7100
rect 14160 6940 14360 7040
rect 14820 7100 15020 7240
rect 14820 7040 14830 7100
rect 15010 7040 15020 7100
rect 14820 6940 15020 7040
rect 15700 7180 15710 7240
rect 15890 7180 15900 7240
rect 15700 6940 15900 7180
rect 16360 7180 16370 7240
rect 16550 7180 16560 7240
rect 16360 6940 16560 7180
rect 17020 7180 17030 7240
rect 17210 7180 17220 7240
rect 17020 6940 17220 7180
rect 17900 7180 17910 7240
rect 18090 7180 18100 7240
rect 17900 6940 18100 7180
rect 18560 7180 18570 7240
rect 18750 7180 18760 7240
rect 18560 6940 18760 7180
rect 19220 7180 19230 7240
rect 19410 7180 19420 7240
rect 27370 7230 27450 7240
rect 19220 6940 19420 7180
rect 27610 7170 27690 7180
rect 27610 7146 27620 7170
rect 27260 7100 27620 7146
rect 27610 7080 27620 7100
rect 27680 7146 27690 7170
rect 27680 7100 27950 7146
rect 27680 7080 27690 7100
rect 27610 7070 27690 7080
rect 27370 7015 27450 7025
rect 27370 6988 27380 7015
rect 27260 6942 27380 6988
rect -90 6930 10 6940
rect -90 6870 -70 6930
rect -10 6870 10 6930
rect -90 6860 10 6870
rect 2110 6930 2210 6940
rect 2110 6870 2130 6930
rect 2190 6870 2210 6930
rect 2110 6860 2210 6870
rect 4310 6930 4410 6940
rect 4310 6870 4330 6930
rect 4390 6870 4410 6930
rect 4310 6860 4410 6870
rect 6510 6930 6610 6940
rect 6510 6870 6530 6930
rect 6590 6870 6610 6930
rect 6510 6860 6610 6870
rect 8710 6930 8810 6940
rect 8710 6870 8730 6930
rect 8790 6870 8810 6930
rect 8710 6860 8810 6870
rect 10910 6930 11010 6940
rect 10910 6870 10930 6930
rect 10990 6870 11010 6930
rect 10910 6860 11010 6870
rect 13110 6930 13210 6940
rect 13110 6870 13130 6930
rect 13190 6870 13210 6930
rect 13110 6860 13210 6870
rect 15310 6930 15410 6940
rect 15310 6870 15330 6930
rect 15390 6870 15410 6930
rect 15310 6860 15410 6870
rect 17510 6930 17610 6940
rect 17510 6870 17530 6930
rect 17590 6870 17610 6930
rect 17510 6860 17610 6870
rect 19710 6930 19810 6940
rect 19710 6870 19730 6930
rect 19790 6870 19810 6930
rect 21910 6930 22010 6940
rect 19710 6860 19810 6870
rect 20230 6900 20310 6910
rect 1410 6810 1490 6820
rect 1410 6660 1420 6810
rect 1480 6710 1490 6810
rect 4100 6760 4510 6820
rect 6300 6760 6420 6820
rect 6480 6760 6710 6820
rect 8500 6760 8840 6820
rect 8900 6760 8910 6820
rect 10700 6760 11040 6820
rect 11100 6760 11110 6820
rect 12900 6760 13240 6820
rect 13300 6760 13310 6820
rect 15100 6760 15440 6820
rect 15500 6760 15510 6820
rect 17300 6760 17420 6820
rect 17480 6760 17710 6820
rect 20230 6800 20240 6900
rect 19500 6750 20240 6800
rect 20300 6750 20310 6900
rect 21910 6870 21930 6930
rect 21990 6870 22010 6930
rect 27370 6925 27380 6942
rect 27440 6988 27450 7015
rect 28770 7020 28810 7240
rect 28870 7080 28950 7090
rect 28870 7020 28880 7080
rect 27440 6942 27950 6988
rect 27440 6925 27450 6942
rect 27370 6915 27450 6925
rect 21910 6860 22010 6870
rect 28770 6910 28880 7020
rect 27610 6855 27690 6865
rect 27610 6830 27620 6855
rect 27260 6784 27620 6830
rect 27610 6765 27620 6784
rect 27680 6830 27690 6855
rect 27680 6784 27950 6830
rect 27680 6765 27690 6784
rect 27610 6755 27690 6765
rect 19500 6740 20310 6750
rect 1480 6660 2420 6710
rect 1410 6650 2420 6660
rect 4210 6650 4220 6710
rect 4280 6650 4620 6710
rect 6410 6650 6640 6710
rect 6700 6650 6820 6710
rect 8610 6650 8840 6710
rect 8900 6650 9020 6710
rect 10810 6650 11040 6710
rect 11100 6650 11220 6710
rect 13010 6650 13240 6710
rect 13300 6650 13420 6710
rect 15210 6650 15220 6710
rect 15280 6650 15620 6710
rect 17410 6650 17820 6710
rect 27370 6700 27450 6710
rect 27370 6672 27380 6700
rect 27260 6626 27380 6672
rect 4700 6610 6220 6622
rect 420 6590 620 6600
rect 420 6510 430 6590
rect 610 6580 620 6590
rect 610 6520 4040 6580
rect 4700 6550 4710 6610
rect 6210 6550 6220 6610
rect 4700 6540 6220 6550
rect 6900 6610 8420 6622
rect 6900 6550 6910 6610
rect 8410 6550 8420 6610
rect 6900 6540 8420 6550
rect 9100 6610 10620 6622
rect 9100 6550 9110 6610
rect 10610 6550 10620 6610
rect 9100 6540 10620 6550
rect 11300 6610 12820 6622
rect 11300 6550 11310 6610
rect 12810 6550 12820 6610
rect 11300 6540 12820 6550
rect 13500 6610 15020 6622
rect 13500 6550 13510 6610
rect 15010 6550 15020 6610
rect 13500 6540 15020 6550
rect 15700 6610 17220 6622
rect 15700 6550 15710 6610
rect 17210 6550 17220 6610
rect 27370 6610 27380 6626
rect 27440 6672 27450 6700
rect 28770 6690 28810 6910
rect 28870 6860 28880 6910
rect 28940 6860 28950 7080
rect 28870 6850 28950 6860
rect 27440 6626 27950 6672
rect 29540 6660 29840 7260
rect 30280 7220 30400 7760
rect 30720 7220 30820 7680
rect 31140 7220 31260 7760
rect 31640 7660 32020 7860
rect 35360 8240 35400 8280
rect 35360 8230 35460 8240
rect 35490 8230 36220 8240
rect 36270 8230 36320 8300
rect 35360 8180 36320 8230
rect 35360 7930 35460 8180
rect 36410 7970 36572 8482
rect 36660 8400 36700 8434
rect 37580 8428 37620 8432
rect 37580 8416 37732 8428
rect 37580 8400 37600 8416
rect 36660 8300 37600 8400
rect 36660 8240 36700 8300
rect 37580 8294 37600 8300
rect 37718 8294 37732 8416
rect 37580 8282 37732 8294
rect 37580 8240 37620 8282
rect 36660 8180 37620 8240
rect 36350 7930 36572 7970
rect 35360 7920 35500 7930
rect 35360 7800 35370 7920
rect 35490 7800 35500 7920
rect 35360 7790 35500 7800
rect 35360 7750 35460 7790
rect 35360 7700 35850 7750
rect 31620 7300 32020 7660
rect 35340 7690 35850 7700
rect 35340 7570 35350 7690
rect 35470 7670 35850 7690
rect 35470 7570 35480 7670
rect 35340 7560 35480 7570
rect 36000 7620 36140 7830
rect 36410 7750 36572 7930
rect 36870 7920 37010 7930
rect 36870 7800 36880 7920
rect 37000 7800 37010 7920
rect 36280 7670 36720 7750
rect 36000 7500 36010 7620
rect 36130 7500 36140 7620
rect 36000 7490 36140 7500
rect 31640 7280 32020 7300
rect 29940 7210 31580 7220
rect 29940 7140 31290 7210
rect 30720 6840 30820 7140
rect 31280 7090 31290 7140
rect 31570 7090 31580 7210
rect 31280 7080 31580 7090
rect 30280 6720 31260 6840
rect 27440 6610 27450 6626
rect 27370 6600 27450 6610
rect 21300 6590 21500 6600
rect 21300 6580 21310 6590
rect 15700 6540 17220 6550
rect 17880 6520 21310 6580
rect 610 6510 620 6520
rect 420 6500 620 6510
rect 21300 6510 21310 6520
rect 21490 6510 21500 6590
rect 29540 6520 29900 6660
rect 21300 6500 21500 6510
rect 2500 6300 2700 6440
rect 2500 6240 2510 6300
rect 2690 6240 2700 6300
rect 2500 6140 2700 6240
rect 3160 6300 3360 6440
rect 3160 6240 3170 6300
rect 3350 6240 3360 6300
rect 3160 6140 3360 6240
rect 3820 6300 4020 6440
rect 3820 6240 3830 6300
rect 4010 6240 4020 6300
rect 3820 6140 4020 6240
rect 4700 6300 4900 6440
rect 4700 6240 4710 6300
rect 4890 6240 4900 6300
rect 4700 6140 4900 6240
rect 5360 6300 5560 6440
rect 5360 6240 5370 6300
rect 5550 6240 5560 6300
rect 5360 6140 5560 6240
rect 6020 6300 6220 6440
rect 6020 6240 6030 6300
rect 6210 6240 6220 6300
rect 6020 6140 6220 6240
rect 6900 6380 6910 6440
rect 7090 6380 7100 6440
rect 6900 6140 7100 6380
rect 7560 6380 7570 6440
rect 7750 6380 7760 6440
rect 7560 6140 7760 6380
rect 8220 6380 8230 6440
rect 8410 6380 8420 6440
rect 8220 6140 8420 6380
rect 9100 6380 9110 6440
rect 9290 6380 9300 6440
rect 9100 6140 9300 6380
rect 9760 6380 9770 6440
rect 9950 6380 9960 6440
rect 9760 6140 9960 6380
rect 10420 6380 10430 6440
rect 10610 6380 10620 6440
rect 10420 6140 10620 6380
rect 11300 6380 11310 6440
rect 11490 6380 11500 6440
rect 11300 6140 11500 6380
rect 11960 6380 11970 6440
rect 12150 6380 12160 6440
rect 11960 6140 12160 6380
rect 12620 6380 12630 6440
rect 12810 6380 12820 6440
rect 12620 6140 12820 6380
rect 13500 6380 13510 6440
rect 13690 6380 13700 6440
rect 13500 6140 13700 6380
rect 14160 6380 14170 6440
rect 14350 6380 14360 6440
rect 14160 6140 14360 6380
rect 14820 6380 14830 6440
rect 15010 6380 15020 6440
rect 14820 6140 15020 6380
rect 15700 6300 15900 6440
rect 15700 6240 15710 6300
rect 15890 6240 15900 6300
rect 15700 6140 15900 6240
rect 16360 6300 16560 6440
rect 16360 6240 16370 6300
rect 16550 6240 16560 6300
rect 16360 6140 16560 6240
rect 17020 6300 17220 6440
rect 17020 6240 17030 6300
rect 17210 6240 17220 6300
rect 17020 6140 17220 6240
rect 17900 6300 18100 6440
rect 17900 6240 17910 6300
rect 18090 6240 18100 6300
rect 17900 6140 18100 6240
rect 18560 6300 18760 6440
rect 18560 6240 18570 6300
rect 18750 6240 18760 6300
rect 18560 6140 18760 6240
rect 19220 6300 19420 6440
rect 27920 6360 29900 6520
rect 19220 6240 19230 6300
rect 19410 6240 19420 6300
rect 27370 6290 27450 6300
rect 27370 6264 27380 6290
rect 19220 6140 19420 6240
rect 27260 6218 27380 6264
rect 27370 6200 27380 6218
rect 27440 6264 27450 6290
rect 27440 6218 27950 6264
rect 27440 6200 27450 6218
rect 27370 6190 27450 6200
rect -90 6130 10 6140
rect -90 6070 -70 6130
rect -10 6070 10 6130
rect -90 6060 10 6070
rect 2110 6130 2210 6140
rect 2110 6070 2130 6130
rect 2190 6070 2210 6130
rect 2110 6060 2210 6070
rect 4310 6130 4410 6140
rect 4310 6070 4330 6130
rect 4390 6070 4410 6130
rect 4310 6060 4410 6070
rect 6510 6130 6610 6140
rect 6510 6070 6530 6130
rect 6590 6070 6610 6130
rect 6510 6060 6610 6070
rect 8710 6130 8810 6140
rect 8710 6070 8730 6130
rect 8790 6070 8810 6130
rect 8710 6060 8810 6070
rect 10910 6130 11010 6140
rect 10910 6070 10930 6130
rect 10990 6070 11010 6130
rect 10910 6060 11010 6070
rect 13110 6130 13210 6140
rect 13110 6070 13130 6130
rect 13190 6070 13210 6130
rect 13110 6060 13210 6070
rect 15310 6130 15410 6140
rect 15310 6070 15330 6130
rect 15390 6070 15410 6130
rect 15310 6060 15410 6070
rect 17510 6130 17610 6140
rect 17510 6070 17530 6130
rect 17590 6070 17610 6130
rect 17510 6060 17610 6070
rect 19710 6130 19810 6140
rect 19710 6070 19730 6130
rect 19790 6070 19810 6130
rect 19710 6060 19810 6070
rect 21910 6130 22010 6140
rect 21910 6070 21930 6130
rect 21990 6070 22010 6130
rect 27490 6130 27570 6140
rect 27490 6106 27500 6130
rect 21910 6060 22010 6070
rect 27260 6060 27500 6106
rect 27490 6040 27500 6060
rect 27560 6106 27570 6130
rect 27560 6060 27950 6106
rect 27560 6040 27570 6060
rect 27490 6030 27570 6040
rect 4100 5960 4440 6020
rect 4500 5960 4510 6020
rect 6300 5960 6640 6020
rect 6700 5960 6710 6020
rect 8500 5960 8620 6020
rect 8680 5960 8910 6020
rect 10700 5960 10820 6020
rect 10880 5960 11110 6020
rect 12900 5960 13020 6020
rect 13080 5960 13310 6020
rect 15100 5960 15220 6020
rect 15280 5960 15510 6020
rect 17300 5960 17640 6020
rect 17700 5960 17710 6020
rect 19500 5940 19840 6000
rect 19900 5940 19910 6000
rect 27370 5975 27450 5985
rect 27370 5948 27380 5975
rect 2010 5850 2240 5910
rect 2300 5850 2420 5910
rect 4210 5850 4440 5910
rect 4500 5850 4620 5910
rect 6410 5850 6420 5910
rect 6480 5850 6820 5910
rect 8610 5850 8620 5910
rect 8680 5850 9020 5910
rect 10810 5850 10820 5910
rect 10880 5850 11220 5910
rect 13010 5850 13020 5910
rect 13080 5850 13420 5910
rect 15210 5850 15440 5910
rect 15500 5850 15620 5910
rect 17410 5850 17640 5910
rect 17700 5850 17820 5910
rect 27260 5902 27380 5948
rect 27370 5885 27380 5902
rect 27440 5948 27450 5975
rect 28770 5970 28810 6200
rect 29000 6040 29080 6050
rect 29000 5970 29010 6040
rect 27440 5902 27950 5948
rect 27440 5885 27450 5902
rect 27370 5875 27450 5885
rect 28760 5860 29010 5970
rect 2500 5810 4020 5822
rect 2500 5750 2510 5810
rect 4010 5750 4020 5810
rect 2500 5740 4020 5750
rect 4700 5810 6220 5822
rect 4700 5750 4710 5810
rect 6210 5750 6220 5810
rect 4700 5740 6220 5750
rect 6900 5810 8420 5822
rect 6900 5750 6910 5810
rect 8410 5750 8420 5810
rect 6900 5740 8420 5750
rect 9100 5810 10620 5822
rect 9100 5750 9110 5810
rect 10610 5750 10620 5810
rect 9100 5740 10620 5750
rect 11300 5810 12820 5822
rect 11300 5750 11310 5810
rect 12810 5750 12820 5810
rect 11300 5740 12820 5750
rect 13500 5810 15020 5822
rect 13500 5750 13510 5810
rect 15010 5750 15020 5810
rect 13500 5740 15020 5750
rect 15700 5810 17220 5822
rect 15700 5750 15710 5810
rect 17210 5750 17220 5810
rect 15700 5740 17220 5750
rect 17900 5810 19420 5822
rect 17900 5750 17910 5810
rect 19410 5750 19420 5810
rect 27490 5815 27570 5825
rect 27490 5790 27500 5815
rect 17900 5740 19420 5750
rect 27260 5744 27500 5790
rect 27490 5725 27500 5744
rect 27560 5790 27570 5815
rect 27560 5744 27950 5790
rect 27560 5725 27570 5744
rect 27490 5715 27570 5725
rect 27370 5660 27450 5670
rect 2500 5580 2510 5640
rect 2690 5580 2700 5640
rect 2500 5340 2700 5580
rect 3160 5580 3170 5640
rect 3350 5580 3360 5640
rect 3160 5340 3360 5580
rect 3820 5580 3830 5640
rect 4010 5580 4020 5640
rect 3820 5340 4020 5580
rect 4700 5580 4710 5640
rect 4890 5580 4900 5640
rect 4700 5340 4900 5580
rect 5360 5580 5370 5640
rect 5550 5580 5560 5640
rect 5360 5340 5560 5580
rect 6020 5580 6030 5640
rect 6210 5580 6220 5640
rect 6020 5340 6220 5580
rect 6900 5500 7100 5640
rect 6900 5440 6910 5500
rect 7090 5440 7100 5500
rect 6900 5340 7100 5440
rect 7560 5500 7760 5640
rect 7560 5440 7570 5500
rect 7750 5440 7760 5500
rect 7560 5340 7760 5440
rect 8220 5500 8420 5640
rect 8220 5440 8230 5500
rect 8410 5440 8420 5500
rect 8220 5340 8420 5440
rect 9100 5500 9300 5640
rect 9100 5440 9110 5500
rect 9290 5440 9300 5500
rect 9100 5340 9300 5440
rect 9760 5500 9960 5640
rect 9760 5440 9770 5500
rect 9950 5440 9960 5500
rect 9760 5340 9960 5440
rect 10420 5500 10620 5640
rect 10420 5440 10430 5500
rect 10610 5440 10620 5500
rect 10420 5340 10620 5440
rect 11300 5500 11500 5640
rect 11300 5440 11310 5500
rect 11490 5440 11500 5500
rect 11300 5340 11500 5440
rect 11960 5500 12160 5640
rect 11960 5440 11970 5500
rect 12150 5440 12160 5500
rect 11960 5340 12160 5440
rect 12620 5500 12820 5640
rect 12620 5440 12630 5500
rect 12810 5440 12820 5500
rect 12620 5340 12820 5440
rect 13500 5500 13700 5640
rect 13500 5440 13510 5500
rect 13690 5440 13700 5500
rect 13500 5340 13700 5440
rect 14160 5500 14360 5640
rect 14160 5440 14170 5500
rect 14350 5440 14360 5500
rect 14160 5340 14360 5440
rect 14820 5500 15020 5640
rect 14820 5440 14830 5500
rect 15010 5440 15020 5500
rect 14820 5340 15020 5440
rect 15700 5580 15710 5640
rect 15890 5580 15900 5640
rect 15700 5340 15900 5580
rect 16360 5580 16370 5640
rect 16550 5580 16560 5640
rect 16360 5340 16560 5580
rect 17020 5580 17030 5640
rect 17210 5580 17220 5640
rect 17020 5340 17220 5580
rect 17900 5580 17910 5640
rect 18090 5580 18100 5640
rect 17900 5340 18100 5580
rect 18560 5580 18570 5640
rect 18750 5580 18760 5640
rect 18560 5340 18760 5580
rect 19220 5580 19230 5640
rect 19410 5580 19420 5640
rect 27370 5632 27380 5660
rect 27260 5586 27380 5632
rect 19220 5340 19420 5580
rect 27370 5570 27380 5586
rect 27440 5632 27450 5660
rect 28770 5650 28810 5860
rect 29000 5820 29010 5860
rect 29070 5820 29080 6040
rect 29000 5810 29080 5820
rect 27440 5586 27950 5632
rect 27440 5570 27450 5586
rect 27370 5560 27450 5570
rect 29540 5580 29900 6360
rect 29540 5500 29670 5580
rect 30280 5560 30400 6720
rect 27920 5340 29670 5500
rect -90 5330 10 5340
rect -90 5270 -70 5330
rect -10 5270 10 5330
rect -90 5260 10 5270
rect 2110 5330 2210 5340
rect 2110 5270 2130 5330
rect 2190 5270 2210 5330
rect 2110 5260 2210 5270
rect 4310 5330 4410 5340
rect 4310 5270 4330 5330
rect 4390 5270 4410 5330
rect 4310 5260 4410 5270
rect 6510 5330 6610 5340
rect 6510 5270 6530 5330
rect 6590 5270 6610 5330
rect 6510 5260 6610 5270
rect 8710 5330 8810 5340
rect 8710 5270 8730 5330
rect 8790 5270 8810 5330
rect 8710 5260 8810 5270
rect 10910 5330 11010 5340
rect 10910 5270 10930 5330
rect 10990 5270 11010 5330
rect 10910 5260 11010 5270
rect 13110 5330 13210 5340
rect 13110 5270 13130 5330
rect 13190 5270 13210 5330
rect 13110 5260 13210 5270
rect 15310 5330 15410 5340
rect 15310 5270 15330 5330
rect 15390 5270 15410 5330
rect 15310 5260 15410 5270
rect 17510 5330 17610 5340
rect 17510 5270 17530 5330
rect 17590 5270 17610 5330
rect 17510 5260 17610 5270
rect 19710 5330 19810 5340
rect 19710 5270 19730 5330
rect 19790 5270 19810 5330
rect 19710 5260 19810 5270
rect 21910 5330 22010 5340
rect 21910 5270 21930 5330
rect 21990 5270 22010 5330
rect 21910 5260 22010 5270
rect 27170 5240 28750 5250
rect 4100 5160 4220 5220
rect 4280 5160 4510 5220
rect 6300 5160 6420 5220
rect 6480 5160 6710 5220
rect 8500 5160 8840 5220
rect 8900 5160 8910 5220
rect 10700 5160 11040 5220
rect 11100 5160 11110 5220
rect 12900 5160 13240 5220
rect 13300 5160 13310 5220
rect 15100 5160 15440 5220
rect 15500 5160 15510 5220
rect 17300 5160 17420 5220
rect 17480 5160 17710 5220
rect 19500 5140 19620 5200
rect 19680 5140 19910 5200
rect 27170 5110 27180 5240
rect 27310 5190 28750 5240
rect 27310 5110 27950 5190
rect 28920 5150 29020 5340
rect 2010 5050 2020 5110
rect 2080 5050 2420 5110
rect 4210 5050 4220 5110
rect 4280 5050 4620 5110
rect 6410 5050 6640 5110
rect 6700 5050 6820 5110
rect 8610 5050 8840 5110
rect 8900 5050 9020 5110
rect 10810 5050 11040 5110
rect 11100 5050 11220 5110
rect 13010 5050 13240 5110
rect 13300 5050 13420 5110
rect 15210 5050 15220 5110
rect 15280 5050 15620 5110
rect 17410 5050 17420 5110
rect 17480 5050 17820 5110
rect 27170 5100 27950 5110
rect 2500 5010 4020 5022
rect 2500 4950 2510 5010
rect 4010 4950 4020 5010
rect 2500 4940 4020 4950
rect 4700 5010 6220 5022
rect 4700 4950 4710 5010
rect 6210 4950 6220 5010
rect 4700 4940 6220 4950
rect 6900 5010 8420 5022
rect 6900 4950 6910 5010
rect 8410 4950 8420 5010
rect 6900 4940 8420 4950
rect 9100 5010 10620 5022
rect 9100 4950 9110 5010
rect 10610 4950 10620 5010
rect 9100 4940 10620 4950
rect 11300 5010 12820 5022
rect 11300 4950 11310 5010
rect 12810 4950 12820 5010
rect 11300 4940 12820 4950
rect 13500 5010 15020 5022
rect 13500 4950 13510 5010
rect 15010 4950 15020 5010
rect 13500 4940 15020 4950
rect 15700 5010 17220 5022
rect 15700 4950 15710 5010
rect 17210 4950 17220 5010
rect 15700 4940 17220 4950
rect 17900 5010 19420 5022
rect 17900 4950 17910 5010
rect 19410 4950 19420 5010
rect 17900 4940 19420 4950
rect 23040 4970 23590 4980
rect 7790 4680 7950 4690
rect 7790 4540 7800 4680
rect 7940 4660 7950 4680
rect 7940 4560 12840 4660
rect 23040 4600 23050 4970
rect 23580 4600 23590 4970
rect 23040 4590 23590 4600
rect 23710 4590 24900 4980
rect 25040 4590 26230 4980
rect 7940 4540 7950 4560
rect 7790 4530 7950 4540
rect 10700 4360 10820 4420
rect 10880 4360 11110 4420
rect 12900 4360 13240 4420
rect 13300 4360 13310 4420
rect 27880 4320 27950 5100
rect 28780 4360 29020 5150
rect 29540 4760 29670 5340
rect 30720 5220 30820 6680
rect 31140 5560 31260 6720
rect 31700 6660 32020 7280
rect 36410 7480 36572 7670
rect 36870 7600 37010 7800
rect 37520 7750 37620 8180
rect 37140 7670 37620 7750
rect 37520 7630 37620 7670
rect 37480 7620 37620 7630
rect 37480 7504 37494 7620
rect 37610 7504 37620 7620
rect 37480 7500 37620 7504
rect 37480 7490 37640 7500
rect 36410 7440 36690 7480
rect 36410 7200 36572 7440
rect 37500 7370 37510 7490
rect 37630 7370 37640 7490
rect 37500 7360 37640 7370
rect 36106 7176 36838 7200
rect 36106 6982 36128 7176
rect 36810 6982 36838 7176
rect 36106 6964 36838 6982
rect 36410 6958 36572 6964
rect 31620 5580 32020 6660
rect 36220 6260 36420 6270
rect 36220 6200 36230 6260
rect 29860 5120 31680 5220
rect 29740 5040 29800 5080
rect 31740 5040 31800 5080
rect 29740 4960 30740 5040
rect 30820 4960 31800 5040
rect 8610 4250 8620 4310
rect 8680 4250 9026 4310
rect 10810 4250 11040 4310
rect 11100 4250 11226 4310
rect 27880 4260 28750 4320
rect 28920 4300 29020 4360
rect 9080 4100 12840 4200
rect 10880 3960 10890 4100
rect 11030 3960 11040 4100
rect 10880 3950 11040 3960
rect 29740 3980 29800 4960
rect 29880 4870 30650 4880
rect 29880 4800 30520 4870
rect 30510 4750 30520 4800
rect 30640 4750 30650 4870
rect 30510 4740 30650 4750
rect 30900 4870 31660 4880
rect 30900 4750 30910 4870
rect 31030 4800 31660 4870
rect 31030 4750 31040 4800
rect 30900 4740 31040 4750
rect 31740 4050 31800 4960
rect 31890 4790 32020 5580
rect 31900 4760 32020 4790
rect 36060 6080 36230 6200
rect 36410 6080 36420 6260
rect 36060 6000 36420 6080
rect 36520 6260 36720 6270
rect 36520 6080 36530 6260
rect 36710 6220 36720 6260
rect 36710 6110 38010 6220
rect 36710 6080 36720 6110
rect 36520 6070 36720 6080
rect 37420 6000 38010 6110
rect 36060 5970 36840 6000
rect 37240 5970 38010 6000
rect 36060 5480 36140 5970
rect 36380 5900 36910 5920
rect 36290 5890 36910 5900
rect 36290 5820 36300 5890
rect 36390 5820 36910 5890
rect 36290 5810 36910 5820
rect 36380 5790 36910 5810
rect 37000 5740 37080 5960
rect 37170 5900 37700 5920
rect 37170 5890 37780 5900
rect 37170 5820 37680 5890
rect 37770 5820 37780 5890
rect 37170 5810 37780 5820
rect 37170 5790 37700 5810
rect 36460 5710 37630 5740
rect 36380 5640 36910 5660
rect 36290 5630 36910 5640
rect 36290 5560 36300 5630
rect 36390 5560 36910 5630
rect 36290 5550 36910 5560
rect 36380 5530 36910 5550
rect 36060 5450 36840 5480
rect 36060 4970 36140 5450
rect 36380 5380 36910 5400
rect 36290 5370 36910 5380
rect 36290 5300 36300 5370
rect 36390 5300 36910 5370
rect 36290 5290 36910 5300
rect 36380 5270 36910 5290
rect 37000 5220 37080 5710
rect 37170 5640 37710 5660
rect 37170 5630 37780 5640
rect 37170 5560 37680 5630
rect 37770 5560 37780 5630
rect 37170 5550 37780 5560
rect 37170 5530 37710 5550
rect 37930 5480 38010 5970
rect 37240 5450 38010 5480
rect 37170 5380 37700 5400
rect 37170 5370 37780 5380
rect 37170 5300 37680 5370
rect 37770 5300 37780 5370
rect 37170 5290 37780 5300
rect 37170 5270 37700 5290
rect 36460 5190 37630 5220
rect 36380 5120 36910 5140
rect 36290 5110 36910 5120
rect 36290 5040 36300 5110
rect 36390 5040 36910 5110
rect 36290 5030 36910 5040
rect 36380 5010 36910 5030
rect 36060 4940 36850 4970
rect 36060 4450 36140 4940
rect 36380 4860 36910 4890
rect 36290 4850 36910 4860
rect 36290 4780 36300 4850
rect 36390 4780 36910 4850
rect 36290 4770 36910 4780
rect 36380 4760 36910 4770
rect 37000 4710 37080 5190
rect 37170 5120 37700 5140
rect 37170 5110 37780 5120
rect 37170 5040 37680 5110
rect 37770 5040 37780 5110
rect 37170 5030 37780 5040
rect 37170 5010 37700 5030
rect 37930 4970 38010 5450
rect 37240 4940 38010 4970
rect 37170 4860 37700 4890
rect 37170 4850 37780 4860
rect 37170 4780 37680 4850
rect 37770 4780 37780 4850
rect 37170 4770 37780 4780
rect 37170 4760 37700 4770
rect 36460 4680 37630 4710
rect 36380 4600 36910 4630
rect 36290 4590 36910 4600
rect 36290 4520 36300 4590
rect 36390 4520 36910 4590
rect 36290 4510 36910 4520
rect 36380 4500 36910 4510
rect 36060 4420 36850 4450
rect 32240 4130 34160 4240
rect 30070 4040 30270 4050
rect 30070 3980 30080 4040
rect 29740 3920 30080 3980
rect 30070 3860 30080 3920
rect 30260 3860 30270 4040
rect 30070 3850 30270 3860
rect 31670 4040 31870 4050
rect 31670 3860 31680 4040
rect 31860 3860 31870 4040
rect 31670 3850 31870 3860
rect 17150 3360 18160 3410
rect 18110 3020 18160 3360
rect 32240 3280 32760 4130
rect 32800 4070 32990 4080
rect 32800 4036 32810 4070
rect 32790 4010 32810 4036
rect 32980 4036 32990 4070
rect 32980 4010 33004 4036
rect 32790 3990 33004 4010
rect 32790 3480 32846 3990
rect 32880 3440 32914 3946
rect 32948 3480 33004 3990
rect 33038 3558 33072 4128
rect 33120 4070 33310 4080
rect 33120 4036 33130 4070
rect 33106 4010 33130 4036
rect 33300 4036 33310 4070
rect 33300 4010 33320 4036
rect 33106 3990 33320 4010
rect 33106 3480 33162 3990
rect 33196 3440 33230 3946
rect 33264 3480 33320 3990
rect 33354 3558 33388 4130
rect 33430 4070 33620 4080
rect 33430 4036 33440 4070
rect 33422 4010 33440 4036
rect 33610 4036 33620 4070
rect 33610 4010 33636 4036
rect 33422 3990 33636 4010
rect 33422 3480 33478 3990
rect 33512 3440 33546 3946
rect 33580 3480 33636 3990
rect 33670 3558 33704 4130
rect 33960 4120 34160 4130
rect 33750 4070 33940 4080
rect 33750 4036 33760 4070
rect 33738 4010 33760 4036
rect 33930 4036 33940 4070
rect 33930 4010 33952 4036
rect 33738 3990 33952 4010
rect 33738 3480 33794 3990
rect 33828 3440 33862 3946
rect 33896 3480 33952 3990
rect 33990 3560 34160 4120
rect 34740 4140 35740 4240
rect 34740 3958 34800 4140
rect 34860 4090 35200 4100
rect 34860 4010 34870 4090
rect 35190 4010 35200 4090
rect 34860 4000 35200 4010
rect 34980 3992 35194 4000
rect 34740 3560 34950 3958
rect 33990 3558 34950 3560
rect 32840 3430 33880 3440
rect 32840 3350 32850 3430
rect 33870 3350 33880 3430
rect 32840 3340 33880 3350
rect 32240 3244 32880 3280
rect 33990 3250 34800 3558
rect 34980 3482 35036 3992
rect 35070 3440 35104 3946
rect 35138 3526 35194 3992
rect 35228 3570 35262 4140
rect 35296 3526 35352 4034
rect 35138 3480 35352 3526
rect 35386 3440 35420 3946
rect 35060 3430 35420 3440
rect 35060 3350 35070 3430
rect 35410 3350 35420 3430
rect 35060 3340 35420 3350
rect 35540 3340 35740 4140
rect 36060 3930 36140 4420
rect 36380 4340 36910 4370
rect 36290 4330 36910 4340
rect 36290 4260 36300 4330
rect 36390 4260 36910 4330
rect 36290 4250 36910 4260
rect 36380 4240 36910 4250
rect 37000 4190 37080 4680
rect 37170 4600 37700 4630
rect 37170 4590 37780 4600
rect 37170 4520 37680 4590
rect 37770 4520 37780 4590
rect 37170 4510 37780 4520
rect 37170 4500 37700 4510
rect 37930 4450 38010 4940
rect 37240 4420 38010 4450
rect 37170 4340 37700 4370
rect 37170 4330 37780 4340
rect 37170 4260 37680 4330
rect 37770 4260 37780 4330
rect 37170 4250 37780 4260
rect 37170 4240 37700 4250
rect 36460 4160 37630 4190
rect 36380 4080 36910 4110
rect 36290 4070 36910 4080
rect 36290 4000 36300 4070
rect 36390 4000 36910 4070
rect 36290 3990 36910 4000
rect 36380 3980 36910 3990
rect 36060 3900 36840 3930
rect 36060 3860 36140 3900
rect 36370 3580 36530 3590
rect 36370 3440 36380 3580
rect 36520 3560 36530 3580
rect 37000 3560 37080 4160
rect 37170 4080 37700 4110
rect 37170 4070 37780 4080
rect 37170 4000 37680 4070
rect 37770 4000 37780 4070
rect 37170 3990 37780 4000
rect 37170 3980 37700 3990
rect 37930 3930 38010 4420
rect 37240 3900 38010 3930
rect 37930 3860 38010 3900
rect 36520 3460 37080 3560
rect 36520 3440 36530 3460
rect 36370 3430 36530 3440
rect 35540 3260 36200 3340
rect 33980 3244 34800 3250
rect 32240 3198 32882 3244
rect 32240 3028 32348 3198
rect 32460 3156 32674 3162
rect 32460 3106 32466 3156
rect 32459 3068 32466 3106
rect 32668 3106 32674 3156
rect 32668 3068 32675 3106
rect 32459 3062 32675 3068
rect 32459 3060 32517 3062
rect 32617 3060 32675 3062
rect 18050 3010 18210 3020
rect 7800 2500 7940 2900
rect 18050 2870 18060 3010
rect 18200 2870 18210 3010
rect 18050 2860 18210 2870
rect 16900 2780 17140 2790
rect 16900 2640 16910 2780
rect 17130 2640 17140 2780
rect 16900 2630 17140 2640
rect 17370 2780 17500 2790
rect 17370 2640 17380 2780
rect 17490 2640 17500 2780
rect 17370 2630 17500 2640
rect 17730 2780 17970 2790
rect 17730 2640 17740 2780
rect 17960 2640 17970 2780
rect 17730 2630 17970 2640
rect 32240 2628 32432 3028
rect -140 2480 14240 2500
rect 17260 2480 17300 2610
rect 17570 2480 17610 2620
rect 32240 2480 32392 2628
rect 32460 2596 32516 3060
rect 32544 2628 32590 3028
rect 32459 2550 32517 2596
rect 32548 2520 32586 2628
rect 32618 2596 32674 3060
rect 32786 3028 32882 3198
rect 32702 2760 32882 3028
rect 33852 3220 34800 3244
rect 33852 3198 34680 3220
rect 33852 3028 33948 3198
rect 34060 3156 34274 3162
rect 34060 3106 34066 3156
rect 34059 3068 34066 3106
rect 34268 3106 34274 3156
rect 34268 3068 34275 3106
rect 34059 3062 34275 3068
rect 34059 3060 34117 3062
rect 34217 3060 34275 3062
rect 33852 2760 34032 3028
rect 32702 2628 34032 2760
rect 32617 2550 32675 2596
rect -140 2380 32392 2480
rect 32440 2510 32700 2520
rect 32440 2430 32450 2510
rect 32690 2430 32700 2510
rect 32440 2420 32700 2430
rect 32742 2380 33992 2628
rect 34060 2596 34116 3060
rect 34144 2628 34190 3028
rect 34059 2550 34117 2596
rect 34148 2520 34186 2628
rect 34218 2596 34274 3060
rect 34386 3028 34680 3198
rect 34302 2628 34680 3028
rect 34217 2550 34275 2596
rect 34040 2510 34300 2520
rect 34040 2430 34050 2510
rect 34290 2430 34300 2510
rect 34040 2420 34300 2430
rect 34342 2380 34680 2628
rect 35360 3198 36200 3260
rect 35360 3028 35548 3198
rect 35660 3156 35874 3162
rect 35660 3068 35666 3156
rect 35868 3068 35874 3156
rect 35660 3062 35874 3068
rect 35360 2628 35632 3028
rect 35360 2380 35592 2628
rect 35660 2552 35716 3062
rect 35748 2520 35786 3026
rect 35818 2552 35874 3062
rect 35986 3028 36200 3198
rect 35902 2628 36200 3028
rect 35640 2510 35900 2520
rect 35640 2430 35650 2510
rect 35890 2430 35900 2510
rect 35640 2420 35900 2430
rect 35942 2380 36200 2628
rect -140 2220 37880 2380
rect -140 2060 480 2220
rect -140 460 0 2060
rect 440 460 480 2060
rect -140 260 480 460
rect -140 -1340 0 260
rect 440 -1340 480 260
rect -140 -1540 480 -1340
rect -140 -3140 0 -1540
rect 440 -3140 480 -1540
rect -140 -3340 480 -3140
rect -140 -4680 0 -3340
rect 440 -4780 480 -3340
rect 660 2180 37880 2220
rect 660 2060 11160 2180
rect 11240 2060 12300 2140
rect 12380 2060 12760 2180
rect 12840 2060 13900 2140
rect 13980 2100 31780 2180
rect 13980 2060 14870 2100
rect 15070 2060 31780 2100
rect 32060 2130 34680 2140
rect 32060 2070 32450 2130
rect 32690 2070 34050 2130
rect 34290 2070 34680 2130
rect 32060 2060 34680 2070
rect 35270 2130 36270 2140
rect 35270 2070 35650 2130
rect 35890 2070 36270 2130
rect 35270 2060 36270 2070
rect 36760 2060 37880 2180
rect 660 460 710 2060
rect 32200 2055 32459 2060
rect 32677 2055 32940 2060
rect 33800 2055 34059 2060
rect 34277 2055 34540 2060
rect 2100 1990 2240 2000
rect 2100 1310 2110 1990
rect 2230 1310 2240 1990
rect 2100 1300 2240 1310
rect 3700 1990 3840 2000
rect 3700 1310 3710 1990
rect 3830 1310 3840 1990
rect 3700 1300 3840 1310
rect 5300 1990 5440 2000
rect 5300 1310 5310 1990
rect 5430 1310 5440 1990
rect 5300 1300 5440 1310
rect 6900 1990 7040 2000
rect 6900 1310 6910 1990
rect 7030 1310 7040 1990
rect 6900 1300 7040 1310
rect 8500 1990 8640 2000
rect 8500 1310 8510 1990
rect 8630 1310 8640 1990
rect 8500 1300 8640 1310
rect 10100 1990 10240 2000
rect 10100 1310 10110 1990
rect 10230 1310 10240 1990
rect 11020 1950 11220 1960
rect 11020 1330 11030 1950
rect 11150 1330 11220 1950
rect 11020 1320 11220 1330
rect 10100 1300 10240 1310
rect 11700 1300 11840 2000
rect 12310 1950 12820 1960
rect 12310 1330 12610 1950
rect 12730 1330 12820 1950
rect 12310 1320 12820 1330
rect 13300 1300 13440 2000
rect 14900 1980 15040 2010
rect 13910 1950 14120 1960
rect 13910 1330 13990 1950
rect 14110 1330 14120 1950
rect 13910 1240 14120 1330
rect 14900 1320 14910 1980
rect 15030 1320 15040 1980
rect 14900 1240 15040 1320
rect 16500 1990 16640 2000
rect 16500 1310 16510 1990
rect 16630 1310 16640 1990
rect 16500 1300 16640 1310
rect 18100 1990 18240 2000
rect 18100 1310 18110 1990
rect 18230 1310 18240 1990
rect 18100 1300 18240 1310
rect 19700 1990 19840 2000
rect 19700 1310 19710 1990
rect 19830 1310 19840 1990
rect 19700 1300 19840 1310
rect 21300 1990 21440 2000
rect 21300 1310 21310 1990
rect 21430 1310 21440 1990
rect 21300 1300 21440 1310
rect 22900 1990 23040 2000
rect 22900 1310 22910 1990
rect 23030 1310 23040 1990
rect 22900 1300 23040 1310
rect 24500 1990 24640 2000
rect 24500 1310 24510 1990
rect 24630 1310 24640 1990
rect 24500 1300 24640 1310
rect 26100 1990 26240 2000
rect 26100 1310 26110 1990
rect 26230 1310 26240 1990
rect 26100 1300 26240 1310
rect 27700 1990 27840 2000
rect 27700 1310 27710 1990
rect 27830 1310 27840 1990
rect 27700 1300 27840 1310
rect 28781 1995 28827 2007
rect 28781 1303 28787 1995
rect 28821 1303 28827 1995
rect 28781 1291 28827 1303
rect 29291 2000 29337 2007
rect 29399 2000 29445 2007
rect 29291 1995 29445 2000
rect 29291 1303 29297 1995
rect 29331 1990 29405 1995
rect 29331 1303 29405 1310
rect 29439 1303 29445 1995
rect 29291 1300 29445 1303
rect 29291 1291 29337 1300
rect 29399 1291 29445 1300
rect 29909 1995 29955 2007
rect 29909 1303 29915 1995
rect 29949 1303 29955 1995
rect 29909 1291 29955 1303
rect 30381 1995 30427 2007
rect 30381 1303 30387 1995
rect 30421 1303 30427 1995
rect 30381 1291 30427 1303
rect 30891 2000 30937 2007
rect 30999 2000 31045 2007
rect 30891 1995 31045 2000
rect 30891 1303 30897 1995
rect 30931 1990 31005 1995
rect 30931 1303 31005 1310
rect 31039 1303 31045 1995
rect 30891 1300 31045 1303
rect 30891 1291 30937 1300
rect 30999 1291 31045 1300
rect 31509 1995 31555 2007
rect 32500 1995 32640 2000
rect 34100 1995 34240 2000
rect 35700 1995 35840 2000
rect 31509 1303 31515 1995
rect 31549 1303 31555 1995
rect 32531 1990 32605 1995
rect 32531 1303 32605 1310
rect 32639 1303 32640 1995
rect 34131 1990 34205 1995
rect 34131 1303 34205 1310
rect 34239 1303 34240 1995
rect 35731 1990 35805 1995
rect 35731 1303 35805 1310
rect 35839 1303 35840 1995
rect 31509 1291 31555 1303
rect 32500 1300 32640 1303
rect 34100 1300 34240 1303
rect 35700 1300 35840 1303
rect 37300 1990 37440 2000
rect 37300 1310 37310 1990
rect 37430 1310 37440 1990
rect 37300 1300 37440 1310
rect 11240 1230 11680 1240
rect 1680 1160 2040 1220
rect 2300 1160 2660 1220
rect 3280 1160 3640 1220
rect 3900 1160 4260 1220
rect 4880 1160 5240 1220
rect 5500 1160 5860 1220
rect 6480 1160 6840 1220
rect 7100 1160 7460 1220
rect 8080 1160 8440 1220
rect 8700 1160 9060 1220
rect 9680 1160 10040 1220
rect 10300 1160 10660 1220
rect 1400 1150 10660 1160
rect 1400 1030 1410 1150
rect 1530 1030 3010 1150
rect 3130 1030 4610 1150
rect 4730 1030 6210 1150
rect 6330 1030 7810 1150
rect 7930 1030 9410 1150
rect 9530 1030 10660 1150
rect 11240 1070 11250 1230
rect 11670 1070 11680 1230
rect 11860 1120 13280 1240
rect 13480 1120 14120 1240
rect 14460 1150 15480 1240
rect 16059 1237 16459 1243
rect 16059 1203 16071 1237
rect 16080 1203 16440 1220
rect 16447 1203 16459 1237
rect 16059 1197 16459 1203
rect 16677 1237 17077 1243
rect 16677 1203 16689 1237
rect 16700 1203 17060 1220
rect 17065 1203 17077 1237
rect 16677 1197 17077 1203
rect 17659 1237 18059 1243
rect 17659 1203 17671 1237
rect 17680 1203 18040 1220
rect 18047 1203 18059 1237
rect 17659 1197 18059 1203
rect 18277 1237 18677 1243
rect 18277 1203 18289 1237
rect 18300 1203 18660 1220
rect 18665 1203 18677 1237
rect 18277 1197 18677 1203
rect 19259 1237 19659 1243
rect 19259 1203 19271 1237
rect 19280 1203 19640 1220
rect 19647 1203 19659 1237
rect 19259 1197 19659 1203
rect 19877 1237 20277 1243
rect 19877 1203 19889 1237
rect 19900 1203 20260 1220
rect 20265 1203 20277 1237
rect 19877 1197 20277 1203
rect 20859 1237 21259 1243
rect 20859 1203 20871 1237
rect 20880 1203 21240 1220
rect 21247 1203 21259 1237
rect 20859 1197 21259 1203
rect 21477 1237 21877 1243
rect 21477 1203 21489 1237
rect 21500 1203 21860 1220
rect 21865 1203 21877 1237
rect 21477 1197 21877 1203
rect 22459 1237 22859 1243
rect 22459 1203 22471 1237
rect 22480 1203 22840 1220
rect 22847 1203 22859 1237
rect 22459 1197 22859 1203
rect 23077 1237 23477 1243
rect 23077 1203 23089 1237
rect 23100 1203 23460 1220
rect 23465 1203 23477 1237
rect 23077 1197 23477 1203
rect 24059 1237 24459 1243
rect 24059 1203 24071 1237
rect 24080 1203 24440 1220
rect 24447 1203 24459 1237
rect 24059 1197 24459 1203
rect 24677 1237 25077 1243
rect 24677 1203 24689 1237
rect 24700 1203 25060 1220
rect 25065 1203 25077 1237
rect 24677 1197 25077 1203
rect 25659 1237 26059 1243
rect 25659 1203 25671 1237
rect 25680 1203 26040 1220
rect 26047 1203 26059 1237
rect 25659 1197 26059 1203
rect 26277 1237 26677 1243
rect 26277 1203 26289 1237
rect 26300 1203 26660 1220
rect 26665 1203 26677 1237
rect 26277 1197 26677 1203
rect 27259 1237 27659 1243
rect 27259 1203 27271 1237
rect 27280 1203 27640 1220
rect 27647 1203 27659 1237
rect 27259 1197 27659 1203
rect 27877 1237 28277 1243
rect 27877 1203 27889 1237
rect 27900 1203 28260 1220
rect 28265 1203 28277 1237
rect 27877 1197 28277 1203
rect 28859 1237 29259 1243
rect 28859 1203 28871 1237
rect 28880 1203 29240 1220
rect 29247 1203 29259 1237
rect 28859 1197 29259 1203
rect 29477 1237 29877 1243
rect 29477 1203 29489 1237
rect 29500 1203 29860 1220
rect 29865 1203 29877 1237
rect 29477 1197 29877 1203
rect 30459 1237 30859 1243
rect 30459 1203 30471 1237
rect 30480 1203 30840 1220
rect 30847 1203 30859 1237
rect 30459 1197 30859 1203
rect 31077 1237 31477 1243
rect 31077 1203 31089 1237
rect 31100 1203 31460 1220
rect 31465 1203 31477 1237
rect 31077 1197 31477 1203
rect 32060 1237 32459 1240
rect 32060 1203 32071 1237
rect 32080 1203 32440 1220
rect 32447 1203 32459 1237
rect 32060 1197 32459 1203
rect 32677 1237 33077 1243
rect 32677 1203 32689 1237
rect 32700 1203 33060 1220
rect 33065 1203 33077 1237
rect 32677 1197 33077 1203
rect 33659 1237 34059 1243
rect 33659 1203 33671 1237
rect 33680 1203 34040 1220
rect 34047 1203 34059 1237
rect 33659 1197 34059 1203
rect 34277 1237 34677 1243
rect 34277 1203 34289 1237
rect 34300 1203 34660 1220
rect 34665 1203 34677 1237
rect 34277 1197 34677 1203
rect 35259 1237 35659 1243
rect 35259 1203 35271 1237
rect 35280 1203 35640 1220
rect 35647 1203 35659 1237
rect 35259 1197 35659 1203
rect 35877 1237 36277 1243
rect 35877 1203 35889 1237
rect 35900 1203 36260 1220
rect 36265 1203 36277 1237
rect 35877 1197 36277 1203
rect 16080 1160 16440 1197
rect 16700 1160 17060 1197
rect 17680 1160 18040 1197
rect 18300 1160 18660 1197
rect 19280 1160 19640 1197
rect 19900 1160 20260 1197
rect 20880 1160 21240 1197
rect 21500 1160 21860 1197
rect 22480 1160 22840 1197
rect 23100 1160 23460 1197
rect 24080 1160 24440 1197
rect 24700 1160 25060 1197
rect 25680 1160 26040 1197
rect 26300 1160 26660 1197
rect 27280 1160 27640 1197
rect 27900 1160 28260 1197
rect 28880 1160 29240 1197
rect 29500 1160 29860 1197
rect 30480 1160 30840 1197
rect 31100 1160 31460 1197
rect 32080 1160 32440 1197
rect 32700 1160 33060 1197
rect 33680 1160 34040 1197
rect 34300 1160 34660 1197
rect 35280 1160 35640 1197
rect 35900 1160 36260 1197
rect 15590 1150 17060 1160
rect 11240 1060 11680 1070
rect 1400 1020 10660 1030
rect 15590 1030 15600 1150
rect 15700 1030 17060 1150
rect 15590 1020 17060 1030
rect 17190 1150 18660 1160
rect 17190 1030 17200 1150
rect 17300 1030 18660 1150
rect 17190 1020 18660 1030
rect 18790 1150 20260 1160
rect 18790 1030 18800 1150
rect 18900 1030 20260 1150
rect 18790 1020 20260 1030
rect 20390 1150 21860 1160
rect 20390 1030 20400 1150
rect 20500 1030 21860 1150
rect 20390 1020 21860 1030
rect 21990 1150 23460 1160
rect 21990 1030 22000 1150
rect 22100 1030 23460 1150
rect 21990 1020 23460 1030
rect 23590 1150 25060 1160
rect 23590 1030 23600 1150
rect 23700 1030 25060 1150
rect 23590 1020 25060 1030
rect 25660 1150 28260 1160
rect 25660 1030 26800 1150
rect 26900 1030 28260 1150
rect 25660 1020 28260 1030
rect 28391 1150 31460 1160
rect 28391 1030 28400 1150
rect 28500 1030 31460 1150
rect 28391 1020 31460 1030
rect 32060 1020 34660 1160
rect 35260 1020 36260 1160
rect 1680 950 2040 1020
rect 2300 950 2660 1020
rect 3280 950 3640 1020
rect 3900 950 4260 1020
rect 4880 950 5240 1020
rect 5500 950 5860 1020
rect 6480 950 6840 1020
rect 7100 950 7460 1020
rect 8080 950 8440 1020
rect 8700 950 9060 1020
rect 9680 950 10040 1020
rect 10300 950 10660 1020
rect 16080 975 16440 1020
rect 16700 975 17060 1020
rect 17680 975 18040 1020
rect 18300 975 18660 1020
rect 19280 975 19640 1020
rect 19900 975 20260 1020
rect 20880 975 21240 1020
rect 21500 975 21860 1020
rect 22480 975 22840 1020
rect 23100 975 23460 1020
rect 24080 975 24440 1020
rect 24700 975 25060 1020
rect 25680 975 26040 1020
rect 26300 975 26660 1020
rect 27280 975 27640 1020
rect 27900 975 28260 1020
rect 28880 975 29240 1020
rect 29500 975 29860 1020
rect 30480 975 30840 1020
rect 31100 975 31460 1020
rect 32080 975 32440 1020
rect 32700 975 33060 1020
rect 33680 975 34040 1020
rect 34300 975 34660 1020
rect 35280 975 35640 1020
rect 35900 975 36260 1020
rect 16059 970 16459 975
rect 11420 870 11500 940
rect 12040 870 12120 940
rect 12320 870 12520 880
rect 13020 870 13100 940
rect 13640 870 13720 940
rect 14620 870 14700 940
rect 15240 870 15320 940
rect 16059 929 16460 970
rect 16677 929 17077 975
rect 17659 970 18059 975
rect 17659 929 18060 970
rect 18277 929 18677 975
rect 19259 970 19659 975
rect 19259 929 19660 970
rect 19877 929 20277 975
rect 20859 970 21259 975
rect 20859 929 21260 970
rect 21477 929 21877 975
rect 22459 970 22859 975
rect 22459 929 22860 970
rect 23077 929 23477 975
rect 24059 970 24459 975
rect 24059 929 24460 970
rect 24677 929 25077 975
rect 25659 970 26059 975
rect 25659 929 26060 970
rect 26277 929 26677 975
rect 27259 970 27659 975
rect 27259 929 27660 970
rect 27877 929 28277 975
rect 28859 970 29259 975
rect 28859 929 29260 970
rect 29477 929 29877 975
rect 30459 970 30859 975
rect 30459 929 30860 970
rect 31077 929 31477 975
rect 32060 970 32459 975
rect 16060 910 16460 929
rect 16680 920 17070 929
rect 16677 909 17077 920
rect 17660 910 18060 929
rect 18280 920 18670 929
rect 18277 909 18677 920
rect 19260 910 19660 929
rect 19880 920 20270 929
rect 19877 909 20277 920
rect 20860 910 21260 929
rect 21480 920 21870 929
rect 21477 909 21877 920
rect 22460 910 22860 929
rect 23080 920 23470 929
rect 23077 909 23477 920
rect 24060 910 24460 929
rect 24680 920 25070 929
rect 24677 909 25077 920
rect 25660 910 26060 929
rect 26280 920 26670 929
rect 26277 909 26677 920
rect 27260 910 27660 929
rect 27880 920 28270 929
rect 27877 909 28277 920
rect 28860 910 29260 929
rect 29480 920 29870 929
rect 29477 909 29877 920
rect 30460 910 30860 929
rect 31080 920 31470 929
rect 31077 909 31477 920
rect 32060 910 32460 970
rect 32677 940 33077 975
rect 33659 970 34059 975
rect 32680 920 33070 940
rect 33659 929 34060 970
rect 34277 929 34677 975
rect 35259 970 35659 975
rect 35259 929 35660 970
rect 35877 929 36277 975
rect 36870 930 37260 1230
rect 37480 930 37870 1230
rect 32677 909 33077 920
rect 33660 910 34060 929
rect 34280 920 34670 929
rect 34277 909 34677 920
rect 35260 910 35660 929
rect 35880 920 36270 929
rect 35877 909 36277 920
rect 1540 750 12390 870
rect 12510 750 37950 870
rect 1540 740 37950 750
rect 1180 680 1320 690
rect 2780 680 2920 690
rect 4380 680 4520 690
rect 5980 680 6120 690
rect 7580 680 7720 690
rect 9180 680 9320 690
rect 11420 680 11500 740
rect 12040 680 12120 740
rect 13020 680 13100 740
rect 13640 680 13720 740
rect 14620 680 14700 740
rect 15240 680 15320 740
rect 30459 691 30859 697
rect 30459 690 30471 691
rect 30847 690 30859 691
rect 31077 691 31477 697
rect 31077 690 31089 691
rect 31465 690 31477 691
rect 15810 680 15930 690
rect 17410 680 17530 690
rect 19010 680 19130 690
rect 20610 680 20730 690
rect 22210 680 22330 690
rect 23810 680 23930 690
rect 27010 680 27130 690
rect 28610 680 31520 690
rect 1180 560 1190 680
rect 1310 560 2790 680
rect 2910 560 4390 680
rect 4510 560 5990 680
rect 6110 560 7590 680
rect 7710 560 9190 680
rect 9310 560 10720 680
rect 15810 560 15820 680
rect 15920 560 17120 680
rect 17410 560 17420 680
rect 17520 560 18720 680
rect 19010 560 19020 680
rect 19120 560 20320 680
rect 20610 560 20620 680
rect 20720 560 21920 680
rect 22210 560 22220 680
rect 22320 560 23520 680
rect 23810 560 23820 680
rect 23920 560 25120 680
rect 25620 560 27020 680
rect 27120 560 28320 680
rect 28610 560 28620 680
rect 28720 560 31520 680
rect 1180 550 1320 560
rect 2780 550 2920 560
rect 4380 550 4520 560
rect 5980 550 6120 560
rect 7580 550 7720 560
rect 9180 550 9320 560
rect 15810 550 15930 560
rect 17410 550 17530 560
rect 19010 550 19130 560
rect 20610 550 20730 560
rect 22210 550 22330 560
rect 23810 550 23930 560
rect 27010 550 27130 560
rect 28610 550 31520 560
rect 31810 680 31930 690
rect 31810 560 31820 680
rect 31920 560 36270 680
rect 36590 670 36730 680
rect 31810 550 31930 560
rect 36590 550 36600 670
rect 36720 660 36730 670
rect 36870 660 37252 690
rect 36720 560 37252 660
rect 37480 660 37870 690
rect 37480 650 37980 660
rect 37480 560 37850 650
rect 36720 550 36730 560
rect 36590 540 36730 550
rect 37840 530 37850 560
rect 37970 530 37980 650
rect 37840 520 37980 530
rect 660 260 38060 460
rect 660 -1340 710 260
rect 2100 190 2240 200
rect 2100 -490 2110 190
rect 2230 -490 2240 190
rect 2100 -500 2240 -490
rect 3700 190 3840 200
rect 3700 -490 3710 190
rect 3830 -490 3840 190
rect 3700 -500 3840 -490
rect 5300 190 5440 200
rect 5300 -490 5310 190
rect 5430 -490 5440 190
rect 5300 -500 5440 -490
rect 6900 190 7040 200
rect 6900 -490 6910 190
rect 7030 -490 7040 190
rect 6900 -500 7040 -490
rect 8500 190 8640 200
rect 8500 -490 8510 190
rect 8630 -490 8640 190
rect 8500 -500 8640 -490
rect 10100 190 10240 200
rect 10100 -490 10110 190
rect 10230 -490 10240 190
rect 10100 -500 10240 -490
rect 11700 190 11840 200
rect 11700 -560 11710 190
rect 11260 -570 11710 -560
rect 11830 -560 11840 190
rect 13300 190 13440 200
rect 13300 -490 13310 190
rect 13430 -490 13440 190
rect 14900 190 15040 200
rect 13300 -500 13440 -490
rect 14380 -560 14430 -490
rect 14900 -560 14910 190
rect 11830 -570 12280 -560
rect 1680 -640 2040 -580
rect 2300 -640 2660 -580
rect 3280 -640 3640 -580
rect 3900 -640 4260 -580
rect 4880 -640 5240 -580
rect 5500 -640 5860 -580
rect 6480 -640 6840 -580
rect 7100 -640 7460 -580
rect 8080 -640 8440 -580
rect 8700 -640 9060 -580
rect 9680 -640 10040 -580
rect 10300 -640 10660 -580
rect 1400 -650 10660 -640
rect 1400 -770 1410 -650
rect 1530 -770 3010 -650
rect 3130 -770 4610 -650
rect 4730 -770 6210 -650
rect 6330 -770 7810 -650
rect 7930 -770 9410 -650
rect 9530 -770 10660 -650
rect 11260 -730 11270 -570
rect 12270 -730 12280 -570
rect 14380 -570 14910 -560
rect 15030 -560 15040 190
rect 16500 190 16640 200
rect 16500 -490 16510 190
rect 16630 -490 16640 190
rect 15510 -560 15560 -490
rect 16500 -500 16640 -490
rect 18100 190 18240 200
rect 18100 -490 18110 190
rect 18230 -490 18240 190
rect 18100 -500 18240 -490
rect 19700 190 19840 200
rect 19700 -490 19710 190
rect 19830 -490 19840 190
rect 19700 -500 19840 -490
rect 21300 190 21440 200
rect 21300 -490 21310 190
rect 21430 -490 21440 190
rect 21300 -500 21440 -490
rect 22900 190 23040 200
rect 22900 -490 22910 190
rect 23030 -490 23040 190
rect 22900 -500 23040 -490
rect 24500 190 24640 200
rect 24500 -490 24510 190
rect 24630 -490 24640 190
rect 24500 -500 24640 -490
rect 26100 190 26240 200
rect 26100 -490 26110 190
rect 26230 -490 26240 190
rect 26100 -500 26240 -490
rect 27700 190 27840 200
rect 27700 -490 27710 190
rect 27830 -490 27840 190
rect 27700 -500 27840 -490
rect 28781 195 28827 207
rect 28781 -497 28787 195
rect 28821 -497 28827 195
rect 28781 -509 28827 -497
rect 29291 200 29337 207
rect 29399 200 29445 207
rect 29291 195 29445 200
rect 29291 -497 29297 195
rect 29331 190 29405 195
rect 29331 -497 29405 -490
rect 29439 -497 29445 195
rect 29291 -500 29445 -497
rect 29291 -509 29337 -500
rect 29399 -509 29445 -500
rect 29909 195 29955 207
rect 29909 -497 29915 195
rect 29949 -497 29955 195
rect 29909 -509 29955 -497
rect 30381 195 30427 207
rect 30381 -497 30387 195
rect 30421 -497 30427 195
rect 30381 -509 30427 -497
rect 30891 200 30937 207
rect 30999 200 31045 207
rect 30891 195 31045 200
rect 30891 -497 30897 195
rect 30931 190 31005 195
rect 30931 -497 31005 -490
rect 31039 -497 31045 195
rect 30891 -500 31045 -497
rect 30891 -509 30937 -500
rect 30999 -509 31045 -500
rect 31509 195 31555 207
rect 32500 195 32640 200
rect 31509 -497 31515 195
rect 31549 -497 31555 195
rect 32531 190 32605 195
rect 32531 -497 32605 -490
rect 32639 -497 32640 195
rect 34100 190 34240 200
rect 35700 195 35840 200
rect 35731 190 35805 195
rect 34100 160 34110 190
rect 34230 160 34240 190
rect 34131 -497 34205 -490
rect 34239 -497 34240 160
rect 35731 -497 35805 -490
rect 35839 -497 35840 195
rect 31509 -509 31555 -497
rect 32500 -500 32640 -497
rect 34100 -500 34240 -497
rect 35700 -500 35840 -497
rect 15030 -570 15560 -560
rect 12880 -597 13240 -580
rect 13247 -597 13259 -580
rect 12880 -603 13259 -597
rect 13477 -597 13489 -580
rect 13500 -597 13860 -580
rect 13477 -603 13860 -597
rect 12880 -640 13240 -603
rect 13500 -640 13860 -603
rect 11260 -740 12280 -730
rect 12380 -650 14300 -640
rect 1400 -780 10660 -770
rect 1680 -850 2040 -780
rect 2300 -850 2660 -780
rect 3280 -850 3640 -780
rect 3900 -850 4260 -780
rect 4880 -850 5240 -780
rect 5500 -850 5860 -780
rect 6480 -850 6840 -780
rect 7100 -850 7460 -780
rect 8080 -850 8440 -780
rect 8700 -850 9060 -780
rect 9680 -850 10040 -780
rect 10300 -850 10660 -780
rect 12380 -810 12390 -650
rect 12510 -780 14300 -650
rect 14380 -730 14470 -570
rect 15470 -730 15560 -570
rect 16059 -563 16459 -557
rect 16059 -597 16071 -563
rect 16080 -597 16440 -580
rect 16447 -597 16459 -563
rect 16059 -603 16459 -597
rect 16677 -563 17077 -557
rect 16677 -597 16689 -563
rect 16700 -597 17060 -580
rect 17065 -597 17077 -563
rect 16677 -603 17077 -597
rect 17659 -563 18059 -557
rect 17659 -597 17671 -563
rect 17680 -597 18040 -580
rect 18047 -597 18059 -563
rect 17659 -603 18059 -597
rect 18277 -563 18677 -557
rect 18277 -597 18289 -563
rect 18300 -597 18660 -580
rect 18665 -597 18677 -563
rect 18277 -603 18677 -597
rect 19259 -563 19659 -557
rect 19259 -597 19271 -563
rect 19280 -597 19640 -580
rect 19647 -597 19659 -563
rect 19259 -603 19659 -597
rect 19877 -563 20277 -557
rect 19877 -597 19889 -563
rect 19900 -597 20260 -580
rect 20265 -597 20277 -563
rect 19877 -603 20277 -597
rect 20859 -563 21259 -557
rect 20859 -597 20871 -563
rect 20880 -597 21240 -580
rect 21247 -597 21259 -563
rect 20859 -603 21259 -597
rect 21477 -563 21877 -557
rect 21477 -597 21489 -563
rect 21500 -597 21860 -580
rect 21865 -597 21877 -563
rect 21477 -603 21877 -597
rect 22459 -563 22859 -557
rect 22459 -597 22471 -563
rect 22480 -597 22840 -580
rect 22847 -597 22859 -563
rect 22459 -603 22859 -597
rect 23077 -563 23477 -557
rect 23077 -597 23089 -563
rect 23100 -597 23460 -580
rect 23465 -597 23477 -563
rect 23077 -603 23477 -597
rect 24059 -563 24459 -557
rect 24059 -597 24071 -563
rect 24080 -597 24440 -580
rect 24447 -597 24459 -563
rect 24059 -603 24459 -597
rect 24677 -563 25077 -557
rect 24677 -597 24689 -563
rect 24700 -597 25060 -580
rect 25065 -597 25077 -563
rect 24677 -603 25077 -597
rect 25659 -563 26059 -557
rect 25659 -597 25671 -563
rect 25680 -597 26040 -580
rect 26047 -597 26059 -563
rect 25659 -603 26059 -597
rect 26277 -563 26677 -557
rect 26277 -597 26289 -563
rect 26300 -597 26660 -580
rect 26665 -597 26677 -563
rect 26277 -603 26677 -597
rect 27259 -563 27659 -557
rect 27259 -597 27271 -563
rect 27280 -597 27640 -580
rect 27647 -597 27659 -563
rect 27259 -603 27659 -597
rect 27877 -563 28277 -557
rect 27877 -597 27889 -563
rect 27900 -597 28260 -580
rect 28265 -597 28277 -563
rect 27877 -603 28277 -597
rect 28859 -563 29259 -557
rect 28859 -597 28871 -563
rect 28880 -597 29240 -580
rect 29247 -597 29259 -563
rect 28859 -603 29259 -597
rect 29477 -563 29877 -557
rect 29477 -597 29489 -563
rect 29500 -597 29860 -580
rect 29865 -597 29877 -563
rect 29477 -603 29877 -597
rect 30459 -563 30859 -557
rect 30459 -597 30471 -563
rect 30480 -597 30840 -580
rect 30847 -597 30859 -563
rect 30459 -603 30859 -597
rect 31077 -563 31477 -557
rect 31077 -597 31089 -563
rect 31100 -597 31460 -580
rect 31465 -597 31477 -563
rect 31077 -603 31477 -597
rect 32060 -563 32459 -560
rect 32060 -597 32071 -563
rect 32080 -597 32440 -580
rect 32447 -597 32459 -563
rect 32060 -603 32459 -597
rect 32677 -563 33077 -557
rect 32677 -597 32689 -563
rect 32700 -597 33060 -580
rect 33065 -597 33077 -563
rect 32677 -603 33077 -597
rect 33659 -563 34059 -557
rect 33659 -597 33671 -563
rect 33680 -597 34040 -580
rect 34047 -597 34059 -563
rect 33659 -603 34059 -597
rect 34277 -563 34677 -557
rect 34277 -597 34289 -563
rect 34300 -597 34660 -580
rect 34665 -597 34677 -563
rect 34277 -603 34677 -597
rect 35259 -563 35659 -557
rect 35259 -597 35271 -563
rect 35280 -597 35640 -580
rect 35647 -597 35659 -563
rect 35259 -603 35659 -597
rect 35877 -563 36277 -557
rect 35877 -597 35889 -563
rect 35900 -597 36260 -580
rect 36265 -597 36277 -563
rect 35877 -603 36277 -597
rect 16080 -640 16440 -603
rect 16700 -640 17060 -603
rect 17680 -640 18040 -603
rect 18300 -640 18660 -603
rect 19280 -640 19640 -603
rect 19900 -640 20260 -603
rect 20880 -640 21240 -603
rect 21500 -640 21860 -603
rect 22480 -640 22840 -603
rect 23100 -640 23460 -603
rect 24080 -640 24440 -603
rect 24700 -640 25060 -603
rect 25680 -640 26040 -603
rect 26300 -640 26660 -603
rect 27280 -640 27640 -603
rect 27900 -640 28260 -603
rect 28880 -640 29240 -603
rect 29500 -640 29860 -603
rect 30480 -640 30840 -603
rect 31100 -640 31460 -603
rect 32080 -640 32440 -603
rect 32700 -640 33060 -603
rect 33680 -640 34040 -603
rect 34300 -640 34660 -603
rect 35280 -640 35640 -603
rect 35900 -640 36260 -603
rect 14380 -740 15560 -730
rect 15590 -650 17060 -640
rect 15590 -770 15600 -650
rect 15700 -770 17060 -650
rect 15590 -780 17060 -770
rect 17190 -650 18660 -640
rect 17190 -770 17200 -650
rect 17300 -770 18660 -650
rect 17190 -780 18660 -770
rect 18790 -650 20260 -640
rect 18790 -770 18800 -650
rect 18900 -770 20260 -650
rect 18790 -780 20260 -770
rect 20390 -650 21860 -640
rect 20390 -770 20400 -650
rect 20500 -770 21860 -650
rect 20390 -780 21860 -770
rect 21990 -650 23460 -640
rect 21990 -770 22000 -650
rect 22100 -770 23460 -650
rect 21990 -780 23460 -770
rect 23590 -650 25060 -640
rect 23590 -770 23600 -650
rect 23700 -770 25060 -650
rect 23590 -780 25060 -770
rect 25660 -650 28260 -640
rect 25660 -770 26800 -650
rect 26900 -770 28260 -650
rect 25660 -780 28260 -770
rect 28390 -650 31460 -640
rect 28390 -770 28400 -650
rect 28500 -770 31460 -650
rect 28390 -780 31460 -770
rect 32060 -780 36260 -640
rect 12510 -810 12520 -780
rect 11400 -930 11480 -860
rect 12020 -930 12100 -860
rect 12380 -910 12520 -810
rect 12880 -880 13240 -780
rect 13500 -880 13860 -780
rect 12310 -930 12520 -910
rect 1540 -980 12520 -930
rect 1540 -1050 12390 -980
rect 12510 -1050 12520 -980
rect 1540 -1060 12520 -1050
rect 12620 -930 12820 -920
rect 1180 -1120 1320 -1110
rect 2780 -1120 2920 -1110
rect 4380 -1120 4520 -1110
rect 5980 -1120 6120 -1110
rect 7580 -1120 7720 -1110
rect 9180 -1120 9320 -1110
rect 11400 -1120 11480 -1060
rect 12020 -1120 12100 -1060
rect 12620 -1070 12630 -930
rect 12750 -1070 12820 -930
rect 12620 -1080 12820 -1070
rect 13920 -930 14100 -920
rect 13920 -1070 13970 -930
rect 14090 -1070 14100 -930
rect 14160 -930 14300 -780
rect 16080 -825 16440 -780
rect 16700 -825 17060 -780
rect 17680 -825 18040 -780
rect 18300 -825 18660 -780
rect 19280 -825 19640 -780
rect 19900 -825 20260 -780
rect 20880 -825 21240 -780
rect 21500 -825 21860 -780
rect 22480 -825 22840 -780
rect 23100 -825 23460 -780
rect 24080 -825 24440 -780
rect 24700 -825 25060 -780
rect 25680 -825 26040 -780
rect 26300 -825 26660 -780
rect 27280 -825 27640 -780
rect 27900 -825 28260 -780
rect 28880 -825 29240 -780
rect 29500 -825 29860 -780
rect 30480 -825 30840 -780
rect 31100 -825 31460 -780
rect 32080 -825 32440 -780
rect 32700 -825 33060 -780
rect 33680 -825 34040 -780
rect 34300 -825 34660 -780
rect 35280 -825 35640 -780
rect 35900 -825 36260 -780
rect 16059 -830 16459 -825
rect 14620 -930 14700 -860
rect 15220 -930 15300 -860
rect 16059 -871 16460 -830
rect 16677 -871 17077 -825
rect 17659 -830 18059 -825
rect 17659 -871 18060 -830
rect 18277 -871 18677 -825
rect 19259 -830 19659 -825
rect 19259 -871 19660 -830
rect 19877 -871 20277 -825
rect 20859 -830 21259 -825
rect 20859 -871 21260 -830
rect 21477 -871 21877 -825
rect 22459 -830 22859 -825
rect 22459 -871 22860 -830
rect 23077 -871 23477 -825
rect 24059 -830 24459 -825
rect 24059 -871 24460 -830
rect 24677 -871 25077 -825
rect 25659 -830 26059 -825
rect 25659 -871 26060 -830
rect 26277 -871 26677 -825
rect 27259 -830 27659 -825
rect 27259 -871 27660 -830
rect 27877 -871 28277 -825
rect 28859 -830 29259 -825
rect 28859 -871 29260 -830
rect 29477 -871 29877 -825
rect 30459 -830 30859 -825
rect 30459 -871 30860 -830
rect 31077 -871 31477 -825
rect 32060 -830 32459 -825
rect 16060 -890 16460 -871
rect 16680 -880 17070 -871
rect 16677 -891 17077 -880
rect 17660 -890 18060 -871
rect 18280 -880 18670 -871
rect 18277 -891 18677 -880
rect 19260 -890 19660 -871
rect 19880 -880 20270 -871
rect 19877 -891 20277 -880
rect 20860 -890 21260 -871
rect 21480 -880 21870 -871
rect 21477 -891 21877 -880
rect 22460 -890 22860 -871
rect 23080 -880 23470 -871
rect 23077 -891 23477 -880
rect 24060 -890 24460 -871
rect 24680 -880 25070 -871
rect 24677 -891 25077 -880
rect 25660 -890 26060 -871
rect 26280 -880 26670 -871
rect 26277 -891 26677 -880
rect 27260 -890 27660 -871
rect 27880 -880 28270 -871
rect 27877 -891 28277 -880
rect 28860 -890 29260 -871
rect 29480 -880 29870 -871
rect 29477 -891 29877 -880
rect 30460 -890 30860 -871
rect 31080 -880 31470 -871
rect 31077 -891 31477 -880
rect 32060 -890 32460 -830
rect 32677 -860 33077 -825
rect 33659 -830 34059 -825
rect 32680 -880 33070 -860
rect 33659 -871 34060 -830
rect 34277 -871 34677 -825
rect 35259 -830 35659 -825
rect 35259 -871 35660 -830
rect 35877 -871 36277 -825
rect 32677 -891 33077 -880
rect 33660 -890 34060 -871
rect 34280 -880 34670 -871
rect 34277 -891 34677 -880
rect 35260 -890 35660 -871
rect 35880 -880 36270 -871
rect 35877 -891 36277 -880
rect 14160 -1060 36400 -930
rect 13920 -1080 14100 -1070
rect 12870 -1110 13250 -1100
rect 1180 -1240 1190 -1120
rect 1310 -1240 2790 -1120
rect 2910 -1240 4390 -1120
rect 4510 -1240 5990 -1120
rect 6110 -1240 7590 -1120
rect 7710 -1240 9190 -1120
rect 9310 -1240 10720 -1120
rect 1180 -1250 1320 -1240
rect 2780 -1250 2920 -1240
rect 4380 -1250 4520 -1240
rect 5980 -1250 6120 -1240
rect 7580 -1250 7720 -1240
rect 9180 -1250 9320 -1240
rect 12870 -1260 12880 -1110
rect 13240 -1120 13250 -1110
rect 14620 -1120 14700 -1060
rect 15220 -1120 15300 -1060
rect 30459 -1109 30859 -1103
rect 30459 -1110 30471 -1109
rect 30847 -1110 30859 -1109
rect 31077 -1109 31477 -1103
rect 31077 -1110 31089 -1109
rect 31465 -1110 31477 -1109
rect 15810 -1120 15930 -1110
rect 17410 -1120 17530 -1110
rect 19010 -1120 19130 -1110
rect 20610 -1120 20730 -1110
rect 22210 -1120 22330 -1110
rect 23810 -1120 23930 -1110
rect 27010 -1120 28270 -1110
rect 13240 -1260 13860 -1120
rect 15810 -1240 15820 -1120
rect 15920 -1240 17120 -1120
rect 17410 -1240 17420 -1120
rect 17520 -1240 18720 -1120
rect 19010 -1240 19020 -1120
rect 19120 -1240 20320 -1120
rect 20610 -1240 20620 -1120
rect 20720 -1240 21920 -1120
rect 22210 -1240 22220 -1120
rect 22320 -1240 23520 -1120
rect 23810 -1240 23820 -1120
rect 23920 -1240 25120 -1120
rect 25620 -1240 27020 -1120
rect 27120 -1240 28270 -1120
rect 15810 -1250 15930 -1240
rect 17410 -1250 17530 -1240
rect 19010 -1250 19130 -1240
rect 20610 -1250 20730 -1240
rect 22210 -1250 22330 -1240
rect 23810 -1250 23930 -1240
rect 27010 -1250 28270 -1240
rect 28610 -1120 31520 -1110
rect 28610 -1240 28620 -1120
rect 28720 -1240 31520 -1120
rect 28610 -1250 31520 -1240
rect 31590 -1120 31710 -1110
rect 31590 -1240 31600 -1120
rect 31700 -1240 36270 -1120
rect 31590 -1250 31710 -1240
rect 12870 -1290 13860 -1260
rect 36660 -1300 36800 260
rect 37300 -1300 37440 260
rect 37920 -1300 38060 260
rect 31760 -1340 38060 -1300
rect 660 -1420 38060 -1340
rect 660 -1540 31780 -1420
rect 32060 -1470 33490 -1460
rect 32060 -1540 33360 -1470
rect 660 -3140 710 -1540
rect 33350 -1590 33360 -1540
rect 33480 -1590 33490 -1470
rect 33660 -1470 35650 -1460
rect 33660 -1540 35020 -1470
rect 2100 -1610 2240 -1600
rect 2100 -2290 2110 -1610
rect 2230 -2290 2240 -1610
rect 2100 -2300 2240 -2290
rect 3700 -1610 3840 -1600
rect 3700 -2290 3710 -1610
rect 3830 -2290 3840 -1610
rect 3700 -2300 3840 -2290
rect 5300 -1610 5440 -1600
rect 5300 -2290 5310 -1610
rect 5430 -2290 5440 -1610
rect 5300 -2300 5440 -2290
rect 6900 -1610 7040 -1600
rect 6900 -2290 6910 -1610
rect 7030 -2290 7040 -1610
rect 6900 -2300 7040 -2290
rect 8500 -1610 8640 -1600
rect 8500 -2290 8510 -1610
rect 8630 -2290 8640 -1610
rect 8500 -2300 8640 -2290
rect 10100 -1610 10240 -1600
rect 10100 -2290 10110 -1610
rect 10230 -2290 10240 -1610
rect 10100 -2300 10240 -2290
rect 11700 -1610 11840 -1600
rect 11700 -2290 11710 -1610
rect 11830 -2290 11840 -1610
rect 11700 -2300 11840 -2290
rect 13300 -1610 13440 -1600
rect 13300 -2290 13310 -1610
rect 13430 -2290 13440 -1610
rect 13300 -2300 13440 -2290
rect 14900 -1610 15040 -1600
rect 14900 -2290 14910 -1610
rect 15030 -2290 15040 -1610
rect 14900 -2300 15040 -2290
rect 16500 -1610 16640 -1600
rect 16500 -2290 16510 -1610
rect 16630 -2290 16640 -1610
rect 16500 -2300 16640 -2290
rect 18100 -1610 18240 -1600
rect 18100 -2290 18110 -1610
rect 18230 -2290 18240 -1610
rect 18100 -2300 18240 -2290
rect 19700 -1610 19840 -1600
rect 19700 -2290 19710 -1610
rect 19830 -2290 19840 -1610
rect 19700 -2300 19840 -2290
rect 21300 -1610 21440 -1600
rect 21300 -2290 21310 -1610
rect 21430 -2290 21440 -1610
rect 21300 -2300 21440 -2290
rect 22900 -1610 23040 -1600
rect 22900 -2290 22910 -1610
rect 23030 -2290 23040 -1610
rect 22900 -2300 23040 -2290
rect 24500 -1610 24640 -1600
rect 24500 -2290 24510 -1610
rect 24630 -2290 24640 -1610
rect 24500 -2300 24640 -2290
rect 26100 -1610 26240 -1600
rect 26100 -2290 26110 -1610
rect 26230 -2290 26240 -1610
rect 26100 -2300 26240 -2290
rect 27700 -1610 27840 -1600
rect 27700 -2290 27710 -1610
rect 27830 -2290 27840 -1610
rect 27700 -2300 27840 -2290
rect 28781 -1605 28827 -1593
rect 28781 -2297 28787 -1605
rect 28821 -2297 28827 -1605
rect 28781 -2309 28827 -2297
rect 29291 -1600 29337 -1593
rect 29399 -1600 29445 -1593
rect 29291 -1605 29445 -1600
rect 29291 -2297 29297 -1605
rect 29331 -1610 29405 -1605
rect 29331 -2297 29405 -2290
rect 29439 -2297 29445 -1605
rect 29291 -2300 29445 -2297
rect 29291 -2309 29337 -2300
rect 29399 -2309 29445 -2300
rect 29909 -1605 29955 -1593
rect 29909 -2297 29915 -1605
rect 29949 -2297 29955 -1605
rect 29909 -2309 29955 -2297
rect 30381 -1605 30427 -1593
rect 30381 -2297 30387 -1605
rect 30421 -2297 30427 -1605
rect 30381 -2309 30427 -2297
rect 30891 -1600 30937 -1593
rect 30999 -1600 31045 -1593
rect 30891 -1605 31045 -1600
rect 30891 -2297 30897 -1605
rect 30931 -1610 31005 -1605
rect 30931 -2297 31005 -2290
rect 31039 -2297 31045 -1605
rect 30891 -2300 31045 -2297
rect 30891 -2309 30937 -2300
rect 30999 -2309 31045 -2300
rect 31509 -1605 31555 -1593
rect 33350 -1600 33490 -1590
rect 35010 -1590 35020 -1540
rect 35140 -1540 35650 -1470
rect 35880 -1540 36270 -1420
rect 35140 -1570 35160 -1540
rect 35140 -1590 35150 -1570
rect 35010 -1600 35150 -1590
rect 35690 -1600 35760 -1590
rect 32500 -1605 32640 -1600
rect 34100 -1605 34240 -1600
rect 31509 -2297 31515 -1605
rect 31549 -2297 31555 -1605
rect 32531 -1610 32605 -1605
rect 32531 -2297 32605 -2290
rect 32639 -2297 32640 -1605
rect 34131 -1610 34205 -1605
rect 34131 -2297 34205 -2290
rect 34239 -2297 34240 -1605
rect 31509 -2309 31555 -2297
rect 32500 -2300 32640 -2297
rect 34100 -2300 34240 -2297
rect 35750 -2310 35760 -1600
rect 36018 -1838 36102 -1540
rect 35818 -2016 36338 -1838
rect 35690 -2320 35760 -2310
rect 11260 -2363 11659 -2360
rect 1680 -2440 2040 -2380
rect 2300 -2440 2660 -2380
rect 3280 -2440 3640 -2380
rect 3900 -2440 4260 -2380
rect 4880 -2440 5240 -2380
rect 5500 -2440 5860 -2380
rect 6480 -2440 6840 -2380
rect 7100 -2440 7460 -2380
rect 8080 -2440 8440 -2380
rect 8700 -2440 9060 -2380
rect 9680 -2440 10040 -2380
rect 10300 -2440 10660 -2380
rect 11260 -2397 11271 -2363
rect 11280 -2397 11640 -2380
rect 11647 -2397 11659 -2363
rect 11260 -2403 11659 -2397
rect 11877 -2363 12277 -2360
rect 11877 -2397 11889 -2363
rect 11900 -2397 12260 -2380
rect 12265 -2397 12277 -2363
rect 11877 -2403 12277 -2397
rect 12860 -2363 13259 -2360
rect 12860 -2397 12871 -2363
rect 12880 -2397 13240 -2380
rect 13247 -2397 13259 -2363
rect 12860 -2403 13259 -2397
rect 13477 -2363 13877 -2360
rect 13477 -2397 13489 -2363
rect 13500 -2397 13860 -2380
rect 13865 -2397 13877 -2363
rect 13477 -2403 13877 -2397
rect 14459 -2363 14859 -2357
rect 14459 -2397 14471 -2363
rect 14480 -2397 14840 -2380
rect 14847 -2397 14859 -2363
rect 14459 -2403 14859 -2397
rect 15077 -2363 15477 -2357
rect 15077 -2397 15089 -2363
rect 15100 -2397 15460 -2380
rect 15465 -2397 15477 -2363
rect 15077 -2403 15477 -2397
rect 16059 -2363 16459 -2357
rect 16059 -2397 16071 -2363
rect 16080 -2397 16440 -2380
rect 16447 -2397 16459 -2363
rect 16059 -2403 16459 -2397
rect 16677 -2363 17077 -2357
rect 16677 -2397 16689 -2363
rect 16700 -2397 17060 -2380
rect 17065 -2397 17077 -2363
rect 16677 -2403 17077 -2397
rect 17659 -2363 18059 -2357
rect 17659 -2397 17671 -2363
rect 17680 -2397 18040 -2380
rect 18047 -2397 18059 -2363
rect 17659 -2403 18059 -2397
rect 18277 -2363 18677 -2357
rect 18277 -2397 18289 -2363
rect 18300 -2397 18660 -2380
rect 18665 -2397 18677 -2363
rect 18277 -2403 18677 -2397
rect 19259 -2363 19659 -2357
rect 19259 -2397 19271 -2363
rect 19280 -2397 19640 -2380
rect 19647 -2397 19659 -2363
rect 19259 -2403 19659 -2397
rect 19877 -2363 20277 -2357
rect 19877 -2397 19889 -2363
rect 19900 -2397 20260 -2380
rect 20265 -2397 20277 -2363
rect 19877 -2403 20277 -2397
rect 20859 -2363 21259 -2357
rect 20859 -2397 20871 -2363
rect 20880 -2397 21240 -2380
rect 21247 -2397 21259 -2363
rect 20859 -2403 21259 -2397
rect 21477 -2363 21877 -2357
rect 21477 -2397 21489 -2363
rect 21500 -2397 21860 -2380
rect 21865 -2397 21877 -2363
rect 21477 -2403 21877 -2397
rect 22459 -2363 22859 -2357
rect 22459 -2397 22471 -2363
rect 22480 -2397 22840 -2380
rect 22847 -2397 22859 -2363
rect 22459 -2403 22859 -2397
rect 23077 -2363 23477 -2357
rect 23077 -2397 23089 -2363
rect 23100 -2397 23460 -2380
rect 23465 -2397 23477 -2363
rect 23077 -2403 23477 -2397
rect 24059 -2363 24459 -2357
rect 24059 -2397 24071 -2363
rect 24080 -2397 24440 -2380
rect 24447 -2397 24459 -2363
rect 24059 -2403 24459 -2397
rect 24677 -2363 25077 -2357
rect 24677 -2397 24689 -2363
rect 24700 -2397 25060 -2380
rect 25065 -2397 25077 -2363
rect 24677 -2403 25077 -2397
rect 25659 -2363 26059 -2357
rect 25659 -2397 25671 -2363
rect 25680 -2397 26040 -2380
rect 26047 -2397 26059 -2363
rect 25659 -2403 26059 -2397
rect 26277 -2363 26677 -2357
rect 26277 -2397 26289 -2363
rect 26300 -2397 26660 -2380
rect 26665 -2397 26677 -2363
rect 26277 -2403 26677 -2397
rect 27259 -2363 27659 -2357
rect 27259 -2397 27271 -2363
rect 27280 -2397 27640 -2380
rect 27647 -2397 27659 -2363
rect 27259 -2403 27659 -2397
rect 27877 -2363 28277 -2357
rect 27877 -2397 27889 -2363
rect 27900 -2397 28260 -2380
rect 28265 -2397 28277 -2363
rect 27877 -2403 28277 -2397
rect 28859 -2363 29259 -2357
rect 28859 -2397 28871 -2363
rect 28880 -2397 29240 -2380
rect 29247 -2397 29259 -2363
rect 28859 -2403 29259 -2397
rect 29477 -2363 29877 -2357
rect 29477 -2397 29489 -2363
rect 29500 -2397 29860 -2380
rect 29865 -2397 29877 -2363
rect 29477 -2403 29877 -2397
rect 30459 -2363 30859 -2357
rect 30459 -2397 30471 -2363
rect 30480 -2397 30840 -2380
rect 30847 -2397 30859 -2363
rect 30459 -2403 30859 -2397
rect 31077 -2363 31477 -2357
rect 31077 -2397 31089 -2363
rect 31100 -2397 31460 -2380
rect 31465 -2397 31477 -2363
rect 31077 -2403 31477 -2397
rect 32060 -2363 32459 -2360
rect 32060 -2397 32071 -2363
rect 32080 -2397 32440 -2380
rect 32447 -2397 32459 -2363
rect 32060 -2403 32459 -2397
rect 32677 -2363 33077 -2357
rect 32677 -2397 32689 -2363
rect 32700 -2397 33060 -2380
rect 33065 -2397 33077 -2363
rect 32677 -2403 33077 -2397
rect 33659 -2363 34059 -2357
rect 33659 -2397 33671 -2363
rect 33680 -2397 34040 -2380
rect 34047 -2397 34059 -2363
rect 33659 -2403 34059 -2397
rect 34277 -2363 34677 -2357
rect 34277 -2397 34289 -2363
rect 34300 -2397 34660 -2380
rect 34665 -2397 34677 -2363
rect 34277 -2403 34677 -2397
rect 35259 -2363 35659 -2357
rect 35259 -2397 35271 -2363
rect 35280 -2397 35640 -2380
rect 35647 -2397 35659 -2363
rect 36018 -2386 36102 -2016
rect 35259 -2403 35659 -2397
rect 11280 -2440 11640 -2403
rect 11900 -2440 12260 -2403
rect 12880 -2440 13240 -2403
rect 13500 -2440 13860 -2403
rect 14480 -2440 14840 -2403
rect 15100 -2440 15460 -2403
rect 16080 -2440 16440 -2403
rect 16700 -2440 17060 -2403
rect 17680 -2440 18040 -2403
rect 18300 -2440 18660 -2403
rect 19280 -2440 19640 -2403
rect 19900 -2440 20260 -2403
rect 20880 -2440 21240 -2403
rect 21500 -2440 21860 -2403
rect 22480 -2440 22840 -2403
rect 23100 -2440 23460 -2403
rect 24080 -2440 24440 -2403
rect 24700 -2440 25060 -2403
rect 25680 -2440 26040 -2403
rect 26300 -2440 26660 -2403
rect 27280 -2440 27640 -2403
rect 27900 -2440 28260 -2403
rect 28880 -2440 29240 -2403
rect 29500 -2440 29860 -2403
rect 30480 -2440 30840 -2403
rect 31100 -2440 31460 -2403
rect 32080 -2440 32440 -2403
rect 32700 -2440 33060 -2403
rect 33680 -2440 34040 -2403
rect 34300 -2440 34660 -2403
rect 35280 -2440 35640 -2403
rect 1400 -2450 10660 -2440
rect 1400 -2570 1410 -2450
rect 1530 -2570 3010 -2450
rect 3130 -2570 4610 -2450
rect 4730 -2570 6210 -2450
rect 6330 -2570 7810 -2450
rect 7930 -2570 9410 -2450
rect 9530 -2570 10660 -2450
rect 1400 -2580 10660 -2570
rect 11260 -2580 12260 -2440
rect 12860 -2580 13860 -2440
rect 14460 -2580 15460 -2440
rect 15590 -2450 17060 -2440
rect 15590 -2570 15600 -2450
rect 15700 -2570 17060 -2450
rect 15590 -2580 17060 -2570
rect 17190 -2450 18660 -2440
rect 17190 -2570 17200 -2450
rect 17300 -2570 18660 -2450
rect 17190 -2580 18660 -2570
rect 18790 -2450 20260 -2440
rect 18790 -2570 18800 -2450
rect 18900 -2570 20260 -2450
rect 18790 -2580 20260 -2570
rect 20390 -2450 21860 -2440
rect 20390 -2570 20400 -2450
rect 20500 -2570 21860 -2450
rect 20390 -2580 21860 -2570
rect 21990 -2450 23460 -2440
rect 21990 -2570 22000 -2450
rect 22100 -2570 23460 -2450
rect 21990 -2580 23460 -2570
rect 23590 -2450 25060 -2440
rect 23590 -2570 23600 -2450
rect 23700 -2570 25060 -2450
rect 23590 -2580 25060 -2570
rect 25190 -2450 26660 -2440
rect 25190 -2570 25200 -2450
rect 25300 -2570 26660 -2450
rect 25190 -2580 26660 -2570
rect 26791 -2450 28260 -2440
rect 26791 -2570 26800 -2450
rect 26900 -2570 28260 -2450
rect 26791 -2580 28260 -2570
rect 28390 -2450 29860 -2440
rect 28390 -2570 28400 -2450
rect 28500 -2570 29860 -2450
rect 28390 -2580 29860 -2570
rect 29990 -2450 31460 -2440
rect 29990 -2570 30000 -2450
rect 30100 -2570 31460 -2450
rect 29990 -2580 31460 -2570
rect 32060 -2450 33310 -2440
rect 32060 -2570 33180 -2450
rect 33300 -2570 33310 -2450
rect 32060 -2580 33310 -2570
rect 33660 -2580 35640 -2440
rect 1680 -2650 2040 -2580
rect 2300 -2650 2660 -2580
rect 3280 -2650 3640 -2580
rect 3900 -2650 4260 -2580
rect 4880 -2650 5240 -2580
rect 5500 -2650 5860 -2580
rect 6480 -2650 6840 -2580
rect 7100 -2650 7460 -2580
rect 8080 -2650 8440 -2580
rect 8700 -2650 9060 -2580
rect 9680 -2650 10040 -2580
rect 10300 -2650 10660 -2580
rect 11280 -2625 11640 -2580
rect 11900 -2625 12260 -2580
rect 12880 -2625 13240 -2580
rect 13500 -2625 13860 -2580
rect 14480 -2625 14840 -2580
rect 15100 -2625 15460 -2580
rect 16080 -2625 16440 -2580
rect 16700 -2625 17060 -2580
rect 17680 -2625 18040 -2580
rect 18300 -2625 18660 -2580
rect 19280 -2625 19640 -2580
rect 19900 -2625 20260 -2580
rect 20880 -2625 21240 -2580
rect 21500 -2625 21860 -2580
rect 22480 -2625 22840 -2580
rect 23100 -2625 23460 -2580
rect 24080 -2625 24440 -2580
rect 24700 -2625 25060 -2580
rect 25680 -2625 26040 -2580
rect 26300 -2625 26660 -2580
rect 27280 -2625 27640 -2580
rect 27900 -2625 28260 -2580
rect 28880 -2625 29240 -2580
rect 29500 -2625 29860 -2580
rect 30480 -2625 30840 -2580
rect 31100 -2625 31460 -2580
rect 32080 -2625 32440 -2580
rect 32700 -2625 33060 -2580
rect 33680 -2625 34040 -2580
rect 34300 -2625 34660 -2580
rect 35280 -2625 35640 -2580
rect 11260 -2671 11659 -2625
rect 11877 -2671 12277 -2625
rect 12860 -2671 13259 -2625
rect 13477 -2671 13877 -2625
rect 14459 -2671 14859 -2625
rect 15077 -2671 15477 -2625
rect 16059 -2630 16459 -2625
rect 16059 -2671 16460 -2630
rect 16677 -2671 17077 -2625
rect 17659 -2630 18059 -2625
rect 17659 -2671 18060 -2630
rect 18277 -2671 18677 -2625
rect 19259 -2630 19659 -2625
rect 19259 -2671 19660 -2630
rect 19877 -2671 20277 -2625
rect 20859 -2630 21259 -2625
rect 20859 -2671 21260 -2630
rect 21477 -2671 21877 -2625
rect 22459 -2630 22859 -2625
rect 22459 -2671 22860 -2630
rect 23077 -2671 23477 -2625
rect 24059 -2630 24459 -2625
rect 24059 -2671 24460 -2630
rect 24677 -2671 25077 -2625
rect 25659 -2630 26059 -2625
rect 25659 -2671 26060 -2630
rect 26277 -2671 26677 -2625
rect 27259 -2630 27659 -2625
rect 27259 -2671 27660 -2630
rect 27877 -2671 28277 -2625
rect 28859 -2630 29259 -2625
rect 28859 -2671 29260 -2630
rect 29477 -2671 29877 -2625
rect 30459 -2630 30859 -2625
rect 30459 -2671 30860 -2630
rect 31077 -2671 31477 -2625
rect 32060 -2630 32459 -2625
rect 16060 -2690 16460 -2671
rect 16680 -2680 17070 -2671
rect 16677 -2691 17077 -2680
rect 17660 -2690 18060 -2671
rect 18280 -2680 18670 -2671
rect 18277 -2691 18677 -2680
rect 19260 -2690 19660 -2671
rect 19880 -2680 20270 -2671
rect 19877 -2691 20277 -2680
rect 20860 -2690 21260 -2671
rect 21480 -2680 21870 -2671
rect 21477 -2691 21877 -2680
rect 22460 -2690 22860 -2671
rect 23080 -2680 23470 -2671
rect 23077 -2691 23477 -2680
rect 24060 -2690 24460 -2671
rect 24680 -2680 25070 -2671
rect 24677 -2691 25077 -2680
rect 25660 -2690 26060 -2671
rect 26280 -2680 26670 -2671
rect 26277 -2691 26677 -2680
rect 27260 -2690 27660 -2671
rect 27880 -2680 28270 -2671
rect 27877 -2691 28277 -2680
rect 28860 -2690 29260 -2671
rect 29480 -2680 29870 -2671
rect 29477 -2691 29877 -2680
rect 30460 -2690 30860 -2671
rect 31080 -2680 31470 -2671
rect 31077 -2691 31477 -2680
rect 32060 -2690 32460 -2630
rect 32677 -2660 33077 -2625
rect 33659 -2630 34059 -2625
rect 32680 -2680 33070 -2660
rect 33659 -2671 34060 -2630
rect 34277 -2671 34677 -2625
rect 35259 -2630 35659 -2625
rect 35259 -2671 35660 -2630
rect 32677 -2691 33077 -2680
rect 33660 -2690 34060 -2671
rect 34280 -2680 34670 -2671
rect 34277 -2691 34677 -2680
rect 35260 -2690 35660 -2671
rect 12320 -2730 12520 -2720
rect 36026 -2730 36116 -2666
rect 1540 -2850 12390 -2730
rect 12510 -2850 36400 -2730
rect 1540 -2860 36400 -2850
rect 1180 -2920 1320 -2910
rect 2780 -2920 2920 -2910
rect 4380 -2920 4520 -2910
rect 5980 -2920 6120 -2910
rect 7580 -2920 7720 -2910
rect 9180 -2920 9320 -2910
rect 11000 -2920 11140 -2910
rect 14200 -2920 14340 -2910
rect 1180 -3040 1190 -2920
rect 1310 -3040 2790 -2920
rect 2910 -3040 4390 -2920
rect 4510 -3040 5990 -2920
rect 6110 -3040 7590 -2920
rect 7710 -3040 9190 -2920
rect 9310 -3040 10720 -2920
rect 11000 -3040 11010 -2920
rect 11130 -3040 12320 -2920
rect 12820 -3040 14210 -2920
rect 14330 -3040 14340 -2920
rect 1180 -3050 1320 -3040
rect 2780 -3050 2920 -3040
rect 4380 -3050 4520 -3040
rect 5980 -3050 6120 -3040
rect 7580 -3050 7720 -3040
rect 9180 -3050 9320 -3040
rect 11000 -3050 11140 -3040
rect 14200 -3050 14340 -3040
rect 14420 -2920 14560 -2910
rect 15810 -2920 15930 -2910
rect 17410 -2920 17530 -2910
rect 19010 -2920 19130 -2910
rect 20610 -2920 20730 -2910
rect 22210 -2920 22330 -2910
rect 23810 -2920 23930 -2910
rect 25410 -2920 25530 -2910
rect 27011 -2920 27130 -2910
rect 28610 -2920 29880 -2910
rect 14420 -3040 14430 -2920
rect 14550 -3040 15520 -2920
rect 15810 -3040 15820 -2920
rect 15920 -3040 17120 -2920
rect 17410 -3040 17420 -2920
rect 17520 -3040 18720 -2920
rect 19010 -3040 19020 -2920
rect 19120 -3040 20320 -2920
rect 20610 -3040 20620 -2920
rect 20720 -3040 21920 -2920
rect 22210 -3040 22220 -2920
rect 22320 -3040 23520 -2920
rect 23810 -3040 23820 -2920
rect 23920 -3040 25120 -2920
rect 25410 -3040 25420 -2920
rect 25520 -3040 26720 -2920
rect 27011 -3040 27020 -2920
rect 27120 -3040 28320 -2920
rect 28610 -3040 28620 -2920
rect 28720 -3040 29880 -2920
rect 14420 -3050 14560 -3040
rect 15810 -3050 15930 -3040
rect 17410 -3050 17530 -3040
rect 19010 -3050 19130 -3040
rect 20610 -3050 20730 -3040
rect 22210 -3050 22330 -3040
rect 23810 -3050 23930 -3040
rect 25410 -3050 25530 -3040
rect 27011 -3050 27130 -3040
rect 28610 -3050 29880 -3040
rect 30210 -2920 30330 -2910
rect 30210 -3040 30220 -2920
rect 30320 -3040 31480 -2920
rect 32060 -2980 35840 -2920
rect 36026 -2930 36116 -2860
rect 36390 -2910 36510 -2900
rect 36390 -2920 36400 -2910
rect 36320 -2980 36400 -2920
rect 32060 -3030 36400 -2980
rect 36500 -3030 36510 -2910
rect 32060 -3040 36510 -3030
rect 30210 -3050 30330 -3040
rect 36660 -3100 36800 -1420
rect 37300 -3100 37440 -1420
rect 37920 -3100 38060 -1420
rect 31720 -3140 38100 -3100
rect 660 -3220 38100 -3140
rect 660 -3240 31960 -3220
rect 660 -3340 12520 -3240
rect 12600 -3290 13260 -3280
rect 660 -4780 710 -3340
rect 12600 -3390 12610 -3290
rect 12730 -3340 13260 -3290
rect 13380 -3340 14120 -3240
rect 14200 -3290 14860 -3280
rect 12730 -3390 12740 -3340
rect 12600 -3400 12740 -3390
rect 2100 -3410 2240 -3400
rect 2100 -4090 2110 -3410
rect 2230 -4090 2240 -3410
rect 2100 -4100 2240 -4090
rect 3700 -3410 3840 -3400
rect 3700 -4090 3710 -3410
rect 3830 -4090 3840 -3410
rect 3700 -4100 3840 -4090
rect 5300 -3410 5440 -3400
rect 5300 -4090 5310 -3410
rect 5430 -4090 5440 -3410
rect 5300 -4100 5440 -4090
rect 6900 -3410 7040 -3400
rect 6900 -4090 6910 -3410
rect 7030 -4090 7040 -3410
rect 6900 -4100 7040 -4090
rect 8500 -3410 8640 -3400
rect 8500 -4090 8510 -3410
rect 8630 -4090 8640 -3410
rect 8500 -4100 8640 -4090
rect 10100 -3410 10240 -3400
rect 10100 -4090 10110 -3410
rect 10230 -4090 10240 -3410
rect 10100 -4100 10240 -4090
rect 11700 -3410 11840 -3400
rect 11700 -4090 11710 -3410
rect 11830 -4090 11840 -3410
rect 11700 -4100 11840 -4090
rect 13300 -3410 13440 -3400
rect 13300 -4090 13310 -3410
rect 13430 -4090 13440 -3410
rect 14200 -3410 14210 -3290
rect 14330 -3340 14860 -3290
rect 14980 -3340 31960 -3240
rect 32060 -3280 36270 -3270
rect 32060 -3340 33400 -3280
rect 14330 -3410 14340 -3340
rect 14200 -3420 14340 -3410
rect 14900 -3410 15040 -3400
rect 13300 -4100 13440 -4090
rect 14900 -4090 14910 -3410
rect 15030 -4090 15040 -3410
rect 14900 -4100 15040 -4090
rect 16500 -3410 16640 -3400
rect 16500 -4090 16510 -3410
rect 16630 -4090 16640 -3410
rect 16500 -4100 16640 -4090
rect 18100 -3410 18240 -3400
rect 18100 -4090 18110 -3410
rect 18230 -4090 18240 -3410
rect 18100 -4100 18240 -4090
rect 19700 -3410 19840 -3400
rect 19700 -4090 19710 -3410
rect 19830 -4090 19840 -3410
rect 19700 -4100 19840 -4090
rect 21300 -3410 21440 -3400
rect 21300 -4090 21310 -3410
rect 21430 -4090 21440 -3410
rect 21300 -4100 21440 -4090
rect 22900 -3410 23040 -3400
rect 22900 -4090 22910 -3410
rect 23030 -4090 23040 -3410
rect 22900 -4100 23040 -4090
rect 24500 -3410 24640 -3400
rect 24500 -4090 24510 -3410
rect 24630 -4090 24640 -3410
rect 24500 -4100 24640 -4090
rect 26100 -3410 26240 -3400
rect 26100 -4090 26110 -3410
rect 26230 -4090 26240 -3410
rect 26100 -4100 26240 -4090
rect 27700 -3410 27840 -3400
rect 27700 -4090 27710 -3410
rect 27830 -4090 27840 -3410
rect 27700 -4100 27840 -4090
rect 28781 -3405 28827 -3393
rect 28781 -4097 28787 -3405
rect 28821 -4097 28827 -3405
rect 28781 -4109 28827 -4097
rect 29291 -3400 29337 -3393
rect 29399 -3400 29445 -3393
rect 29291 -3405 29445 -3400
rect 29291 -4097 29297 -3405
rect 29331 -3410 29405 -3405
rect 29331 -4097 29405 -4090
rect 29439 -4097 29445 -3405
rect 29291 -4100 29445 -4097
rect 29291 -4109 29337 -4100
rect 29399 -4109 29445 -4100
rect 29909 -3405 29955 -3393
rect 29909 -4097 29915 -3405
rect 29949 -4097 29955 -3405
rect 29909 -4109 29955 -4097
rect 30381 -3405 30427 -3393
rect 30381 -4097 30387 -3405
rect 30421 -4097 30427 -3405
rect 30381 -4109 30427 -4097
rect 30891 -3400 30937 -3393
rect 30999 -3400 31045 -3393
rect 30891 -3405 31045 -3400
rect 30891 -4097 30897 -3405
rect 30931 -3410 31005 -3405
rect 30931 -4097 31005 -4090
rect 31039 -4097 31045 -3405
rect 30891 -4100 31045 -4097
rect 30891 -4109 30937 -4100
rect 30999 -4109 31045 -4100
rect 31509 -3405 31555 -3393
rect 33390 -3400 33400 -3340
rect 33530 -3340 36270 -3280
rect 36530 -3340 38100 -3220
rect 31509 -4097 31515 -3405
rect 31549 -4097 31555 -3405
rect 31509 -4109 31555 -4097
rect 32500 -3410 32640 -3400
rect 33390 -3410 33530 -3400
rect 34100 -3405 34240 -3400
rect 35700 -3405 35840 -3400
rect 34131 -3410 34205 -3405
rect 32500 -4090 32510 -3410
rect 32630 -4090 32640 -3410
rect 32500 -4100 32640 -4090
rect 34131 -4097 34205 -4090
rect 34239 -4097 34240 -3405
rect 35731 -3410 35805 -3405
rect 35731 -4097 35805 -4090
rect 35839 -4097 35840 -3405
rect 34100 -4100 34240 -4097
rect 35700 -4100 35840 -4097
rect 11260 -4163 11659 -4160
rect 1680 -4240 2040 -4180
rect 2300 -4240 2660 -4180
rect 3280 -4240 3640 -4180
rect 3900 -4240 4260 -4180
rect 4880 -4240 5240 -4180
rect 5500 -4240 5860 -4180
rect 6480 -4240 6840 -4180
rect 7100 -4240 7460 -4180
rect 8080 -4240 8440 -4180
rect 8700 -4240 9060 -4180
rect 9680 -4240 10040 -4180
rect 10300 -4240 10660 -4180
rect 11260 -4197 11271 -4163
rect 11280 -4197 11640 -4180
rect 11647 -4197 11659 -4163
rect 11260 -4203 11659 -4197
rect 11877 -4163 12277 -4160
rect 11877 -4197 11889 -4163
rect 11900 -4197 12260 -4180
rect 12265 -4197 12277 -4163
rect 12860 -4163 13259 -4160
rect 12860 -4180 12871 -4163
rect 13247 -4180 13259 -4163
rect 13477 -4163 13877 -4160
rect 13477 -4180 13489 -4163
rect 13865 -4180 13877 -4163
rect 16059 -4163 16459 -4157
rect 11877 -4203 12277 -4197
rect 11280 -4240 11640 -4203
rect 11900 -4240 12260 -4203
rect 1400 -4250 10660 -4240
rect 1400 -4370 1410 -4250
rect 1530 -4370 3010 -4250
rect 3130 -4370 4610 -4250
rect 4730 -4370 6210 -4250
rect 6330 -4370 7810 -4250
rect 7930 -4370 9410 -4250
rect 9530 -4370 10660 -4250
rect 1400 -4380 10660 -4370
rect 11260 -4380 12260 -4240
rect 12840 -4260 13880 -4180
rect 14440 -4260 15480 -4180
rect 16059 -4197 16071 -4163
rect 16080 -4197 16440 -4180
rect 16447 -4197 16459 -4163
rect 16059 -4203 16459 -4197
rect 16677 -4163 17077 -4157
rect 16677 -4197 16689 -4163
rect 16700 -4197 17060 -4180
rect 17065 -4197 17077 -4163
rect 16677 -4203 17077 -4197
rect 17659 -4163 18059 -4157
rect 17659 -4197 17671 -4163
rect 17680 -4197 18040 -4180
rect 18047 -4197 18059 -4163
rect 17659 -4203 18059 -4197
rect 18277 -4163 18677 -4157
rect 18277 -4197 18289 -4163
rect 18300 -4197 18660 -4180
rect 18665 -4197 18677 -4163
rect 18277 -4203 18677 -4197
rect 19259 -4163 19659 -4157
rect 19259 -4197 19271 -4163
rect 19280 -4197 19640 -4180
rect 19647 -4197 19659 -4163
rect 19259 -4203 19659 -4197
rect 19877 -4163 20277 -4157
rect 19877 -4197 19889 -4163
rect 19900 -4197 20260 -4180
rect 20265 -4197 20277 -4163
rect 19877 -4203 20277 -4197
rect 20859 -4163 21259 -4157
rect 20859 -4197 20871 -4163
rect 20880 -4197 21240 -4180
rect 21247 -4197 21259 -4163
rect 20859 -4203 21259 -4197
rect 21477 -4163 21877 -4157
rect 21477 -4197 21489 -4163
rect 21500 -4197 21860 -4180
rect 21865 -4197 21877 -4163
rect 21477 -4203 21877 -4197
rect 22459 -4163 22859 -4157
rect 22459 -4197 22471 -4163
rect 22480 -4197 22840 -4180
rect 22847 -4197 22859 -4163
rect 22459 -4203 22859 -4197
rect 23077 -4163 23477 -4157
rect 23077 -4197 23089 -4163
rect 23100 -4197 23460 -4180
rect 23465 -4197 23477 -4163
rect 23077 -4203 23477 -4197
rect 24059 -4163 24459 -4157
rect 24059 -4197 24071 -4163
rect 24080 -4197 24440 -4180
rect 24447 -4197 24459 -4163
rect 24059 -4203 24459 -4197
rect 24677 -4163 25077 -4157
rect 24677 -4197 24689 -4163
rect 24700 -4197 25060 -4180
rect 25065 -4197 25077 -4163
rect 24677 -4203 25077 -4197
rect 25659 -4163 26059 -4157
rect 25659 -4197 25671 -4163
rect 25680 -4197 26040 -4180
rect 26047 -4197 26059 -4163
rect 25659 -4203 26059 -4197
rect 26277 -4163 26677 -4157
rect 26277 -4197 26289 -4163
rect 26300 -4197 26660 -4180
rect 26665 -4197 26677 -4163
rect 26277 -4203 26677 -4197
rect 27259 -4163 27659 -4157
rect 27259 -4197 27271 -4163
rect 27280 -4197 27640 -4180
rect 27647 -4197 27659 -4163
rect 27259 -4203 27659 -4197
rect 27877 -4163 28277 -4157
rect 27877 -4197 27889 -4163
rect 27900 -4197 28260 -4180
rect 28265 -4197 28277 -4163
rect 27877 -4203 28277 -4197
rect 28859 -4163 29259 -4157
rect 28859 -4197 28871 -4163
rect 28880 -4197 29240 -4180
rect 29247 -4197 29259 -4163
rect 28859 -4203 29259 -4197
rect 29477 -4163 29877 -4157
rect 29477 -4197 29489 -4163
rect 29500 -4197 29860 -4180
rect 29865 -4197 29877 -4163
rect 29477 -4203 29877 -4197
rect 30459 -4163 30859 -4157
rect 30459 -4197 30471 -4163
rect 30480 -4197 30840 -4180
rect 30847 -4197 30859 -4163
rect 30459 -4203 30859 -4197
rect 31077 -4163 31477 -4157
rect 31077 -4197 31089 -4163
rect 31100 -4197 31460 -4180
rect 31465 -4197 31477 -4163
rect 31077 -4203 31477 -4197
rect 32060 -4163 32459 -4160
rect 32060 -4197 32071 -4163
rect 32080 -4197 32440 -4180
rect 32447 -4197 32459 -4163
rect 32060 -4203 32459 -4197
rect 32677 -4163 33077 -4157
rect 32677 -4197 32689 -4163
rect 32700 -4197 33060 -4180
rect 33065 -4197 33077 -4163
rect 32677 -4203 33077 -4197
rect 33659 -4163 34059 -4157
rect 33659 -4197 33671 -4163
rect 33680 -4197 34040 -4180
rect 34047 -4197 34059 -4163
rect 33659 -4203 34059 -4197
rect 34277 -4163 34677 -4157
rect 34277 -4197 34289 -4163
rect 34300 -4197 34660 -4180
rect 34665 -4197 34677 -4163
rect 34277 -4203 34677 -4197
rect 35259 -4163 35659 -4157
rect 35259 -4197 35271 -4163
rect 35280 -4197 35640 -4180
rect 35647 -4197 35659 -4163
rect 35259 -4203 35659 -4197
rect 35877 -4163 36277 -4157
rect 35877 -4197 35889 -4163
rect 35900 -4197 36260 -4180
rect 36265 -4197 36277 -4163
rect 35877 -4203 36277 -4197
rect 16080 -4240 16440 -4203
rect 16700 -4240 17060 -4203
rect 17680 -4240 18040 -4203
rect 18300 -4240 18660 -4203
rect 19280 -4240 19640 -4203
rect 19900 -4240 20260 -4203
rect 20880 -4240 21240 -4203
rect 21500 -4240 21860 -4203
rect 22480 -4240 22840 -4203
rect 23100 -4240 23460 -4203
rect 24080 -4240 24440 -4203
rect 24700 -4240 25060 -4203
rect 25680 -4240 26040 -4203
rect 26300 -4240 26660 -4203
rect 27280 -4240 27640 -4203
rect 27900 -4240 28260 -4203
rect 28880 -4240 29240 -4203
rect 29500 -4240 29860 -4203
rect 30480 -4240 30840 -4203
rect 31100 -4240 31460 -4203
rect 32080 -4240 32440 -4203
rect 32700 -4240 33060 -4203
rect 33680 -4240 34040 -4203
rect 34300 -4240 34660 -4203
rect 35280 -4240 35640 -4203
rect 35900 -4240 36260 -4203
rect 15590 -4250 17060 -4240
rect 15590 -4370 15600 -4250
rect 15700 -4370 17060 -4250
rect 1680 -4450 2040 -4380
rect 2300 -4450 2660 -4380
rect 3280 -4450 3640 -4380
rect 3900 -4450 4260 -4380
rect 4880 -4450 5240 -4380
rect 5500 -4450 5860 -4380
rect 6480 -4450 6840 -4380
rect 7100 -4450 7460 -4380
rect 8080 -4450 8440 -4380
rect 8700 -4450 9060 -4380
rect 9680 -4450 10040 -4380
rect 10300 -4450 10660 -4380
rect 11280 -4425 11640 -4380
rect 11900 -4425 12260 -4380
rect 11260 -4430 11659 -4425
rect 11260 -4490 11660 -4430
rect 11877 -4460 12277 -4425
rect 12850 -4460 13880 -4370
rect 14450 -4460 15480 -4370
rect 15590 -4380 17060 -4370
rect 17190 -4250 18660 -4240
rect 17190 -4370 17200 -4250
rect 17300 -4370 18660 -4250
rect 17190 -4380 18660 -4370
rect 18790 -4250 20260 -4240
rect 18790 -4370 18800 -4250
rect 18900 -4370 20260 -4250
rect 18790 -4380 20260 -4370
rect 20390 -4250 21860 -4240
rect 20390 -4370 20400 -4250
rect 20500 -4370 21860 -4250
rect 20390 -4380 21860 -4370
rect 21990 -4250 23460 -4240
rect 21990 -4370 22000 -4250
rect 22100 -4370 23460 -4250
rect 21990 -4380 23460 -4370
rect 23590 -4250 25060 -4240
rect 23590 -4370 23600 -4250
rect 23700 -4370 25060 -4250
rect 23590 -4380 25060 -4370
rect 25190 -4250 26660 -4240
rect 25190 -4370 25200 -4250
rect 25300 -4370 26660 -4250
rect 25190 -4380 26660 -4370
rect 26791 -4250 28260 -4240
rect 26791 -4370 26800 -4250
rect 26900 -4370 28260 -4250
rect 26791 -4380 28260 -4370
rect 28391 -4250 29860 -4240
rect 28391 -4370 28400 -4250
rect 28500 -4370 29860 -4250
rect 28391 -4380 29860 -4370
rect 29990 -4250 31460 -4240
rect 29990 -4370 30000 -4250
rect 30100 -4370 31460 -4250
rect 29990 -4380 31460 -4370
rect 32060 -4250 36260 -4240
rect 32060 -4370 33180 -4250
rect 33300 -4370 36260 -4250
rect 36660 -4320 36800 -3340
rect 37300 -4320 37440 -3340
rect 37920 -4320 38060 -3340
rect 32060 -4380 36260 -4370
rect 16080 -4425 16440 -4380
rect 16700 -4425 17060 -4380
rect 17680 -4425 18040 -4380
rect 18300 -4425 18660 -4380
rect 19280 -4425 19640 -4380
rect 19900 -4425 20260 -4380
rect 20880 -4425 21240 -4380
rect 21500 -4425 21860 -4380
rect 22480 -4425 22840 -4380
rect 23100 -4425 23460 -4380
rect 24080 -4425 24440 -4380
rect 24700 -4425 25060 -4380
rect 25680 -4425 26040 -4380
rect 26300 -4425 26660 -4380
rect 27280 -4425 27640 -4380
rect 27900 -4425 28260 -4380
rect 28880 -4425 29240 -4380
rect 29500 -4425 29860 -4380
rect 30480 -4425 30840 -4380
rect 31100 -4425 31460 -4380
rect 32080 -4425 32440 -4380
rect 32700 -4425 33060 -4380
rect 33680 -4425 34040 -4380
rect 34300 -4425 34660 -4380
rect 35280 -4425 35640 -4380
rect 35900 -4425 36260 -4380
rect 16059 -4430 16459 -4425
rect 16059 -4460 16460 -4430
rect 16677 -4460 17077 -4425
rect 17659 -4430 18059 -4425
rect 17659 -4460 18060 -4430
rect 18277 -4460 18677 -4425
rect 19259 -4430 19659 -4425
rect 19259 -4460 19660 -4430
rect 19877 -4460 20277 -4425
rect 20859 -4430 21259 -4425
rect 20859 -4460 21260 -4430
rect 21477 -4460 21877 -4425
rect 22459 -4430 22859 -4425
rect 22459 -4460 22860 -4430
rect 23077 -4460 23477 -4425
rect 24059 -4430 24459 -4425
rect 24059 -4460 24460 -4430
rect 24677 -4460 25077 -4425
rect 25659 -4430 26059 -4425
rect 25659 -4460 26060 -4430
rect 26277 -4460 26677 -4425
rect 27259 -4430 27659 -4425
rect 27259 -4460 27660 -4430
rect 27877 -4460 28277 -4425
rect 28859 -4430 29259 -4425
rect 28859 -4460 29260 -4430
rect 29477 -4460 29877 -4425
rect 30459 -4430 30859 -4425
rect 30459 -4460 30860 -4430
rect 31077 -4460 31477 -4425
rect 32060 -4430 32459 -4425
rect 11880 -4480 12270 -4460
rect 16060 -4480 16460 -4460
rect 16680 -4480 17070 -4460
rect 17660 -4480 18060 -4460
rect 18280 -4480 18670 -4460
rect 19260 -4480 19660 -4460
rect 19880 -4480 20270 -4460
rect 20860 -4480 21260 -4460
rect 21480 -4480 21870 -4460
rect 22460 -4480 22860 -4460
rect 23080 -4480 23470 -4460
rect 24060 -4480 24460 -4460
rect 24680 -4480 25070 -4460
rect 25660 -4480 26060 -4460
rect 26280 -4480 26670 -4460
rect 27260 -4480 27660 -4460
rect 27880 -4480 28270 -4460
rect 28860 -4480 29260 -4460
rect 29480 -4480 29870 -4460
rect 30460 -4480 30860 -4460
rect 31080 -4480 31470 -4460
rect 11260 -4491 11659 -4490
rect 11877 -4491 12277 -4480
rect 16059 -4490 16460 -4480
rect 16059 -4491 16459 -4490
rect 16677 -4491 17077 -4480
rect 17659 -4490 18060 -4480
rect 17659 -4491 18059 -4490
rect 18277 -4491 18677 -4480
rect 19259 -4490 19660 -4480
rect 19259 -4491 19659 -4490
rect 19877 -4491 20277 -4480
rect 20859 -4490 21260 -4480
rect 20859 -4491 21259 -4490
rect 21477 -4491 21877 -4480
rect 22459 -4490 22860 -4480
rect 22459 -4491 22859 -4490
rect 23077 -4491 23477 -4480
rect 24059 -4490 24460 -4480
rect 24059 -4491 24459 -4490
rect 24677 -4491 25077 -4480
rect 25659 -4490 26060 -4480
rect 25659 -4491 26059 -4490
rect 26277 -4491 26677 -4480
rect 27259 -4490 27660 -4480
rect 27259 -4491 27659 -4490
rect 27877 -4491 28277 -4480
rect 28859 -4490 29260 -4480
rect 28859 -4491 29259 -4490
rect 29477 -4491 29877 -4480
rect 30459 -4490 30860 -4480
rect 30459 -4491 30859 -4490
rect 31077 -4491 31477 -4480
rect 32060 -4490 32460 -4430
rect 32677 -4460 33077 -4425
rect 33659 -4430 34059 -4425
rect 33659 -4460 34060 -4430
rect 34277 -4460 34677 -4425
rect 35259 -4430 35659 -4425
rect 35259 -4460 35660 -4430
rect 35877 -4460 36277 -4425
rect 32680 -4480 33070 -4460
rect 33660 -4480 34060 -4460
rect 34280 -4480 34670 -4460
rect 35260 -4480 35660 -4460
rect 35880 -4480 36270 -4460
rect 32677 -4491 33077 -4480
rect 33659 -4490 34060 -4480
rect 33659 -4491 34059 -4490
rect 34277 -4491 34677 -4480
rect 35259 -4490 35660 -4480
rect 35259 -4491 35659 -4490
rect 35877 -4491 36277 -4480
rect 12320 -4530 12520 -4520
rect 1540 -4650 12390 -4530
rect 12510 -4650 36400 -4530
rect 1540 -4660 36400 -4650
rect 30459 -4709 30859 -4703
rect 440 -4800 710 -4780
rect 1180 -4720 1320 -4710
rect 2780 -4720 2920 -4710
rect 4380 -4720 4520 -4710
rect 5980 -4720 6120 -4710
rect 7580 -4720 7720 -4710
rect 9180 -4720 9320 -4710
rect 15810 -4720 15930 -4710
rect 17410 -4720 17530 -4710
rect 19010 -4720 19130 -4710
rect 20610 -4720 20730 -4710
rect 22210 -4720 22330 -4710
rect 23810 -4720 23930 -4710
rect 25410 -4720 25530 -4710
rect 27011 -4720 27130 -4710
rect 28611 -4720 28730 -4710
rect 30211 -4720 30330 -4710
rect 30459 -4720 30471 -4709
rect 30847 -4720 30859 -4709
rect 31077 -4709 31477 -4703
rect 31077 -4720 31089 -4709
rect 1180 -4840 1190 -4720
rect 1310 -4840 2790 -4720
rect 2910 -4840 4390 -4720
rect 4510 -4840 5990 -4720
rect 6110 -4840 7590 -4720
rect 7710 -4840 9190 -4720
rect 9310 -4840 10720 -4720
rect 11220 -4810 12350 -4720
rect 11220 -4840 11710 -4810
rect 1180 -4850 1320 -4840
rect 2780 -4850 2920 -4840
rect 4380 -4850 4520 -4840
rect 5980 -4850 6120 -4840
rect 7580 -4850 7720 -4840
rect 9180 -4850 9320 -4840
rect 11700 -4930 11710 -4840
rect 11830 -4840 12350 -4810
rect 12600 -4730 12740 -4720
rect 11830 -4930 11840 -4840
rect 12600 -4850 12610 -4730
rect 12730 -4740 12740 -4730
rect 12730 -4840 13260 -4740
rect 13470 -4790 13890 -4720
rect 13470 -4840 13630 -4790
rect 12730 -4850 12740 -4840
rect 12600 -4860 12740 -4850
rect 13620 -4910 13630 -4840
rect 13750 -4840 13890 -4790
rect 14200 -4730 14340 -4720
rect 13750 -4910 13760 -4840
rect 14200 -4850 14210 -4730
rect 14330 -4740 14340 -4730
rect 14330 -4840 14860 -4740
rect 15070 -4790 15490 -4720
rect 15070 -4840 15230 -4790
rect 14330 -4850 14340 -4840
rect 14200 -4860 14340 -4850
rect 13620 -4920 13760 -4910
rect 15220 -4910 15230 -4840
rect 15350 -4840 15490 -4790
rect 15810 -4840 15820 -4720
rect 15920 -4840 17120 -4720
rect 17410 -4840 17420 -4720
rect 17520 -4840 18720 -4720
rect 19010 -4840 19020 -4720
rect 19120 -4840 20320 -4720
rect 20610 -4840 20620 -4720
rect 20720 -4840 21920 -4720
rect 22210 -4840 22220 -4720
rect 22320 -4840 23520 -4720
rect 23810 -4840 23820 -4720
rect 23920 -4840 25120 -4720
rect 25410 -4840 25420 -4720
rect 25520 -4840 26720 -4720
rect 27011 -4840 27020 -4720
rect 27120 -4840 28320 -4720
rect 28611 -4840 28620 -4720
rect 28720 -4840 29920 -4720
rect 30211 -4840 30220 -4720
rect 30320 -4743 31089 -4720
rect 31465 -4720 31477 -4709
rect 36390 -4710 36510 -4700
rect 36390 -4720 36400 -4710
rect 31465 -4743 31520 -4720
rect 30320 -4840 31520 -4743
rect 32060 -4830 36400 -4720
rect 36500 -4830 36510 -4710
rect 32060 -4840 36510 -4830
rect 15350 -4910 15360 -4840
rect 15810 -4850 15930 -4840
rect 17410 -4850 17530 -4840
rect 19010 -4850 19130 -4840
rect 20610 -4850 20730 -4840
rect 22210 -4850 22330 -4840
rect 23810 -4850 23930 -4840
rect 25410 -4850 25530 -4840
rect 27011 -4850 27130 -4840
rect 28611 -4850 28730 -4840
rect 30211 -4850 30330 -4840
rect 15220 -4920 15360 -4910
rect 11700 -4940 11840 -4930
rect 11700 -5830 11840 -5820
rect 11700 -5950 11710 -5830
rect 11830 -5840 11840 -5830
rect 13300 -5830 13440 -5820
rect 13300 -5840 13310 -5830
rect 11830 -5940 13310 -5840
rect 11830 -5950 11840 -5940
rect 11700 -5960 11840 -5950
rect 13300 -5950 13310 -5940
rect 13430 -5950 13440 -5830
rect 13300 -5960 13440 -5950
rect 11700 -6050 11840 -6040
rect 11700 -6170 11710 -6050
rect 11830 -6060 11840 -6050
rect 13620 -6050 13760 -6040
rect 13620 -6060 13630 -6050
rect 11830 -6160 13630 -6060
rect 11830 -6170 11840 -6160
rect 11700 -6180 11840 -6170
rect 13620 -6170 13630 -6160
rect 13750 -6170 13760 -6050
rect 13620 -6180 13760 -6170
rect 14220 -6050 14360 -6040
rect 14220 -6170 14230 -6050
rect 14350 -6060 14360 -6050
rect 15220 -6050 15360 -6040
rect 15220 -6060 15230 -6050
rect 14350 -6160 15230 -6060
rect 14350 -6170 14360 -6160
rect 14220 -6180 14360 -6170
rect 15220 -6170 15230 -6160
rect 15350 -6170 15360 -6050
rect 15220 -6180 15360 -6170
rect 12620 -6270 12760 -6260
rect 12620 -6390 12630 -6270
rect 12750 -6280 12760 -6270
rect 16500 -6270 16640 -6260
rect 16500 -6280 16510 -6270
rect 12750 -6380 16510 -6280
rect 12750 -6390 12760 -6380
rect 12620 -6400 12760 -6390
rect 16500 -6390 16510 -6380
rect 16630 -6390 16640 -6270
rect 16500 -6400 16640 -6390
rect 12400 -6490 12540 -6480
rect 12400 -6610 12410 -6490
rect 12530 -6500 12540 -6490
rect 14900 -6490 15040 -6480
rect 14900 -6500 14910 -6490
rect 12530 -6600 14910 -6500
rect 12530 -6610 12540 -6600
rect 12400 -6620 12540 -6610
rect 14900 -6610 14910 -6600
rect 15030 -6610 15040 -6490
rect 14900 -6620 15040 -6610
rect 12940 -6830 13120 -6820
rect 12940 -6900 12950 -6830
rect 440 -6990 12950 -6900
rect 13110 -6990 13120 -6830
rect 440 -8090 720 -6990
rect 12940 -7000 13120 -6990
rect 7800 -7870 7940 -7860
rect 7800 -7990 7810 -7870
rect 7930 -7880 7940 -7870
rect 14900 -7880 15050 -7870
rect 7930 -7990 14910 -7880
rect 7800 -8000 14910 -7990
rect 15040 -8000 15050 -7880
rect 14900 -8010 15050 -8000
rect 440 -9580 490 -8090
rect 0 -9600 490 -9580
rect -1349 -9800 490 -9600
rect -1349 -11400 -1300 -9800
rect 0 -9820 490 -9800
rect 440 -11360 490 -9820
rect 20 -11400 490 -11360
rect -1349 -11600 490 -11400
rect -1349 -13200 -1300 -11600
rect 0 -11620 490 -11600
rect 440 -13180 490 -11620
rect 0 -13200 490 -13180
rect -1349 -13400 490 -13200
rect -1349 -15000 -1300 -13400
rect 0 -13420 490 -13400
rect 440 -14980 490 -13420
rect 0 -15000 490 -14980
rect -1349 -15200 490 -15000
rect -1349 -16800 -1300 -15200
rect 0 -15220 490 -15200
rect 440 -16760 490 -15220
rect 0 -16800 490 -16760
rect -1349 -17000 490 -16800
rect -1349 -18600 -1300 -17000
rect 0 -17020 490 -17000
rect 440 -18560 490 -17020
rect 0 -18600 490 -18560
rect -1349 -18800 490 -18600
rect -1349 -20400 -1300 -18800
rect 0 -18820 490 -18800
rect 440 -20380 490 -18820
rect 0 -20400 490 -20380
rect -1349 -20600 490 -20400
rect -1349 -22200 -1300 -20600
rect 0 -20620 490 -20600
rect 440 -22160 490 -20620
rect 0 -22200 490 -22160
rect -1349 -22380 490 -22200
rect 670 -9580 720 -8090
rect 1200 -8070 1340 -8060
rect 1200 -8190 1210 -8070
rect 1330 -8080 1340 -8070
rect 2800 -8070 2940 -8060
rect 2800 -8080 2810 -8070
rect 1330 -8180 2810 -8080
rect 1330 -8190 1340 -8180
rect 1200 -8200 1340 -8190
rect 2800 -8190 2810 -8180
rect 2930 -8080 2940 -8070
rect 4400 -8070 4540 -8060
rect 4400 -8080 4410 -8070
rect 2930 -8180 4410 -8080
rect 2930 -8190 2940 -8180
rect 2800 -8200 2940 -8190
rect 4400 -8190 4410 -8180
rect 4530 -8080 4540 -8070
rect 6000 -8070 6140 -8060
rect 6000 -8080 6010 -8070
rect 4530 -8180 6010 -8080
rect 4530 -8190 4540 -8180
rect 4400 -8200 4540 -8190
rect 6000 -8190 6010 -8180
rect 6130 -8080 6140 -8070
rect 7600 -8070 7740 -8060
rect 7600 -8080 7610 -8070
rect 6130 -8180 7610 -8080
rect 6130 -8190 6140 -8180
rect 6000 -8200 6140 -8190
rect 7600 -8190 7610 -8180
rect 7730 -8080 7740 -8070
rect 9200 -8070 9340 -8060
rect 9200 -8080 9210 -8070
rect 7730 -8180 9210 -8080
rect 7730 -8190 7740 -8180
rect 7600 -8200 7740 -8190
rect 9200 -8190 9210 -8180
rect 9330 -8080 9340 -8070
rect 15820 -8070 15960 -8060
rect 9330 -8180 10700 -8080
rect 11270 -8110 15480 -8100
rect 9330 -8190 9340 -8180
rect 9200 -8200 9340 -8190
rect 11270 -8200 11710 -8110
rect 11690 -8230 11710 -8200
rect 11840 -8200 15480 -8110
rect 15820 -8190 15830 -8070
rect 15950 -8100 15960 -8070
rect 17420 -8070 17560 -8060
rect 15950 -8190 17090 -8100
rect 15820 -8200 17090 -8190
rect 17420 -8190 17430 -8070
rect 17550 -8100 17560 -8070
rect 19020 -8070 19160 -8060
rect 17550 -8190 18690 -8100
rect 17420 -8200 18690 -8190
rect 19020 -8190 19030 -8070
rect 19150 -8100 19160 -8070
rect 20620 -8070 20760 -8060
rect 19150 -8190 20290 -8100
rect 19020 -8200 20290 -8190
rect 20620 -8190 20630 -8070
rect 20750 -8100 20760 -8070
rect 22220 -8070 22360 -8060
rect 20750 -8190 21890 -8100
rect 20620 -8200 21890 -8190
rect 22220 -8190 22230 -8070
rect 22350 -8100 22360 -8070
rect 23820 -8070 23960 -8060
rect 22350 -8190 23490 -8100
rect 22220 -8200 23490 -8190
rect 23820 -8190 23830 -8070
rect 23950 -8100 23960 -8070
rect 25420 -8070 25560 -8060
rect 23950 -8190 25090 -8100
rect 23820 -8200 25090 -8190
rect 25420 -8190 25430 -8070
rect 25550 -8100 25560 -8070
rect 27020 -8070 27160 -8060
rect 25550 -8190 26680 -8100
rect 25420 -8200 26680 -8190
rect 27020 -8190 27030 -8070
rect 27150 -8100 27160 -8070
rect 28620 -8070 28760 -8060
rect 27150 -8190 28290 -8100
rect 27020 -8200 28290 -8190
rect 28620 -8190 28630 -8070
rect 28750 -8100 28760 -8070
rect 30220 -8070 30360 -8060
rect 28750 -8190 29890 -8100
rect 28620 -8200 29890 -8190
rect 30220 -8190 30230 -8070
rect 30350 -8100 30360 -8070
rect 31820 -8070 31960 -8060
rect 30350 -8164 31490 -8100
rect 30350 -8190 31493 -8164
rect 30220 -8200 31493 -8190
rect 31820 -8190 31830 -8070
rect 31950 -8100 31960 -8070
rect 34800 -8070 34940 -8060
rect 34800 -8100 34810 -8070
rect 31950 -8190 34810 -8100
rect 34930 -8100 34940 -8070
rect 34930 -8190 36280 -8100
rect 31820 -8200 36280 -8190
rect 11840 -8230 11860 -8200
rect 11690 -8240 11860 -8230
rect 13290 -8240 13460 -8200
rect 14890 -8240 15060 -8200
rect 30457 -8204 30469 -8200
rect 30845 -8204 30857 -8200
rect 30457 -8210 30857 -8204
rect 31093 -8204 31105 -8200
rect 31481 -8204 31493 -8200
rect 31093 -8210 31493 -8204
rect 32057 -8204 32069 -8200
rect 32057 -8210 32140 -8204
rect 10750 -8260 10940 -8250
rect 1560 -8380 10810 -8260
rect 10930 -8380 10940 -8260
rect 10750 -8390 10940 -8380
rect 11180 -8390 15570 -8240
rect 30370 -8249 30416 -8237
rect 16500 -8260 16650 -8250
rect 30370 -8260 30376 -8249
rect 30410 -8260 30416 -8249
rect 30898 -8249 30944 -8237
rect 30898 -8260 30904 -8249
rect 30938 -8260 30944 -8249
rect 31006 -8249 31052 -8237
rect 31006 -8260 31012 -8249
rect 31046 -8260 31052 -8249
rect 31534 -8260 31540 -8257
rect 15970 -8380 16510 -8260
rect 16640 -8380 36380 -8260
rect 16500 -8390 16650 -8380
rect 30370 -8383 30376 -8380
rect 30410 -8383 30416 -8380
rect 30370 -8395 30416 -8383
rect 30898 -8383 30904 -8380
rect 30938 -8383 30944 -8380
rect 30898 -8395 30944 -8383
rect 31006 -8383 31012 -8380
rect 31046 -8383 31052 -8380
rect 31006 -8395 31052 -8383
rect 30457 -8428 30857 -8422
rect 30457 -8430 30469 -8428
rect 30845 -8430 30857 -8428
rect 1420 -8510 1560 -8500
rect 1420 -8630 1430 -8510
rect 1550 -8520 1560 -8510
rect 1660 -8520 2060 -8430
rect 2290 -8520 2690 -8430
rect 3020 -8510 3160 -8500
rect 3020 -8520 3030 -8510
rect 1550 -8620 3030 -8520
rect 1550 -8630 1560 -8620
rect 1420 -8640 1560 -8630
rect 1660 -8640 2690 -8620
rect 3020 -8630 3030 -8620
rect 3150 -8520 3160 -8510
rect 3260 -8520 3660 -8430
rect 3890 -8520 4290 -8430
rect 4620 -8510 4760 -8500
rect 4620 -8520 4630 -8510
rect 3150 -8620 4630 -8520
rect 3150 -8630 3160 -8620
rect 3020 -8640 3160 -8630
rect 3260 -8640 4290 -8620
rect 4620 -8630 4630 -8620
rect 4750 -8520 4760 -8510
rect 4860 -8520 5260 -8430
rect 5490 -8520 5890 -8430
rect 6220 -8510 6360 -8500
rect 6220 -8520 6230 -8510
rect 4750 -8620 6230 -8520
rect 4750 -8630 4760 -8620
rect 4620 -8640 4760 -8630
rect 4860 -8640 5890 -8620
rect 6220 -8630 6230 -8620
rect 6350 -8520 6360 -8510
rect 6460 -8520 6860 -8430
rect 7090 -8520 7490 -8430
rect 7820 -8510 7960 -8500
rect 7820 -8520 7830 -8510
rect 6350 -8620 7830 -8520
rect 6350 -8630 6360 -8620
rect 6220 -8640 6360 -8630
rect 6460 -8640 7490 -8620
rect 7820 -8630 7830 -8620
rect 7950 -8520 7960 -8510
rect 8060 -8520 8460 -8430
rect 8690 -8520 9090 -8430
rect 9420 -8510 9560 -8500
rect 9420 -8520 9430 -8510
rect 7950 -8620 9430 -8520
rect 7950 -8630 7960 -8620
rect 7820 -8640 7960 -8630
rect 8060 -8640 9090 -8620
rect 9420 -8630 9430 -8620
rect 9550 -8520 9560 -8510
rect 9660 -8520 10060 -8430
rect 10290 -8520 10690 -8430
rect 11260 -8490 15490 -8430
rect 9550 -8620 10690 -8520
rect 9550 -8630 9560 -8620
rect 9420 -8640 9560 -8630
rect 9660 -8640 10690 -8620
rect 1660 -8730 2060 -8640
rect 2290 -8730 2690 -8640
rect 3260 -8730 3660 -8640
rect 3890 -8730 4290 -8640
rect 4860 -8730 5260 -8640
rect 5490 -8730 5890 -8640
rect 6460 -8730 6860 -8640
rect 7090 -8730 7490 -8640
rect 8060 -8730 8460 -8640
rect 8690 -8730 9090 -8640
rect 9660 -8730 10060 -8640
rect 10290 -8730 10690 -8640
rect 11420 -8650 11480 -8490
rect 12070 -8650 12130 -8490
rect 11260 -8730 12290 -8650
rect 2120 -8810 2240 -8800
rect 2120 -9470 2130 -8810
rect 2230 -9470 2240 -8810
rect 2120 -9480 2240 -9470
rect 3720 -8810 3840 -8800
rect 3720 -9470 3730 -8810
rect 3830 -9470 3840 -8810
rect 3720 -9480 3840 -9470
rect 5320 -8810 5440 -8800
rect 5320 -9470 5330 -8810
rect 5430 -9470 5440 -8810
rect 5320 -9480 5440 -9470
rect 6920 -8810 7040 -8800
rect 6920 -9470 6930 -8810
rect 7030 -9470 7040 -8810
rect 6920 -9480 7040 -9470
rect 8520 -8810 8640 -8800
rect 8520 -9470 8530 -8810
rect 8630 -9470 8640 -8810
rect 8520 -9480 8640 -9470
rect 10120 -8810 10240 -8800
rect 10120 -9470 10130 -8810
rect 10230 -9470 10240 -8810
rect 10120 -9480 10240 -9470
rect 11710 -8810 11840 -8800
rect 11710 -9470 11720 -8810
rect 11830 -9470 11840 -8810
rect 11710 -9480 11840 -9470
rect 12480 -9550 12680 -8490
rect 15600 -8520 15740 -8510
rect 12860 -8730 15490 -8630
rect 15600 -8640 15610 -8520
rect 15730 -8530 15740 -8520
rect 16060 -8530 16450 -8430
rect 16700 -8530 17090 -8430
rect 15730 -8630 17090 -8530
rect 15730 -8640 15740 -8630
rect 15600 -8650 15740 -8640
rect 16060 -8730 16450 -8630
rect 16700 -8730 17090 -8630
rect 17200 -8520 17340 -8510
rect 17200 -8640 17210 -8520
rect 17330 -8530 17340 -8520
rect 17660 -8530 18050 -8430
rect 18300 -8530 18690 -8430
rect 17330 -8630 18690 -8530
rect 17330 -8640 17340 -8630
rect 17200 -8650 17340 -8640
rect 17660 -8730 18050 -8630
rect 18300 -8730 18690 -8630
rect 18800 -8520 18940 -8510
rect 18800 -8640 18810 -8520
rect 18930 -8530 18940 -8520
rect 19260 -8530 19650 -8430
rect 19900 -8530 20290 -8430
rect 18930 -8630 20290 -8530
rect 18930 -8640 18940 -8630
rect 18800 -8650 18940 -8640
rect 19260 -8730 19650 -8630
rect 19900 -8730 20290 -8630
rect 20400 -8520 20540 -8510
rect 20400 -8640 20410 -8520
rect 20530 -8530 20540 -8520
rect 20860 -8530 21250 -8430
rect 21500 -8530 21890 -8430
rect 20530 -8630 21890 -8530
rect 20530 -8640 20540 -8630
rect 20400 -8650 20540 -8640
rect 20860 -8730 21250 -8630
rect 21500 -8730 21890 -8630
rect 22000 -8520 22140 -8510
rect 22000 -8640 22010 -8520
rect 22130 -8530 22140 -8520
rect 22460 -8530 22850 -8430
rect 23100 -8530 23490 -8430
rect 22130 -8630 23490 -8530
rect 22130 -8640 22140 -8630
rect 22000 -8650 22140 -8640
rect 22460 -8730 22850 -8630
rect 23100 -8730 23490 -8630
rect 23600 -8520 23740 -8510
rect 23600 -8640 23610 -8520
rect 23730 -8530 23740 -8520
rect 24060 -8530 24450 -8430
rect 24700 -8530 25090 -8430
rect 23730 -8630 25090 -8530
rect 23730 -8640 23740 -8630
rect 23600 -8650 23740 -8640
rect 24060 -8730 24450 -8630
rect 24700 -8730 25090 -8630
rect 25200 -8520 25340 -8510
rect 25200 -8640 25210 -8520
rect 25330 -8530 25340 -8520
rect 25660 -8530 26050 -8430
rect 26300 -8530 26690 -8430
rect 27260 -8468 27657 -8430
rect 27893 -8468 28290 -8430
rect 25330 -8630 26690 -8530
rect 25330 -8640 25340 -8630
rect 25200 -8650 25340 -8640
rect 25660 -8730 26050 -8630
rect 26300 -8730 26690 -8630
rect 26800 -8520 26940 -8510
rect 26800 -8640 26810 -8520
rect 26930 -8530 26940 -8520
rect 27260 -8530 27650 -8468
rect 27900 -8530 28290 -8468
rect 28860 -8468 29257 -8430
rect 29493 -8468 29890 -8430
rect 30457 -8468 30857 -8430
rect 31093 -8428 31493 -8422
rect 31093 -8430 31105 -8428
rect 31481 -8430 31493 -8428
rect 31093 -8468 31493 -8430
rect 32060 -8468 32457 -8430
rect 32693 -8468 33090 -8430
rect 26930 -8630 28290 -8530
rect 26930 -8640 26940 -8630
rect 26800 -8650 26940 -8640
rect 27260 -8690 27650 -8630
rect 27900 -8690 28290 -8630
rect 28400 -8520 28540 -8510
rect 28400 -8640 28410 -8520
rect 28530 -8530 28540 -8520
rect 28860 -8530 29250 -8468
rect 29500 -8530 29890 -8468
rect 28530 -8630 29890 -8530
rect 28530 -8640 28540 -8630
rect 28400 -8650 28540 -8640
rect 27260 -8730 27657 -8690
rect 27893 -8730 28290 -8690
rect 28860 -8690 29250 -8630
rect 29500 -8690 29890 -8630
rect 30000 -8520 30140 -8510
rect 30000 -8640 30010 -8520
rect 30130 -8530 30140 -8520
rect 30460 -8530 30850 -8468
rect 31100 -8530 31490 -8468
rect 30130 -8630 31490 -8530
rect 30130 -8640 30140 -8630
rect 30000 -8650 30140 -8640
rect 28860 -8730 29257 -8690
rect 29493 -8730 29890 -8690
rect 30460 -8690 30850 -8630
rect 31100 -8690 31490 -8630
rect 30460 -8730 30857 -8690
rect 31093 -8730 31490 -8690
rect 32060 -8530 32450 -8468
rect 32700 -8530 33090 -8468
rect 33660 -8468 34057 -8430
rect 34293 -8468 34690 -8430
rect 33660 -8530 34050 -8468
rect 34300 -8530 34690 -8468
rect 35260 -8468 35657 -8430
rect 35893 -8468 36290 -8430
rect 35260 -8530 35650 -8468
rect 35900 -8530 36290 -8468
rect 32060 -8630 36290 -8530
rect 32060 -8690 32450 -8630
rect 32700 -8690 33090 -8630
rect 33660 -8690 34050 -8630
rect 34300 -8690 34690 -8630
rect 35260 -8690 35650 -8630
rect 35900 -8690 36290 -8630
rect 32060 -8730 32457 -8690
rect 13310 -8810 13440 -8730
rect 13310 -9470 13320 -8810
rect 13430 -9470 13440 -8810
rect 13310 -9480 13440 -9470
rect 14910 -9480 15040 -8730
rect 32340 -8736 32457 -8730
rect 32693 -8736 33093 -8690
rect 33657 -8736 34057 -8690
rect 34293 -8736 34693 -8690
rect 35257 -8736 35657 -8690
rect 35893 -8730 36290 -8690
rect 35893 -8736 36030 -8730
rect 32498 -8790 32544 -8784
rect 32606 -8790 32652 -8784
rect 16510 -8800 16640 -8790
rect 16510 -9480 16520 -8800
rect 16630 -9480 16640 -8800
rect 16510 -9490 16640 -9480
rect 18110 -8800 18240 -8790
rect 18110 -9480 18120 -8800
rect 18230 -9480 18240 -8800
rect 18110 -9490 18240 -9480
rect 19710 -8800 19840 -8790
rect 19710 -9480 19720 -8800
rect 19830 -9480 19840 -8800
rect 19710 -9490 19840 -9480
rect 21310 -8800 21440 -8790
rect 21310 -9480 21320 -8800
rect 21430 -9480 21440 -8800
rect 21310 -9490 21440 -9480
rect 22910 -8800 23040 -8790
rect 22910 -9480 22920 -8800
rect 23030 -9480 23040 -8800
rect 22910 -9490 23040 -9480
rect 24510 -8800 24640 -8790
rect 24510 -9480 24520 -8800
rect 24630 -9480 24640 -8800
rect 24510 -9490 24640 -9480
rect 26110 -8800 26240 -8790
rect 26110 -9480 26120 -8800
rect 26230 -9480 26240 -8800
rect 26110 -9490 26240 -9480
rect 27710 -8800 27840 -8790
rect 27710 -9480 27720 -8800
rect 27830 -9480 27840 -8800
rect 27710 -9490 27840 -9480
rect 29310 -8800 29440 -8790
rect 29310 -9480 29320 -8800
rect 29430 -9480 29440 -8800
rect 29310 -9490 29440 -9480
rect 30910 -8800 31040 -8790
rect 30910 -9480 30920 -8800
rect 31030 -9480 31040 -8800
rect 32498 -8796 32652 -8790
rect 32498 -9360 32504 -8796
rect 32510 -8800 32640 -8796
rect 32510 -9360 32520 -8800
rect 32630 -9360 32640 -8800
rect 32646 -9360 32652 -8796
rect 33134 -8796 33180 -8784
rect 33134 -9360 33140 -8796
rect 33174 -9360 33180 -8796
rect 33570 -8796 33616 -8784
rect 33570 -9360 33576 -8796
rect 33610 -9360 33616 -8796
rect 34098 -8790 34144 -8784
rect 34206 -8790 34252 -8784
rect 34098 -8796 34252 -8790
rect 34098 -9360 34104 -8796
rect 34110 -8800 34240 -8796
rect 34110 -9360 34120 -8800
rect 34230 -9360 34240 -8800
rect 34246 -9360 34252 -8796
rect 34734 -8796 34780 -8784
rect 34734 -9360 34740 -8796
rect 34774 -9360 34780 -8796
rect 35170 -8796 35216 -8784
rect 35170 -9360 35176 -8796
rect 35210 -9360 35216 -8796
rect 35698 -8790 35744 -8784
rect 35806 -8790 35852 -8784
rect 35698 -8796 35852 -8790
rect 35698 -9360 35704 -8796
rect 35710 -8800 35840 -8796
rect 35710 -9360 35720 -8800
rect 35830 -9360 35840 -8800
rect 35846 -9360 35852 -8796
rect 39100 -9400 39229 8940
rect 30910 -9490 31040 -9480
rect 33400 -9510 33540 -9500
rect 33400 -9550 33410 -9510
rect 670 -9700 12420 -9580
rect 12480 -9620 15490 -9550
rect 15700 -9700 31760 -9580
rect 32060 -9630 33410 -9550
rect 33530 -9550 33540 -9510
rect 33530 -9630 36290 -9550
rect 32060 -9640 36290 -9630
rect 36700 -9700 39229 -9400
rect 670 -9800 39229 -9700
rect 670 -9820 37940 -9800
rect 670 -11360 720 -9820
rect 1200 -9870 1340 -9860
rect 1200 -9990 1210 -9870
rect 1330 -9880 1340 -9870
rect 2800 -9870 2940 -9860
rect 2800 -9880 2810 -9870
rect 1330 -9980 2810 -9880
rect 1330 -9990 1340 -9980
rect 1200 -10000 1340 -9990
rect 2800 -9990 2810 -9980
rect 2930 -9880 2940 -9870
rect 4400 -9870 4540 -9860
rect 4400 -9880 4410 -9870
rect 2930 -9980 4410 -9880
rect 2930 -9990 2940 -9980
rect 2800 -10000 2940 -9990
rect 4400 -9990 4410 -9980
rect 4530 -9880 4540 -9870
rect 6000 -9870 6140 -9860
rect 6000 -9880 6010 -9870
rect 4530 -9980 6010 -9880
rect 4530 -9990 4540 -9980
rect 4400 -10000 4540 -9990
rect 6000 -9990 6010 -9980
rect 6130 -9880 6140 -9870
rect 7600 -9870 7740 -9860
rect 7600 -9880 7610 -9870
rect 6130 -9980 7610 -9880
rect 6130 -9990 6140 -9980
rect 6000 -10000 6140 -9990
rect 7600 -9990 7610 -9980
rect 7730 -9880 7740 -9870
rect 9200 -9870 9340 -9860
rect 9200 -9880 9210 -9870
rect 7730 -9980 9210 -9880
rect 7730 -9990 7740 -9980
rect 7600 -10000 7740 -9990
rect 9200 -9990 9210 -9980
rect 9330 -9880 9340 -9870
rect 15820 -9870 15960 -9860
rect 9330 -9980 10700 -9880
rect 9330 -9990 9340 -9980
rect 9200 -10000 9340 -9990
rect 10750 -10060 10940 -10050
rect 11400 -10060 11520 -9980
rect 12040 -10060 12160 -9980
rect 13000 -10060 13120 -9980
rect 13640 -10060 13760 -9980
rect 14600 -10060 14720 -9980
rect 15240 -10060 15360 -9980
rect 15820 -9990 15830 -9870
rect 15950 -9900 15960 -9870
rect 17420 -9870 17560 -9860
rect 15950 -9990 17090 -9900
rect 15820 -10000 17090 -9990
rect 17420 -9990 17430 -9870
rect 17550 -9900 17560 -9870
rect 19020 -9870 19160 -9860
rect 17550 -9990 18690 -9900
rect 17420 -10000 18690 -9990
rect 19020 -9990 19030 -9870
rect 19150 -9900 19160 -9870
rect 20620 -9870 20760 -9860
rect 19150 -9990 20290 -9900
rect 19020 -10000 20290 -9990
rect 20620 -9990 20630 -9870
rect 20750 -9900 20760 -9870
rect 22220 -9870 22360 -9860
rect 20750 -9990 21890 -9900
rect 20620 -10000 21890 -9990
rect 22220 -9990 22230 -9870
rect 22350 -9900 22360 -9870
rect 23820 -9870 23960 -9860
rect 22350 -9990 23490 -9900
rect 22220 -10000 23490 -9990
rect 23820 -9990 23830 -9870
rect 23950 -9900 23960 -9870
rect 25420 -9870 25560 -9860
rect 23950 -9990 25090 -9900
rect 23820 -10000 25090 -9990
rect 25420 -9990 25430 -9870
rect 25550 -9900 25560 -9870
rect 27020 -9870 27160 -9860
rect 25550 -9990 26680 -9900
rect 25420 -10000 26680 -9990
rect 27020 -9990 27030 -9870
rect 27150 -9900 27160 -9870
rect 28620 -9870 28760 -9860
rect 27150 -9990 28290 -9900
rect 27020 -10000 28290 -9990
rect 28620 -9990 28630 -9870
rect 28750 -9900 28760 -9870
rect 30220 -9870 30360 -9860
rect 28750 -9990 29890 -9900
rect 28620 -10000 29890 -9990
rect 30220 -9990 30230 -9870
rect 30350 -9900 30360 -9870
rect 31820 -9870 31960 -9860
rect 30350 -9964 31490 -9900
rect 30350 -9990 31493 -9964
rect 30220 -10000 31493 -9990
rect 31820 -9990 31830 -9870
rect 31950 -9900 31960 -9870
rect 34800 -9870 34940 -9860
rect 34800 -9900 34810 -9870
rect 31950 -9990 34810 -9900
rect 34930 -9900 34940 -9870
rect 34930 -9990 36280 -9900
rect 31820 -10000 36280 -9990
rect 30457 -10004 30469 -10000
rect 30845 -10004 30857 -10000
rect 30457 -10010 30857 -10004
rect 31093 -10004 31105 -10000
rect 31481 -10004 31493 -10000
rect 31093 -10010 31493 -10004
rect 32057 -10004 32069 -10000
rect 32057 -10010 32140 -10004
rect 30370 -10049 30416 -10037
rect 30370 -10060 30376 -10049
rect 30410 -10060 30416 -10049
rect 30898 -10049 30944 -10037
rect 30898 -10060 30904 -10049
rect 30938 -10060 30944 -10049
rect 31006 -10049 31052 -10037
rect 31006 -10060 31012 -10049
rect 31046 -10060 31052 -10049
rect 1560 -10180 10810 -10060
rect 10930 -10180 36380 -10060
rect 10750 -10190 10940 -10180
rect 1420 -10310 1560 -10300
rect 1420 -10430 1430 -10310
rect 1550 -10320 1560 -10310
rect 1660 -10320 2060 -10230
rect 2290 -10320 2690 -10230
rect 3020 -10310 3160 -10300
rect 3020 -10320 3030 -10310
rect 1550 -10420 3030 -10320
rect 1550 -10430 1560 -10420
rect 1420 -10440 1560 -10430
rect 1660 -10440 2690 -10420
rect 3020 -10430 3030 -10420
rect 3150 -10320 3160 -10310
rect 3260 -10320 3660 -10230
rect 3890 -10320 4290 -10230
rect 4620 -10310 4760 -10300
rect 4620 -10320 4630 -10310
rect 3150 -10420 4630 -10320
rect 3150 -10430 3160 -10420
rect 3020 -10440 3160 -10430
rect 3260 -10440 4290 -10420
rect 4620 -10430 4630 -10420
rect 4750 -10320 4760 -10310
rect 4860 -10320 5260 -10230
rect 5490 -10320 5890 -10230
rect 6220 -10310 6360 -10300
rect 6220 -10320 6230 -10310
rect 4750 -10420 6230 -10320
rect 4750 -10430 4760 -10420
rect 4620 -10440 4760 -10430
rect 4860 -10440 5890 -10420
rect 6220 -10430 6230 -10420
rect 6350 -10320 6360 -10310
rect 6460 -10320 6860 -10230
rect 7090 -10320 7490 -10230
rect 7820 -10310 7960 -10300
rect 7820 -10320 7830 -10310
rect 6350 -10420 7830 -10320
rect 6350 -10430 6360 -10420
rect 6220 -10440 6360 -10430
rect 6460 -10440 7490 -10420
rect 7820 -10430 7830 -10420
rect 7950 -10320 7960 -10310
rect 8060 -10320 8460 -10230
rect 8690 -10320 9090 -10230
rect 9420 -10310 9560 -10300
rect 9420 -10320 9430 -10310
rect 7950 -10420 9430 -10320
rect 7950 -10430 7960 -10420
rect 7820 -10440 7960 -10430
rect 8060 -10440 9090 -10420
rect 9420 -10430 9430 -10420
rect 9550 -10320 9560 -10310
rect 9660 -10320 10060 -10230
rect 10290 -10320 10690 -10230
rect 11400 -10260 11520 -10180
rect 12040 -10260 12160 -10180
rect 13000 -10260 13120 -10180
rect 13640 -10260 13760 -10180
rect 14600 -10260 14720 -10180
rect 15240 -10260 15360 -10180
rect 30370 -10183 30376 -10180
rect 30410 -10183 30416 -10180
rect 30370 -10195 30416 -10183
rect 30898 -10183 30904 -10180
rect 30938 -10183 30944 -10180
rect 30898 -10195 30944 -10183
rect 31006 -10183 31012 -10180
rect 31046 -10183 31052 -10180
rect 31006 -10195 31052 -10183
rect 30457 -10228 30857 -10222
rect 30457 -10230 30469 -10228
rect 30845 -10230 30857 -10228
rect 9550 -10420 10690 -10320
rect 15600 -10320 15740 -10310
rect 9550 -10430 9560 -10420
rect 9420 -10440 9560 -10430
rect 9660 -10440 10690 -10420
rect 1660 -10530 2060 -10440
rect 2290 -10530 2690 -10440
rect 3260 -10530 3660 -10440
rect 3890 -10530 4290 -10440
rect 4860 -10530 5260 -10440
rect 5490 -10530 5890 -10440
rect 6460 -10530 6860 -10440
rect 7090 -10530 7490 -10440
rect 8060 -10530 8460 -10440
rect 8690 -10530 9090 -10440
rect 9660 -10530 10060 -10440
rect 10290 -10530 10690 -10440
rect 11020 -10410 11160 -10400
rect 11020 -10530 11030 -10410
rect 11150 -10530 13890 -10410
rect 15600 -10440 15610 -10320
rect 15730 -10330 15740 -10320
rect 16060 -10330 16450 -10230
rect 16700 -10330 17090 -10230
rect 15730 -10430 17090 -10330
rect 15730 -10440 15740 -10430
rect 15600 -10450 15740 -10440
rect 11020 -10540 11160 -10530
rect 2120 -10610 2240 -10600
rect 2120 -11270 2130 -10610
rect 2230 -11270 2240 -10610
rect 2120 -11280 2240 -11270
rect 3720 -10610 3840 -10600
rect 3720 -11270 3730 -10610
rect 3830 -11270 3840 -10610
rect 3720 -11280 3840 -11270
rect 5320 -10610 5440 -10600
rect 5320 -11270 5330 -10610
rect 5430 -11270 5440 -10610
rect 5320 -11280 5440 -11270
rect 6920 -10610 7040 -10600
rect 6920 -11270 6930 -10610
rect 7030 -11270 7040 -10610
rect 6920 -11280 7040 -11270
rect 8520 -10610 8640 -10600
rect 8520 -11270 8530 -10610
rect 8630 -11270 8640 -10610
rect 8520 -11280 8640 -11270
rect 10120 -10610 10240 -10600
rect 10120 -11270 10130 -10610
rect 10230 -11270 10240 -10610
rect 10120 -11280 10240 -11270
rect 11710 -10610 11840 -10530
rect 11710 -11270 11720 -10610
rect 11830 -11270 11840 -10610
rect 11710 -11280 11840 -11270
rect 13310 -10610 13440 -10530
rect 13310 -11270 13320 -10610
rect 13430 -11270 13440 -10610
rect 14610 -10880 14740 -10510
rect 15220 -10880 15350 -10500
rect 16060 -10530 16450 -10430
rect 16700 -10530 17090 -10430
rect 17200 -10320 17340 -10310
rect 17200 -10440 17210 -10320
rect 17330 -10330 17340 -10320
rect 17660 -10330 18050 -10230
rect 18300 -10330 18690 -10230
rect 17330 -10430 18690 -10330
rect 17330 -10440 17340 -10430
rect 17200 -10450 17340 -10440
rect 17660 -10530 18050 -10430
rect 18300 -10530 18690 -10430
rect 18800 -10320 18940 -10310
rect 18800 -10440 18810 -10320
rect 18930 -10330 18940 -10320
rect 19260 -10330 19650 -10230
rect 19900 -10330 20290 -10230
rect 18930 -10430 20290 -10330
rect 18930 -10440 18940 -10430
rect 18800 -10450 18940 -10440
rect 19260 -10530 19650 -10430
rect 19900 -10530 20290 -10430
rect 20400 -10320 20540 -10310
rect 20400 -10440 20410 -10320
rect 20530 -10330 20540 -10320
rect 20860 -10330 21250 -10230
rect 21500 -10330 21890 -10230
rect 20530 -10430 21890 -10330
rect 20530 -10440 20540 -10430
rect 20400 -10450 20540 -10440
rect 20860 -10530 21250 -10430
rect 21500 -10530 21890 -10430
rect 22000 -10320 22140 -10310
rect 22000 -10440 22010 -10320
rect 22130 -10330 22140 -10320
rect 22460 -10330 22850 -10230
rect 23100 -10330 23490 -10230
rect 22130 -10430 23490 -10330
rect 22130 -10440 22140 -10430
rect 22000 -10450 22140 -10440
rect 22460 -10530 22850 -10430
rect 23100 -10530 23490 -10430
rect 23600 -10320 23740 -10310
rect 23600 -10440 23610 -10320
rect 23730 -10330 23740 -10320
rect 24060 -10330 24450 -10230
rect 24700 -10330 25090 -10230
rect 23730 -10430 25090 -10330
rect 23730 -10440 23740 -10430
rect 23600 -10450 23740 -10440
rect 24060 -10530 24450 -10430
rect 24700 -10530 25090 -10430
rect 25200 -10320 25340 -10310
rect 25200 -10440 25210 -10320
rect 25330 -10330 25340 -10320
rect 25660 -10330 26050 -10230
rect 26300 -10330 26690 -10230
rect 27260 -10268 27657 -10230
rect 27893 -10268 28290 -10230
rect 25330 -10430 26690 -10330
rect 25330 -10440 25340 -10430
rect 25200 -10450 25340 -10440
rect 25660 -10530 26050 -10430
rect 26300 -10530 26690 -10430
rect 26800 -10320 26940 -10310
rect 26800 -10440 26810 -10320
rect 26930 -10330 26940 -10320
rect 27260 -10330 27650 -10268
rect 27900 -10330 28290 -10268
rect 28860 -10268 29257 -10230
rect 29493 -10268 29890 -10230
rect 30457 -10268 30857 -10230
rect 31093 -10228 31493 -10222
rect 31093 -10230 31105 -10228
rect 31481 -10230 31493 -10228
rect 31093 -10268 31493 -10230
rect 32060 -10268 32457 -10230
rect 32693 -10268 33090 -10230
rect 26930 -10430 28290 -10330
rect 26930 -10440 26940 -10430
rect 26800 -10450 26940 -10440
rect 27260 -10490 27650 -10430
rect 27900 -10490 28290 -10430
rect 28400 -10320 28540 -10310
rect 28400 -10440 28410 -10320
rect 28530 -10330 28540 -10320
rect 28860 -10330 29250 -10268
rect 29500 -10330 29890 -10268
rect 28530 -10430 29890 -10330
rect 28530 -10440 28540 -10430
rect 28400 -10450 28540 -10440
rect 27260 -10530 27657 -10490
rect 27893 -10530 28290 -10490
rect 28860 -10490 29250 -10430
rect 29500 -10490 29890 -10430
rect 30000 -10320 30140 -10310
rect 30000 -10440 30010 -10320
rect 30130 -10330 30140 -10320
rect 30460 -10330 30850 -10268
rect 31100 -10330 31490 -10268
rect 30130 -10430 31490 -10330
rect 30130 -10440 30140 -10430
rect 30000 -10450 30140 -10440
rect 28860 -10530 29257 -10490
rect 29493 -10530 29890 -10490
rect 30460 -10490 30850 -10430
rect 31100 -10490 31490 -10430
rect 31600 -10320 31740 -10310
rect 31600 -10440 31610 -10320
rect 31730 -10330 31740 -10320
rect 32060 -10330 32450 -10268
rect 32700 -10330 33090 -10268
rect 33660 -10268 34057 -10230
rect 34293 -10268 34690 -10230
rect 33660 -10330 34050 -10268
rect 34300 -10330 34690 -10268
rect 35260 -10268 35657 -10230
rect 35893 -10268 36290 -10230
rect 35260 -10330 35650 -10268
rect 35900 -10330 36290 -10268
rect 31730 -10430 36290 -10330
rect 31730 -10440 31740 -10430
rect 31600 -10450 31740 -10440
rect 30460 -10530 30857 -10490
rect 31093 -10530 31490 -10490
rect 32060 -10490 32450 -10430
rect 32700 -10490 33090 -10430
rect 33660 -10490 34050 -10430
rect 34300 -10490 34690 -10430
rect 35260 -10490 35650 -10430
rect 35900 -10490 36290 -10430
rect 32060 -10530 32457 -10490
rect 32340 -10536 32457 -10530
rect 32693 -10536 33093 -10490
rect 33657 -10536 34057 -10490
rect 34293 -10536 34693 -10490
rect 35257 -10536 35657 -10490
rect 35893 -10530 36290 -10490
rect 35893 -10536 36030 -10530
rect 32498 -10590 32544 -10584
rect 32606 -10590 32652 -10584
rect 16510 -10600 16640 -10590
rect 14400 -11030 15570 -10880
rect 13310 -11280 13440 -11270
rect 14610 -11360 14740 -11030
rect 15220 -11360 15350 -11030
rect 16510 -11280 16520 -10600
rect 16630 -11280 16640 -10600
rect 16510 -11290 16640 -11280
rect 18110 -10600 18240 -10590
rect 18110 -11280 18120 -10600
rect 18230 -11280 18240 -10600
rect 18110 -11290 18240 -11280
rect 19710 -10600 19840 -10590
rect 19710 -11280 19720 -10600
rect 19830 -11280 19840 -10600
rect 19710 -11290 19840 -11280
rect 21310 -10600 21440 -10590
rect 21310 -11280 21320 -10600
rect 21430 -11280 21440 -10600
rect 21310 -11290 21440 -11280
rect 22910 -10600 23040 -10590
rect 22910 -11280 22920 -10600
rect 23030 -11280 23040 -10600
rect 22910 -11290 23040 -11280
rect 24510 -10600 24640 -10590
rect 24510 -11280 24520 -10600
rect 24630 -11280 24640 -10600
rect 24510 -11290 24640 -11280
rect 26110 -10600 26240 -10590
rect 26110 -11280 26120 -10600
rect 26230 -11280 26240 -10600
rect 26110 -11290 26240 -11280
rect 27710 -10600 27840 -10590
rect 27710 -11280 27720 -10600
rect 27830 -11280 27840 -10600
rect 27710 -11290 27840 -11280
rect 29310 -10600 29440 -10590
rect 29310 -11280 29320 -10600
rect 29430 -11280 29440 -10600
rect 29310 -11290 29440 -11280
rect 30910 -10600 31040 -10590
rect 30910 -11280 30920 -10600
rect 31030 -11280 31040 -10600
rect 32498 -10596 32652 -10590
rect 32498 -11110 32504 -10596
rect 32510 -10600 32640 -10596
rect 32510 -11110 32520 -10600
rect 32630 -11110 32640 -10600
rect 32646 -11110 32652 -10596
rect 33134 -10596 33180 -10584
rect 33134 -11110 33140 -10596
rect 33174 -11110 33180 -10596
rect 33570 -10596 33616 -10584
rect 33570 -11110 33576 -10596
rect 33610 -11110 33616 -10596
rect 34098 -10590 34144 -10584
rect 34206 -10590 34252 -10584
rect 34098 -10596 34252 -10590
rect 34098 -11110 34104 -10596
rect 34110 -10600 34240 -10596
rect 34110 -11110 34120 -10600
rect 34230 -11110 34240 -10600
rect 34246 -11110 34252 -10596
rect 34734 -10596 34780 -10584
rect 34734 -11110 34740 -10596
rect 34774 -11110 34780 -10596
rect 35170 -10596 35216 -10584
rect 35170 -11110 35176 -10596
rect 35210 -11110 35216 -10596
rect 35698 -10590 35744 -10584
rect 35806 -10590 35852 -10584
rect 35698 -10596 35852 -10590
rect 35698 -11110 35704 -10596
rect 35710 -10600 35840 -10596
rect 35710 -11110 35720 -10600
rect 35830 -11110 35840 -10600
rect 35846 -11110 35852 -10596
rect 30910 -11290 31040 -11280
rect 35000 -11310 35140 -11300
rect 35000 -11350 35010 -11310
rect 670 -11500 31880 -11360
rect 32060 -11430 35010 -11350
rect 35130 -11350 35140 -11310
rect 35130 -11430 36290 -11350
rect 32060 -11440 36290 -11430
rect 39100 -11500 39229 -9800
rect 670 -11600 39229 -11500
rect 670 -11620 37940 -11600
rect 670 -13180 720 -11620
rect 1200 -11670 1340 -11660
rect 1200 -11790 1210 -11670
rect 1330 -11680 1340 -11670
rect 2800 -11670 2940 -11660
rect 2800 -11680 2810 -11670
rect 1330 -11780 2810 -11680
rect 1330 -11790 1340 -11780
rect 1200 -11800 1340 -11790
rect 2800 -11790 2810 -11780
rect 2930 -11680 2940 -11670
rect 4400 -11670 4540 -11660
rect 4400 -11680 4410 -11670
rect 2930 -11780 4410 -11680
rect 2930 -11790 2940 -11780
rect 2800 -11800 2940 -11790
rect 4400 -11790 4410 -11780
rect 4530 -11680 4540 -11670
rect 6000 -11670 6140 -11660
rect 6000 -11680 6010 -11670
rect 4530 -11780 6010 -11680
rect 4530 -11790 4540 -11780
rect 4400 -11800 4540 -11790
rect 6000 -11790 6010 -11780
rect 6130 -11680 6140 -11670
rect 7600 -11670 7740 -11660
rect 7600 -11680 7610 -11670
rect 6130 -11780 7610 -11680
rect 6130 -11790 6140 -11780
rect 6000 -11800 6140 -11790
rect 7600 -11790 7610 -11780
rect 7730 -11680 7740 -11670
rect 9200 -11670 9340 -11660
rect 13300 -11670 13440 -11660
rect 14220 -11670 14360 -11660
rect 15820 -11670 15960 -11660
rect 9200 -11680 9210 -11670
rect 7730 -11780 9210 -11680
rect 7730 -11790 7740 -11780
rect 7600 -11800 7740 -11790
rect 9200 -11790 9210 -11780
rect 9330 -11680 9340 -11670
rect 9330 -11780 10700 -11680
rect 9330 -11790 9340 -11780
rect 9200 -11800 9340 -11790
rect 10750 -11860 10940 -11850
rect 11400 -11860 11520 -11780
rect 12040 -11860 12160 -11780
rect 12860 -11790 13310 -11670
rect 13430 -11790 14230 -11670
rect 14350 -11790 15490 -11670
rect 12860 -11800 15490 -11790
rect 15820 -11790 15830 -11670
rect 15950 -11700 15960 -11670
rect 17420 -11670 17560 -11660
rect 15950 -11790 17090 -11700
rect 15820 -11800 17090 -11790
rect 17420 -11790 17430 -11670
rect 17550 -11700 17560 -11670
rect 19020 -11670 19160 -11660
rect 17550 -11790 18690 -11700
rect 17420 -11800 18690 -11790
rect 19020 -11790 19030 -11670
rect 19150 -11700 19160 -11670
rect 20620 -11670 20760 -11660
rect 19150 -11790 20290 -11700
rect 19020 -11800 20290 -11790
rect 20620 -11790 20630 -11670
rect 20750 -11700 20760 -11670
rect 22220 -11670 22360 -11660
rect 20750 -11790 21890 -11700
rect 20620 -11800 21890 -11790
rect 22220 -11790 22230 -11670
rect 22350 -11700 22360 -11670
rect 23820 -11670 23960 -11660
rect 22350 -11790 23490 -11700
rect 22220 -11800 23490 -11790
rect 23820 -11790 23830 -11670
rect 23950 -11700 23960 -11670
rect 25420 -11670 25560 -11660
rect 23950 -11790 25090 -11700
rect 23820 -11800 25090 -11790
rect 25420 -11790 25430 -11670
rect 25550 -11700 25560 -11670
rect 27020 -11670 27160 -11660
rect 25550 -11790 26680 -11700
rect 25420 -11800 26680 -11790
rect 27020 -11790 27030 -11670
rect 27150 -11700 27160 -11670
rect 28620 -11670 28760 -11660
rect 27150 -11790 28290 -11700
rect 27020 -11800 28290 -11790
rect 28620 -11790 28630 -11670
rect 28750 -11700 28760 -11670
rect 30220 -11670 30360 -11660
rect 28750 -11790 29890 -11700
rect 28620 -11800 29890 -11790
rect 30220 -11790 30230 -11670
rect 30350 -11700 30360 -11670
rect 31820 -11670 31960 -11660
rect 30350 -11764 31490 -11700
rect 30350 -11790 31493 -11764
rect 30220 -11800 31493 -11790
rect 31820 -11790 31830 -11670
rect 31950 -11700 31960 -11670
rect 34800 -11670 34940 -11660
rect 34800 -11700 34810 -11670
rect 31950 -11790 34810 -11700
rect 34930 -11700 34940 -11670
rect 34930 -11790 36280 -11700
rect 31820 -11800 36280 -11790
rect 30457 -11804 30469 -11800
rect 30845 -11804 30857 -11800
rect 30457 -11810 30857 -11804
rect 31093 -11804 31105 -11800
rect 31481 -11804 31493 -11800
rect 31093 -11810 31493 -11804
rect 32057 -11804 32069 -11800
rect 32057 -11810 32140 -11804
rect 30370 -11849 30416 -11837
rect 30370 -11860 30376 -11849
rect 30410 -11860 30416 -11849
rect 30898 -11849 30944 -11837
rect 30898 -11860 30904 -11849
rect 30938 -11860 30944 -11849
rect 31006 -11849 31052 -11837
rect 31006 -11860 31012 -11849
rect 31046 -11860 31052 -11849
rect 1560 -11980 10810 -11860
rect 10930 -11980 36380 -11860
rect 10750 -11990 10940 -11980
rect 1420 -12110 1560 -12100
rect 1420 -12230 1430 -12110
rect 1550 -12120 1560 -12110
rect 1660 -12120 2060 -12030
rect 2290 -12120 2690 -12030
rect 3020 -12110 3160 -12100
rect 3020 -12120 3030 -12110
rect 1550 -12220 3030 -12120
rect 1550 -12230 1560 -12220
rect 1420 -12240 1560 -12230
rect 1660 -12240 2690 -12220
rect 3020 -12230 3030 -12220
rect 3150 -12120 3160 -12110
rect 3260 -12120 3660 -12030
rect 3890 -12120 4290 -12030
rect 4620 -12110 4760 -12100
rect 4620 -12120 4630 -12110
rect 3150 -12220 4630 -12120
rect 3150 -12230 3160 -12220
rect 3020 -12240 3160 -12230
rect 3260 -12240 4290 -12220
rect 4620 -12230 4630 -12220
rect 4750 -12120 4760 -12110
rect 4860 -12120 5260 -12030
rect 5490 -12120 5890 -12030
rect 6220 -12110 6360 -12100
rect 6220 -12120 6230 -12110
rect 4750 -12220 6230 -12120
rect 4750 -12230 4760 -12220
rect 4620 -12240 4760 -12230
rect 4860 -12240 5890 -12220
rect 6220 -12230 6230 -12220
rect 6350 -12120 6360 -12110
rect 6460 -12120 6860 -12030
rect 7090 -12120 7490 -12030
rect 7820 -12110 7960 -12100
rect 7820 -12120 7830 -12110
rect 6350 -12220 7830 -12120
rect 6350 -12230 6360 -12220
rect 6220 -12240 6360 -12230
rect 6460 -12240 7490 -12220
rect 7820 -12230 7830 -12220
rect 7950 -12120 7960 -12110
rect 8060 -12120 8460 -12030
rect 8690 -12120 9090 -12030
rect 9420 -12110 9560 -12100
rect 9420 -12120 9430 -12110
rect 7950 -12220 9430 -12120
rect 7950 -12230 7960 -12220
rect 7820 -12240 7960 -12230
rect 8060 -12240 9090 -12220
rect 9420 -12230 9430 -12220
rect 9550 -12120 9560 -12110
rect 9660 -12120 10060 -12030
rect 10290 -12120 10690 -12030
rect 11400 -12060 11520 -11980
rect 12040 -12060 12160 -11980
rect 30370 -11983 30376 -11980
rect 30410 -11983 30416 -11980
rect 30370 -11995 30416 -11983
rect 30898 -11983 30904 -11980
rect 30938 -11983 30944 -11980
rect 30898 -11995 30944 -11983
rect 31006 -11983 31012 -11980
rect 31046 -11983 31052 -11980
rect 31006 -11995 31052 -11983
rect 30457 -12028 30857 -12022
rect 30457 -12030 30469 -12028
rect 30845 -12030 30857 -12028
rect 12857 -12068 13260 -12030
rect 12860 -12120 13260 -12068
rect 13490 -12068 13893 -12030
rect 14457 -12068 14860 -12030
rect 13490 -12120 13890 -12068
rect 14460 -12120 14860 -12068
rect 15090 -12068 15493 -12030
rect 14900 -12100 15050 -12090
rect 14900 -12120 14910 -12100
rect 9550 -12220 10690 -12120
rect 9550 -12230 9560 -12220
rect 9420 -12240 9560 -12230
rect 9660 -12240 10690 -12220
rect 1660 -12330 2060 -12240
rect 2290 -12330 2690 -12240
rect 3260 -12330 3660 -12240
rect 3890 -12330 4290 -12240
rect 4860 -12330 5260 -12240
rect 5490 -12330 5890 -12240
rect 6460 -12330 6860 -12240
rect 7090 -12330 7490 -12240
rect 8060 -12330 8460 -12240
rect 8690 -12330 9090 -12240
rect 9660 -12330 10060 -12240
rect 10290 -12330 10690 -12240
rect 11260 -12230 14910 -12120
rect 15040 -12120 15050 -12100
rect 15090 -12120 15490 -12068
rect 15040 -12230 15490 -12120
rect 11260 -12240 15490 -12230
rect 11260 -12330 12290 -12240
rect 12860 -12290 13260 -12240
rect 12857 -12330 13260 -12290
rect 13490 -12290 13890 -12240
rect 14460 -12290 14860 -12240
rect 13490 -12330 13893 -12290
rect 14457 -12330 14860 -12290
rect 15090 -12290 15490 -12240
rect 15600 -12120 15740 -12110
rect 15600 -12240 15610 -12120
rect 15730 -12130 15740 -12120
rect 16060 -12130 16450 -12030
rect 16700 -12130 17090 -12030
rect 15730 -12230 17090 -12130
rect 15730 -12240 15740 -12230
rect 15600 -12250 15740 -12240
rect 15090 -12330 15493 -12290
rect 16060 -12330 16450 -12230
rect 16700 -12330 17090 -12230
rect 17200 -12120 17340 -12110
rect 17200 -12240 17210 -12120
rect 17330 -12130 17340 -12120
rect 17660 -12130 18050 -12030
rect 18300 -12130 18690 -12030
rect 17330 -12230 18690 -12130
rect 17330 -12240 17340 -12230
rect 17200 -12250 17340 -12240
rect 17660 -12330 18050 -12230
rect 18300 -12330 18690 -12230
rect 18800 -12120 18940 -12110
rect 18800 -12240 18810 -12120
rect 18930 -12130 18940 -12120
rect 19260 -12130 19650 -12030
rect 19900 -12130 20290 -12030
rect 18930 -12230 20290 -12130
rect 18930 -12240 18940 -12230
rect 18800 -12250 18940 -12240
rect 19260 -12330 19650 -12230
rect 19900 -12330 20290 -12230
rect 20400 -12120 20540 -12110
rect 20400 -12240 20410 -12120
rect 20530 -12130 20540 -12120
rect 20860 -12130 21250 -12030
rect 21500 -12130 21890 -12030
rect 20530 -12230 21890 -12130
rect 20530 -12240 20540 -12230
rect 20400 -12250 20540 -12240
rect 20860 -12330 21250 -12230
rect 21500 -12330 21890 -12230
rect 22000 -12120 22140 -12110
rect 22000 -12240 22010 -12120
rect 22130 -12130 22140 -12120
rect 22460 -12130 22850 -12030
rect 23100 -12130 23490 -12030
rect 22130 -12230 23490 -12130
rect 22130 -12240 22140 -12230
rect 22000 -12250 22140 -12240
rect 22460 -12330 22850 -12230
rect 23100 -12330 23490 -12230
rect 23600 -12120 23740 -12110
rect 23600 -12240 23610 -12120
rect 23730 -12130 23740 -12120
rect 24060 -12130 24450 -12030
rect 24700 -12130 25090 -12030
rect 23730 -12230 25090 -12130
rect 23730 -12240 23740 -12230
rect 23600 -12250 23740 -12240
rect 24060 -12330 24450 -12230
rect 24700 -12330 25090 -12230
rect 25200 -12120 25340 -12110
rect 25200 -12240 25210 -12120
rect 25330 -12130 25340 -12120
rect 25660 -12130 26050 -12030
rect 26300 -12130 26690 -12030
rect 27260 -12068 27657 -12030
rect 27893 -12068 28290 -12030
rect 25330 -12230 26690 -12130
rect 25330 -12240 25340 -12230
rect 25200 -12250 25340 -12240
rect 25660 -12330 26050 -12230
rect 26300 -12330 26690 -12230
rect 26800 -12120 26940 -12110
rect 26800 -12240 26810 -12120
rect 26930 -12130 26940 -12120
rect 27260 -12130 27650 -12068
rect 27900 -12130 28290 -12068
rect 28860 -12068 29257 -12030
rect 29493 -12068 29890 -12030
rect 30457 -12068 30857 -12030
rect 31093 -12028 31493 -12022
rect 31093 -12030 31105 -12028
rect 31481 -12030 31493 -12028
rect 31093 -12068 31493 -12030
rect 32060 -12068 32457 -12030
rect 32693 -12068 33090 -12030
rect 26930 -12230 28290 -12130
rect 26930 -12240 26940 -12230
rect 26800 -12250 26940 -12240
rect 27260 -12290 27650 -12230
rect 27900 -12290 28290 -12230
rect 28400 -12120 28540 -12110
rect 28400 -12240 28410 -12120
rect 28530 -12130 28540 -12120
rect 28860 -12130 29250 -12068
rect 29500 -12130 29890 -12068
rect 28530 -12230 29890 -12130
rect 28530 -12240 28540 -12230
rect 28400 -12250 28540 -12240
rect 27260 -12330 27657 -12290
rect 27893 -12330 28290 -12290
rect 28860 -12290 29250 -12230
rect 29500 -12290 29890 -12230
rect 30000 -12120 30140 -12110
rect 30000 -12240 30010 -12120
rect 30130 -12130 30140 -12120
rect 30460 -12130 30850 -12068
rect 31100 -12130 31490 -12068
rect 30130 -12230 31490 -12130
rect 30130 -12240 30140 -12230
rect 30000 -12250 30140 -12240
rect 28860 -12330 29257 -12290
rect 29493 -12330 29890 -12290
rect 30460 -12290 30850 -12230
rect 31100 -12290 31490 -12230
rect 31600 -12120 31740 -12110
rect 31600 -12240 31610 -12120
rect 31730 -12130 31740 -12120
rect 32060 -12130 32450 -12068
rect 32700 -12130 33090 -12068
rect 33660 -12068 34057 -12030
rect 34293 -12068 34690 -12030
rect 33660 -12130 34050 -12068
rect 34300 -12130 34690 -12068
rect 35260 -12068 35657 -12030
rect 35893 -12068 36290 -12030
rect 35260 -12130 35650 -12068
rect 35900 -12130 36290 -12068
rect 31730 -12230 36290 -12130
rect 31730 -12240 31740 -12230
rect 31600 -12250 31740 -12240
rect 30460 -12330 30857 -12290
rect 31093 -12330 31490 -12290
rect 32060 -12290 32450 -12230
rect 32700 -12290 33090 -12230
rect 33660 -12290 34050 -12230
rect 34300 -12290 34690 -12230
rect 35260 -12290 35650 -12230
rect 35900 -12290 36290 -12230
rect 32060 -12330 32457 -12290
rect 32340 -12336 32457 -12330
rect 32693 -12336 33093 -12290
rect 33657 -12336 34057 -12290
rect 34293 -12336 34693 -12290
rect 35257 -12336 35657 -12290
rect 35893 -12330 36290 -12290
rect 35893 -12336 36030 -12330
rect 32498 -12390 32544 -12384
rect 32606 -12390 32652 -12384
rect 16510 -12400 16640 -12390
rect 2120 -12410 2240 -12400
rect 2120 -13070 2130 -12410
rect 2230 -13070 2240 -12410
rect 2120 -13080 2240 -13070
rect 3720 -12410 3840 -12400
rect 3720 -13070 3730 -12410
rect 3830 -13070 3840 -12410
rect 3720 -13080 3840 -13070
rect 5320 -12410 5440 -12400
rect 5320 -13070 5330 -12410
rect 5430 -13070 5440 -12410
rect 5320 -13080 5440 -13070
rect 6920 -12410 7040 -12400
rect 6920 -13070 6930 -12410
rect 7030 -13070 7040 -12410
rect 6920 -13080 7040 -13070
rect 8520 -12410 8640 -12400
rect 8520 -13070 8530 -12410
rect 8630 -13070 8640 -12410
rect 8520 -13080 8640 -13070
rect 10120 -12410 10240 -12400
rect 10120 -13070 10130 -12410
rect 10230 -13070 10240 -12410
rect 10120 -13080 10240 -13070
rect 11710 -12410 11840 -12400
rect 11710 -13070 11720 -12410
rect 11830 -13070 11840 -12410
rect 11710 -13080 11840 -13070
rect 13310 -12410 13440 -12400
rect 13310 -13070 13320 -12410
rect 13430 -13070 13440 -12410
rect 13310 -13080 13440 -13070
rect 14910 -12410 15040 -12400
rect 14910 -13070 14920 -12410
rect 15030 -13070 15040 -12410
rect 14910 -13080 15040 -13070
rect 16510 -13080 16520 -12400
rect 16630 -13080 16640 -12400
rect 16510 -13090 16640 -13080
rect 18110 -12400 18240 -12390
rect 18110 -13080 18120 -12400
rect 18230 -13080 18240 -12400
rect 18110 -13090 18240 -13080
rect 19710 -12400 19840 -12390
rect 19710 -13080 19720 -12400
rect 19830 -13080 19840 -12400
rect 19710 -13090 19840 -13080
rect 21310 -12400 21440 -12390
rect 21310 -13080 21320 -12400
rect 21430 -13080 21440 -12400
rect 21310 -13090 21440 -13080
rect 22910 -12400 23040 -12390
rect 22910 -13080 22920 -12400
rect 23030 -13080 23040 -12400
rect 22910 -13090 23040 -13080
rect 24510 -12400 24640 -12390
rect 24510 -13080 24520 -12400
rect 24630 -13080 24640 -12400
rect 24510 -13090 24640 -13080
rect 26110 -12400 26240 -12390
rect 26110 -13080 26120 -12400
rect 26230 -13080 26240 -12400
rect 26110 -13090 26240 -13080
rect 27710 -12400 27840 -12390
rect 27710 -13080 27720 -12400
rect 27830 -13080 27840 -12400
rect 27710 -13090 27840 -13080
rect 29310 -12400 29440 -12390
rect 29310 -13080 29320 -12400
rect 29430 -13080 29440 -12400
rect 29310 -13090 29440 -13080
rect 30910 -12400 31040 -12390
rect 30910 -13080 30920 -12400
rect 31030 -13080 31040 -12400
rect 32498 -12396 32652 -12390
rect 32498 -12910 32504 -12396
rect 32510 -12400 32640 -12396
rect 32510 -12910 32520 -12400
rect 32630 -12910 32640 -12400
rect 32646 -12910 32652 -12396
rect 33134 -12396 33180 -12384
rect 33134 -12910 33140 -12396
rect 33174 -12910 33180 -12396
rect 33570 -12396 33616 -12384
rect 33570 -12910 33576 -12396
rect 33610 -12910 33616 -12396
rect 34098 -12390 34144 -12384
rect 34206 -12390 34252 -12384
rect 34098 -12396 34252 -12390
rect 34098 -12910 34104 -12396
rect 34110 -12400 34240 -12396
rect 34110 -12910 34120 -12400
rect 34230 -12910 34240 -12400
rect 34246 -12910 34252 -12396
rect 34734 -12396 34780 -12384
rect 34734 -12910 34740 -12396
rect 34774 -12910 34780 -12396
rect 35170 -12396 35216 -12384
rect 35170 -12910 35176 -12396
rect 35210 -12910 35216 -12396
rect 35698 -12390 35744 -12384
rect 35806 -12390 35852 -12384
rect 35698 -12396 35852 -12390
rect 35698 -12910 35704 -12396
rect 35710 -12400 35840 -12396
rect 35710 -12910 35720 -12400
rect 35830 -12910 35840 -12400
rect 35846 -12910 35852 -12396
rect 30910 -13090 31040 -13080
rect 35000 -13110 35140 -13100
rect 35000 -13150 35010 -13110
rect 670 -13300 11080 -13180
rect 11260 -13210 11270 -13150
rect 11650 -13210 12300 -13150
rect 12720 -13300 31860 -13180
rect 32060 -13230 35010 -13150
rect 35130 -13150 35140 -13110
rect 35130 -13230 36290 -13150
rect 32060 -13240 36290 -13230
rect 39100 -13300 39229 -11600
rect 670 -13400 39229 -13300
rect 670 -13420 37940 -13400
rect 670 -14980 720 -13420
rect 1200 -13470 1340 -13460
rect 1200 -13590 1210 -13470
rect 1330 -13480 1340 -13470
rect 2800 -13470 2940 -13460
rect 2800 -13480 2810 -13470
rect 1330 -13580 2810 -13480
rect 1330 -13590 1340 -13580
rect 1200 -13600 1340 -13590
rect 2800 -13590 2810 -13580
rect 2930 -13480 2940 -13470
rect 4400 -13470 4540 -13460
rect 4400 -13480 4410 -13470
rect 2930 -13580 4410 -13480
rect 2930 -13590 2940 -13580
rect 2800 -13600 2940 -13590
rect 4400 -13590 4410 -13580
rect 4530 -13480 4540 -13470
rect 6000 -13470 6140 -13460
rect 6000 -13480 6010 -13470
rect 4530 -13580 6010 -13480
rect 4530 -13590 4540 -13580
rect 4400 -13600 4540 -13590
rect 6000 -13590 6010 -13580
rect 6130 -13480 6140 -13470
rect 7600 -13470 7740 -13460
rect 7600 -13480 7610 -13470
rect 6130 -13580 7610 -13480
rect 6130 -13590 6140 -13580
rect 6000 -13600 6140 -13590
rect 7600 -13590 7610 -13580
rect 7730 -13480 7740 -13470
rect 9200 -13470 9340 -13460
rect 15820 -13470 15960 -13460
rect 9200 -13480 9210 -13470
rect 7730 -13580 9210 -13480
rect 7730 -13590 7740 -13580
rect 7600 -13600 7740 -13590
rect 9200 -13590 9210 -13580
rect 9330 -13480 9340 -13470
rect 14000 -13480 14140 -13470
rect 9330 -13580 10700 -13480
rect 14000 -13520 14010 -13480
rect 9330 -13590 9340 -13580
rect 9200 -13600 9340 -13590
rect 10750 -13660 10940 -13650
rect 11400 -13660 11520 -13580
rect 12040 -13660 12160 -13580
rect 12860 -13600 14010 -13520
rect 14130 -13520 14140 -13480
rect 14130 -13600 15490 -13520
rect 15820 -13590 15830 -13470
rect 15950 -13500 15960 -13470
rect 17420 -13470 17560 -13460
rect 15950 -13590 17090 -13500
rect 15820 -13600 17090 -13590
rect 17420 -13590 17430 -13470
rect 17550 -13500 17560 -13470
rect 19020 -13470 19160 -13460
rect 17550 -13590 18690 -13500
rect 17420 -13600 18690 -13590
rect 19020 -13590 19030 -13470
rect 19150 -13500 19160 -13470
rect 20620 -13470 20760 -13460
rect 19150 -13590 20290 -13500
rect 19020 -13600 20290 -13590
rect 20620 -13590 20630 -13470
rect 20750 -13500 20760 -13470
rect 22220 -13470 22360 -13460
rect 20750 -13590 21890 -13500
rect 20620 -13600 21890 -13590
rect 22220 -13590 22230 -13470
rect 22350 -13500 22360 -13470
rect 23820 -13470 23960 -13460
rect 22350 -13590 23490 -13500
rect 22220 -13600 23490 -13590
rect 23820 -13590 23830 -13470
rect 23950 -13500 23960 -13470
rect 25420 -13470 25560 -13460
rect 23950 -13590 25090 -13500
rect 23820 -13600 25090 -13590
rect 25420 -13590 25430 -13470
rect 25550 -13500 25560 -13470
rect 27020 -13470 27160 -13460
rect 25550 -13590 26680 -13500
rect 25420 -13600 26680 -13590
rect 27020 -13590 27030 -13470
rect 27150 -13500 27160 -13470
rect 28620 -13470 28760 -13460
rect 27150 -13590 28290 -13500
rect 27020 -13600 28290 -13590
rect 28620 -13590 28630 -13470
rect 28750 -13500 28760 -13470
rect 30220 -13470 30360 -13460
rect 28750 -13590 29890 -13500
rect 28620 -13600 29890 -13590
rect 30220 -13590 30230 -13470
rect 30350 -13500 30360 -13470
rect 31820 -13470 31960 -13460
rect 30350 -13564 31490 -13500
rect 30350 -13590 31493 -13564
rect 30220 -13600 31493 -13590
rect 31820 -13590 31830 -13470
rect 31950 -13500 31960 -13470
rect 34800 -13470 34940 -13460
rect 34800 -13500 34810 -13470
rect 31950 -13590 34810 -13500
rect 34930 -13500 34940 -13470
rect 34930 -13590 36280 -13500
rect 31820 -13600 36280 -13590
rect 14000 -13610 14140 -13600
rect 30457 -13604 30469 -13600
rect 30845 -13604 30857 -13600
rect 30457 -13610 30857 -13604
rect 31093 -13604 31105 -13600
rect 31481 -13604 31493 -13600
rect 31093 -13610 31493 -13604
rect 32057 -13604 32069 -13600
rect 32057 -13610 32140 -13604
rect 30370 -13649 30416 -13637
rect 30370 -13660 30376 -13649
rect 30410 -13660 30416 -13649
rect 30898 -13649 30944 -13637
rect 30898 -13660 30904 -13649
rect 30938 -13660 30944 -13649
rect 31006 -13649 31052 -13637
rect 31006 -13660 31012 -13649
rect 31046 -13660 31052 -13649
rect 1560 -13780 10810 -13660
rect 10930 -13780 36380 -13660
rect 10750 -13790 10940 -13780
rect 1420 -13910 1560 -13900
rect 1420 -14030 1430 -13910
rect 1550 -13920 1560 -13910
rect 1660 -13920 2060 -13830
rect 2290 -13920 2690 -13830
rect 3020 -13910 3160 -13900
rect 3020 -13920 3030 -13910
rect 1550 -14020 3030 -13920
rect 1550 -14030 1560 -14020
rect 1420 -14040 1560 -14030
rect 1660 -14040 2690 -14020
rect 3020 -14030 3030 -14020
rect 3150 -13920 3160 -13910
rect 3260 -13920 3660 -13830
rect 3890 -13920 4290 -13830
rect 4620 -13910 4760 -13900
rect 4620 -13920 4630 -13910
rect 3150 -14020 4630 -13920
rect 3150 -14030 3160 -14020
rect 3020 -14040 3160 -14030
rect 3260 -14040 4290 -14020
rect 4620 -14030 4630 -14020
rect 4750 -13920 4760 -13910
rect 4860 -13920 5260 -13830
rect 5490 -13920 5890 -13830
rect 6220 -13910 6360 -13900
rect 6220 -13920 6230 -13910
rect 4750 -14020 6230 -13920
rect 4750 -14030 4760 -14020
rect 4620 -14040 4760 -14030
rect 4860 -14040 5890 -14020
rect 6220 -14030 6230 -14020
rect 6350 -13920 6360 -13910
rect 6460 -13920 6860 -13830
rect 7090 -13920 7490 -13830
rect 7820 -13910 7960 -13900
rect 7820 -13920 7830 -13910
rect 6350 -14020 7830 -13920
rect 6350 -14030 6360 -14020
rect 6220 -14040 6360 -14030
rect 6460 -14040 7490 -14020
rect 7820 -14030 7830 -14020
rect 7950 -13920 7960 -13910
rect 8060 -13920 8460 -13830
rect 8690 -13920 9090 -13830
rect 9420 -13910 9560 -13900
rect 9420 -13920 9430 -13910
rect 7950 -14020 9430 -13920
rect 7950 -14030 7960 -14020
rect 7820 -14040 7960 -14030
rect 8060 -14040 9090 -14020
rect 9420 -14030 9430 -14020
rect 9550 -13920 9560 -13910
rect 9660 -13920 10060 -13830
rect 10290 -13920 10690 -13830
rect 11400 -13860 11520 -13780
rect 12040 -13860 12160 -13780
rect 30370 -13783 30376 -13780
rect 30410 -13783 30416 -13780
rect 30370 -13795 30416 -13783
rect 30898 -13783 30904 -13780
rect 30938 -13783 30944 -13780
rect 30898 -13795 30944 -13783
rect 31006 -13783 31012 -13780
rect 31046 -13783 31052 -13780
rect 31006 -13795 31052 -13783
rect 30457 -13828 30857 -13822
rect 30457 -13830 30469 -13828
rect 30845 -13830 30857 -13828
rect 9550 -14020 10690 -13920
rect 9550 -14030 9560 -14020
rect 9420 -14040 9560 -14030
rect 9660 -14040 10690 -14020
rect 1660 -14130 2060 -14040
rect 2290 -14130 2690 -14040
rect 3260 -14130 3660 -14040
rect 3890 -14130 4290 -14040
rect 4860 -14130 5260 -14040
rect 5490 -14130 5890 -14040
rect 6460 -14130 6860 -14040
rect 7090 -14130 7490 -14040
rect 8060 -14130 8460 -14040
rect 8690 -14130 9090 -14040
rect 9660 -14130 10060 -14040
rect 10290 -14130 10690 -14040
rect 12860 -13920 13260 -13830
rect 13490 -13920 13890 -13830
rect 14460 -13920 14860 -13830
rect 15090 -13920 15490 -13830
rect 12860 -14040 15490 -13920
rect 11260 -14060 12290 -14050
rect 11260 -14120 11270 -14060
rect 11650 -14120 12290 -14060
rect 11260 -14130 11660 -14120
rect 12860 -14130 13260 -14040
rect 13490 -14130 13890 -14040
rect 14460 -14130 14860 -14040
rect 15090 -14130 15490 -14040
rect 15600 -13920 15740 -13910
rect 15600 -14040 15610 -13920
rect 15730 -13930 15740 -13920
rect 16060 -13930 16450 -13830
rect 16700 -13930 17090 -13830
rect 15730 -14030 17090 -13930
rect 15730 -14040 15740 -14030
rect 15600 -14050 15740 -14040
rect 16060 -14130 16450 -14030
rect 16700 -14130 17090 -14030
rect 17200 -13920 17340 -13910
rect 17200 -14040 17210 -13920
rect 17330 -13930 17340 -13920
rect 17660 -13930 18050 -13830
rect 18300 -13930 18690 -13830
rect 17330 -14030 18690 -13930
rect 17330 -14040 17340 -14030
rect 17200 -14050 17340 -14040
rect 17660 -14130 18050 -14030
rect 18300 -14130 18690 -14030
rect 18800 -13920 18940 -13910
rect 18800 -14040 18810 -13920
rect 18930 -13930 18940 -13920
rect 19260 -13930 19650 -13830
rect 19900 -13930 20290 -13830
rect 18930 -14030 20290 -13930
rect 18930 -14040 18940 -14030
rect 18800 -14050 18940 -14040
rect 19260 -14130 19650 -14030
rect 19900 -14130 20290 -14030
rect 20400 -13920 20540 -13910
rect 20400 -14040 20410 -13920
rect 20530 -13930 20540 -13920
rect 20860 -13930 21250 -13830
rect 21500 -13930 21890 -13830
rect 20530 -14030 21890 -13930
rect 20530 -14040 20540 -14030
rect 20400 -14050 20540 -14040
rect 20860 -14130 21250 -14030
rect 21500 -14130 21890 -14030
rect 22000 -13920 22140 -13910
rect 22000 -14040 22010 -13920
rect 22130 -13930 22140 -13920
rect 22460 -13930 22850 -13830
rect 23100 -13930 23490 -13830
rect 22130 -14030 23490 -13930
rect 22130 -14040 22140 -14030
rect 22000 -14050 22140 -14040
rect 22460 -14130 22850 -14030
rect 23100 -14130 23490 -14030
rect 23600 -13920 23740 -13910
rect 23600 -14040 23610 -13920
rect 23730 -13930 23740 -13920
rect 24060 -13930 24450 -13830
rect 24700 -13930 25090 -13830
rect 23730 -14030 25090 -13930
rect 23730 -14040 23740 -14030
rect 23600 -14050 23740 -14040
rect 24060 -14130 24450 -14030
rect 24700 -14130 25090 -14030
rect 25200 -13920 25340 -13910
rect 25200 -14040 25210 -13920
rect 25330 -13930 25340 -13920
rect 25660 -13930 26050 -13830
rect 26300 -13930 26690 -13830
rect 27260 -13868 27657 -13830
rect 27893 -13868 28290 -13830
rect 25330 -14030 26690 -13930
rect 25330 -14040 25340 -14030
rect 25200 -14050 25340 -14040
rect 25660 -14130 26050 -14030
rect 26300 -14130 26690 -14030
rect 26800 -13920 26940 -13910
rect 26800 -14040 26810 -13920
rect 26930 -13930 26940 -13920
rect 27260 -13930 27650 -13868
rect 27900 -13930 28290 -13868
rect 28860 -13868 29257 -13830
rect 29493 -13868 29890 -13830
rect 30457 -13868 30857 -13830
rect 31093 -13828 31493 -13822
rect 31093 -13830 31105 -13828
rect 31481 -13830 31493 -13828
rect 31093 -13868 31493 -13830
rect 32060 -13868 32457 -13830
rect 32693 -13868 33090 -13830
rect 26930 -14030 28290 -13930
rect 26930 -14040 26940 -14030
rect 26800 -14050 26940 -14040
rect 27260 -14090 27650 -14030
rect 27900 -14090 28290 -14030
rect 28400 -13920 28540 -13910
rect 28400 -14040 28410 -13920
rect 28530 -13930 28540 -13920
rect 28860 -13930 29250 -13868
rect 29500 -13930 29890 -13868
rect 28530 -14030 29890 -13930
rect 28530 -14040 28540 -14030
rect 28400 -14050 28540 -14040
rect 27260 -14130 27657 -14090
rect 27893 -14130 28290 -14090
rect 28860 -14090 29250 -14030
rect 29500 -14090 29890 -14030
rect 30000 -13920 30140 -13910
rect 30000 -14040 30010 -13920
rect 30130 -13930 30140 -13920
rect 30460 -13930 30850 -13868
rect 31100 -13930 31490 -13868
rect 30130 -14030 31490 -13930
rect 30130 -14040 30140 -14030
rect 30000 -14050 30140 -14040
rect 28860 -14130 29257 -14090
rect 29493 -14130 29890 -14090
rect 30460 -14090 30850 -14030
rect 31100 -14090 31490 -14030
rect 31600 -13920 31740 -13910
rect 31600 -14040 31610 -13920
rect 31730 -13930 31740 -13920
rect 32060 -13930 32450 -13868
rect 32700 -13930 33090 -13868
rect 33660 -13868 34057 -13830
rect 34293 -13868 34690 -13830
rect 33660 -13930 34050 -13868
rect 34300 -13930 34690 -13868
rect 35260 -13868 35657 -13830
rect 35893 -13868 36290 -13830
rect 35260 -13930 35650 -13868
rect 35900 -13930 36290 -13868
rect 31730 -14030 36290 -13930
rect 31730 -14040 31740 -14030
rect 31600 -14050 31740 -14040
rect 30460 -14130 30857 -14090
rect 31093 -14130 31490 -14090
rect 32060 -14090 32450 -14030
rect 32700 -14090 33090 -14030
rect 33660 -14090 34050 -14030
rect 34300 -14090 34690 -14030
rect 35260 -14090 35650 -14030
rect 35900 -14090 36290 -14030
rect 32060 -14130 32457 -14090
rect 32340 -14136 32457 -14130
rect 32693 -14136 33093 -14090
rect 33657 -14136 34057 -14090
rect 34293 -14136 34693 -14090
rect 35257 -14136 35657 -14090
rect 35893 -14130 36290 -14090
rect 35893 -14136 36030 -14130
rect 32498 -14190 32544 -14184
rect 32606 -14190 32652 -14184
rect 16510 -14200 16640 -14190
rect 2120 -14210 2240 -14200
rect 2120 -14870 2130 -14210
rect 2230 -14870 2240 -14210
rect 2120 -14880 2240 -14870
rect 3720 -14210 3840 -14200
rect 3720 -14870 3730 -14210
rect 3830 -14870 3840 -14210
rect 3720 -14880 3840 -14870
rect 5320 -14210 5440 -14200
rect 5320 -14870 5330 -14210
rect 5430 -14870 5440 -14210
rect 5320 -14880 5440 -14870
rect 6920 -14210 7040 -14200
rect 6920 -14870 6930 -14210
rect 7030 -14870 7040 -14210
rect 6920 -14880 7040 -14870
rect 8520 -14210 8640 -14200
rect 8520 -14870 8530 -14210
rect 8630 -14870 8640 -14210
rect 8520 -14880 8640 -14870
rect 10120 -14210 10240 -14200
rect 10120 -14870 10130 -14210
rect 10230 -14870 10240 -14210
rect 10120 -14880 10240 -14870
rect 11710 -14210 11840 -14200
rect 11710 -14870 11720 -14210
rect 11830 -14870 11840 -14210
rect 11710 -14880 11840 -14870
rect 13310 -14210 13440 -14200
rect 13310 -14870 13320 -14210
rect 13430 -14870 13440 -14210
rect 13310 -14880 13440 -14870
rect 14910 -14210 15040 -14200
rect 14910 -14870 14920 -14210
rect 15030 -14870 15040 -14210
rect 14910 -14880 15040 -14870
rect 16510 -14880 16520 -14200
rect 16630 -14880 16640 -14200
rect 16510 -14890 16640 -14880
rect 18110 -14200 18240 -14190
rect 18110 -14880 18120 -14200
rect 18230 -14880 18240 -14200
rect 18110 -14890 18240 -14880
rect 19710 -14200 19840 -14190
rect 19710 -14880 19720 -14200
rect 19830 -14880 19840 -14200
rect 19710 -14890 19840 -14880
rect 21310 -14200 21440 -14190
rect 21310 -14880 21320 -14200
rect 21430 -14880 21440 -14200
rect 21310 -14890 21440 -14880
rect 22910 -14200 23040 -14190
rect 22910 -14880 22920 -14200
rect 23030 -14880 23040 -14200
rect 22910 -14890 23040 -14880
rect 24510 -14200 24640 -14190
rect 24510 -14880 24520 -14200
rect 24630 -14880 24640 -14200
rect 24510 -14890 24640 -14880
rect 26110 -14200 26240 -14190
rect 26110 -14880 26120 -14200
rect 26230 -14880 26240 -14200
rect 26110 -14890 26240 -14880
rect 27710 -14200 27840 -14190
rect 27710 -14880 27720 -14200
rect 27830 -14880 27840 -14200
rect 27710 -14890 27840 -14880
rect 29310 -14200 29440 -14190
rect 29310 -14880 29320 -14200
rect 29430 -14880 29440 -14200
rect 29310 -14890 29440 -14880
rect 30910 -14200 31040 -14190
rect 30910 -14880 30920 -14200
rect 31030 -14880 31040 -14200
rect 32498 -14196 32652 -14190
rect 32498 -14710 32504 -14196
rect 32510 -14200 32640 -14196
rect 32510 -14710 32520 -14200
rect 32630 -14710 32640 -14200
rect 32646 -14710 32652 -14196
rect 33134 -14196 33180 -14184
rect 33134 -14710 33140 -14196
rect 33174 -14710 33180 -14196
rect 33570 -14196 33616 -14184
rect 33570 -14710 33576 -14196
rect 33610 -14710 33616 -14196
rect 34098 -14190 34144 -14184
rect 34206 -14190 34252 -14184
rect 34098 -14196 34252 -14190
rect 34098 -14710 34104 -14196
rect 34110 -14200 34240 -14196
rect 34110 -14710 34120 -14200
rect 34230 -14710 34240 -14200
rect 34246 -14710 34252 -14196
rect 34734 -14196 34780 -14184
rect 34734 -14710 34740 -14196
rect 34774 -14710 34780 -14196
rect 35170 -14196 35216 -14184
rect 35170 -14710 35176 -14196
rect 35210 -14710 35216 -14196
rect 35698 -14190 35744 -14184
rect 35806 -14190 35852 -14184
rect 35698 -14196 35852 -14190
rect 35698 -14710 35704 -14196
rect 35710 -14200 35840 -14196
rect 35710 -14710 35720 -14200
rect 35830 -14710 35840 -14200
rect 35846 -14710 35852 -14196
rect 30910 -14890 31040 -14880
rect 35000 -14910 35140 -14900
rect 35000 -14950 35010 -14910
rect 670 -15100 31800 -14980
rect 32060 -15030 35010 -14950
rect 35130 -14950 35140 -14910
rect 35130 -15030 36290 -14950
rect 32060 -15040 36290 -15030
rect 39100 -15100 39229 -13400
rect 670 -15200 39229 -15100
rect 670 -15220 37940 -15200
rect 670 -16760 720 -15220
rect 1200 -15270 1340 -15260
rect 1200 -15390 1210 -15270
rect 1330 -15280 1340 -15270
rect 2800 -15270 2940 -15260
rect 2800 -15280 2810 -15270
rect 1330 -15380 2810 -15280
rect 1330 -15390 1340 -15380
rect 1200 -15400 1340 -15390
rect 2800 -15390 2810 -15380
rect 2930 -15280 2940 -15270
rect 4400 -15270 4540 -15260
rect 4400 -15280 4410 -15270
rect 2930 -15380 4410 -15280
rect 2930 -15390 2940 -15380
rect 2800 -15400 2940 -15390
rect 4400 -15390 4410 -15380
rect 4530 -15280 4540 -15270
rect 6000 -15270 6140 -15260
rect 6000 -15280 6010 -15270
rect 4530 -15380 6010 -15280
rect 4530 -15390 4540 -15380
rect 4400 -15400 4540 -15390
rect 6000 -15390 6010 -15380
rect 6130 -15280 6140 -15270
rect 7600 -15270 7740 -15260
rect 7600 -15280 7610 -15270
rect 6130 -15380 7610 -15280
rect 6130 -15390 6140 -15380
rect 6000 -15400 6140 -15390
rect 7600 -15390 7610 -15380
rect 7730 -15280 7740 -15270
rect 9200 -15270 9340 -15260
rect 9200 -15280 9210 -15270
rect 7730 -15380 9210 -15280
rect 7730 -15390 7740 -15380
rect 7600 -15400 7740 -15390
rect 9200 -15390 9210 -15380
rect 9330 -15280 9340 -15270
rect 15820 -15270 15960 -15260
rect 9330 -15380 10700 -15280
rect 13320 -15290 13440 -15280
rect 13320 -15320 13330 -15290
rect 9330 -15390 9340 -15380
rect 9200 -15400 9340 -15390
rect 10750 -15460 10940 -15450
rect 11400 -15460 11520 -15380
rect 12040 -15460 12160 -15380
rect 12860 -15390 13330 -15320
rect 13430 -15320 13440 -15290
rect 14920 -15290 15040 -15280
rect 14010 -15310 14130 -15300
rect 14010 -15320 14020 -15310
rect 13430 -15390 14020 -15320
rect 12860 -15400 14020 -15390
rect 14010 -15410 14020 -15400
rect 14120 -15320 14130 -15310
rect 14920 -15320 14930 -15290
rect 14120 -15390 14930 -15320
rect 15030 -15320 15040 -15290
rect 15030 -15390 15490 -15320
rect 14120 -15400 15490 -15390
rect 15820 -15390 15830 -15270
rect 15950 -15300 15960 -15270
rect 17420 -15270 17560 -15260
rect 15950 -15390 17090 -15300
rect 15820 -15400 17090 -15390
rect 17420 -15390 17430 -15270
rect 17550 -15300 17560 -15270
rect 19020 -15270 19160 -15260
rect 17550 -15390 18690 -15300
rect 17420 -15400 18690 -15390
rect 19020 -15390 19030 -15270
rect 19150 -15300 19160 -15270
rect 20620 -15270 20760 -15260
rect 19150 -15390 20290 -15300
rect 19020 -15400 20290 -15390
rect 20620 -15390 20630 -15270
rect 20750 -15300 20760 -15270
rect 22220 -15270 22360 -15260
rect 20750 -15390 21890 -15300
rect 20620 -15400 21890 -15390
rect 22220 -15390 22230 -15270
rect 22350 -15300 22360 -15270
rect 23820 -15270 23960 -15260
rect 22350 -15390 23490 -15300
rect 22220 -15400 23490 -15390
rect 23820 -15390 23830 -15270
rect 23950 -15300 23960 -15270
rect 27020 -15270 27160 -15260
rect 27020 -15300 27030 -15270
rect 23950 -15390 25090 -15300
rect 23820 -15400 25090 -15390
rect 25660 -15390 27030 -15300
rect 27150 -15300 27160 -15270
rect 28620 -15270 28760 -15260
rect 27150 -15390 28290 -15300
rect 25660 -15400 28290 -15390
rect 28620 -15390 28630 -15270
rect 28750 -15300 28760 -15270
rect 31840 -15280 31980 -15270
rect 28750 -15390 31490 -15300
rect 28620 -15400 31490 -15390
rect 31840 -15400 31850 -15280
rect 31970 -15300 31980 -15280
rect 31970 -15400 36290 -15300
rect 14120 -15410 14130 -15400
rect 31840 -15410 31980 -15400
rect 14010 -15420 14130 -15410
rect 1560 -15580 10810 -15460
rect 10930 -15580 36380 -15460
rect 10750 -15590 10940 -15580
rect 1420 -15710 1560 -15700
rect 1420 -15830 1430 -15710
rect 1550 -15720 1560 -15710
rect 1660 -15720 2060 -15630
rect 2290 -15720 2690 -15630
rect 3020 -15710 3160 -15700
rect 3020 -15720 3030 -15710
rect 1550 -15820 3030 -15720
rect 1550 -15830 1560 -15820
rect 1420 -15840 1560 -15830
rect 1660 -15840 2690 -15820
rect 3020 -15830 3030 -15820
rect 3150 -15720 3160 -15710
rect 3260 -15720 3660 -15630
rect 3890 -15720 4290 -15630
rect 4620 -15710 4760 -15700
rect 4620 -15720 4630 -15710
rect 3150 -15820 4630 -15720
rect 3150 -15830 3160 -15820
rect 3020 -15840 3160 -15830
rect 3260 -15840 4290 -15820
rect 4620 -15830 4630 -15820
rect 4750 -15720 4760 -15710
rect 4860 -15720 5260 -15630
rect 5490 -15720 5890 -15630
rect 6220 -15710 6360 -15700
rect 6220 -15720 6230 -15710
rect 4750 -15820 6230 -15720
rect 4750 -15830 4760 -15820
rect 4620 -15840 4760 -15830
rect 4860 -15840 5890 -15820
rect 6220 -15830 6230 -15820
rect 6350 -15720 6360 -15710
rect 6460 -15720 6860 -15630
rect 7090 -15720 7490 -15630
rect 7820 -15710 7960 -15700
rect 7820 -15720 7830 -15710
rect 6350 -15820 7830 -15720
rect 6350 -15830 6360 -15820
rect 6220 -15840 6360 -15830
rect 6460 -15840 7490 -15820
rect 7820 -15830 7830 -15820
rect 7950 -15720 7960 -15710
rect 8060 -15720 8460 -15630
rect 8690 -15720 9090 -15630
rect 9420 -15710 9560 -15700
rect 9420 -15720 9430 -15710
rect 7950 -15820 9430 -15720
rect 7950 -15830 7960 -15820
rect 7820 -15840 7960 -15830
rect 8060 -15840 9090 -15820
rect 9420 -15830 9430 -15820
rect 9550 -15720 9560 -15710
rect 9660 -15720 10060 -15630
rect 10290 -15720 10690 -15630
rect 11400 -15660 11520 -15580
rect 12040 -15660 12160 -15580
rect 9550 -15820 10690 -15720
rect 9550 -15830 9560 -15820
rect 9420 -15840 9560 -15830
rect 9660 -15840 10690 -15820
rect 1660 -15930 2060 -15840
rect 2290 -15930 2690 -15840
rect 3260 -15930 3660 -15840
rect 3890 -15930 4290 -15840
rect 4860 -15930 5260 -15840
rect 5490 -15930 5890 -15840
rect 6460 -15930 6860 -15840
rect 7090 -15930 7490 -15840
rect 8060 -15930 8460 -15840
rect 8690 -15930 9090 -15840
rect 9660 -15930 10060 -15840
rect 10290 -15930 10690 -15840
rect 12860 -15710 13260 -15630
rect 13490 -15710 13890 -15630
rect 14460 -15710 14860 -15630
rect 12860 -15720 15050 -15710
rect 15090 -15720 15490 -15630
rect 12860 -15830 15490 -15720
rect 12860 -15840 13890 -15830
rect 2120 -16010 2240 -16000
rect 2120 -16430 2130 -16010
rect 2120 -16670 2130 -16630
rect 2230 -16430 2240 -16010
rect 3720 -16010 3840 -16000
rect 3720 -16430 3730 -16010
rect 2230 -16670 2240 -16630
rect 2120 -16680 2240 -16670
rect 3720 -16670 3730 -16630
rect 3830 -16430 3840 -16010
rect 5320 -16010 5440 -16000
rect 5320 -16430 5330 -16010
rect 3830 -16670 3840 -16630
rect 3720 -16680 3840 -16670
rect 5320 -16670 5330 -16630
rect 5430 -16430 5440 -16010
rect 6920 -16010 7040 -16000
rect 6920 -16430 6930 -16010
rect 5430 -16670 5440 -16630
rect 5320 -16680 5440 -16670
rect 6920 -16670 6930 -16630
rect 7030 -16430 7040 -16010
rect 8520 -16010 8640 -16000
rect 7030 -16670 7040 -16630
rect 6920 -16680 7040 -16670
rect 8520 -16670 8530 -16010
rect 8630 -16670 8640 -16010
rect 8520 -16680 8640 -16670
rect 10120 -16010 10240 -16000
rect 10120 -16670 10130 -16010
rect 10230 -16670 10240 -16010
rect 11420 -16290 11500 -15900
rect 12040 -16290 12120 -15900
rect 12860 -15930 13260 -15840
rect 13490 -15930 13890 -15840
rect 14460 -15840 15490 -15830
rect 14460 -15930 14860 -15840
rect 15090 -15930 15490 -15840
rect 15600 -15720 15740 -15710
rect 15600 -15840 15610 -15720
rect 15730 -15730 15740 -15720
rect 16060 -15730 16450 -15630
rect 16700 -15730 17090 -15630
rect 15730 -15830 17090 -15730
rect 15730 -15840 15740 -15830
rect 15600 -15850 15740 -15840
rect 16060 -15930 16450 -15830
rect 16700 -15930 17090 -15830
rect 17200 -15720 17340 -15710
rect 17200 -15840 17210 -15720
rect 17330 -15730 17340 -15720
rect 17660 -15730 18050 -15630
rect 18300 -15730 18690 -15630
rect 17330 -15830 18690 -15730
rect 17330 -15840 17340 -15830
rect 17200 -15850 17340 -15840
rect 17660 -15930 18050 -15830
rect 18300 -15930 18690 -15830
rect 18800 -15720 18940 -15710
rect 18800 -15840 18810 -15720
rect 18930 -15730 18940 -15720
rect 19260 -15730 19650 -15630
rect 19900 -15730 20290 -15630
rect 18930 -15830 20290 -15730
rect 18930 -15840 18940 -15830
rect 18800 -15850 18940 -15840
rect 19260 -15930 19650 -15830
rect 19900 -15930 20290 -15830
rect 20400 -15720 20540 -15710
rect 20400 -15840 20410 -15720
rect 20530 -15730 20540 -15720
rect 20860 -15730 21250 -15630
rect 21500 -15730 21890 -15630
rect 20530 -15830 21890 -15730
rect 20530 -15840 20540 -15830
rect 20400 -15850 20540 -15840
rect 20860 -15930 21250 -15830
rect 21500 -15930 21890 -15830
rect 22000 -15720 22140 -15710
rect 22000 -15840 22010 -15720
rect 22130 -15730 22140 -15720
rect 22460 -15730 22850 -15630
rect 23100 -15730 23490 -15630
rect 22130 -15830 23490 -15730
rect 22130 -15840 22140 -15830
rect 22000 -15850 22140 -15840
rect 22460 -15930 22850 -15830
rect 23100 -15930 23490 -15830
rect 23600 -15720 23740 -15710
rect 23600 -15840 23610 -15720
rect 23730 -15730 23740 -15720
rect 24060 -15730 24450 -15630
rect 24700 -15730 25090 -15630
rect 23730 -15830 25090 -15730
rect 23730 -15840 23740 -15830
rect 23600 -15850 23740 -15840
rect 24060 -15930 24450 -15830
rect 24700 -15930 25090 -15830
rect 25660 -15730 26050 -15630
rect 26300 -15730 26690 -15630
rect 27260 -15668 27657 -15630
rect 27893 -15668 28290 -15630
rect 26800 -15720 26940 -15710
rect 26800 -15730 26810 -15720
rect 25660 -15830 26810 -15730
rect 25660 -15930 26050 -15830
rect 26300 -15930 26690 -15830
rect 26800 -15840 26810 -15830
rect 26930 -15730 26940 -15720
rect 27260 -15730 27650 -15668
rect 27900 -15730 28290 -15668
rect 28860 -15668 29257 -15630
rect 29493 -15668 29890 -15630
rect 26930 -15830 28290 -15730
rect 26930 -15840 26940 -15830
rect 26800 -15850 26940 -15840
rect 27260 -15890 27650 -15830
rect 27900 -15890 28290 -15830
rect 28400 -15720 28540 -15710
rect 28400 -15840 28410 -15720
rect 28530 -15730 28540 -15720
rect 28860 -15730 29250 -15668
rect 29500 -15730 29890 -15668
rect 30460 -15668 30857 -15630
rect 31093 -15668 31490 -15630
rect 30460 -15730 30850 -15668
rect 31100 -15730 31490 -15668
rect 32060 -15668 32457 -15630
rect 32693 -15668 33090 -15630
rect 28530 -15830 31490 -15730
rect 28530 -15840 28540 -15830
rect 28400 -15850 28540 -15840
rect 27260 -15930 27657 -15890
rect 27893 -15930 28290 -15890
rect 28860 -15890 29250 -15830
rect 29500 -15890 29890 -15830
rect 28860 -15930 29257 -15890
rect 29493 -15930 29890 -15890
rect 30460 -15890 30850 -15830
rect 31100 -15890 31490 -15830
rect 31580 -15720 31720 -15710
rect 31580 -15840 31590 -15720
rect 31710 -15730 31720 -15720
rect 32060 -15730 32450 -15668
rect 32700 -15730 33090 -15668
rect 33660 -15668 34057 -15630
rect 34293 -15668 34690 -15630
rect 33660 -15730 34050 -15668
rect 34300 -15730 34690 -15668
rect 35260 -15668 35657 -15630
rect 35893 -15668 36290 -15630
rect 35260 -15730 35650 -15668
rect 35900 -15730 36290 -15668
rect 31710 -15830 36290 -15730
rect 31710 -15840 31720 -15830
rect 31580 -15850 31720 -15840
rect 30460 -15930 30857 -15890
rect 31093 -15930 31490 -15890
rect 32060 -15890 32450 -15830
rect 32700 -15890 33090 -15830
rect 33660 -15890 34050 -15830
rect 34300 -15890 34690 -15830
rect 35260 -15890 35650 -15830
rect 35900 -15890 36290 -15830
rect 32060 -15930 32457 -15890
rect 32340 -15936 32457 -15930
rect 32693 -15936 33093 -15890
rect 33657 -15936 34057 -15890
rect 34293 -15936 34693 -15890
rect 35257 -15936 35657 -15890
rect 35893 -15930 36290 -15890
rect 35893 -15936 36030 -15930
rect 32498 -15990 32544 -15984
rect 32606 -15990 32652 -15984
rect 16510 -16000 16640 -15990
rect 13310 -16010 13440 -16000
rect 11180 -16410 12360 -16290
rect 10120 -16680 10240 -16670
rect 11420 -16760 11500 -16410
rect 12040 -16760 12120 -16410
rect 13310 -16670 13320 -16010
rect 13430 -16670 13440 -16010
rect 13310 -16680 13440 -16670
rect 14910 -16010 15040 -16000
rect 14910 -16670 14920 -16010
rect 15030 -16670 15040 -16010
rect 14910 -16680 15040 -16670
rect 16510 -16680 16520 -16000
rect 16630 -16680 16640 -16000
rect 16510 -16690 16640 -16680
rect 18110 -16000 18240 -15990
rect 18110 -16680 18120 -16000
rect 18230 -16680 18240 -16000
rect 18110 -16690 18240 -16680
rect 19710 -16000 19840 -15990
rect 19710 -16680 19720 -16000
rect 19830 -16680 19840 -16000
rect 19710 -16690 19840 -16680
rect 21310 -16000 21440 -15990
rect 21310 -16680 21320 -16000
rect 21430 -16680 21440 -16000
rect 21310 -16690 21440 -16680
rect 22910 -16000 23040 -15990
rect 22910 -16680 22920 -16000
rect 23030 -16680 23040 -16000
rect 22910 -16690 23040 -16680
rect 24510 -16000 24640 -15990
rect 24510 -16680 24520 -16000
rect 24630 -16680 24640 -16000
rect 24510 -16690 24640 -16680
rect 26110 -16000 26240 -15990
rect 26110 -16680 26120 -16000
rect 26230 -16680 26240 -16000
rect 26110 -16690 26240 -16680
rect 27710 -16000 27840 -15990
rect 27710 -16680 27720 -16000
rect 27830 -16680 27840 -16000
rect 27710 -16690 27840 -16680
rect 29310 -16000 29440 -15990
rect 29310 -16680 29320 -16000
rect 29430 -16680 29440 -16000
rect 29310 -16690 29440 -16680
rect 30910 -16000 31040 -15990
rect 30910 -16680 30920 -16000
rect 31030 -16680 31040 -16000
rect 30910 -16690 31040 -16680
rect 32498 -15996 32652 -15990
rect 32498 -16688 32504 -15996
rect 32510 -16000 32640 -15996
rect 32510 -16680 32520 -16000
rect 32630 -16680 32640 -16000
rect 32510 -16688 32640 -16680
rect 32646 -16688 32652 -15996
rect 32498 -16690 32652 -16688
rect 32498 -16700 32544 -16690
rect 32606 -16700 32652 -16690
rect 33134 -15996 33180 -15984
rect 33134 -16688 33140 -15996
rect 33174 -16688 33180 -15996
rect 33134 -16700 33180 -16688
rect 33570 -15996 33616 -15984
rect 33570 -16688 33576 -15996
rect 33610 -16688 33616 -15996
rect 33570 -16700 33616 -16688
rect 34098 -15990 34144 -15984
rect 34206 -15990 34252 -15984
rect 34098 -15996 34252 -15990
rect 34098 -16688 34104 -15996
rect 34110 -16000 34240 -15996
rect 34110 -16680 34120 -16000
rect 34230 -16680 34240 -16000
rect 34110 -16688 34240 -16680
rect 34246 -16688 34252 -15996
rect 34098 -16690 34252 -16688
rect 34098 -16700 34144 -16690
rect 34206 -16700 34252 -16690
rect 34734 -15996 34780 -15984
rect 34734 -16688 34740 -15996
rect 34774 -16688 34780 -15996
rect 34734 -16700 34780 -16688
rect 35170 -15996 35216 -15984
rect 35170 -16688 35176 -15996
rect 35210 -16688 35216 -15996
rect 35170 -16700 35216 -16688
rect 35698 -15990 35744 -15984
rect 35806 -15990 35852 -15984
rect 35698 -15996 35852 -15990
rect 35698 -16688 35704 -15996
rect 35710 -16000 35840 -15996
rect 35710 -16680 35720 -16000
rect 35830 -16680 35840 -16000
rect 35710 -16688 35840 -16680
rect 35846 -16688 35852 -15996
rect 39100 -16600 39229 -15200
rect 35698 -16690 35852 -16688
rect 35698 -16700 35744 -16690
rect 35806 -16700 35852 -16690
rect 36700 -16760 39229 -16600
rect 670 -17000 39229 -16760
rect 670 -17020 37940 -17000
rect 670 -18560 720 -17020
rect 1200 -17070 1340 -17060
rect 1200 -17190 1210 -17070
rect 1330 -17080 1340 -17070
rect 2800 -17070 2940 -17060
rect 2800 -17080 2810 -17070
rect 1330 -17180 2810 -17080
rect 1330 -17190 1340 -17180
rect 1200 -17200 1340 -17190
rect 2800 -17190 2810 -17180
rect 2930 -17080 2940 -17070
rect 4400 -17070 4540 -17060
rect 4400 -17080 4410 -17070
rect 2930 -17180 4410 -17080
rect 2930 -17190 2940 -17180
rect 2800 -17200 2940 -17190
rect 4400 -17190 4410 -17180
rect 4530 -17080 4540 -17070
rect 6000 -17070 6140 -17060
rect 6000 -17080 6010 -17070
rect 4530 -17180 6010 -17080
rect 4530 -17190 4540 -17180
rect 4400 -17200 4540 -17190
rect 6000 -17190 6010 -17180
rect 6130 -17080 6140 -17070
rect 7600 -17070 7740 -17060
rect 7600 -17080 7610 -17070
rect 6130 -17180 7610 -17080
rect 6130 -17190 6140 -17180
rect 6000 -17200 6140 -17190
rect 7600 -17190 7610 -17180
rect 7730 -17080 7740 -17070
rect 9200 -17070 9340 -17060
rect 15820 -17070 15960 -17060
rect 9200 -17080 9210 -17070
rect 7730 -17180 9210 -17080
rect 7730 -17190 7740 -17180
rect 7600 -17200 7740 -17190
rect 9200 -17190 9210 -17180
rect 9330 -17080 9340 -17070
rect 12620 -17080 12760 -17070
rect 9330 -17180 10700 -17080
rect 9330 -17190 9340 -17180
rect 9200 -17200 9340 -17190
rect 10750 -17260 10940 -17250
rect 11380 -17260 11500 -17180
rect 12040 -17260 12160 -17180
rect 12620 -17200 12630 -17080
rect 12750 -17110 12760 -17080
rect 12750 -17200 15490 -17110
rect 15820 -17190 15830 -17070
rect 15950 -17100 15960 -17070
rect 17420 -17070 17560 -17060
rect 15950 -17190 17090 -17100
rect 15820 -17200 17090 -17190
rect 17420 -17190 17430 -17070
rect 17550 -17100 17560 -17070
rect 19020 -17070 19160 -17060
rect 17550 -17190 18690 -17100
rect 17420 -17200 18690 -17190
rect 19020 -17190 19030 -17070
rect 19150 -17100 19160 -17070
rect 20620 -17070 20760 -17060
rect 19150 -17190 20290 -17100
rect 19020 -17200 20290 -17190
rect 20620 -17190 20630 -17070
rect 20750 -17100 20760 -17070
rect 22220 -17070 22360 -17060
rect 20750 -17190 21890 -17100
rect 20620 -17200 21890 -17190
rect 22220 -17190 22230 -17070
rect 22350 -17100 22360 -17070
rect 23820 -17070 23960 -17060
rect 22350 -17190 23490 -17100
rect 22220 -17200 23490 -17190
rect 23820 -17190 23830 -17070
rect 23950 -17100 23960 -17070
rect 27020 -17070 27160 -17060
rect 27020 -17100 27030 -17070
rect 23950 -17190 25090 -17100
rect 23820 -17200 25090 -17190
rect 25660 -17190 27030 -17100
rect 27150 -17100 27160 -17070
rect 28620 -17070 28760 -17060
rect 27150 -17190 28290 -17100
rect 25660 -17200 28290 -17190
rect 28620 -17190 28630 -17070
rect 28750 -17100 28760 -17070
rect 31840 -17080 31980 -17070
rect 28750 -17190 31490 -17100
rect 28620 -17200 31490 -17190
rect 31840 -17200 31850 -17080
rect 31970 -17100 31980 -17080
rect 31970 -17200 36290 -17100
rect 12620 -17210 12760 -17200
rect 31840 -17210 31980 -17200
rect 1560 -17380 10810 -17260
rect 10930 -17380 36380 -17260
rect 10750 -17390 10940 -17380
rect 1420 -17510 1560 -17500
rect 1420 -17630 1430 -17510
rect 1550 -17520 1560 -17510
rect 1660 -17520 2060 -17430
rect 2290 -17520 2690 -17430
rect 3020 -17510 3160 -17500
rect 3020 -17520 3030 -17510
rect 1550 -17620 3030 -17520
rect 1550 -17630 1560 -17620
rect 1420 -17640 1560 -17630
rect 1660 -17640 2690 -17620
rect 3020 -17630 3030 -17620
rect 3150 -17520 3160 -17510
rect 3260 -17520 3660 -17430
rect 3890 -17520 4290 -17430
rect 4620 -17510 4760 -17500
rect 4620 -17520 4630 -17510
rect 3150 -17620 4630 -17520
rect 3150 -17630 3160 -17620
rect 3020 -17640 3160 -17630
rect 3260 -17640 4290 -17620
rect 4620 -17630 4630 -17620
rect 4750 -17520 4760 -17510
rect 4860 -17520 5260 -17430
rect 5490 -17520 5890 -17430
rect 6220 -17510 6360 -17500
rect 6220 -17520 6230 -17510
rect 4750 -17620 6230 -17520
rect 4750 -17630 4760 -17620
rect 4620 -17640 4760 -17630
rect 4860 -17640 5890 -17620
rect 6220 -17630 6230 -17620
rect 6350 -17520 6360 -17510
rect 6460 -17520 6860 -17430
rect 7090 -17520 7490 -17430
rect 7820 -17510 7960 -17500
rect 7820 -17520 7830 -17510
rect 6350 -17620 7830 -17520
rect 6350 -17630 6360 -17620
rect 6220 -17640 6360 -17630
rect 6460 -17640 7490 -17620
rect 7820 -17630 7830 -17620
rect 7950 -17520 7960 -17510
rect 8060 -17520 8460 -17430
rect 8690 -17520 9090 -17430
rect 9420 -17510 9560 -17500
rect 9420 -17520 9430 -17510
rect 7950 -17620 9430 -17520
rect 7950 -17630 7960 -17620
rect 7820 -17640 7960 -17630
rect 8060 -17640 9090 -17620
rect 9420 -17630 9430 -17620
rect 9550 -17520 9560 -17510
rect 9660 -17520 10060 -17430
rect 10290 -17520 10690 -17430
rect 11380 -17460 11500 -17380
rect 12040 -17460 12160 -17380
rect 9550 -17620 10690 -17520
rect 9550 -17630 9560 -17620
rect 9420 -17640 9560 -17630
rect 9660 -17640 10690 -17620
rect 1660 -17730 2060 -17640
rect 2290 -17730 2690 -17640
rect 3260 -17730 3660 -17640
rect 3890 -17730 4290 -17640
rect 4860 -17730 5260 -17640
rect 5490 -17730 5890 -17640
rect 6460 -17730 6860 -17640
rect 7090 -17730 7490 -17640
rect 8060 -17730 8460 -17640
rect 8690 -17730 9090 -17640
rect 9660 -17730 10060 -17640
rect 10290 -17730 10690 -17640
rect 12860 -17520 13260 -17430
rect 13490 -17520 13890 -17430
rect 14460 -17520 14860 -17430
rect 15090 -17520 15490 -17430
rect 12860 -17640 15490 -17520
rect 2120 -17810 2240 -17800
rect 2120 -17970 2130 -17810
rect 2120 -18470 2130 -18170
rect 2230 -17970 2240 -17810
rect 3720 -17810 3840 -17800
rect 3720 -17970 3730 -17810
rect 2230 -18470 2240 -18170
rect 2120 -18480 2240 -18470
rect 3720 -18470 3730 -18170
rect 3830 -17970 3840 -17810
rect 5320 -17810 5440 -17800
rect 5320 -17970 5330 -17810
rect 3830 -18470 3840 -18170
rect 3720 -18480 3840 -18470
rect 5320 -18470 5330 -18170
rect 5430 -17970 5440 -17810
rect 6920 -17810 7040 -17800
rect 6920 -17970 6930 -17810
rect 5430 -18470 5440 -18170
rect 5320 -18480 5440 -18470
rect 6920 -18470 6930 -18170
rect 7030 -17970 7040 -17810
rect 8520 -17810 8640 -17800
rect 7030 -18470 7040 -18170
rect 6920 -18480 7040 -18470
rect 8520 -18470 8530 -17810
rect 8630 -18470 8640 -17810
rect 8520 -18480 8640 -18470
rect 10120 -17810 10240 -17800
rect 10120 -18470 10130 -17810
rect 10230 -18470 10240 -17810
rect 11400 -18070 11510 -17700
rect 12040 -18070 12150 -17710
rect 12860 -17730 13260 -17640
rect 13490 -17730 13890 -17640
rect 14460 -17730 14860 -17640
rect 15090 -17730 15490 -17640
rect 15600 -17520 15740 -17510
rect 15600 -17640 15610 -17520
rect 15730 -17530 15740 -17520
rect 16060 -17530 16450 -17430
rect 16700 -17530 17090 -17430
rect 15730 -17630 17090 -17530
rect 15730 -17640 15740 -17630
rect 15600 -17650 15740 -17640
rect 16060 -17730 16450 -17630
rect 16700 -17730 17090 -17630
rect 17200 -17520 17340 -17510
rect 17200 -17640 17210 -17520
rect 17330 -17530 17340 -17520
rect 17660 -17530 18050 -17430
rect 18300 -17530 18690 -17430
rect 17330 -17630 18690 -17530
rect 17330 -17640 17340 -17630
rect 17200 -17650 17340 -17640
rect 17660 -17730 18050 -17630
rect 18300 -17730 18690 -17630
rect 18800 -17520 18940 -17510
rect 18800 -17640 18810 -17520
rect 18930 -17530 18940 -17520
rect 19260 -17530 19650 -17430
rect 19900 -17530 20290 -17430
rect 18930 -17630 20290 -17530
rect 18930 -17640 18940 -17630
rect 18800 -17650 18940 -17640
rect 19260 -17730 19650 -17630
rect 19900 -17730 20290 -17630
rect 20400 -17520 20540 -17510
rect 20400 -17640 20410 -17520
rect 20530 -17530 20540 -17520
rect 20860 -17530 21250 -17430
rect 21500 -17530 21890 -17430
rect 20530 -17630 21890 -17530
rect 20530 -17640 20540 -17630
rect 20400 -17650 20540 -17640
rect 20860 -17730 21250 -17630
rect 21500 -17730 21890 -17630
rect 22000 -17520 22140 -17510
rect 22000 -17640 22010 -17520
rect 22130 -17530 22140 -17520
rect 22460 -17530 22850 -17430
rect 23100 -17530 23490 -17430
rect 22130 -17630 23490 -17530
rect 22130 -17640 22140 -17630
rect 22000 -17650 22140 -17640
rect 22460 -17730 22850 -17630
rect 23100 -17730 23490 -17630
rect 23600 -17520 23740 -17510
rect 23600 -17640 23610 -17520
rect 23730 -17530 23740 -17520
rect 24060 -17530 24450 -17430
rect 24700 -17530 25090 -17430
rect 23730 -17630 25090 -17530
rect 23730 -17640 23740 -17630
rect 23600 -17650 23740 -17640
rect 24060 -17730 24450 -17630
rect 24700 -17730 25090 -17630
rect 25660 -17530 26050 -17430
rect 26300 -17530 26690 -17430
rect 27260 -17468 27657 -17430
rect 27893 -17468 28290 -17430
rect 26800 -17520 26940 -17510
rect 26800 -17530 26810 -17520
rect 25660 -17630 26810 -17530
rect 25660 -17730 26050 -17630
rect 26300 -17730 26690 -17630
rect 26800 -17640 26810 -17630
rect 26930 -17530 26940 -17520
rect 27260 -17530 27650 -17468
rect 27900 -17530 28290 -17468
rect 28860 -17468 29257 -17430
rect 29493 -17468 29890 -17430
rect 26930 -17630 28290 -17530
rect 26930 -17640 26940 -17630
rect 26800 -17650 26940 -17640
rect 27260 -17690 27650 -17630
rect 27900 -17690 28290 -17630
rect 28400 -17520 28540 -17510
rect 28400 -17640 28410 -17520
rect 28530 -17530 28540 -17520
rect 28860 -17530 29250 -17468
rect 29500 -17530 29890 -17468
rect 30460 -17468 30857 -17430
rect 31093 -17468 31490 -17430
rect 30460 -17530 30850 -17468
rect 31100 -17530 31490 -17468
rect 32060 -17468 32457 -17430
rect 32693 -17468 33090 -17430
rect 28530 -17630 31490 -17530
rect 28530 -17640 28540 -17630
rect 28400 -17650 28540 -17640
rect 27260 -17730 27657 -17690
rect 27893 -17730 28290 -17690
rect 28860 -17690 29250 -17630
rect 29500 -17690 29890 -17630
rect 28860 -17730 29257 -17690
rect 29493 -17730 29890 -17690
rect 30460 -17690 30850 -17630
rect 31100 -17690 31490 -17630
rect 31580 -17520 31720 -17510
rect 31580 -17640 31590 -17520
rect 31710 -17540 31720 -17520
rect 32060 -17530 32450 -17468
rect 32700 -17530 33090 -17468
rect 33660 -17468 34057 -17430
rect 34293 -17468 34690 -17430
rect 33660 -17530 34050 -17468
rect 34300 -17530 34690 -17468
rect 35260 -17468 35657 -17430
rect 35893 -17468 36290 -17430
rect 35260 -17530 35650 -17468
rect 35900 -17530 36290 -17468
rect 32060 -17540 36290 -17530
rect 31710 -17630 36290 -17540
rect 31710 -17640 31720 -17630
rect 31580 -17650 31720 -17640
rect 30460 -17730 30857 -17690
rect 31093 -17730 31490 -17690
rect 32060 -17690 32450 -17630
rect 32700 -17690 33090 -17630
rect 32060 -17730 32457 -17690
rect 32693 -17730 33090 -17690
rect 33660 -17690 34050 -17630
rect 34300 -17690 34690 -17630
rect 33660 -17730 34057 -17690
rect 34293 -17730 34690 -17690
rect 35260 -17690 35650 -17630
rect 35900 -17690 36290 -17630
rect 35260 -17730 35657 -17690
rect 35893 -17730 36290 -17690
rect 16510 -17800 16640 -17790
rect 13310 -17810 13440 -17800
rect 11200 -18220 12360 -18070
rect 10120 -18480 10240 -18470
rect 11400 -18560 11510 -18220
rect 12040 -18560 12150 -18220
rect 13310 -18470 13320 -17810
rect 13430 -18470 13440 -17810
rect 13310 -18480 13440 -18470
rect 14910 -17810 15040 -17800
rect 14910 -18470 14920 -17810
rect 15030 -18470 15040 -17810
rect 14910 -18480 15040 -18470
rect 16510 -18480 16520 -17800
rect 16630 -18480 16640 -17800
rect 16510 -18490 16640 -18480
rect 18110 -17800 18240 -17790
rect 18110 -18480 18120 -17800
rect 18230 -18480 18240 -17800
rect 18110 -18490 18240 -18480
rect 19710 -17800 19840 -17790
rect 19710 -18480 19720 -17800
rect 19830 -18480 19840 -17800
rect 19710 -18490 19840 -18480
rect 21310 -17800 21440 -17790
rect 21310 -18480 21320 -17800
rect 21430 -18480 21440 -17800
rect 21310 -18490 21440 -18480
rect 22910 -17800 23040 -17790
rect 22910 -18480 22920 -17800
rect 23030 -18480 23040 -17800
rect 22910 -18490 23040 -18480
rect 24510 -17800 24640 -17790
rect 24510 -18480 24520 -17800
rect 24630 -18480 24640 -17800
rect 24510 -18490 24640 -18480
rect 26110 -17800 26240 -17790
rect 26110 -18480 26120 -17800
rect 26230 -18480 26240 -17800
rect 26110 -18490 26240 -18480
rect 27710 -17800 27840 -17790
rect 27710 -18480 27720 -17800
rect 27830 -18480 27840 -17800
rect 27710 -18490 27840 -18480
rect 29310 -17800 29440 -17790
rect 29310 -18480 29320 -17800
rect 29430 -18480 29440 -17800
rect 29310 -18490 29440 -18480
rect 30910 -17800 31040 -17790
rect 30910 -18480 30920 -17800
rect 31030 -18480 31040 -17800
rect 30910 -18490 31040 -18480
rect 32510 -17800 32640 -17790
rect 32510 -18480 32520 -17800
rect 32630 -18480 32640 -17800
rect 32510 -18490 32640 -18480
rect 34110 -17800 34240 -17790
rect 34110 -18480 34120 -17800
rect 34230 -18480 34240 -17800
rect 34110 -18490 34240 -18480
rect 35710 -17800 35840 -17790
rect 35710 -18480 35720 -17800
rect 35830 -18480 35840 -17800
rect 35710 -18490 35840 -18480
rect 670 -18700 37880 -18560
rect 39100 -18700 39229 -17000
rect 670 -18800 39229 -18700
rect 670 -18820 37940 -18800
rect 670 -20380 720 -18820
rect 1200 -18870 1340 -18860
rect 1200 -18990 1210 -18870
rect 1330 -18880 1340 -18870
rect 2800 -18870 2940 -18860
rect 2800 -18880 2810 -18870
rect 1330 -18980 2810 -18880
rect 1330 -18990 1340 -18980
rect 1200 -19000 1340 -18990
rect 2800 -18990 2810 -18980
rect 2930 -18880 2940 -18870
rect 4400 -18870 4540 -18860
rect 4400 -18880 4410 -18870
rect 2930 -18980 4410 -18880
rect 2930 -18990 2940 -18980
rect 2800 -19000 2940 -18990
rect 4400 -18990 4410 -18980
rect 4530 -18880 4540 -18870
rect 6000 -18870 6140 -18860
rect 6000 -18880 6010 -18870
rect 4530 -18980 6010 -18880
rect 4530 -18990 4540 -18980
rect 4400 -19000 4540 -18990
rect 6000 -18990 6010 -18980
rect 6130 -18880 6140 -18870
rect 7600 -18870 7740 -18860
rect 7600 -18880 7610 -18870
rect 6130 -18980 7610 -18880
rect 6130 -18990 6140 -18980
rect 6000 -19000 6140 -18990
rect 7600 -18990 7610 -18980
rect 7730 -18880 7740 -18870
rect 9200 -18870 9340 -18860
rect 15820 -18870 15960 -18860
rect 9200 -18880 9210 -18870
rect 7730 -18980 9210 -18880
rect 7730 -18990 7740 -18980
rect 7600 -19000 7740 -18990
rect 9200 -18990 9210 -18980
rect 9330 -18880 9340 -18870
rect 12400 -18880 12540 -18870
rect 9330 -18980 10700 -18880
rect 9330 -18990 9340 -18980
rect 9200 -19000 9340 -18990
rect 10750 -19060 10940 -19050
rect 11400 -19060 11520 -18980
rect 12040 -19060 12160 -18980
rect 12400 -19000 12410 -18880
rect 12530 -18910 12540 -18880
rect 12530 -19000 15490 -18910
rect 15820 -18990 15830 -18870
rect 15950 -18900 15960 -18870
rect 17420 -18870 17560 -18860
rect 15950 -18990 17090 -18900
rect 15820 -19000 17090 -18990
rect 17420 -18990 17430 -18870
rect 17550 -18900 17560 -18870
rect 19020 -18870 19160 -18860
rect 17550 -18990 18690 -18900
rect 17420 -19000 18690 -18990
rect 19020 -18990 19030 -18870
rect 19150 -18900 19160 -18870
rect 20620 -18870 20760 -18860
rect 19150 -18990 20290 -18900
rect 19020 -19000 20290 -18990
rect 20620 -18990 20630 -18870
rect 20750 -18900 20760 -18870
rect 22220 -18870 22360 -18860
rect 20750 -18990 21890 -18900
rect 20620 -19000 21890 -18990
rect 22220 -18990 22230 -18870
rect 22350 -18900 22360 -18870
rect 23820 -18870 23960 -18860
rect 22350 -18990 23490 -18900
rect 22220 -19000 23490 -18990
rect 23820 -18990 23830 -18870
rect 23950 -18900 23960 -18870
rect 27020 -18870 27160 -18860
rect 27020 -18900 27030 -18870
rect 23950 -18990 25090 -18900
rect 23820 -19000 25090 -18990
rect 25660 -18990 27030 -18900
rect 27150 -18900 27160 -18870
rect 28620 -18870 28760 -18860
rect 27150 -18990 28290 -18900
rect 25660 -19000 28290 -18990
rect 28620 -18990 28630 -18870
rect 28750 -18900 28760 -18870
rect 31580 -18880 31720 -18870
rect 28750 -18990 31490 -18900
rect 28620 -19000 31490 -18990
rect 31580 -19000 31590 -18880
rect 31710 -18900 31720 -18880
rect 31710 -19000 36280 -18900
rect 12400 -19010 12540 -19000
rect 31580 -19010 31720 -19000
rect 1560 -19180 10810 -19060
rect 10930 -19180 36380 -19060
rect 10750 -19190 10940 -19180
rect 1420 -19310 1560 -19300
rect 1420 -19430 1430 -19310
rect 1550 -19320 1560 -19310
rect 1660 -19320 2060 -19230
rect 2290 -19320 2690 -19230
rect 3020 -19310 3160 -19300
rect 3020 -19320 3030 -19310
rect 1550 -19420 3030 -19320
rect 1550 -19430 1560 -19420
rect 1420 -19440 1560 -19430
rect 1660 -19440 2690 -19420
rect 3020 -19430 3030 -19420
rect 3150 -19320 3160 -19310
rect 3260 -19320 3660 -19230
rect 3890 -19320 4290 -19230
rect 4620 -19310 4760 -19300
rect 4620 -19320 4630 -19310
rect 3150 -19420 4630 -19320
rect 3150 -19430 3160 -19420
rect 3020 -19440 3160 -19430
rect 3260 -19440 4290 -19420
rect 4620 -19430 4630 -19420
rect 4750 -19320 4760 -19310
rect 4860 -19320 5260 -19230
rect 5490 -19320 5890 -19230
rect 6220 -19310 6360 -19300
rect 6220 -19320 6230 -19310
rect 4750 -19420 6230 -19320
rect 4750 -19430 4760 -19420
rect 4620 -19440 4760 -19430
rect 4860 -19440 5890 -19420
rect 6220 -19430 6230 -19420
rect 6350 -19320 6360 -19310
rect 6460 -19320 6860 -19230
rect 7090 -19320 7490 -19230
rect 7820 -19310 7960 -19300
rect 7820 -19320 7830 -19310
rect 6350 -19420 7830 -19320
rect 6350 -19430 6360 -19420
rect 6220 -19440 6360 -19430
rect 6460 -19440 7490 -19420
rect 7820 -19430 7830 -19420
rect 7950 -19320 7960 -19310
rect 8060 -19320 8460 -19230
rect 8690 -19320 9090 -19230
rect 9420 -19310 9560 -19300
rect 9420 -19320 9430 -19310
rect 7950 -19420 9430 -19320
rect 7950 -19430 7960 -19420
rect 7820 -19440 7960 -19430
rect 8060 -19440 9090 -19420
rect 9420 -19430 9430 -19420
rect 9550 -19320 9560 -19310
rect 9660 -19320 10060 -19230
rect 10290 -19320 10690 -19230
rect 11400 -19260 11520 -19180
rect 12040 -19260 12160 -19180
rect 9550 -19420 10690 -19320
rect 9550 -19430 9560 -19420
rect 9420 -19440 9560 -19430
rect 9660 -19440 10690 -19420
rect 1660 -19530 2060 -19440
rect 2290 -19530 2690 -19440
rect 3260 -19530 3660 -19440
rect 3890 -19530 4290 -19440
rect 4860 -19530 5260 -19440
rect 5490 -19530 5890 -19440
rect 6460 -19530 6860 -19440
rect 7090 -19530 7490 -19440
rect 8060 -19530 8460 -19440
rect 8690 -19530 9090 -19440
rect 9660 -19530 10060 -19440
rect 10290 -19530 10690 -19440
rect 12860 -19320 13260 -19230
rect 13490 -19320 13890 -19230
rect 14460 -19320 14860 -19230
rect 15090 -19320 15490 -19230
rect 12860 -19440 15490 -19320
rect 2120 -19610 2240 -19600
rect 2120 -20170 2130 -19610
rect 2230 -20170 2240 -19610
rect 3720 -19610 3840 -19600
rect 3720 -20170 3730 -19610
rect 3830 -20170 3840 -19610
rect 5320 -19610 5440 -19600
rect 5320 -20170 5330 -19610
rect 5430 -20170 5440 -19610
rect 6920 -19610 7040 -19600
rect 6920 -20170 6930 -19610
rect 7030 -20170 7040 -19610
rect 8520 -19610 8640 -19600
rect 8520 -20270 8530 -19610
rect 8630 -20270 8640 -19610
rect 8520 -20280 8640 -20270
rect 10120 -19610 10240 -19600
rect 10120 -20270 10130 -19610
rect 10230 -20270 10240 -19610
rect 11370 -19840 11510 -19510
rect 12030 -19840 12140 -19510
rect 12860 -19530 13260 -19440
rect 13490 -19530 13890 -19440
rect 14460 -19530 14860 -19440
rect 15090 -19530 15490 -19440
rect 15600 -19320 15740 -19310
rect 15600 -19440 15610 -19320
rect 15730 -19330 15740 -19320
rect 16060 -19330 16450 -19230
rect 16700 -19330 17090 -19230
rect 15730 -19430 17090 -19330
rect 15730 -19440 15740 -19430
rect 15600 -19450 15740 -19440
rect 16060 -19530 16450 -19430
rect 16700 -19530 17090 -19430
rect 17200 -19320 17340 -19310
rect 17200 -19440 17210 -19320
rect 17330 -19330 17340 -19320
rect 17660 -19330 18050 -19230
rect 18300 -19330 18690 -19230
rect 17330 -19430 18690 -19330
rect 17330 -19440 17340 -19430
rect 17200 -19450 17340 -19440
rect 17660 -19530 18050 -19430
rect 18300 -19530 18690 -19430
rect 18800 -19320 18940 -19310
rect 18800 -19440 18810 -19320
rect 18930 -19330 18940 -19320
rect 19260 -19330 19650 -19230
rect 19900 -19330 20290 -19230
rect 18930 -19430 20290 -19330
rect 18930 -19440 18940 -19430
rect 18800 -19450 18940 -19440
rect 19260 -19530 19650 -19430
rect 19900 -19530 20290 -19430
rect 20400 -19320 20540 -19310
rect 20400 -19440 20410 -19320
rect 20530 -19330 20540 -19320
rect 20860 -19330 21250 -19230
rect 21500 -19330 21890 -19230
rect 20530 -19430 21890 -19330
rect 20530 -19440 20540 -19430
rect 20400 -19450 20540 -19440
rect 20860 -19530 21250 -19430
rect 21500 -19530 21890 -19430
rect 22000 -19320 22140 -19310
rect 22000 -19440 22010 -19320
rect 22130 -19330 22140 -19320
rect 22460 -19330 22850 -19230
rect 23100 -19330 23490 -19230
rect 22130 -19430 23490 -19330
rect 22130 -19440 22140 -19430
rect 22000 -19450 22140 -19440
rect 22460 -19530 22850 -19430
rect 23100 -19530 23490 -19430
rect 23600 -19320 23740 -19310
rect 23600 -19440 23610 -19320
rect 23730 -19330 23740 -19320
rect 24060 -19330 24450 -19230
rect 24700 -19330 25090 -19230
rect 23730 -19430 25090 -19330
rect 23730 -19440 23740 -19430
rect 23600 -19450 23740 -19440
rect 24060 -19530 24450 -19430
rect 24700 -19530 25090 -19430
rect 25660 -19330 26050 -19230
rect 26300 -19330 26690 -19230
rect 27260 -19268 27657 -19230
rect 27893 -19268 28290 -19230
rect 26800 -19320 26940 -19310
rect 26800 -19330 26810 -19320
rect 25660 -19430 26810 -19330
rect 25660 -19530 26050 -19430
rect 26300 -19530 26690 -19430
rect 26800 -19440 26810 -19430
rect 26930 -19330 26940 -19320
rect 27260 -19330 27650 -19268
rect 27900 -19330 28290 -19268
rect 28860 -19268 29257 -19230
rect 29493 -19268 29890 -19230
rect 26930 -19430 28290 -19330
rect 26930 -19440 26940 -19430
rect 26800 -19450 26940 -19440
rect 27260 -19490 27650 -19430
rect 27900 -19490 28290 -19430
rect 28400 -19320 28540 -19310
rect 28400 -19440 28410 -19320
rect 28530 -19330 28540 -19320
rect 28860 -19330 29250 -19268
rect 29500 -19330 29890 -19268
rect 30460 -19268 30857 -19230
rect 31093 -19268 31490 -19230
rect 30460 -19330 30850 -19268
rect 31100 -19330 31490 -19268
rect 28530 -19430 31490 -19330
rect 28530 -19440 28540 -19430
rect 28400 -19450 28540 -19440
rect 27260 -19530 27657 -19490
rect 27893 -19530 28290 -19490
rect 28860 -19490 29250 -19430
rect 29500 -19490 29890 -19430
rect 28860 -19530 29257 -19490
rect 29493 -19530 29890 -19490
rect 30460 -19490 30850 -19430
rect 31100 -19490 31490 -19430
rect 30460 -19530 30857 -19490
rect 31093 -19530 31490 -19490
rect 31740 -19240 31820 -19230
rect 31740 -19520 31750 -19240
rect 31810 -19330 31820 -19240
rect 32060 -19268 32457 -19230
rect 32693 -19268 33090 -19230
rect 32060 -19330 32450 -19268
rect 32700 -19330 33090 -19268
rect 33660 -19268 34057 -19230
rect 34293 -19268 34690 -19230
rect 33660 -19330 34050 -19268
rect 34300 -19330 34690 -19268
rect 35260 -19268 35657 -19230
rect 35893 -19268 36290 -19230
rect 35260 -19330 35650 -19268
rect 35900 -19330 36290 -19268
rect 31810 -19430 36290 -19330
rect 31810 -19520 31820 -19430
rect 31740 -19530 31820 -19520
rect 32060 -19490 32450 -19430
rect 32700 -19490 33090 -19430
rect 32060 -19530 32457 -19490
rect 32693 -19530 33090 -19490
rect 33660 -19490 34050 -19430
rect 34300 -19490 34690 -19430
rect 33660 -19530 34057 -19490
rect 34293 -19530 34690 -19490
rect 35260 -19490 35650 -19430
rect 35900 -19490 36290 -19430
rect 35260 -19530 35657 -19490
rect 35893 -19530 36290 -19490
rect 16510 -19600 16640 -19590
rect 13310 -19610 13440 -19600
rect 11200 -20030 12370 -19840
rect 10120 -20280 10240 -20270
rect 11370 -20380 11510 -20030
rect 12030 -20380 12140 -20030
rect 13310 -20270 13320 -19610
rect 13430 -20270 13440 -19610
rect 13310 -20280 13440 -20270
rect 14910 -19610 15040 -19600
rect 14910 -20270 14920 -19610
rect 15030 -20270 15040 -19610
rect 14910 -20280 15040 -20270
rect 16510 -20280 16520 -19600
rect 16630 -20280 16640 -19600
rect 16510 -20290 16640 -20280
rect 18110 -19600 18240 -19590
rect 18110 -20280 18120 -19600
rect 18230 -20280 18240 -19600
rect 18110 -20290 18240 -20280
rect 19710 -19600 19840 -19590
rect 19710 -20280 19720 -19600
rect 19830 -20280 19840 -19600
rect 19710 -20290 19840 -20280
rect 21310 -19600 21440 -19590
rect 21310 -20280 21320 -19600
rect 21430 -20280 21440 -19600
rect 21310 -20290 21440 -20280
rect 22910 -19600 23040 -19590
rect 22910 -20280 22920 -19600
rect 23030 -20280 23040 -19600
rect 22910 -20290 23040 -20280
rect 24510 -19600 24640 -19590
rect 24510 -20280 24520 -19600
rect 24630 -20280 24640 -19600
rect 24510 -20290 24640 -20280
rect 26110 -19600 26240 -19590
rect 26110 -20280 26120 -19600
rect 26230 -20280 26240 -19600
rect 26110 -20290 26240 -20280
rect 27710 -19600 27840 -19590
rect 27710 -20280 27720 -19600
rect 27830 -20280 27840 -19600
rect 27710 -20290 27840 -20280
rect 29310 -19600 29440 -19590
rect 29310 -20280 29320 -19600
rect 29430 -20280 29440 -19600
rect 29310 -20290 29440 -20280
rect 30910 -19600 31040 -19590
rect 30910 -20280 30920 -19600
rect 31030 -20280 31040 -19600
rect 30910 -20290 31040 -20280
rect 32510 -19600 32640 -19590
rect 32510 -20280 32520 -19600
rect 32630 -20280 32640 -19600
rect 32510 -20290 32640 -20280
rect 34110 -19600 34240 -19590
rect 34110 -20280 34120 -19600
rect 34230 -20280 34240 -19600
rect 34110 -20290 34240 -20280
rect 35710 -19600 35840 -19590
rect 35710 -20280 35720 -19600
rect 35830 -20280 35840 -19600
rect 35710 -20290 35840 -20280
rect 33180 -20340 33320 -20330
rect 32060 -20360 32330 -20350
rect 33180 -20360 33190 -20340
rect 670 -20500 31480 -20380
rect 32060 -20450 33190 -20360
rect 33180 -20460 33190 -20450
rect 33310 -20360 33320 -20340
rect 33310 -20450 36280 -20360
rect 33310 -20460 33320 -20450
rect 33180 -20470 33320 -20460
rect 39100 -20500 39229 -18800
rect 670 -20600 39229 -20500
rect 670 -20620 37940 -20600
rect 670 -22160 720 -20620
rect 1200 -20670 1340 -20660
rect 1200 -20790 1210 -20670
rect 1330 -20680 1340 -20670
rect 2800 -20670 2940 -20660
rect 2800 -20680 2810 -20670
rect 1330 -20780 2810 -20680
rect 1330 -20790 1340 -20780
rect 1200 -20800 1340 -20790
rect 2800 -20790 2810 -20780
rect 2930 -20680 2940 -20670
rect 4400 -20670 4540 -20660
rect 4400 -20680 4410 -20670
rect 2930 -20780 4410 -20680
rect 2930 -20790 2940 -20780
rect 2800 -20800 2940 -20790
rect 4400 -20790 4410 -20780
rect 4530 -20680 4540 -20670
rect 6000 -20670 6140 -20660
rect 6000 -20680 6010 -20670
rect 4530 -20780 6010 -20680
rect 4530 -20790 4540 -20780
rect 4400 -20800 4540 -20790
rect 6000 -20790 6010 -20780
rect 6130 -20680 6140 -20670
rect 7600 -20670 7740 -20660
rect 7600 -20680 7610 -20670
rect 6130 -20780 7610 -20680
rect 6130 -20790 6140 -20780
rect 6000 -20800 6140 -20790
rect 7600 -20790 7610 -20780
rect 7730 -20680 7740 -20670
rect 9200 -20670 9340 -20660
rect 15820 -20670 15960 -20660
rect 9200 -20680 9210 -20670
rect 7730 -20780 9210 -20680
rect 7730 -20790 7740 -20780
rect 7600 -20800 7740 -20790
rect 9200 -20790 9210 -20780
rect 9330 -20680 9340 -20670
rect 12400 -20680 12540 -20670
rect 9330 -20780 10700 -20680
rect 12400 -20700 12410 -20680
rect 9330 -20790 9340 -20780
rect 9200 -20800 9340 -20790
rect 11260 -20800 12410 -20700
rect 12530 -20800 12540 -20680
rect 12400 -20810 12540 -20800
rect 10750 -20860 10940 -20850
rect 13000 -20860 13120 -20780
rect 13640 -20860 13760 -20780
rect 14600 -20860 14720 -20780
rect 15240 -20860 15360 -20780
rect 15820 -20790 15830 -20670
rect 15950 -20700 15960 -20670
rect 17420 -20670 17560 -20660
rect 15950 -20790 17090 -20700
rect 15820 -20800 17090 -20790
rect 17420 -20790 17430 -20670
rect 17550 -20700 17560 -20670
rect 19020 -20670 19160 -20660
rect 17550 -20790 18690 -20700
rect 17420 -20800 18690 -20790
rect 19020 -20790 19030 -20670
rect 19150 -20700 19160 -20670
rect 20620 -20670 20760 -20660
rect 19150 -20790 20290 -20700
rect 19020 -20800 20290 -20790
rect 20620 -20790 20630 -20670
rect 20750 -20700 20760 -20670
rect 22220 -20670 22360 -20660
rect 20750 -20790 21890 -20700
rect 20620 -20800 21890 -20790
rect 22220 -20790 22230 -20670
rect 22350 -20700 22360 -20670
rect 23820 -20670 23960 -20660
rect 22350 -20790 23490 -20700
rect 22220 -20800 23490 -20790
rect 23820 -20790 23830 -20670
rect 23950 -20700 23960 -20670
rect 27020 -20670 27160 -20660
rect 27020 -20700 27030 -20670
rect 23950 -20790 25090 -20700
rect 23820 -20800 25090 -20790
rect 25660 -20790 27030 -20700
rect 27150 -20700 27160 -20670
rect 28620 -20670 28760 -20660
rect 27150 -20790 28290 -20700
rect 25660 -20800 28290 -20790
rect 28620 -20790 28630 -20670
rect 28750 -20700 28760 -20670
rect 31580 -20680 31720 -20670
rect 28750 -20790 31490 -20700
rect 28620 -20800 31490 -20790
rect 31580 -20800 31590 -20680
rect 31710 -20700 31720 -20680
rect 31710 -20800 36280 -20700
rect 31580 -20810 31720 -20800
rect 1560 -20980 10810 -20860
rect 10930 -20980 36380 -20860
rect 10750 -20990 10940 -20980
rect 1420 -21110 1560 -21100
rect 1420 -21230 1430 -21110
rect 1550 -21120 1560 -21110
rect 1660 -21120 2060 -21030
rect 2290 -21120 2690 -21030
rect 3020 -21110 3160 -21100
rect 3020 -21120 3030 -21110
rect 1550 -21220 3030 -21120
rect 1550 -21230 1560 -21220
rect 1420 -21240 1560 -21230
rect 1660 -21240 2690 -21220
rect 3020 -21230 3030 -21220
rect 3150 -21120 3160 -21110
rect 3260 -21120 3660 -21030
rect 3890 -21120 4290 -21030
rect 4620 -21110 4760 -21100
rect 4620 -21120 4630 -21110
rect 3150 -21220 4630 -21120
rect 3150 -21230 3160 -21220
rect 3020 -21240 3160 -21230
rect 3260 -21240 4290 -21220
rect 4620 -21230 4630 -21220
rect 4750 -21120 4760 -21110
rect 4860 -21120 5260 -21030
rect 5490 -21120 5890 -21030
rect 6220 -21110 6360 -21100
rect 6220 -21120 6230 -21110
rect 4750 -21220 6230 -21120
rect 4750 -21230 4760 -21220
rect 4620 -21240 4760 -21230
rect 4860 -21240 5890 -21220
rect 6220 -21230 6230 -21220
rect 6350 -21120 6360 -21110
rect 6460 -21120 6860 -21030
rect 7090 -21120 7490 -21030
rect 7820 -21110 7960 -21100
rect 7820 -21120 7830 -21110
rect 6350 -21220 7830 -21120
rect 6350 -21230 6360 -21220
rect 6220 -21240 6360 -21230
rect 6460 -21240 7490 -21220
rect 7820 -21230 7830 -21220
rect 7950 -21120 7960 -21110
rect 8060 -21120 8460 -21030
rect 8690 -21120 9090 -21030
rect 9420 -21110 9560 -21100
rect 9420 -21120 9430 -21110
rect 7950 -21220 9430 -21120
rect 7950 -21230 7960 -21220
rect 7820 -21240 7960 -21230
rect 8060 -21240 9090 -21220
rect 9420 -21230 9430 -21220
rect 9550 -21120 9560 -21110
rect 9660 -21120 10060 -21030
rect 10290 -21120 10690 -21030
rect 9550 -21220 10690 -21120
rect 9550 -21230 9560 -21220
rect 9420 -21240 9560 -21230
rect 9660 -21240 10690 -21220
rect 1660 -21330 2060 -21240
rect 2290 -21330 2690 -21240
rect 3260 -21330 3660 -21240
rect 3890 -21330 4290 -21240
rect 4860 -21330 5260 -21240
rect 5490 -21330 5890 -21240
rect 6460 -21330 6860 -21240
rect 7090 -21330 7490 -21240
rect 8060 -21330 8460 -21240
rect 8690 -21330 9090 -21240
rect 9660 -21330 10060 -21240
rect 10290 -21330 10690 -21240
rect 11260 -21120 11660 -21030
rect 11890 -21120 12290 -21030
rect 13000 -21060 13120 -20980
rect 13640 -21060 13760 -20980
rect 14600 -21060 14720 -20980
rect 15240 -21060 15360 -20980
rect 11260 -21240 12290 -21120
rect 11260 -21330 11660 -21240
rect 11890 -21330 12290 -21240
rect 15600 -21120 15740 -21110
rect 15600 -21240 15610 -21120
rect 15730 -21130 15740 -21120
rect 16060 -21130 16450 -21030
rect 16700 -21130 17090 -21030
rect 15730 -21230 17090 -21130
rect 15730 -21240 15740 -21230
rect 15600 -21250 15740 -21240
rect 11700 -21400 11850 -21390
rect 2120 -21410 2240 -21400
rect 2120 -21490 2130 -21410
rect 2120 -22070 2130 -21690
rect 2230 -21490 2240 -21410
rect 3720 -21410 3840 -21400
rect 3720 -21490 3730 -21410
rect 2230 -22070 2240 -21690
rect 2120 -22080 2240 -22070
rect 3720 -22070 3730 -21690
rect 3830 -21490 3840 -21410
rect 5320 -21410 5440 -21400
rect 5320 -21490 5330 -21410
rect 3830 -22070 3840 -21690
rect 3720 -22080 3840 -22070
rect 5320 -22070 5330 -21690
rect 5430 -21490 5440 -21410
rect 6920 -21410 7040 -21400
rect 6920 -21490 6930 -21410
rect 5430 -22070 5440 -21690
rect 5320 -22080 5440 -22070
rect 6920 -22070 6930 -21690
rect 7030 -21490 7040 -21410
rect 8520 -21410 8640 -21400
rect 7030 -22070 7040 -21690
rect 6920 -22080 7040 -22070
rect 8520 -22070 8530 -21410
rect 8630 -22070 8640 -21410
rect 8520 -22080 8640 -22070
rect 10120 -21410 10240 -21400
rect 10120 -22070 10130 -21410
rect 10230 -22070 10240 -21410
rect 10120 -22080 10240 -22070
rect 11700 -22080 11710 -21400
rect 11840 -22080 11850 -21400
rect 13010 -21650 13110 -21320
rect 13640 -21650 13740 -21300
rect 14630 -21640 14700 -21310
rect 15260 -21640 15330 -21300
rect 16060 -21330 16450 -21230
rect 16700 -21330 17090 -21230
rect 17200 -21120 17340 -21110
rect 17200 -21240 17210 -21120
rect 17330 -21130 17340 -21120
rect 17660 -21130 18050 -21030
rect 18300 -21130 18690 -21030
rect 17330 -21230 18690 -21130
rect 17330 -21240 17340 -21230
rect 17200 -21250 17340 -21240
rect 17660 -21330 18050 -21230
rect 18300 -21330 18690 -21230
rect 18800 -21120 18940 -21110
rect 18800 -21240 18810 -21120
rect 18930 -21130 18940 -21120
rect 19260 -21130 19650 -21030
rect 19900 -21130 20290 -21030
rect 18930 -21230 20290 -21130
rect 18930 -21240 18940 -21230
rect 18800 -21250 18940 -21240
rect 19260 -21330 19650 -21230
rect 19900 -21330 20290 -21230
rect 20400 -21120 20540 -21110
rect 20400 -21240 20410 -21120
rect 20530 -21130 20540 -21120
rect 20860 -21130 21250 -21030
rect 21500 -21130 21890 -21030
rect 20530 -21230 21890 -21130
rect 20530 -21240 20540 -21230
rect 20400 -21250 20540 -21240
rect 20860 -21330 21250 -21230
rect 21500 -21330 21890 -21230
rect 22000 -21120 22140 -21110
rect 22000 -21240 22010 -21120
rect 22130 -21130 22140 -21120
rect 22460 -21130 22850 -21030
rect 23100 -21130 23490 -21030
rect 22130 -21230 23490 -21130
rect 22130 -21240 22140 -21230
rect 22000 -21250 22140 -21240
rect 22460 -21330 22850 -21230
rect 23100 -21330 23490 -21230
rect 23600 -21120 23740 -21110
rect 23600 -21240 23610 -21120
rect 23730 -21130 23740 -21120
rect 24060 -21130 24450 -21030
rect 24700 -21130 25090 -21030
rect 23730 -21230 25090 -21130
rect 23730 -21240 23740 -21230
rect 23600 -21250 23740 -21240
rect 24060 -21330 24450 -21230
rect 24700 -21330 25090 -21230
rect 25660 -21130 26050 -21030
rect 26300 -21130 26690 -21030
rect 27260 -21068 27657 -21030
rect 27893 -21068 28290 -21030
rect 26800 -21120 26940 -21110
rect 26800 -21130 26810 -21120
rect 25660 -21230 26810 -21130
rect 25660 -21330 26050 -21230
rect 26300 -21330 26690 -21230
rect 26800 -21240 26810 -21230
rect 26930 -21130 26940 -21120
rect 27260 -21130 27650 -21068
rect 27900 -21130 28290 -21068
rect 28860 -21068 29257 -21030
rect 29493 -21068 29890 -21030
rect 26930 -21230 28290 -21130
rect 26930 -21240 26940 -21230
rect 26800 -21250 26940 -21240
rect 27260 -21290 27650 -21230
rect 27900 -21290 28290 -21230
rect 28400 -21120 28540 -21110
rect 28400 -21240 28410 -21120
rect 28530 -21130 28540 -21120
rect 28860 -21130 29250 -21068
rect 29500 -21130 29890 -21068
rect 30460 -21068 30857 -21030
rect 31093 -21068 31490 -21030
rect 30460 -21130 30850 -21068
rect 31100 -21130 31490 -21068
rect 28530 -21230 31490 -21130
rect 28530 -21240 28540 -21230
rect 28400 -21250 28540 -21240
rect 27260 -21330 27657 -21290
rect 27893 -21330 28290 -21290
rect 28860 -21290 29250 -21230
rect 29500 -21290 29890 -21230
rect 28860 -21330 29257 -21290
rect 29493 -21330 29890 -21290
rect 30460 -21290 30850 -21230
rect 31100 -21290 31490 -21230
rect 30460 -21330 30857 -21290
rect 31093 -21330 31490 -21290
rect 31740 -21040 31820 -21030
rect 31740 -21320 31750 -21040
rect 31810 -21130 31820 -21040
rect 32060 -21068 32457 -21030
rect 32693 -21068 33090 -21030
rect 32060 -21130 32450 -21068
rect 32700 -21130 33090 -21068
rect 31810 -21230 33090 -21130
rect 31810 -21320 31820 -21230
rect 31740 -21330 31820 -21320
rect 32060 -21290 32450 -21230
rect 32700 -21290 33090 -21230
rect 33660 -21068 34057 -21030
rect 34293 -21068 34690 -21030
rect 33660 -21130 34050 -21068
rect 34300 -21130 34690 -21068
rect 35260 -21068 35657 -21030
rect 35893 -21068 36290 -21030
rect 35260 -21130 35650 -21068
rect 35900 -21130 36290 -21068
rect 33660 -21230 36290 -21130
rect 33660 -21290 34050 -21230
rect 34300 -21290 34690 -21230
rect 35260 -21290 35650 -21230
rect 35900 -21290 36290 -21230
rect 32060 -21330 32457 -21290
rect 32340 -21336 32457 -21330
rect 32693 -21336 33093 -21290
rect 33657 -21336 34057 -21290
rect 34293 -21336 34693 -21290
rect 35257 -21336 35657 -21290
rect 35893 -21330 36290 -21290
rect 35893 -21336 36030 -21330
rect 32498 -21390 32544 -21384
rect 32606 -21390 32652 -21384
rect 16510 -21400 16640 -21390
rect 12800 -21810 13960 -21650
rect 14390 -21780 15560 -21640
rect 11700 -22090 11850 -22080
rect 13010 -22160 13110 -21810
rect 13640 -22160 13740 -21810
rect 14630 -22160 14700 -21780
rect 15260 -22160 15330 -21780
rect 16510 -22080 16520 -21400
rect 16630 -22080 16640 -21400
rect 16510 -22090 16640 -22080
rect 18110 -21400 18240 -21390
rect 18110 -22080 18120 -21400
rect 18230 -22080 18240 -21400
rect 18110 -22090 18240 -22080
rect 19710 -21400 19840 -21390
rect 19710 -22080 19720 -21400
rect 19830 -22080 19840 -21400
rect 19710 -22090 19840 -22080
rect 21310 -21400 21440 -21390
rect 21310 -22080 21320 -21400
rect 21430 -22080 21440 -21400
rect 21310 -22090 21440 -22080
rect 22910 -21400 23040 -21390
rect 22910 -22080 22920 -21400
rect 23030 -22080 23040 -21400
rect 22910 -22090 23040 -22080
rect 24510 -21400 24640 -21390
rect 24510 -22080 24520 -21400
rect 24630 -22080 24640 -21400
rect 24510 -22090 24640 -22080
rect 26110 -21400 26240 -21390
rect 26110 -22080 26120 -21400
rect 26230 -22080 26240 -21400
rect 26110 -22090 26240 -22080
rect 27710 -21400 27840 -21390
rect 27710 -22080 27720 -21400
rect 27830 -22080 27840 -21400
rect 27710 -22090 27840 -22080
rect 29310 -21400 29440 -21390
rect 29310 -22080 29320 -21400
rect 29430 -22080 29440 -21400
rect 29310 -22090 29440 -22080
rect 30910 -21400 31040 -21390
rect 30910 -22080 30920 -21400
rect 31030 -22080 31040 -21400
rect 30910 -22090 31040 -22080
rect 32498 -21396 32652 -21390
rect 32498 -22088 32504 -21396
rect 32510 -21400 32640 -21396
rect 32510 -22080 32520 -21400
rect 32630 -22080 32640 -21400
rect 32510 -22088 32640 -22080
rect 32646 -22088 32652 -21396
rect 32498 -22090 32652 -22088
rect 32498 -22100 32544 -22090
rect 32606 -22100 32652 -22090
rect 33134 -21396 33180 -21384
rect 33134 -22088 33140 -21396
rect 33174 -22088 33180 -21396
rect 33134 -22100 33180 -22088
rect 33570 -21396 33616 -21384
rect 33570 -22088 33576 -21396
rect 33610 -22088 33616 -21396
rect 33570 -22100 33616 -22088
rect 34098 -21390 34144 -21384
rect 34206 -21390 34252 -21384
rect 34098 -21396 34252 -21390
rect 34098 -22088 34104 -21396
rect 34110 -21400 34240 -21396
rect 34110 -22080 34120 -21400
rect 34230 -22080 34240 -21400
rect 34110 -22088 34240 -22080
rect 34246 -22088 34252 -21396
rect 34098 -22090 34252 -22088
rect 34098 -22100 34144 -22090
rect 34206 -22100 34252 -22090
rect 34734 -21396 34780 -21384
rect 34734 -22088 34740 -21396
rect 34774 -22088 34780 -21396
rect 34734 -22100 34780 -22088
rect 35170 -21396 35216 -21384
rect 35170 -22088 35176 -21396
rect 35210 -22088 35216 -21396
rect 35170 -22100 35216 -22088
rect 35698 -21390 35744 -21384
rect 35806 -21390 35852 -21384
rect 35698 -21396 35852 -21390
rect 35698 -22088 35704 -21396
rect 35710 -21400 35840 -21396
rect 35710 -22080 35720 -21400
rect 35830 -22080 35840 -21400
rect 35710 -22088 35840 -22080
rect 35846 -22088 35852 -21396
rect 35698 -22090 35852 -22088
rect 35698 -22100 35744 -22090
rect 35806 -22100 35852 -22090
rect 33200 -22140 33300 -22130
rect 33200 -22150 33210 -22140
rect 33070 -22160 33210 -22150
rect 670 -22300 31480 -22160
rect 32060 -22240 33210 -22160
rect 33290 -22240 33300 -22140
rect 32060 -22250 33300 -22240
rect 33660 -22170 36290 -22160
rect 33660 -22240 34020 -22170
rect 34360 -22240 36290 -22170
rect 33660 -22250 34000 -22240
rect 34320 -22250 36290 -22240
rect 39100 -22300 39229 -20600
rect 670 -22380 39229 -22300
rect -1349 -22390 39229 -22380
rect -1349 -22400 32490 -22390
rect -1349 -33000 -1300 -22400
rect 0 -22420 32490 -22400
rect 36180 -22400 39229 -22390
rect 36180 -22420 37940 -22400
rect 28140 -22730 28380 -22720
rect 28140 -22870 28150 -22730
rect 28370 -22870 28380 -22730
rect 28500 -22760 28540 -22420
rect 28620 -22740 28750 -22730
rect 28140 -22880 28380 -22870
rect 28620 -22870 28630 -22740
rect 28740 -22870 28750 -22740
rect 28820 -22760 28860 -22420
rect 28990 -22730 29230 -22720
rect 28620 -22880 28750 -22870
rect 28990 -22870 29000 -22730
rect 29220 -22870 29230 -22730
rect 28990 -22880 29230 -22870
rect 31890 -23240 32390 -22420
rect 32620 -22430 33310 -22420
rect 32620 -22490 32630 -22430
rect 33300 -22490 33310 -22430
rect 32620 -22500 33310 -22490
rect 34030 -22430 34320 -22420
rect 34030 -22490 34040 -22430
rect 34310 -22490 34320 -22430
rect 34030 -22500 34320 -22490
rect 32620 -23240 32660 -22840
rect 32710 -23060 32750 -22550
rect 32790 -22640 32820 -22500
rect 32870 -23060 32910 -22550
rect 32690 -23070 32920 -23060
rect 32690 -23150 32700 -23070
rect 32910 -23150 32920 -23070
rect 32690 -23160 32920 -23150
rect 32950 -23240 32980 -22970
rect 33030 -23060 33070 -22550
rect 33110 -22640 33140 -22500
rect 33180 -23060 33220 -22550
rect 33010 -23070 33240 -23060
rect 33010 -23150 33020 -23070
rect 33230 -23150 33240 -23070
rect 33010 -23160 33240 -23150
rect 33290 -23240 33330 -22630
rect 34000 -23240 34030 -22980
rect 34080 -23090 34120 -22560
rect 34160 -22770 34190 -22500
rect 34240 -23090 34280 -22560
rect 34060 -23100 34310 -23090
rect 34060 -23160 34070 -23100
rect 34300 -23160 34310 -23100
rect 34060 -23170 34310 -23160
rect 34350 -23240 34380 -22960
rect 31890 -23370 34480 -23240
rect 32300 -23460 34480 -23370
rect 29740 -23520 29890 -23510
rect 28370 -23590 29750 -23520
rect 29880 -23590 29890 -23520
rect 29740 -23600 29890 -23590
rect 32540 -24360 33040 -23460
rect 33400 -23560 33920 -23550
rect 33400 -23590 33410 -23560
rect 33170 -23620 33410 -23590
rect 33910 -23590 33920 -23560
rect 34620 -23560 37030 -23550
rect 33910 -23620 34150 -23590
rect 33170 -23630 34150 -23620
rect 34620 -23620 35000 -23560
rect 37020 -23620 37030 -23560
rect 34620 -23630 35180 -23620
rect 35210 -23630 37030 -23620
rect 33170 -23830 33200 -23630
rect 33250 -24210 33290 -23690
rect 33160 -24220 33290 -24210
rect 33160 -24280 33170 -24220
rect 33280 -24280 33290 -24220
rect 33160 -24290 33290 -24280
rect 33330 -24360 33360 -23950
rect 33410 -24210 33440 -23680
rect 33490 -23890 33520 -23630
rect 33570 -24210 33600 -23680
rect 33400 -24220 33610 -24210
rect 33400 -24280 33410 -24220
rect 33600 -24280 33610 -24220
rect 33400 -24290 33610 -24280
rect 33650 -24360 33680 -23940
rect 33730 -24210 33760 -23680
rect 33810 -23890 33840 -23630
rect 33890 -24210 33920 -23680
rect 34042 -23690 34074 -23688
rect 33720 -24220 33930 -24210
rect 33720 -24280 33730 -24220
rect 33920 -24280 33930 -24220
rect 33720 -24290 33930 -24280
rect 33960 -24360 33990 -23950
rect 34040 -24210 34080 -23690
rect 34120 -23840 34150 -23630
rect 34030 -24220 34150 -24210
rect 34030 -24280 34040 -24220
rect 34140 -24280 34150 -24220
rect 34030 -24290 34150 -24280
rect 34540 -24360 34570 -23930
rect 34620 -24210 34650 -23680
rect 34700 -23810 34730 -23630
rect 34780 -24210 34810 -23680
rect 34610 -24220 34820 -24210
rect 34610 -24280 34620 -24220
rect 34770 -24280 34820 -24220
rect 34610 -24290 34820 -24280
rect 34860 -24360 34890 -23930
rect 34940 -24210 34970 -23680
rect 35020 -23800 35050 -23630
rect 35100 -24210 35130 -23680
rect 34930 -24220 35140 -24210
rect 34930 -24280 34990 -24220
rect 35130 -24280 35140 -24220
rect 34930 -24290 35140 -24280
rect 35180 -24360 35210 -23930
rect 35250 -24210 35280 -23680
rect 35330 -23810 35360 -23630
rect 35410 -24210 35440 -23680
rect 35250 -24220 35460 -24210
rect 35250 -24280 35260 -24220
rect 35450 -24280 35460 -24220
rect 35250 -24290 35460 -24280
rect 35490 -24360 35520 -23940
rect 35570 -24210 35600 -23680
rect 35650 -23800 35680 -23630
rect 35730 -24210 35760 -23680
rect 35560 -24220 35770 -24210
rect 35560 -24280 35570 -24220
rect 35760 -24280 35770 -24220
rect 35560 -24290 35770 -24280
rect 35810 -24360 35840 -23960
rect 35890 -24210 35920 -23680
rect 35970 -23810 36000 -23630
rect 36050 -24210 36080 -23680
rect 35880 -24220 36090 -24210
rect 35880 -24280 35890 -24220
rect 36080 -24280 36090 -24220
rect 35880 -24290 36090 -24280
rect 36120 -24360 36150 -23940
rect 36200 -24210 36230 -23680
rect 36280 -23800 36310 -23630
rect 36360 -24210 36390 -23680
rect 36190 -24220 36400 -24210
rect 36190 -24280 36200 -24220
rect 36390 -24280 36400 -24220
rect 36190 -24290 36400 -24280
rect 36440 -24360 36470 -23960
rect 36520 -24210 36550 -23680
rect 36600 -23790 36630 -23630
rect 36680 -24210 36710 -23680
rect 36510 -24220 36720 -24210
rect 36510 -24280 36520 -24220
rect 36710 -24280 36720 -24220
rect 36510 -24290 36720 -24280
rect 36750 -24360 36780 -23930
rect 36830 -24210 36860 -23680
rect 36910 -23800 36940 -23630
rect 36990 -24210 37020 -23680
rect 36820 -24220 37030 -24210
rect 36820 -24280 36830 -24220
rect 37020 -24280 37030 -24220
rect 36820 -24290 37030 -24280
rect 37070 -24360 37100 -23940
rect 27940 -24520 29990 -24390
rect 32540 -24410 37260 -24360
rect 32980 -24420 37260 -24410
rect 27870 -24680 28760 -24630
rect 23030 -24690 23570 -24680
rect 2500 -25070 4020 -25060
rect 2500 -25130 2510 -25070
rect 4010 -25130 4020 -25070
rect 2500 -25142 4020 -25130
rect 4700 -25070 6220 -25060
rect 4700 -25130 4710 -25070
rect 6210 -25130 6220 -25070
rect 4700 -25142 6220 -25130
rect 6900 -25070 8420 -25060
rect 6900 -25130 6910 -25070
rect 8410 -25130 8420 -25070
rect 6900 -25142 8420 -25130
rect 9100 -25070 10620 -25060
rect 9100 -25130 9110 -25070
rect 10610 -25130 10620 -25070
rect 9100 -25142 10620 -25130
rect 11300 -25070 12820 -25060
rect 11300 -25130 11310 -25070
rect 12810 -25130 12820 -25070
rect 11300 -25142 12820 -25130
rect 13500 -25070 15020 -25060
rect 13500 -25130 13510 -25070
rect 15010 -25130 15020 -25070
rect 13500 -25142 15020 -25130
rect 15700 -25070 17220 -25060
rect 15700 -25130 15710 -25070
rect 17210 -25130 17220 -25070
rect 15700 -25142 17220 -25130
rect 17900 -25070 19420 -25060
rect 17900 -25130 17910 -25070
rect 19410 -25130 19420 -25070
rect 23030 -25070 23040 -24690
rect 23560 -25070 23570 -24690
rect 23030 -25080 23570 -25070
rect 23690 -25080 24900 -24680
rect 25020 -25080 26230 -24680
rect 27870 -24720 27970 -24680
rect 27870 -24810 27960 -24720
rect 27250 -24910 27960 -24810
rect 17900 -25142 19420 -25130
rect 4100 -25230 4440 -25170
rect 4500 -25230 4510 -25170
rect 6300 -25230 6640 -25170
rect 6700 -25230 6710 -25170
rect 8500 -25230 8620 -25170
rect 8680 -25230 8910 -25170
rect 10700 -25230 10820 -25170
rect 10880 -25230 11110 -25170
rect 12900 -25230 13020 -25170
rect 13080 -25230 13310 -25170
rect 15100 -25230 15220 -25170
rect 15280 -25230 15510 -25170
rect 17300 -25230 17640 -25170
rect 17700 -25230 17710 -25170
rect 19500 -25230 19840 -25170
rect 19900 -25230 19910 -25170
rect 2010 -25320 2240 -25260
rect 2300 -25320 2420 -25260
rect 4210 -25340 4440 -25280
rect 4500 -25340 4620 -25280
rect 6410 -25340 6420 -25280
rect 6480 -25340 6820 -25280
rect 8610 -25340 8620 -25280
rect 8680 -25340 9020 -25280
rect 10810 -25340 10820 -25280
rect 10880 -25340 11220 -25280
rect 13010 -25340 13020 -25280
rect 13080 -25340 13420 -25280
rect 15210 -25340 15440 -25280
rect 15500 -25340 15620 -25280
rect 17410 -25340 17640 -25280
rect 17700 -25340 17820 -25280
rect 2500 -25700 2700 -25460
rect 2500 -25760 2510 -25700
rect 2690 -25760 2700 -25700
rect 3160 -25700 3360 -25460
rect 3160 -25760 3170 -25700
rect 3350 -25760 3360 -25700
rect 3820 -25700 4020 -25460
rect 3820 -25760 3830 -25700
rect 4010 -25760 4020 -25700
rect 4700 -25700 4900 -25460
rect 4700 -25760 4710 -25700
rect 4890 -25760 4900 -25700
rect 5360 -25700 5560 -25460
rect 5360 -25760 5370 -25700
rect 5550 -25760 5560 -25700
rect 6020 -25700 6220 -25460
rect 6020 -25760 6030 -25700
rect 6210 -25760 6220 -25700
rect 6900 -25560 7100 -25460
rect 6900 -25620 6910 -25560
rect 7090 -25620 7100 -25560
rect 6900 -25760 7100 -25620
rect 7560 -25560 7760 -25460
rect 7560 -25620 7570 -25560
rect 7750 -25620 7760 -25560
rect 7560 -25760 7760 -25620
rect 8220 -25560 8420 -25460
rect 8220 -25620 8230 -25560
rect 8410 -25620 8420 -25560
rect 8220 -25760 8420 -25620
rect 9100 -25560 9300 -25460
rect 9100 -25620 9110 -25560
rect 9290 -25620 9300 -25560
rect 9100 -25760 9300 -25620
rect 9760 -25560 9960 -25460
rect 9760 -25620 9770 -25560
rect 9950 -25620 9960 -25560
rect 9760 -25760 9960 -25620
rect 10420 -25560 10620 -25460
rect 10420 -25620 10430 -25560
rect 10610 -25620 10620 -25560
rect 10420 -25760 10620 -25620
rect 11300 -25560 11500 -25460
rect 11300 -25620 11310 -25560
rect 11490 -25620 11500 -25560
rect 11300 -25760 11500 -25620
rect 11960 -25560 12160 -25460
rect 11960 -25620 11970 -25560
rect 12150 -25620 12160 -25560
rect 11960 -25760 12160 -25620
rect 12620 -25560 12820 -25460
rect 12620 -25620 12630 -25560
rect 12810 -25620 12820 -25560
rect 12620 -25760 12820 -25620
rect 13500 -25560 13700 -25460
rect 13500 -25620 13510 -25560
rect 13690 -25620 13700 -25560
rect 13500 -25760 13700 -25620
rect 14160 -25560 14360 -25460
rect 14160 -25620 14170 -25560
rect 14350 -25620 14360 -25560
rect 14160 -25760 14360 -25620
rect 14820 -25560 15020 -25460
rect 14820 -25620 14830 -25560
rect 15010 -25620 15020 -25560
rect 14820 -25760 15020 -25620
rect 15700 -25700 15900 -25460
rect 15700 -25760 15710 -25700
rect 15890 -25760 15900 -25700
rect 16360 -25700 16560 -25460
rect 16360 -25760 16370 -25700
rect 16550 -25760 16560 -25700
rect 17020 -25700 17220 -25460
rect 17020 -25760 17030 -25700
rect 17210 -25760 17220 -25700
rect 17900 -25700 18100 -25460
rect 17900 -25760 17910 -25700
rect 18090 -25760 18100 -25700
rect 18560 -25700 18760 -25460
rect 18560 -25760 18570 -25700
rect 18750 -25760 18760 -25700
rect 19220 -25700 19420 -25460
rect 27250 -25510 27330 -24910
rect 27870 -25110 27960 -24910
rect 28780 -25110 28940 -24720
rect 27870 -25150 27990 -25110
rect 27870 -25200 28760 -25150
rect 29790 -25300 29990 -24520
rect 34800 -24490 34940 -24480
rect 35960 -24490 36140 -24460
rect 34800 -24610 34810 -24490
rect 34930 -24610 36140 -24490
rect 34800 -24620 34940 -24610
rect 27930 -25402 29990 -25300
rect 27910 -25408 29990 -25402
rect 27910 -25442 27922 -25408
rect 27930 -25430 29990 -25408
rect 28802 -25442 28814 -25430
rect 27910 -25448 28814 -25442
rect 27250 -25600 27260 -25510
rect 27320 -25536 27330 -25510
rect 27320 -25542 28726 -25536
rect 27320 -25576 27950 -25542
rect 28714 -25576 28726 -25542
rect 27320 -25582 28726 -25576
rect 27320 -25600 27330 -25582
rect 27250 -25610 27330 -25600
rect 27730 -25670 27810 -25660
rect 27730 -25694 27740 -25670
rect 19220 -25760 19230 -25700
rect 19410 -25760 19420 -25700
rect 27260 -25740 27740 -25694
rect 27730 -25760 27740 -25740
rect 27800 -25694 27810 -25670
rect 28767 -25677 28814 -25599
rect 27800 -25700 28726 -25694
rect 27800 -25734 27950 -25700
rect 28714 -25734 28726 -25700
rect 27800 -25740 28726 -25734
rect 27800 -25760 27810 -25740
rect 28770 -25757 28810 -25677
rect 27730 -25770 27810 -25760
rect 27250 -25830 27330 -25820
rect 2500 -25870 4020 -25860
rect 2500 -25930 2510 -25870
rect 4010 -25930 4020 -25870
rect 2500 -25942 4020 -25930
rect 4700 -25870 6220 -25860
rect 4700 -25930 4710 -25870
rect 6210 -25930 6220 -25870
rect 4700 -25942 6220 -25930
rect 6900 -25870 8420 -25860
rect 6900 -25930 6910 -25870
rect 8410 -25930 8420 -25870
rect 6900 -25942 8420 -25930
rect 9100 -25870 10620 -25860
rect 9100 -25930 9110 -25870
rect 10610 -25930 10620 -25870
rect 9100 -25942 10620 -25930
rect 11300 -25870 12820 -25860
rect 11300 -25930 11310 -25870
rect 12810 -25930 12820 -25870
rect 11300 -25942 12820 -25930
rect 13500 -25870 15020 -25860
rect 13500 -25930 13510 -25870
rect 15010 -25930 15020 -25870
rect 13500 -25942 15020 -25930
rect 15700 -25870 17220 -25860
rect 15700 -25930 15710 -25870
rect 17210 -25930 17220 -25870
rect 15700 -25942 17220 -25930
rect 17900 -25870 19420 -25860
rect 17900 -25930 17910 -25870
rect 19410 -25930 19420 -25870
rect 27250 -25920 27260 -25830
rect 27320 -25852 27330 -25830
rect 28767 -25830 28814 -25757
rect 29370 -25770 29450 -25760
rect 29370 -25830 29380 -25770
rect 28767 -25835 29380 -25830
rect 27320 -25858 28726 -25852
rect 27320 -25892 27950 -25858
rect 28714 -25892 28726 -25858
rect 27320 -25898 28726 -25892
rect 27320 -25920 27330 -25898
rect 28770 -25915 29380 -25835
rect 27250 -25930 27330 -25920
rect 28767 -25920 29380 -25915
rect 17900 -25942 19420 -25930
rect 4100 -26030 4220 -25970
rect 4280 -26030 4510 -25970
rect 6300 -26030 6420 -25970
rect 6480 -26030 6710 -25970
rect 8500 -26030 8840 -25970
rect 8900 -26030 8910 -25970
rect 10700 -26030 11040 -25970
rect 11100 -26030 11110 -25970
rect 12900 -26030 13240 -25970
rect 13300 -26030 13310 -25970
rect 15100 -26030 15440 -25970
rect 15500 -26030 15510 -25970
rect 17300 -26030 17420 -25970
rect 17480 -26030 17710 -25970
rect 19500 -26030 19620 -25970
rect 19680 -26030 19910 -25970
rect 27730 -25985 27810 -25975
rect 27730 -26010 27740 -25985
rect 27260 -26056 27740 -26010
rect 2010 -26120 2020 -26060
rect 2080 -26120 2420 -26060
rect 27730 -26075 27740 -26056
rect 27800 -26010 27810 -25985
rect 28767 -25993 28814 -25920
rect 29370 -25970 29380 -25920
rect 29440 -25970 29450 -25770
rect 29370 -25980 29450 -25970
rect 27800 -26016 28726 -26010
rect 27800 -26050 27950 -26016
rect 28714 -26050 28726 -26016
rect 27800 -26056 28726 -26050
rect 27800 -26075 27810 -26056
rect 28770 -26073 28810 -25993
rect 4210 -26140 4220 -26080
rect 4280 -26140 4620 -26080
rect 6410 -26140 6640 -26080
rect 6700 -26140 6820 -26080
rect 8610 -26140 8840 -26080
rect 8900 -26140 9020 -26080
rect 10810 -26140 11040 -26080
rect 11100 -26140 11220 -26080
rect 13010 -26140 13240 -26080
rect 13300 -26140 13420 -26080
rect 15210 -26140 15220 -26080
rect 15280 -26140 15620 -26080
rect 17410 -26140 17420 -26080
rect 17480 -26140 17820 -26080
rect 27730 -26085 27810 -26075
rect 27250 -26145 27330 -26135
rect 27250 -26235 27260 -26145
rect 27320 -26168 27330 -26145
rect 28767 -26151 28814 -26073
rect 27320 -26174 28726 -26168
rect 27320 -26208 27950 -26174
rect 28714 -26208 28726 -26174
rect 27320 -26214 28726 -26208
rect 27320 -26235 27330 -26214
rect 27250 -26245 27330 -26235
rect 2500 -26360 2700 -26260
rect 2500 -26420 2510 -26360
rect 2690 -26420 2700 -26360
rect 2500 -26560 2700 -26420
rect 3160 -26360 3360 -26260
rect 3160 -26420 3170 -26360
rect 3350 -26420 3360 -26360
rect 3160 -26560 3360 -26420
rect 3820 -26360 4020 -26260
rect 3820 -26420 3830 -26360
rect 4010 -26420 4020 -26360
rect 3820 -26560 4020 -26420
rect 4700 -26360 4900 -26260
rect 4700 -26420 4710 -26360
rect 4890 -26420 4900 -26360
rect 4700 -26560 4900 -26420
rect 5360 -26360 5560 -26260
rect 5360 -26420 5370 -26360
rect 5550 -26420 5560 -26360
rect 5360 -26560 5560 -26420
rect 6020 -26360 6220 -26260
rect 6020 -26420 6030 -26360
rect 6210 -26420 6220 -26360
rect 6020 -26560 6220 -26420
rect 6900 -26500 7100 -26260
rect 6900 -26560 6910 -26500
rect 7090 -26560 7100 -26500
rect 7560 -26500 7760 -26260
rect 7560 -26560 7570 -26500
rect 7750 -26560 7760 -26500
rect 8220 -26500 8420 -26260
rect 8220 -26560 8230 -26500
rect 8410 -26560 8420 -26500
rect 9100 -26500 9300 -26260
rect 9100 -26560 9110 -26500
rect 9290 -26560 9300 -26500
rect 9760 -26500 9960 -26260
rect 9760 -26560 9770 -26500
rect 9950 -26560 9960 -26500
rect 10420 -26500 10620 -26260
rect 10420 -26560 10430 -26500
rect 10610 -26560 10620 -26500
rect 11300 -26500 11500 -26260
rect 11300 -26560 11310 -26500
rect 11490 -26560 11500 -26500
rect 11960 -26500 12160 -26260
rect 11960 -26560 11970 -26500
rect 12150 -26560 12160 -26500
rect 12620 -26500 12820 -26260
rect 12620 -26560 12630 -26500
rect 12810 -26560 12820 -26500
rect 13500 -26500 13700 -26260
rect 13500 -26560 13510 -26500
rect 13690 -26560 13700 -26500
rect 14160 -26500 14360 -26260
rect 14160 -26560 14170 -26500
rect 14350 -26560 14360 -26500
rect 14820 -26500 15020 -26260
rect 14820 -26560 14830 -26500
rect 15010 -26560 15020 -26500
rect 15700 -26360 15900 -26260
rect 15700 -26420 15710 -26360
rect 15890 -26420 15900 -26360
rect 15700 -26560 15900 -26420
rect 16360 -26360 16560 -26260
rect 16360 -26420 16370 -26360
rect 16550 -26420 16560 -26360
rect 16360 -26560 16560 -26420
rect 17020 -26360 17220 -26260
rect 17020 -26420 17030 -26360
rect 17210 -26420 17220 -26360
rect 17020 -26560 17220 -26420
rect 17900 -26360 18100 -26260
rect 17900 -26420 17910 -26360
rect 18090 -26420 18100 -26360
rect 17900 -26560 18100 -26420
rect 18560 -26360 18760 -26260
rect 18560 -26420 18570 -26360
rect 18750 -26420 18760 -26360
rect 18560 -26560 18760 -26420
rect 19220 -26360 19420 -26260
rect 27910 -26308 28814 -26302
rect 27910 -26342 27922 -26308
rect 28802 -26330 28814 -26308
rect 29790 -26330 29990 -25430
rect 27930 -26342 29990 -26330
rect 27910 -26348 29990 -26342
rect 19220 -26420 19230 -26360
rect 19410 -26420 19420 -26360
rect 19220 -26560 19420 -26420
rect 27930 -26442 29990 -26348
rect 27910 -26448 29990 -26442
rect 27910 -26482 27922 -26448
rect 27930 -26460 29990 -26448
rect 28802 -26482 28814 -26460
rect 27910 -26488 28814 -26482
rect 27730 -26550 27810 -26540
rect 27730 -26576 27740 -26550
rect 420 -26630 620 -26620
rect 420 -26710 430 -26630
rect 610 -26640 620 -26630
rect 21300 -26630 21500 -26620
rect 27260 -26622 27740 -26576
rect 21300 -26640 21310 -26630
rect 610 -26700 4040 -26640
rect 4700 -26670 6220 -26660
rect 610 -26710 620 -26700
rect 420 -26720 620 -26710
rect 4700 -26730 4710 -26670
rect 6210 -26730 6220 -26670
rect 4700 -26742 6220 -26730
rect 6900 -26670 8420 -26660
rect 6900 -26730 6910 -26670
rect 8410 -26730 8420 -26670
rect 6900 -26742 8420 -26730
rect 9100 -26670 10620 -26660
rect 9100 -26730 9110 -26670
rect 10610 -26730 10620 -26670
rect 9100 -26742 10620 -26730
rect 11300 -26670 12820 -26660
rect 11300 -26730 11310 -26670
rect 12810 -26730 12820 -26670
rect 11300 -26742 12820 -26730
rect 13500 -26670 15020 -26660
rect 13500 -26730 13510 -26670
rect 15010 -26730 15020 -26670
rect 13500 -26742 15020 -26730
rect 15700 -26670 17220 -26660
rect 15700 -26730 15710 -26670
rect 17210 -26730 17220 -26670
rect 17880 -26700 21310 -26640
rect 21300 -26710 21310 -26700
rect 21490 -26710 21500 -26630
rect 27730 -26640 27740 -26622
rect 27800 -26576 27810 -26550
rect 27800 -26582 28726 -26576
rect 27800 -26616 27950 -26582
rect 28714 -26616 28726 -26582
rect 27800 -26622 28726 -26616
rect 27800 -26640 27810 -26622
rect 27730 -26650 27810 -26640
rect 21300 -26720 21500 -26710
rect 27370 -26710 27450 -26700
rect 15700 -26742 17220 -26730
rect 27370 -26734 27380 -26710
rect 4100 -26830 4510 -26770
rect 6300 -26830 6640 -26770
rect 6700 -26830 6710 -26770
rect 8500 -26830 8620 -26770
rect 8680 -26830 8910 -26770
rect 10700 -26830 10820 -26770
rect 10880 -26830 11110 -26770
rect 12900 -26830 13020 -26770
rect 13080 -26830 13310 -26770
rect 15100 -26830 15220 -26770
rect 15280 -26830 15510 -26770
rect 17300 -26830 17640 -26770
rect 17700 -26830 17710 -26770
rect 19500 -26780 20310 -26770
rect 27260 -26780 27380 -26734
rect 19500 -26830 20240 -26780
rect 1410 -26870 2420 -26860
rect 1410 -27020 1420 -26870
rect 1480 -26920 2420 -26870
rect 1480 -27020 1490 -26920
rect 4210 -26940 4440 -26880
rect 4500 -26940 4620 -26880
rect 6410 -26940 6420 -26880
rect 6480 -26940 6820 -26880
rect 8610 -26940 8620 -26880
rect 8680 -26940 9020 -26880
rect 10810 -26940 10820 -26880
rect 10880 -26940 11220 -26880
rect 13010 -26940 13020 -26880
rect 13080 -26940 13420 -26880
rect 15210 -26940 15440 -26880
rect 15500 -26940 15620 -26880
rect 17410 -26940 17820 -26880
rect 20230 -26930 20240 -26830
rect 20300 -26930 20310 -26780
rect 27370 -26800 27380 -26780
rect 27440 -26734 27450 -26710
rect 28767 -26717 28813 -26639
rect 27440 -26740 28726 -26734
rect 27440 -26774 27950 -26740
rect 28714 -26774 28726 -26740
rect 27440 -26780 28726 -26774
rect 27440 -26800 27450 -26780
rect 28770 -26797 28810 -26717
rect 27370 -26810 27450 -26800
rect 27730 -26870 27810 -26860
rect 27730 -26892 27740 -26870
rect 20230 -26940 20310 -26930
rect 27260 -26938 27740 -26892
rect 27730 -26960 27740 -26938
rect 27800 -26892 27810 -26870
rect 28767 -26870 28813 -26797
rect 29520 -26810 29600 -26800
rect 29520 -26870 29530 -26810
rect 28767 -26875 29530 -26870
rect 27800 -26898 28726 -26892
rect 27800 -26932 27950 -26898
rect 28714 -26932 28726 -26898
rect 27800 -26938 28726 -26932
rect 27800 -26960 27810 -26938
rect 28770 -26955 29530 -26875
rect 27730 -26970 27810 -26960
rect 28767 -26960 29530 -26955
rect 1410 -27030 1490 -27020
rect 27370 -27025 27450 -27015
rect 27370 -27050 27380 -27025
rect 2500 -27300 2700 -27060
rect 2500 -27360 2510 -27300
rect 2690 -27360 2700 -27300
rect 3160 -27300 3360 -27060
rect 3160 -27360 3170 -27300
rect 3350 -27360 3360 -27300
rect 3820 -27300 4020 -27060
rect 3820 -27360 3830 -27300
rect 4010 -27360 4020 -27300
rect 4700 -27300 4900 -27060
rect 4700 -27360 4710 -27300
rect 4890 -27360 4900 -27300
rect 5360 -27300 5560 -27060
rect 5360 -27360 5370 -27300
rect 5550 -27360 5560 -27300
rect 6020 -27300 6220 -27060
rect 6020 -27360 6030 -27300
rect 6210 -27360 6220 -27300
rect 6900 -27160 7100 -27060
rect 6900 -27220 6910 -27160
rect 7090 -27220 7100 -27160
rect 6900 -27360 7100 -27220
rect 7560 -27160 7760 -27060
rect 7560 -27220 7570 -27160
rect 7750 -27220 7760 -27160
rect 7560 -27360 7760 -27220
rect 8220 -27160 8420 -27060
rect 8220 -27220 8230 -27160
rect 8410 -27220 8420 -27160
rect 8220 -27360 8420 -27220
rect 9100 -27160 9300 -27060
rect 9100 -27220 9110 -27160
rect 9290 -27220 9300 -27160
rect 9100 -27360 9300 -27220
rect 9760 -27160 9960 -27060
rect 9760 -27220 9770 -27160
rect 9950 -27220 9960 -27160
rect 9760 -27360 9960 -27220
rect 10420 -27160 10620 -27060
rect 10420 -27220 10430 -27160
rect 10610 -27220 10620 -27160
rect 10420 -27360 10620 -27220
rect 11300 -27160 11500 -27060
rect 11300 -27220 11310 -27160
rect 11490 -27220 11500 -27160
rect 11300 -27360 11500 -27220
rect 11960 -27160 12160 -27060
rect 11960 -27220 11970 -27160
rect 12150 -27220 12160 -27160
rect 11960 -27360 12160 -27220
rect 12620 -27160 12820 -27060
rect 12620 -27220 12630 -27160
rect 12810 -27220 12820 -27160
rect 12620 -27360 12820 -27220
rect 13500 -27160 13700 -27060
rect 13500 -27220 13510 -27160
rect 13690 -27220 13700 -27160
rect 13500 -27360 13700 -27220
rect 14160 -27160 14360 -27060
rect 14160 -27220 14170 -27160
rect 14350 -27220 14360 -27160
rect 14160 -27360 14360 -27220
rect 14820 -27160 15020 -27060
rect 14820 -27220 14830 -27160
rect 15010 -27220 15020 -27160
rect 14820 -27360 15020 -27220
rect 15700 -27300 15900 -27060
rect 15700 -27360 15710 -27300
rect 15890 -27360 15900 -27300
rect 16360 -27300 16560 -27060
rect 16360 -27360 16370 -27300
rect 16550 -27360 16560 -27300
rect 17020 -27300 17220 -27060
rect 17020 -27360 17030 -27300
rect 17210 -27360 17220 -27300
rect 17900 -27300 18100 -27060
rect 17900 -27360 17910 -27300
rect 18090 -27360 18100 -27300
rect 18560 -27300 18760 -27060
rect 18560 -27360 18570 -27300
rect 18750 -27360 18760 -27300
rect 19220 -27300 19420 -27060
rect 27260 -27096 27380 -27050
rect 27370 -27115 27380 -27096
rect 27440 -27050 27450 -27025
rect 28767 -27033 28813 -26960
rect 29520 -27010 29530 -26960
rect 29590 -27010 29600 -26810
rect 29520 -27020 29600 -27010
rect 27440 -27056 28726 -27050
rect 27440 -27090 27950 -27056
rect 28714 -27090 28726 -27056
rect 27440 -27096 28726 -27090
rect 27440 -27115 27450 -27096
rect 28770 -27113 28810 -27033
rect 27370 -27125 27450 -27115
rect 27730 -27185 27810 -27175
rect 27730 -27208 27740 -27185
rect 27260 -27254 27740 -27208
rect 27730 -27275 27740 -27254
rect 27800 -27208 27810 -27185
rect 28767 -27191 28813 -27113
rect 27800 -27214 28726 -27208
rect 27800 -27248 27950 -27214
rect 28714 -27248 28726 -27214
rect 27800 -27254 28726 -27248
rect 27800 -27275 27810 -27254
rect 27730 -27285 27810 -27275
rect 19220 -27360 19230 -27300
rect 19410 -27360 19420 -27300
rect 27910 -27348 28814 -27342
rect 27910 -27382 27922 -27348
rect 28802 -27370 28814 -27348
rect 29790 -27370 29990 -26460
rect 34630 -24830 34730 -24700
rect 34630 -24860 35000 -24830
rect 34630 -25350 34730 -24860
rect 34800 -24940 35850 -24930
rect 34800 -25010 34810 -24940
rect 34900 -25010 35850 -24940
rect 34800 -25020 35850 -25010
rect 34800 -25190 34900 -25020
rect 35960 -25090 36140 -24610
rect 37330 -24830 37430 -24710
rect 37070 -24860 37430 -24830
rect 36250 -24940 37290 -24930
rect 36250 -25010 37190 -24940
rect 37280 -25010 37290 -24940
rect 36250 -25020 37290 -25010
rect 35740 -25120 36370 -25090
rect 34800 -25200 35850 -25190
rect 34800 -25270 34810 -25200
rect 34900 -25270 35850 -25200
rect 34800 -25280 35850 -25270
rect 34630 -25380 35030 -25350
rect 34630 -25860 34730 -25380
rect 34800 -25460 35850 -25450
rect 34800 -25530 34810 -25460
rect 34900 -25530 35850 -25460
rect 34800 -25540 35850 -25530
rect 34800 -25710 34900 -25540
rect 35960 -25610 36140 -25120
rect 37180 -25190 37290 -25020
rect 36250 -25200 37290 -25190
rect 36250 -25270 37190 -25200
rect 37280 -25270 37290 -25200
rect 36250 -25280 37290 -25270
rect 37330 -25350 37430 -24860
rect 37070 -25380 37430 -25350
rect 36250 -25460 37290 -25450
rect 36250 -25530 37190 -25460
rect 37280 -25530 37290 -25460
rect 36250 -25540 37290 -25530
rect 35740 -25640 36370 -25610
rect 34800 -25720 35850 -25710
rect 34800 -25790 34810 -25720
rect 34900 -25790 35850 -25720
rect 34800 -25800 35850 -25790
rect 34630 -25890 35020 -25860
rect 34630 -26380 34730 -25890
rect 34800 -25980 35850 -25970
rect 34800 -26050 34810 -25980
rect 34900 -26050 35850 -25980
rect 34800 -26060 35850 -26050
rect 34800 -26230 34900 -26060
rect 35960 -26120 36140 -25640
rect 37180 -25710 37290 -25540
rect 36250 -25720 37290 -25710
rect 36250 -25790 37190 -25720
rect 37280 -25790 37290 -25720
rect 36250 -25800 37290 -25790
rect 37330 -25860 37430 -25380
rect 37080 -25890 37430 -25860
rect 36250 -25980 37290 -25970
rect 36250 -26050 37190 -25980
rect 37280 -26050 37290 -25980
rect 36250 -26060 37290 -26050
rect 35740 -26150 36370 -26120
rect 34800 -26240 35850 -26230
rect 34800 -26310 34810 -26240
rect 34900 -26310 35850 -26240
rect 34800 -26320 35850 -26310
rect 34630 -26410 35030 -26380
rect 34630 -26900 34730 -26410
rect 34800 -26500 35850 -26490
rect 34800 -26570 34810 -26500
rect 34900 -26570 35850 -26500
rect 34800 -26580 35850 -26570
rect 34800 -26750 34900 -26580
rect 35960 -26640 36140 -26150
rect 37180 -26230 37290 -26060
rect 36250 -26240 37290 -26230
rect 36250 -26310 37190 -26240
rect 37280 -26310 37290 -26240
rect 36250 -26320 37290 -26310
rect 37330 -26380 37430 -25890
rect 37090 -26410 37430 -26380
rect 36250 -26500 37290 -26490
rect 36250 -26570 37190 -26500
rect 37280 -26570 37290 -26500
rect 36250 -26580 37290 -26570
rect 35740 -26670 36370 -26640
rect 34800 -26760 35850 -26750
rect 34800 -26830 34810 -26760
rect 34900 -26830 35850 -26760
rect 34800 -26840 35850 -26830
rect 34630 -26930 35020 -26900
rect 35960 -26910 36140 -26670
rect 37180 -26750 37290 -26580
rect 36250 -26760 37290 -26750
rect 36250 -26830 37190 -26760
rect 37280 -26830 37290 -26760
rect 36250 -26840 37290 -26830
rect 37330 -26900 37430 -26410
rect 37080 -26930 37430 -26900
rect 34630 -27020 34730 -26930
rect 36020 -27010 36420 -27000
rect 36020 -27020 36030 -27010
rect 34630 -27130 36030 -27020
rect 36020 -27140 36030 -27130
rect 36410 -27140 36420 -27010
rect 36020 -27150 36420 -27140
rect 36520 -27010 36920 -27000
rect 36520 -27140 36530 -27010
rect 36910 -27020 36920 -27010
rect 37330 -27020 37430 -26930
rect 36910 -27130 37430 -27020
rect 36910 -27140 36920 -27130
rect 36520 -27150 36920 -27140
rect 27930 -27382 29990 -27370
rect 27910 -27388 29990 -27382
rect 420 -27430 620 -27420
rect 420 -27510 430 -27430
rect 610 -27440 620 -27430
rect 21300 -27430 21500 -27420
rect 21300 -27440 21310 -27430
rect 610 -27500 4040 -27440
rect 4700 -27470 6220 -27460
rect 610 -27510 620 -27500
rect 420 -27520 620 -27510
rect 4700 -27530 4710 -27470
rect 6210 -27530 6220 -27470
rect 4700 -27542 6220 -27530
rect 6900 -27470 8420 -27460
rect 6900 -27530 6910 -27470
rect 8410 -27530 8420 -27470
rect 6900 -27542 8420 -27530
rect 9100 -27470 10620 -27460
rect 9100 -27530 9110 -27470
rect 10610 -27530 10620 -27470
rect 9100 -27542 10620 -27530
rect 11300 -27470 12820 -27460
rect 11300 -27530 11310 -27470
rect 12810 -27530 12820 -27470
rect 11300 -27542 12820 -27530
rect 13500 -27470 15020 -27460
rect 13500 -27530 13510 -27470
rect 15010 -27530 15020 -27470
rect 13500 -27542 15020 -27530
rect 15700 -27470 17220 -27460
rect 15700 -27530 15710 -27470
rect 17210 -27530 17220 -27470
rect 17880 -27500 21310 -27440
rect 21300 -27510 21310 -27500
rect 21490 -27510 21500 -27430
rect 27930 -27482 29990 -27388
rect 21300 -27520 21500 -27510
rect 27910 -27488 29990 -27482
rect 27910 -27522 27922 -27488
rect 27930 -27500 29990 -27488
rect 28802 -27522 28814 -27500
rect 27910 -27528 28814 -27522
rect 29790 -27520 29990 -27500
rect 15700 -27542 17220 -27530
rect 29790 -27540 37700 -27520
rect 4100 -27630 4510 -27570
rect 6300 -27630 6420 -27570
rect 6480 -27630 6710 -27570
rect 8500 -27630 8840 -27570
rect 8900 -27630 8910 -27570
rect 10700 -27630 11040 -27570
rect 11100 -27630 11110 -27570
rect 12900 -27630 13240 -27570
rect 13300 -27630 13310 -27570
rect 15100 -27630 15440 -27570
rect 15500 -27630 15510 -27570
rect 17300 -27630 17420 -27570
rect 17480 -27630 17710 -27570
rect 19500 -27580 20510 -27570
rect 19500 -27630 20440 -27580
rect 1610 -27670 2420 -27660
rect 1610 -27820 1620 -27670
rect 1680 -27720 2420 -27670
rect 1680 -27820 1690 -27720
rect 4210 -27740 4220 -27680
rect 4280 -27740 4620 -27680
rect 6410 -27740 6640 -27680
rect 6700 -27740 6820 -27680
rect 8610 -27740 8840 -27680
rect 8900 -27740 9020 -27680
rect 10810 -27740 11040 -27680
rect 11100 -27740 11220 -27680
rect 13010 -27740 13240 -27680
rect 13300 -27740 13420 -27680
rect 15210 -27740 15220 -27680
rect 15280 -27740 15620 -27680
rect 17410 -27740 17820 -27680
rect 20430 -27730 20440 -27630
rect 20500 -27730 20510 -27580
rect 27250 -27595 27330 -27585
rect 27250 -27685 27260 -27595
rect 27320 -27616 27330 -27595
rect 27320 -27622 28726 -27616
rect 27320 -27656 27950 -27622
rect 28714 -27656 28726 -27622
rect 27320 -27662 28726 -27656
rect 27320 -27685 27330 -27662
rect 27250 -27695 27330 -27685
rect 20430 -27740 20510 -27730
rect 27490 -27750 27570 -27740
rect 27490 -27774 27500 -27750
rect 27260 -27820 27500 -27774
rect 1610 -27830 1690 -27820
rect 27490 -27840 27500 -27820
rect 27560 -27774 27570 -27750
rect 28767 -27757 28813 -27679
rect 27560 -27780 28726 -27774
rect 27560 -27814 27950 -27780
rect 28714 -27814 28726 -27780
rect 27560 -27820 28726 -27814
rect 27560 -27840 27570 -27820
rect 28770 -27837 28810 -27757
rect 27490 -27850 27570 -27840
rect 2500 -27960 2700 -27860
rect 2500 -28020 2510 -27960
rect 2690 -28020 2700 -27960
rect 2500 -28160 2700 -28020
rect 3160 -27960 3360 -27860
rect 3160 -28020 3170 -27960
rect 3350 -28020 3360 -27960
rect 3160 -28160 3360 -28020
rect 3820 -27960 4020 -27860
rect 3820 -28020 3830 -27960
rect 4010 -28020 4020 -27960
rect 3820 -28160 4020 -28020
rect 4700 -27960 4900 -27860
rect 4700 -28020 4710 -27960
rect 4890 -28020 4900 -27960
rect 4700 -28160 4900 -28020
rect 5360 -27960 5560 -27860
rect 5360 -28020 5370 -27960
rect 5550 -28020 5560 -27960
rect 5360 -28160 5560 -28020
rect 6020 -27960 6220 -27860
rect 6020 -28020 6030 -27960
rect 6210 -28020 6220 -27960
rect 6020 -28160 6220 -28020
rect 6900 -28100 7100 -27860
rect 6900 -28160 6910 -28100
rect 7090 -28160 7100 -28100
rect 7560 -28100 7760 -27860
rect 7560 -28160 7570 -28100
rect 7750 -28160 7760 -28100
rect 8220 -28100 8420 -27860
rect 8220 -28160 8230 -28100
rect 8410 -28160 8420 -28100
rect 9100 -28100 9300 -27860
rect 9100 -28160 9110 -28100
rect 9290 -28160 9300 -28100
rect 9760 -28100 9960 -27860
rect 9760 -28160 9770 -28100
rect 9950 -28160 9960 -28100
rect 10420 -28100 10620 -27860
rect 10420 -28160 10430 -28100
rect 10610 -28160 10620 -28100
rect 11300 -28100 11500 -27860
rect 11300 -28160 11310 -28100
rect 11490 -28160 11500 -28100
rect 11960 -28100 12160 -27860
rect 11960 -28160 11970 -28100
rect 12150 -28160 12160 -28100
rect 12620 -28100 12820 -27860
rect 12620 -28160 12630 -28100
rect 12810 -28160 12820 -28100
rect 13500 -28100 13700 -27860
rect 13500 -28160 13510 -28100
rect 13690 -28160 13700 -28100
rect 14160 -28100 14360 -27860
rect 14160 -28160 14170 -28100
rect 14350 -28160 14360 -28100
rect 14820 -28100 15020 -27860
rect 14820 -28160 14830 -28100
rect 15010 -28160 15020 -28100
rect 15700 -27960 15900 -27860
rect 15700 -28020 15710 -27960
rect 15890 -28020 15900 -27960
rect 15700 -28160 15900 -28020
rect 16360 -27960 16560 -27860
rect 16360 -28020 16370 -27960
rect 16550 -28020 16560 -27960
rect 16360 -28160 16560 -28020
rect 17020 -27960 17220 -27860
rect 17020 -28020 17030 -27960
rect 17210 -28020 17220 -27960
rect 17020 -28160 17220 -28020
rect 17900 -27960 18100 -27860
rect 17900 -28020 17910 -27960
rect 18090 -28020 18100 -27960
rect 17900 -28160 18100 -28020
rect 18560 -27960 18760 -27860
rect 18560 -28020 18570 -27960
rect 18750 -28020 18760 -27960
rect 18560 -28160 18760 -28020
rect 19220 -27960 19420 -27860
rect 19220 -28020 19230 -27960
rect 19410 -28020 19420 -27960
rect 27250 -27910 27330 -27900
rect 27250 -28000 27260 -27910
rect 27320 -27932 27330 -27910
rect 28767 -27910 28813 -27837
rect 29070 -27850 29150 -27840
rect 29070 -27910 29080 -27850
rect 28767 -27915 29080 -27910
rect 27320 -27938 28726 -27932
rect 27320 -27972 27950 -27938
rect 28714 -27972 28726 -27938
rect 27320 -27978 28726 -27972
rect 27320 -28000 27330 -27978
rect 28770 -27995 29080 -27915
rect 27250 -28010 27330 -28000
rect 28767 -28000 29080 -27995
rect 19220 -28160 19420 -28020
rect 27490 -28065 27570 -28055
rect 27490 -28090 27500 -28065
rect 27260 -28136 27500 -28090
rect 27490 -28155 27500 -28136
rect 27560 -28090 27570 -28065
rect 28767 -28073 28813 -28000
rect 29070 -28050 29080 -28000
rect 29140 -28050 29150 -27850
rect 29070 -28060 29150 -28050
rect 29790 -27900 36920 -27540
rect 37680 -27900 37700 -27540
rect 29790 -27920 37700 -27900
rect 27560 -28096 28726 -28090
rect 27560 -28130 27950 -28096
rect 28714 -28130 28726 -28096
rect 27560 -28136 28726 -28130
rect 27560 -28155 27570 -28136
rect 28770 -28153 28810 -28073
rect 27490 -28165 27570 -28155
rect 420 -28230 620 -28220
rect 420 -28310 430 -28230
rect 610 -28240 620 -28230
rect 21300 -28230 21500 -28220
rect 21300 -28240 21310 -28230
rect 610 -28300 4040 -28240
rect 4700 -28270 6220 -28260
rect 610 -28310 620 -28300
rect 420 -28320 620 -28310
rect 4700 -28330 4710 -28270
rect 6210 -28330 6220 -28270
rect 4700 -28342 6220 -28330
rect 6900 -28270 8420 -28260
rect 6900 -28330 6910 -28270
rect 8410 -28330 8420 -28270
rect 6900 -28342 8420 -28330
rect 9100 -28270 10620 -28260
rect 9100 -28330 9110 -28270
rect 10610 -28330 10620 -28270
rect 9100 -28342 10620 -28330
rect 11300 -28270 12820 -28260
rect 11300 -28330 11310 -28270
rect 12810 -28330 12820 -28270
rect 11300 -28342 12820 -28330
rect 13500 -28270 15020 -28260
rect 13500 -28330 13510 -28270
rect 15010 -28330 15020 -28270
rect 13500 -28342 15020 -28330
rect 15700 -28270 17220 -28260
rect 15700 -28330 15710 -28270
rect 17210 -28330 17220 -28270
rect 17880 -28300 21310 -28240
rect 21300 -28310 21310 -28300
rect 21490 -28310 21500 -28230
rect 21300 -28320 21500 -28310
rect 27250 -28225 27330 -28215
rect 27250 -28315 27260 -28225
rect 27320 -28248 27330 -28225
rect 28767 -28231 28813 -28153
rect 27320 -28254 28726 -28248
rect 27320 -28288 27950 -28254
rect 28714 -28288 28726 -28254
rect 27320 -28294 28726 -28288
rect 27320 -28315 27330 -28294
rect 27250 -28325 27330 -28315
rect 15700 -28342 17220 -28330
rect 4100 -28430 4510 -28370
rect 6300 -28430 6420 -28370
rect 6480 -28430 6710 -28370
rect 8500 -28430 8840 -28370
rect 8900 -28430 8910 -28370
rect 10700 -28430 11040 -28370
rect 11100 -28430 11110 -28370
rect 12900 -28430 13240 -28370
rect 13300 -28430 13310 -28370
rect 15100 -28430 15440 -28370
rect 15500 -28430 15510 -28370
rect 17300 -28430 17420 -28370
rect 17480 -28430 17710 -28370
rect 19500 -28380 20510 -28370
rect 19500 -28430 20440 -28380
rect 1610 -28470 2420 -28460
rect 1610 -28620 1620 -28470
rect 1680 -28520 2420 -28470
rect 1680 -28620 1690 -28520
rect 4210 -28540 4220 -28480
rect 4280 -28540 4620 -28480
rect 6410 -28540 6640 -28480
rect 6700 -28540 6820 -28480
rect 8610 -28540 8840 -28480
rect 8900 -28540 9020 -28480
rect 10810 -28540 11040 -28480
rect 11100 -28540 11220 -28480
rect 13010 -28540 13240 -28480
rect 13300 -28540 13420 -28480
rect 15210 -28540 15220 -28480
rect 15280 -28540 15620 -28480
rect 17410 -28540 17820 -28480
rect 20430 -28530 20440 -28430
rect 20500 -28530 20510 -28380
rect 27910 -28388 28814 -28382
rect 27910 -28422 27922 -28388
rect 28802 -28410 28814 -28388
rect 29790 -28410 29990 -27920
rect 39100 -28140 39229 -22400
rect 27930 -28422 29990 -28410
rect 27910 -28428 29990 -28422
rect 27930 -28522 29990 -28428
rect 20430 -28540 20510 -28530
rect 27910 -28528 29990 -28522
rect 27910 -28562 27922 -28528
rect 27930 -28540 29990 -28528
rect 36900 -28160 39229 -28140
rect 36900 -28520 36920 -28160
rect 37680 -28520 39229 -28160
rect 36900 -28540 39229 -28520
rect 28802 -28562 28814 -28540
rect 27910 -28568 28814 -28562
rect 1610 -28630 1690 -28620
rect 27250 -28630 27330 -28620
rect 2500 -28760 2700 -28660
rect 2500 -28820 2510 -28760
rect 2690 -28820 2700 -28760
rect 2500 -28960 2700 -28820
rect 3160 -28760 3360 -28660
rect 3160 -28820 3170 -28760
rect 3350 -28820 3360 -28760
rect 3160 -28960 3360 -28820
rect 3820 -28760 4020 -28660
rect 3820 -28820 3830 -28760
rect 4010 -28820 4020 -28760
rect 3820 -28960 4020 -28820
rect 4700 -28760 4900 -28660
rect 4700 -28820 4710 -28760
rect 4890 -28820 4900 -28760
rect 4700 -28960 4900 -28820
rect 5360 -28760 5560 -28660
rect 5360 -28820 5370 -28760
rect 5550 -28820 5560 -28760
rect 5360 -28960 5560 -28820
rect 6020 -28760 6220 -28660
rect 6020 -28820 6030 -28760
rect 6210 -28820 6220 -28760
rect 6020 -28960 6220 -28820
rect 6900 -28900 7100 -28660
rect 6900 -28960 6910 -28900
rect 7090 -28960 7100 -28900
rect 7560 -28900 7760 -28660
rect 7560 -28960 7570 -28900
rect 7750 -28960 7760 -28900
rect 8220 -28900 8420 -28660
rect 8220 -28960 8230 -28900
rect 8410 -28960 8420 -28900
rect 9100 -28900 9300 -28660
rect 9100 -28960 9110 -28900
rect 9290 -28960 9300 -28900
rect 9760 -28900 9960 -28660
rect 9760 -28960 9770 -28900
rect 9950 -28960 9960 -28900
rect 10420 -28900 10620 -28660
rect 10420 -28960 10430 -28900
rect 10610 -28960 10620 -28900
rect 11300 -28900 11500 -28660
rect 11300 -28960 11310 -28900
rect 11490 -28960 11500 -28900
rect 11960 -28900 12160 -28660
rect 11960 -28960 11970 -28900
rect 12150 -28960 12160 -28900
rect 12620 -28900 12820 -28660
rect 12620 -28960 12630 -28900
rect 12810 -28960 12820 -28900
rect 13500 -28900 13700 -28660
rect 13500 -28960 13510 -28900
rect 13690 -28960 13700 -28900
rect 14160 -28900 14360 -28660
rect 14160 -28960 14170 -28900
rect 14350 -28960 14360 -28900
rect 14820 -28900 15020 -28660
rect 14820 -28960 14830 -28900
rect 15010 -28960 15020 -28900
rect 15700 -28760 15900 -28660
rect 15700 -28820 15710 -28760
rect 15890 -28820 15900 -28760
rect 15700 -28960 15900 -28820
rect 16360 -28760 16560 -28660
rect 16360 -28820 16370 -28760
rect 16550 -28820 16560 -28760
rect 16360 -28960 16560 -28820
rect 17020 -28760 17220 -28660
rect 17020 -28820 17030 -28760
rect 17210 -28820 17220 -28760
rect 17020 -28960 17220 -28820
rect 17900 -28760 18100 -28660
rect 17900 -28820 17910 -28760
rect 18090 -28820 18100 -28760
rect 17900 -28960 18100 -28820
rect 18560 -28760 18760 -28660
rect 18560 -28820 18570 -28760
rect 18750 -28820 18760 -28760
rect 18560 -28960 18760 -28820
rect 19220 -28760 19420 -28660
rect 27250 -28720 27260 -28630
rect 27320 -28656 27330 -28630
rect 27320 -28662 28726 -28656
rect 27320 -28696 27950 -28662
rect 28714 -28696 28726 -28662
rect 27320 -28702 28726 -28696
rect 27320 -28720 27330 -28702
rect 27250 -28730 27330 -28720
rect 19220 -28820 19230 -28760
rect 19410 -28820 19420 -28760
rect 27610 -28790 27690 -28780
rect 27610 -28814 27620 -28790
rect 19220 -28960 19420 -28820
rect 27260 -28860 27620 -28814
rect 27610 -28880 27620 -28860
rect 27680 -28814 27690 -28790
rect 28767 -28797 28813 -28719
rect 27680 -28820 28726 -28814
rect 27680 -28854 27950 -28820
rect 28714 -28854 28726 -28820
rect 27680 -28860 28726 -28854
rect 27680 -28880 27690 -28860
rect 28770 -28877 28810 -28797
rect 27610 -28890 27690 -28880
rect 27250 -28950 27330 -28940
rect 420 -29030 620 -29020
rect 420 -29110 430 -29030
rect 610 -29040 620 -29030
rect 21300 -29030 21500 -29020
rect 21300 -29040 21310 -29030
rect 610 -29100 4040 -29040
rect 4700 -29070 6220 -29060
rect 610 -29110 620 -29100
rect 420 -29120 620 -29110
rect 4700 -29130 4710 -29070
rect 6210 -29130 6220 -29070
rect 4700 -29142 6220 -29130
rect 6900 -29070 8420 -29060
rect 6900 -29130 6910 -29070
rect 8410 -29130 8420 -29070
rect 6900 -29142 8420 -29130
rect 9100 -29070 10620 -29060
rect 9100 -29130 9110 -29070
rect 10610 -29130 10620 -29070
rect 9100 -29142 10620 -29130
rect 11300 -29070 12820 -29060
rect 11300 -29130 11310 -29070
rect 12810 -29130 12820 -29070
rect 11300 -29142 12820 -29130
rect 13500 -29070 15020 -29060
rect 13500 -29130 13510 -29070
rect 15010 -29130 15020 -29070
rect 13500 -29142 15020 -29130
rect 15700 -29070 17220 -29060
rect 15700 -29130 15710 -29070
rect 17210 -29130 17220 -29070
rect 17880 -29100 21310 -29040
rect 21300 -29110 21310 -29100
rect 21490 -29110 21500 -29030
rect 27250 -29040 27260 -28950
rect 27320 -28972 27330 -28950
rect 28767 -28950 28813 -28877
rect 29220 -28890 29300 -28880
rect 29220 -28950 29230 -28890
rect 28767 -28955 29230 -28950
rect 27320 -28978 28726 -28972
rect 27320 -29012 27950 -28978
rect 28714 -29012 28726 -28978
rect 27320 -29018 28726 -29012
rect 27320 -29040 27330 -29018
rect 28770 -29035 29230 -28955
rect 27250 -29050 27330 -29040
rect 28767 -29040 29230 -29035
rect 21300 -29120 21500 -29110
rect 27610 -29110 27690 -29100
rect 27610 -29130 27620 -29110
rect 15700 -29142 17220 -29130
rect 4100 -29230 4510 -29170
rect 6300 -29230 6640 -29170
rect 6700 -29230 6710 -29170
rect 8500 -29230 8620 -29170
rect 8680 -29230 8910 -29170
rect 10700 -29230 10820 -29170
rect 10880 -29230 11110 -29170
rect 12900 -29230 13020 -29170
rect 13080 -29230 13310 -29170
rect 15100 -29230 15220 -29170
rect 15280 -29230 15510 -29170
rect 17300 -29230 17640 -29170
rect 17700 -29230 17710 -29170
rect 19500 -29180 20310 -29170
rect 27260 -29176 27620 -29130
rect 19500 -29230 20240 -29180
rect 1410 -29270 2420 -29260
rect 1410 -29420 1420 -29270
rect 1480 -29320 2420 -29270
rect 1480 -29420 1490 -29320
rect 4210 -29340 4440 -29280
rect 4500 -29340 4620 -29280
rect 6410 -29340 6420 -29280
rect 6480 -29340 6820 -29280
rect 8610 -29340 8620 -29280
rect 8680 -29340 9020 -29280
rect 10810 -29340 10820 -29280
rect 10880 -29340 11220 -29280
rect 13010 -29340 13020 -29280
rect 13080 -29340 13420 -29280
rect 15210 -29340 15440 -29280
rect 15500 -29340 15620 -29280
rect 17410 -29340 17820 -29280
rect 20230 -29330 20240 -29230
rect 20300 -29330 20310 -29180
rect 27610 -29200 27620 -29176
rect 27680 -29130 27690 -29110
rect 28767 -29113 28813 -29040
rect 29220 -29090 29230 -29040
rect 29290 -29090 29300 -28890
rect 29220 -29100 29300 -29090
rect 27680 -29136 28726 -29130
rect 27680 -29170 27950 -29136
rect 28714 -29170 28726 -29136
rect 27680 -29176 28726 -29170
rect 27680 -29200 27690 -29176
rect 28770 -29193 28810 -29113
rect 27610 -29210 27690 -29200
rect 20230 -29340 20310 -29330
rect 27250 -29260 27330 -29250
rect 27250 -29350 27260 -29260
rect 27320 -29288 27330 -29260
rect 28767 -29271 28813 -29193
rect 27320 -29294 28726 -29288
rect 27320 -29328 27950 -29294
rect 28714 -29328 28726 -29294
rect 27320 -29334 28726 -29328
rect 27320 -29350 27330 -29334
rect 27250 -29360 27330 -29350
rect 1410 -29430 1490 -29420
rect 27910 -29428 28814 -29422
rect 27910 -29450 27922 -29428
rect 28802 -29450 28814 -29428
rect 29790 -29450 29990 -28540
rect 37220 -29060 37420 -28540
rect 32620 -29360 38320 -29060
rect 2500 -29700 2700 -29460
rect 2500 -29760 2510 -29700
rect 2690 -29760 2700 -29700
rect 3160 -29700 3360 -29460
rect 3160 -29760 3170 -29700
rect 3350 -29760 3360 -29700
rect 3820 -29700 4020 -29460
rect 3820 -29760 3830 -29700
rect 4010 -29760 4020 -29700
rect 4700 -29700 4900 -29460
rect 4700 -29760 4710 -29700
rect 4890 -29760 4900 -29700
rect 5360 -29700 5560 -29460
rect 5360 -29760 5370 -29700
rect 5550 -29760 5560 -29700
rect 6020 -29700 6220 -29460
rect 6020 -29760 6030 -29700
rect 6210 -29760 6220 -29700
rect 6900 -29560 7100 -29460
rect 6900 -29620 6910 -29560
rect 7090 -29620 7100 -29560
rect 6900 -29760 7100 -29620
rect 7560 -29560 7760 -29460
rect 7560 -29620 7570 -29560
rect 7750 -29620 7760 -29560
rect 7560 -29760 7760 -29620
rect 8220 -29560 8420 -29460
rect 8220 -29620 8230 -29560
rect 8410 -29620 8420 -29560
rect 8220 -29760 8420 -29620
rect 9100 -29560 9300 -29460
rect 9100 -29620 9110 -29560
rect 9290 -29620 9300 -29560
rect 9100 -29760 9300 -29620
rect 9760 -29560 9960 -29460
rect 9760 -29620 9770 -29560
rect 9950 -29620 9960 -29560
rect 9760 -29760 9960 -29620
rect 10420 -29560 10620 -29460
rect 10420 -29620 10430 -29560
rect 10610 -29620 10620 -29560
rect 10420 -29760 10620 -29620
rect 11300 -29560 11500 -29460
rect 11300 -29620 11310 -29560
rect 11490 -29620 11500 -29560
rect 11300 -29760 11500 -29620
rect 11960 -29560 12160 -29460
rect 11960 -29620 11970 -29560
rect 12150 -29620 12160 -29560
rect 11960 -29760 12160 -29620
rect 12620 -29560 12820 -29460
rect 12620 -29620 12630 -29560
rect 12810 -29620 12820 -29560
rect 12620 -29760 12820 -29620
rect 13500 -29560 13700 -29460
rect 13500 -29620 13510 -29560
rect 13690 -29620 13700 -29560
rect 13500 -29760 13700 -29620
rect 14160 -29560 14360 -29460
rect 14160 -29620 14170 -29560
rect 14350 -29620 14360 -29560
rect 14160 -29760 14360 -29620
rect 14820 -29560 15020 -29460
rect 14820 -29620 14830 -29560
rect 15010 -29620 15020 -29560
rect 14820 -29760 15020 -29620
rect 15700 -29700 15900 -29460
rect 15700 -29760 15710 -29700
rect 15890 -29760 15900 -29700
rect 16360 -29700 16560 -29460
rect 16360 -29760 16370 -29700
rect 16550 -29760 16560 -29700
rect 17020 -29700 17220 -29460
rect 17020 -29760 17030 -29700
rect 17210 -29760 17220 -29700
rect 17900 -29700 18100 -29460
rect 17900 -29760 17910 -29700
rect 18090 -29760 18100 -29700
rect 18560 -29700 18760 -29460
rect 18560 -29760 18570 -29700
rect 18750 -29760 18760 -29700
rect 19220 -29700 19420 -29460
rect 27910 -29468 29990 -29450
rect 27920 -29562 29990 -29468
rect 27910 -29580 29990 -29562
rect 27910 -29602 27922 -29580
rect 28802 -29602 28814 -29580
rect 27910 -29608 28814 -29602
rect 27370 -29670 27450 -29660
rect 27370 -29696 27380 -29670
rect 19220 -29760 19230 -29700
rect 19410 -29760 19420 -29700
rect 27260 -29742 27380 -29696
rect 27370 -29760 27380 -29742
rect 27440 -29696 27450 -29670
rect 27440 -29702 28726 -29696
rect 27440 -29736 27950 -29702
rect 28714 -29736 28726 -29702
rect 27440 -29742 28726 -29736
rect 27440 -29760 27450 -29742
rect 27370 -29770 27450 -29760
rect 27610 -29830 27690 -29820
rect 27610 -29854 27620 -29830
rect 2500 -29870 4020 -29860
rect 2500 -29930 2510 -29870
rect 4010 -29930 4020 -29870
rect 2500 -29942 4020 -29930
rect 4700 -29870 6220 -29860
rect 4700 -29930 4710 -29870
rect 6210 -29930 6220 -29870
rect 4700 -29942 6220 -29930
rect 6900 -29870 8420 -29860
rect 6900 -29930 6910 -29870
rect 8410 -29930 8420 -29870
rect 6900 -29942 8420 -29930
rect 9100 -29870 10620 -29860
rect 9100 -29930 9110 -29870
rect 10610 -29930 10620 -29870
rect 9100 -29942 10620 -29930
rect 11300 -29870 12820 -29860
rect 11300 -29930 11310 -29870
rect 12810 -29930 12820 -29870
rect 11300 -29942 12820 -29930
rect 13500 -29870 15020 -29860
rect 13500 -29930 13510 -29870
rect 15010 -29930 15020 -29870
rect 13500 -29942 15020 -29930
rect 15700 -29870 17220 -29860
rect 15700 -29930 15710 -29870
rect 17210 -29930 17220 -29870
rect 15700 -29942 17220 -29930
rect 17900 -29870 19420 -29860
rect 17900 -29930 17910 -29870
rect 19410 -29930 19420 -29870
rect 27260 -29900 27620 -29854
rect 27610 -29920 27620 -29900
rect 27680 -29854 27690 -29830
rect 28767 -29837 28813 -29759
rect 29790 -29800 29990 -29580
rect 27680 -29860 28726 -29854
rect 27680 -29894 27950 -29860
rect 28714 -29894 28726 -29860
rect 27680 -29900 28726 -29894
rect 27680 -29920 27690 -29900
rect 28770 -29917 28810 -29837
rect 27610 -29930 27690 -29920
rect 17900 -29942 19420 -29930
rect 4100 -30030 4220 -29970
rect 4280 -30030 4510 -29970
rect 6300 -30030 6420 -29970
rect 6480 -30030 6710 -29970
rect 8500 -30030 8840 -29970
rect 8900 -30030 8910 -29970
rect 10700 -30030 11040 -29970
rect 11100 -30030 11110 -29970
rect 12900 -30030 13240 -29970
rect 13300 -30030 13310 -29970
rect 15100 -30030 15440 -29970
rect 15500 -30030 15510 -29970
rect 17300 -30030 17420 -29970
rect 17480 -30030 17710 -29970
rect 19500 -30030 19620 -29970
rect 19680 -30030 19910 -29970
rect 27370 -29985 27450 -29975
rect 27370 -30012 27380 -29985
rect 27260 -30058 27380 -30012
rect 2010 -30120 2020 -30060
rect 2080 -30120 2420 -30060
rect 27370 -30075 27380 -30058
rect 27440 -30012 27450 -29985
rect 28767 -29990 28813 -29917
rect 29070 -29930 29150 -29920
rect 29070 -29990 29080 -29930
rect 28767 -29995 29080 -29990
rect 27440 -30018 28726 -30012
rect 27440 -30052 27950 -30018
rect 28714 -30052 28726 -30018
rect 27440 -30058 28726 -30052
rect 27440 -30075 27450 -30058
rect 28770 -30075 29080 -29995
rect 4210 -30140 4220 -30080
rect 4280 -30140 4620 -30080
rect 6410 -30140 6640 -30080
rect 6700 -30140 6820 -30080
rect 8610 -30140 8840 -30080
rect 8900 -30140 9020 -30080
rect 10810 -30140 11040 -30080
rect 11100 -30140 11220 -30080
rect 13010 -30140 13240 -30080
rect 13300 -30140 13420 -30080
rect 15210 -30140 15220 -30080
rect 15280 -30140 15620 -30080
rect 17410 -30140 17420 -30080
rect 17480 -30140 17820 -30080
rect 27370 -30085 27450 -30075
rect 28767 -30080 29080 -30075
rect 27610 -30145 27690 -30135
rect 27610 -30170 27620 -30145
rect 27260 -30216 27620 -30170
rect 27610 -30235 27620 -30216
rect 27680 -30170 27690 -30145
rect 28767 -30153 28813 -30080
rect 29070 -30130 29080 -30080
rect 29140 -30130 29150 -29930
rect 29070 -30140 29150 -30130
rect 27680 -30176 28726 -30170
rect 27680 -30210 27950 -30176
rect 28714 -30210 28726 -30176
rect 27680 -30216 28726 -30210
rect 27680 -30235 27690 -30216
rect 28770 -30233 28810 -30153
rect 29790 -30220 29980 -29800
rect 38260 -30140 38294 -30100
rect 27610 -30245 27690 -30235
rect 2500 -30360 2700 -30260
rect 2500 -30420 2510 -30360
rect 2690 -30420 2700 -30360
rect 2500 -30560 2700 -30420
rect 3160 -30360 3360 -30260
rect 3160 -30420 3170 -30360
rect 3350 -30420 3360 -30360
rect 3160 -30560 3360 -30420
rect 3820 -30360 4020 -30260
rect 3820 -30420 3830 -30360
rect 4010 -30420 4020 -30360
rect 3820 -30560 4020 -30420
rect 4700 -30360 4900 -30260
rect 4700 -30420 4710 -30360
rect 4890 -30420 4900 -30360
rect 4700 -30560 4900 -30420
rect 5360 -30360 5560 -30260
rect 5360 -30420 5370 -30360
rect 5550 -30420 5560 -30360
rect 5360 -30560 5560 -30420
rect 6020 -30360 6220 -30260
rect 6020 -30420 6030 -30360
rect 6210 -30420 6220 -30360
rect 6020 -30560 6220 -30420
rect 6900 -30500 7100 -30260
rect 6900 -30560 6910 -30500
rect 7090 -30560 7100 -30500
rect 7560 -30500 7760 -30260
rect 7560 -30560 7570 -30500
rect 7750 -30560 7760 -30500
rect 8220 -30500 8420 -30260
rect 8220 -30560 8230 -30500
rect 8410 -30560 8420 -30500
rect 9100 -30500 9300 -30260
rect 9100 -30560 9110 -30500
rect 9290 -30560 9300 -30500
rect 9760 -30500 9960 -30260
rect 9760 -30560 9770 -30500
rect 9950 -30560 9960 -30500
rect 10420 -30500 10620 -30260
rect 10420 -30560 10430 -30500
rect 10610 -30560 10620 -30500
rect 11300 -30500 11500 -30260
rect 11300 -30560 11310 -30500
rect 11490 -30560 11500 -30500
rect 11960 -30500 12160 -30260
rect 11960 -30560 11970 -30500
rect 12150 -30560 12160 -30500
rect 12620 -30500 12820 -30260
rect 12620 -30560 12630 -30500
rect 12810 -30560 12820 -30500
rect 13500 -30500 13700 -30260
rect 13500 -30560 13510 -30500
rect 13690 -30560 13700 -30500
rect 14160 -30500 14360 -30260
rect 14160 -30560 14170 -30500
rect 14350 -30560 14360 -30500
rect 14820 -30500 15020 -30260
rect 14820 -30560 14830 -30500
rect 15010 -30560 15020 -30500
rect 15700 -30360 15900 -30260
rect 15700 -30420 15710 -30360
rect 15890 -30420 15900 -30360
rect 15700 -30560 15900 -30420
rect 16360 -30360 16560 -30260
rect 16360 -30420 16370 -30360
rect 16550 -30420 16560 -30360
rect 16360 -30560 16560 -30420
rect 17020 -30360 17220 -30260
rect 17020 -30420 17030 -30360
rect 17210 -30420 17220 -30360
rect 17020 -30560 17220 -30420
rect 17900 -30360 18100 -30260
rect 17900 -30420 17910 -30360
rect 18090 -30420 18100 -30360
rect 17900 -30560 18100 -30420
rect 18560 -30360 18760 -30260
rect 18560 -30420 18570 -30360
rect 18750 -30420 18760 -30360
rect 18560 -30560 18760 -30420
rect 19220 -30360 19420 -30260
rect 27370 -30300 27450 -30290
rect 27370 -30328 27380 -30300
rect 19220 -30420 19230 -30360
rect 19410 -30420 19420 -30360
rect 27260 -30374 27380 -30328
rect 27370 -30390 27380 -30374
rect 27440 -30328 27450 -30300
rect 28767 -30311 28813 -30233
rect 27440 -30334 28726 -30328
rect 27440 -30368 27950 -30334
rect 28714 -30368 28726 -30334
rect 27440 -30374 28726 -30368
rect 27440 -30390 27450 -30374
rect 27370 -30400 27450 -30390
rect 19220 -30560 19420 -30420
rect 27910 -30468 28814 -30462
rect 27910 -30502 27922 -30468
rect 28802 -30480 28814 -30468
rect 29790 -30480 29990 -30220
rect 27930 -30502 29990 -30480
rect 27910 -30508 29990 -30502
rect 27930 -30602 29990 -30508
rect 27910 -30608 29990 -30602
rect 27910 -30642 27922 -30608
rect 27930 -30610 29990 -30608
rect 28802 -30642 28814 -30610
rect 27910 -30648 28814 -30642
rect 2500 -30670 4020 -30660
rect 2500 -30730 2510 -30670
rect 4010 -30730 4020 -30670
rect 2500 -30742 4020 -30730
rect 4700 -30670 6220 -30660
rect 4700 -30730 4710 -30670
rect 6210 -30730 6220 -30670
rect 4700 -30742 6220 -30730
rect 6900 -30670 8420 -30660
rect 6900 -30730 6910 -30670
rect 8410 -30730 8420 -30670
rect 6900 -30742 8420 -30730
rect 9100 -30670 10620 -30660
rect 9100 -30730 9110 -30670
rect 10610 -30730 10620 -30670
rect 9100 -30742 10620 -30730
rect 11300 -30670 12820 -30660
rect 11300 -30730 11310 -30670
rect 12810 -30730 12820 -30670
rect 11300 -30742 12820 -30730
rect 13500 -30670 15020 -30660
rect 13500 -30730 13510 -30670
rect 15010 -30730 15020 -30670
rect 13500 -30742 15020 -30730
rect 15700 -30670 17220 -30660
rect 15700 -30730 15710 -30670
rect 17210 -30730 17220 -30670
rect 15700 -30742 17220 -30730
rect 17900 -30670 19420 -30660
rect 17900 -30730 17910 -30670
rect 19410 -30730 19420 -30670
rect 17900 -30740 19420 -30730
rect 27370 -30710 27450 -30700
rect 27370 -30736 27380 -30710
rect 4100 -30830 4440 -30770
rect 4500 -30830 4510 -30770
rect 6300 -30830 6640 -30770
rect 6700 -30830 6710 -30770
rect 8500 -30830 8620 -30770
rect 8680 -30830 8910 -30770
rect 10700 -30830 10820 -30770
rect 10880 -30830 11110 -30770
rect 12900 -30830 13020 -30770
rect 13080 -30830 13310 -30770
rect 15100 -30830 15220 -30770
rect 15280 -30830 15510 -30770
rect 17300 -30830 17640 -30770
rect 17700 -30830 17710 -30770
rect 19500 -30830 19840 -30770
rect 19900 -30830 19910 -30770
rect 27260 -30782 27380 -30736
rect 27370 -30800 27380 -30782
rect 27440 -30736 27450 -30710
rect 27440 -30742 28726 -30736
rect 27440 -30776 27950 -30742
rect 28714 -30776 28726 -30742
rect 27440 -30782 28726 -30776
rect 27440 -30800 27450 -30782
rect 27370 -30810 27450 -30800
rect 2010 -30920 2240 -30860
rect 2300 -30920 2420 -30860
rect 27490 -30870 27570 -30860
rect 4210 -30940 4440 -30880
rect 4500 -30940 4620 -30880
rect 6410 -30940 6420 -30880
rect 6480 -30940 6820 -30880
rect 8610 -30940 8620 -30880
rect 8680 -30940 9020 -30880
rect 10810 -30940 10820 -30880
rect 10880 -30940 11220 -30880
rect 13010 -30940 13020 -30880
rect 13080 -30940 13420 -30880
rect 15210 -30940 15440 -30880
rect 15500 -30940 15620 -30880
rect 17410 -30940 17640 -30880
rect 17700 -30940 17820 -30880
rect 27490 -30894 27500 -30870
rect 27260 -30940 27500 -30894
rect 27490 -30960 27500 -30940
rect 27560 -30894 27570 -30870
rect 28767 -30877 28813 -30799
rect 27560 -30900 28726 -30894
rect 27560 -30934 27950 -30900
rect 28714 -30934 28726 -30900
rect 27560 -30940 28726 -30934
rect 27560 -30960 27570 -30940
rect 28770 -30957 28810 -30877
rect 27490 -30970 27570 -30960
rect 28767 -30960 28813 -30957
rect 29060 -30960 29300 -30950
rect 27370 -31025 27450 -31015
rect 27370 -31052 27380 -31025
rect 2500 -31300 2700 -31060
rect 2500 -31360 2510 -31300
rect 2690 -31360 2700 -31300
rect 3160 -31300 3360 -31060
rect 3160 -31360 3170 -31300
rect 3350 -31360 3360 -31300
rect 3820 -31300 4020 -31060
rect 3820 -31360 3830 -31300
rect 4010 -31360 4020 -31300
rect 4700 -31300 4900 -31060
rect 4700 -31360 4710 -31300
rect 4890 -31360 4900 -31300
rect 5360 -31300 5560 -31060
rect 5360 -31360 5370 -31300
rect 5550 -31360 5560 -31300
rect 6020 -31300 6220 -31060
rect 6020 -31360 6030 -31300
rect 6210 -31360 6220 -31300
rect 6900 -31160 7100 -31060
rect 6900 -31220 6910 -31160
rect 7090 -31220 7100 -31160
rect 6900 -31360 7100 -31220
rect 7560 -31160 7760 -31060
rect 7560 -31220 7570 -31160
rect 7750 -31220 7760 -31160
rect 7560 -31360 7760 -31220
rect 8220 -31160 8420 -31060
rect 8220 -31220 8230 -31160
rect 8410 -31220 8420 -31160
rect 8220 -31360 8420 -31220
rect 9100 -31160 9300 -31060
rect 9100 -31220 9110 -31160
rect 9290 -31220 9300 -31160
rect 9100 -31360 9300 -31220
rect 9760 -31160 9960 -31060
rect 9760 -31220 9770 -31160
rect 9950 -31220 9960 -31160
rect 9760 -31360 9960 -31220
rect 10420 -31160 10620 -31060
rect 10420 -31220 10430 -31160
rect 10610 -31220 10620 -31160
rect 10420 -31360 10620 -31220
rect 11300 -31160 11500 -31060
rect 11300 -31220 11310 -31160
rect 11490 -31220 11500 -31160
rect 11300 -31360 11500 -31220
rect 11960 -31160 12160 -31060
rect 11960 -31220 11970 -31160
rect 12150 -31220 12160 -31160
rect 11960 -31360 12160 -31220
rect 12620 -31160 12820 -31060
rect 12620 -31220 12630 -31160
rect 12810 -31220 12820 -31160
rect 12620 -31360 12820 -31220
rect 13500 -31160 13700 -31060
rect 13500 -31220 13510 -31160
rect 13690 -31220 13700 -31160
rect 13500 -31360 13700 -31220
rect 14160 -31160 14360 -31060
rect 14160 -31220 14170 -31160
rect 14350 -31220 14360 -31160
rect 14160 -31360 14360 -31220
rect 14820 -31160 15020 -31060
rect 14820 -31220 14830 -31160
rect 15010 -31220 15020 -31160
rect 14820 -31360 15020 -31220
rect 15700 -31300 15900 -31060
rect 15700 -31360 15710 -31300
rect 15890 -31360 15900 -31300
rect 16360 -31300 16560 -31060
rect 16360 -31360 16370 -31300
rect 16550 -31360 16560 -31300
rect 17020 -31300 17220 -31060
rect 17020 -31360 17030 -31300
rect 17210 -31360 17220 -31300
rect 17900 -31300 18100 -31060
rect 17900 -31360 17910 -31300
rect 18090 -31360 18100 -31300
rect 18560 -31300 18760 -31060
rect 18560 -31360 18570 -31300
rect 18750 -31360 18760 -31300
rect 19220 -31300 19420 -31060
rect 27260 -31098 27380 -31052
rect 27370 -31115 27380 -31098
rect 27440 -31052 27450 -31025
rect 28767 -31030 29070 -30960
rect 29290 -31030 29300 -30960
rect 28767 -31035 28813 -31030
rect 27440 -31058 28726 -31052
rect 27440 -31092 27950 -31058
rect 28714 -31092 28726 -31058
rect 27440 -31098 28726 -31092
rect 27440 -31115 27450 -31098
rect 28770 -31115 28810 -31035
rect 29060 -31040 29300 -31030
rect 27370 -31125 27450 -31115
rect 27490 -31185 27570 -31175
rect 27490 -31210 27500 -31185
rect 27260 -31256 27500 -31210
rect 27490 -31275 27500 -31256
rect 27560 -31210 27570 -31185
rect 28767 -31193 28813 -31115
rect 27560 -31216 28726 -31210
rect 27560 -31250 27950 -31216
rect 28714 -31250 28726 -31216
rect 27560 -31256 28726 -31250
rect 27560 -31275 27570 -31256
rect 28770 -31273 28810 -31193
rect 27490 -31285 27570 -31275
rect 19220 -31360 19230 -31300
rect 19410 -31360 19420 -31300
rect 27370 -31340 27450 -31330
rect 27370 -31368 27380 -31340
rect 27260 -31414 27380 -31368
rect 27370 -31430 27380 -31414
rect 27440 -31368 27450 -31340
rect 28767 -31351 28813 -31273
rect 27440 -31374 28726 -31368
rect 27440 -31408 27950 -31374
rect 28714 -31408 28726 -31374
rect 27440 -31414 28726 -31408
rect 27440 -31430 27450 -31414
rect 27370 -31440 27450 -31430
rect 23030 -31900 24240 -31500
rect 24360 -31900 25570 -31500
rect 25690 -31510 26230 -31500
rect 25690 -31880 25700 -31510
rect 26220 -31880 26230 -31510
rect 27910 -31508 28814 -31502
rect 27910 -31542 27922 -31508
rect 28802 -31520 28814 -31508
rect 29790 -31520 29990 -30610
rect 32600 -30690 32700 -30140
rect 32786 -30336 32854 -30326
rect 32786 -30488 32794 -30336
rect 32846 -30488 32854 -30336
rect 32786 -30498 32854 -30488
rect 33118 -30342 33186 -30330
rect 33118 -30494 33126 -30342
rect 33178 -30494 33186 -30342
rect 33118 -30502 33186 -30494
rect 33280 -30690 33700 -30140
rect 33780 -30336 33854 -30326
rect 34130 -30330 34190 -30328
rect 33780 -30488 33794 -30336
rect 33846 -30488 33854 -30336
rect 33780 -30498 33854 -30488
rect 34118 -30342 34190 -30330
rect 34118 -30494 34126 -30342
rect 34178 -30494 34190 -30342
rect 34118 -30500 34190 -30494
rect 34280 -30690 34700 -30140
rect 34780 -30336 34854 -30326
rect 35130 -30330 35190 -30328
rect 34780 -30488 34794 -30336
rect 34846 -30488 34854 -30336
rect 34780 -30498 34854 -30488
rect 35118 -30342 35190 -30330
rect 35118 -30494 35126 -30342
rect 35178 -30494 35190 -30342
rect 35118 -30500 35190 -30494
rect 35280 -30690 35700 -30140
rect 35780 -30336 35854 -30326
rect 36130 -30330 36190 -30328
rect 35780 -30488 35794 -30336
rect 35846 -30488 35854 -30336
rect 35780 -30498 35854 -30488
rect 36118 -30342 36190 -30330
rect 36118 -30494 36126 -30342
rect 36178 -30494 36190 -30342
rect 36118 -30500 36190 -30494
rect 36280 -30690 36700 -30140
rect 36780 -30336 36854 -30326
rect 37130 -30330 37190 -30328
rect 36780 -30488 36794 -30336
rect 36846 -30488 36854 -30336
rect 36780 -30498 36854 -30488
rect 37118 -30342 37190 -30330
rect 37118 -30494 37126 -30342
rect 37178 -30494 37190 -30342
rect 37118 -30500 37190 -30494
rect 37280 -30690 37700 -30140
rect 38260 -30154 38612 -30140
rect 37780 -30336 37854 -30326
rect 38130 -30330 38190 -30328
rect 37780 -30488 37794 -30336
rect 37846 -30488 37854 -30336
rect 37780 -30498 37854 -30488
rect 38118 -30342 38190 -30330
rect 38118 -30494 38126 -30342
rect 38178 -30494 38190 -30342
rect 38118 -30500 38190 -30494
rect 38260 -30690 38410 -30154
rect 32580 -30730 38410 -30690
rect 38588 -30730 38612 -30154
rect 32580 -30742 38612 -30730
rect 27940 -31542 29990 -31520
rect 27910 -31548 29990 -31542
rect 27940 -31650 29990 -31548
rect 25690 -31890 26230 -31880
rect 29790 -31940 29990 -31650
rect 31500 -31002 31800 -31000
rect 39150 -31002 39229 -28540
rect 31500 -31083 39229 -31002
rect 39263 -31002 39350 8958
rect 39263 -31083 39351 -31002
rect 31500 -31142 39351 -31083
rect 31500 -31206 31742 -31142
rect 39152 -31206 39351 -31142
rect 31500 -31249 39351 -31206
rect 31500 -31660 31636 -31249
rect 30780 -31680 31636 -31660
rect 30780 -32060 30840 -31680
rect 30820 -32440 30840 -32060
rect 31240 -32060 31636 -31680
rect 31240 -32440 31260 -32060
rect 30820 -32460 31260 -32440
rect 31500 -33000 31636 -32060
rect -1349 -33123 31636 -33000
rect 31670 -31292 39351 -31249
rect 31670 -33123 31800 -31292
rect 39500 -31400 39566 9820
rect 32600 -31580 39566 -31400
rect 32600 -31980 32700 -31580
rect 33280 -31980 33700 -31580
rect 34280 -31980 34700 -31580
rect 35280 -31980 35700 -31580
rect 36280 -31980 36700 -31580
rect 37280 -31980 37700 -31580
rect 38260 -32000 39566 -31580
rect 33128 -32592 33202 -32370
rect 33280 -32680 33680 -32170
rect 34128 -32592 34202 -32370
rect 34290 -32680 34690 -32170
rect 35128 -32592 35202 -32370
rect 35280 -32680 35680 -32170
rect 36128 -32592 36202 -32370
rect 36290 -32680 36690 -32170
rect 37128 -32592 37202 -32370
rect 37290 -32680 37690 -32170
rect 38270 -32180 38540 -32160
rect 38270 -32314 38406 -32180
rect 38128 -32592 38202 -32370
rect 38270 -32680 38320 -32314
rect 32660 -32690 38320 -32680
rect 38520 -32690 38540 -32180
rect 32660 -32910 38310 -32690
rect 38530 -32910 38540 -32690
rect 32660 -32920 38540 -32910
rect -1500 -33189 31800 -33123
rect -1500 -33223 -1283 -33189
rect 31570 -33223 31800 -33189
rect -1500 -33300 31800 -33223
rect 39500 -33500 39566 -32000
rect -1766 -33504 39566 -33500
rect 39600 -33504 39700 13504
rect -1900 -33566 39700 -33504
rect -1900 -33600 -1704 -33566
rect 39504 -33600 39700 -33566
rect -1900 -33700 39700 -33600
<< via1 >>
rect 25720 11410 26240 11780
rect 27260 11400 27320 11490
rect 27740 11240 27800 11330
rect 2510 11180 2690 11240
rect 3170 11180 3350 11240
rect 3830 11180 4010 11240
rect 4710 11180 4890 11240
rect 5370 11180 5550 11240
rect 6030 11180 6210 11240
rect 6910 11040 7090 11100
rect 7570 11040 7750 11100
rect 8230 11040 8410 11100
rect 9110 11040 9290 11100
rect 9770 11040 9950 11100
rect 10430 11040 10610 11100
rect 11310 11040 11490 11100
rect 11970 11040 12150 11100
rect 12630 11040 12810 11100
rect 13510 11040 13690 11100
rect 14170 11040 14350 11100
rect 14830 11040 15010 11100
rect 15710 11180 15890 11240
rect 16370 11180 16550 11240
rect 17030 11180 17210 11240
rect 17910 11180 18090 11240
rect 18570 11180 18750 11240
rect 19230 11180 19410 11240
rect 27260 11080 27320 11170
rect -70 10870 -10 10930
rect 2130 10870 2190 10930
rect 4330 10870 4390 10930
rect 6530 10870 6590 10930
rect 8730 10870 8790 10930
rect 10930 10870 10990 10930
rect 13130 10870 13190 10930
rect 15330 10870 15390 10930
rect 17530 10870 17590 10930
rect 19730 10870 19790 10930
rect 21930 10870 21990 10930
rect 27740 10925 27800 11015
rect 4220 10760 4280 10820
rect 6420 10760 6480 10820
rect 8840 10760 8900 10820
rect 11040 10760 11100 10820
rect 13240 10760 13300 10820
rect 15440 10760 15500 10820
rect 17420 10760 17480 10820
rect 19620 10740 19680 10800
rect 27260 10765 27320 10855
rect 29270 11060 29330 11280
rect 2020 10650 2080 10710
rect 4220 10650 4280 10710
rect 6640 10650 6700 10710
rect 8840 10650 8900 10710
rect 11040 10650 11100 10710
rect 13240 10650 13300 10710
rect 15220 10650 15280 10710
rect 17420 10650 17480 10710
rect 2510 10550 4010 10610
rect 4710 10550 6210 10610
rect 6910 10550 8410 10610
rect 9110 10550 10610 10610
rect 11310 10550 12810 10610
rect 13510 10550 15010 10610
rect 15710 10550 17210 10610
rect 17910 10550 19410 10610
rect 2510 10240 2690 10300
rect 3170 10240 3350 10300
rect 3830 10240 4010 10300
rect 4710 10240 4890 10300
rect 5370 10240 5550 10300
rect 6030 10240 6210 10300
rect 6910 10380 7090 10440
rect 7570 10380 7750 10440
rect 8230 10380 8410 10440
rect 9110 10380 9290 10440
rect 9770 10380 9950 10440
rect 10430 10380 10610 10440
rect 11310 10380 11490 10440
rect 11970 10380 12150 10440
rect 12630 10380 12810 10440
rect 13510 10380 13690 10440
rect 14170 10380 14350 10440
rect 14830 10380 15010 10440
rect 15710 10240 15890 10300
rect 16370 10240 16550 10300
rect 17030 10240 17210 10300
rect 17910 10240 18090 10300
rect 18570 10240 18750 10300
rect 27740 10360 27800 10450
rect 19230 10240 19410 10300
rect 27380 10200 27440 10290
rect -70 10070 -10 10130
rect 2130 10070 2190 10130
rect 4330 10070 4390 10130
rect 6530 10070 6590 10130
rect 8730 10070 8790 10130
rect 10930 10070 10990 10130
rect 13130 10070 13190 10130
rect 15330 10070 15390 10130
rect 17530 10070 17590 10130
rect 19730 10070 19790 10130
rect 21930 10070 21990 10130
rect 27740 10040 27800 10130
rect 4440 9960 4500 10020
rect 6640 9960 6700 10020
rect 8620 9960 8680 10020
rect 10820 9960 10880 10020
rect 13020 9960 13080 10020
rect 15220 9960 15280 10020
rect 17640 9960 17700 10020
rect 19840 9940 19900 10000
rect 2240 9850 2300 9910
rect 4440 9850 4500 9910
rect 6420 9850 6480 9910
rect 8620 9850 8680 9910
rect 10820 9850 10880 9910
rect 13020 9850 13080 9910
rect 15440 9850 15500 9910
rect 17640 9850 17700 9910
rect 27380 9885 27440 9975
rect 2510 9750 4010 9810
rect 4710 9750 6210 9810
rect 6910 9750 8410 9810
rect 9110 9750 10610 9810
rect 11310 9750 12810 9810
rect 13510 9750 15010 9810
rect 15710 9750 17210 9810
rect 17910 9750 19410 9810
rect 27740 9725 27800 9815
rect 29140 9970 29200 10190
rect 36920 12280 38280 12540
rect 30826 10346 31190 10876
rect 31422 10082 31494 10262
rect 31756 10082 31828 10262
rect 32556 10082 32628 10262
rect 33356 10082 33428 10262
rect 2510 9580 2690 9640
rect 3170 9580 3350 9640
rect 3830 9580 4010 9640
rect 4710 9580 4890 9640
rect 5370 9580 5550 9640
rect 6030 9580 6210 9640
rect 6910 9440 7090 9500
rect 7570 9440 7750 9500
rect 8230 9440 8410 9500
rect 9110 9440 9290 9500
rect 9770 9440 9950 9500
rect 10430 9440 10610 9500
rect 11310 9440 11490 9500
rect 11970 9440 12150 9500
rect 12630 9440 12810 9500
rect 13510 9440 13690 9500
rect 14170 9440 14350 9500
rect 14830 9440 15010 9500
rect 15710 9580 15890 9640
rect 16370 9580 16550 9640
rect 17030 9580 17210 9640
rect 17910 9580 18090 9640
rect 18570 9580 18750 9640
rect 19230 9580 19410 9640
rect -70 9270 -10 9330
rect 2130 9270 2190 9330
rect 4330 9270 4390 9330
rect 6530 9270 6590 9330
rect 8730 9270 8790 9330
rect 10930 9270 10990 9330
rect 13130 9270 13190 9330
rect 15330 9270 15390 9330
rect 17530 9270 17590 9330
rect 19730 9270 19790 9330
rect 1420 9060 1480 9210
rect 6420 9160 6480 9220
rect 8840 9160 8900 9220
rect 11040 9160 11100 9220
rect 13240 9160 13300 9220
rect 15440 9160 15500 9220
rect 17420 9160 17480 9220
rect 20240 9150 20300 9300
rect 21930 9270 21990 9330
rect 27260 9315 27320 9405
rect 27500 9160 27560 9250
rect 4220 9050 4280 9110
rect 6640 9050 6700 9110
rect 8840 9050 8900 9110
rect 11040 9050 11100 9110
rect 13240 9050 13300 9110
rect 15220 9050 15280 9110
rect 430 8910 610 8990
rect 4710 8950 6210 9010
rect 6910 8950 8410 9010
rect 9110 8950 10610 9010
rect 11310 8950 12810 9010
rect 13510 8950 15010 9010
rect 15710 8950 17210 9010
rect 27260 9000 27320 9090
rect 21310 8910 21490 8990
rect 27500 8845 27560 8935
rect 2510 8640 2690 8700
rect 3170 8640 3350 8700
rect 3830 8640 4010 8700
rect 4710 8640 4890 8700
rect 5370 8640 5550 8700
rect 6030 8640 6210 8700
rect 6910 8780 7090 8840
rect 7570 8780 7750 8840
rect 8230 8780 8410 8840
rect 9110 8780 9290 8840
rect 9770 8780 9950 8840
rect 10430 8780 10610 8840
rect 11310 8780 11490 8840
rect 11970 8780 12150 8840
rect 12630 8780 12810 8840
rect 13510 8780 13690 8840
rect 14170 8780 14350 8840
rect 14830 8780 15010 8840
rect 15710 8640 15890 8700
rect 16370 8640 16550 8700
rect 17030 8640 17210 8700
rect 17910 8640 18090 8700
rect 18570 8640 18750 8700
rect 19230 8640 19410 8700
rect 27260 8685 27320 8775
rect 28880 8940 28940 9160
rect 34490 10846 34848 11022
rect 36940 11850 37070 12030
rect 37360 11850 37490 12030
rect 37780 11850 37910 12030
rect 36990 11300 37050 11680
rect 35820 10070 36010 10140
rect 36140 10070 36330 10140
rect 37410 11300 37470 11680
rect 37190 10860 37340 11010
rect 36990 10320 37050 10500
rect 37830 11300 37890 11680
rect 37610 10600 37760 10750
rect 37410 10320 37470 10500
rect 37990 10780 38120 10960
rect 37830 10320 37890 10500
rect 36950 9980 37080 10160
rect 37370 9980 37500 10160
rect 37790 9980 37920 10160
rect 35266 9542 35384 9664
rect 36430 9434 36542 9924
rect 38298 9848 39274 10406
rect 37584 9542 37702 9664
rect -70 8470 -10 8530
rect 2130 8470 2190 8530
rect 4330 8470 4390 8530
rect 6530 8470 6590 8530
rect 8730 8470 8790 8530
rect 10930 8470 10990 8530
rect 13130 8470 13190 8530
rect 15330 8470 15390 8530
rect 17530 8470 17590 8530
rect 19730 8470 19790 8530
rect 1620 8260 1680 8410
rect 6640 8360 6700 8420
rect 8620 8360 8680 8420
rect 10820 8360 10880 8420
rect 13020 8360 13080 8420
rect 15220 8360 15280 8420
rect 17640 8360 17700 8420
rect 20440 8350 20500 8500
rect 21930 8470 21990 8530
rect 4440 8250 4500 8310
rect 6420 8250 6480 8310
rect 8620 8250 8680 8310
rect 10820 8250 10880 8310
rect 13020 8250 13080 8310
rect 15440 8250 15500 8310
rect 27260 8280 27320 8370
rect 430 8110 610 8190
rect 4710 8150 6210 8210
rect 6910 8150 8410 8210
rect 9110 8150 10610 8210
rect 11310 8150 12810 8210
rect 13510 8150 15010 8210
rect 15710 8150 17210 8210
rect 21310 8110 21490 8190
rect 27620 8120 27680 8210
rect 2510 7840 2690 7900
rect 3170 7840 3350 7900
rect 3830 7840 4010 7900
rect 4710 7840 4890 7900
rect 5370 7840 5550 7900
rect 6030 7840 6210 7900
rect 6910 7980 7090 8040
rect 7570 7980 7750 8040
rect 8230 7980 8410 8040
rect 9110 7980 9290 8040
rect 9770 7980 9950 8040
rect 10430 7980 10610 8040
rect 11310 7980 11490 8040
rect 11970 7980 12150 8040
rect 12630 7980 12810 8040
rect 13510 7980 13690 8040
rect 14170 7980 14350 8040
rect 14830 7980 15010 8040
rect 15710 7840 15890 7900
rect 16370 7840 16550 7900
rect 17030 7840 17210 7900
rect 17910 7840 18090 7900
rect 18570 7840 18750 7900
rect 27260 7960 27320 8050
rect 19230 7840 19410 7900
rect 27620 7800 27680 7890
rect -70 7670 -10 7730
rect 2130 7670 2190 7730
rect 4330 7670 4390 7730
rect 6530 7670 6590 7730
rect 8730 7670 8790 7730
rect 10930 7670 10990 7730
rect 13130 7670 13190 7730
rect 15330 7670 15390 7730
rect 17530 7670 17590 7730
rect 19730 7670 19790 7730
rect 1620 7460 1680 7610
rect 6640 7560 6700 7620
rect 8620 7560 8680 7620
rect 10820 7560 10880 7620
rect 13020 7560 13080 7620
rect 15220 7560 15280 7620
rect 17640 7560 17700 7620
rect 20440 7550 20500 7700
rect 21930 7670 21990 7730
rect 27260 7650 27320 7740
rect 29010 7890 29070 8110
rect 35254 8292 35372 8414
rect 4440 7450 4500 7510
rect 6420 7450 6480 7510
rect 8620 7450 8680 7510
rect 10820 7450 10880 7510
rect 13020 7450 13080 7510
rect 15440 7450 15500 7510
rect 430 7310 610 7390
rect 4710 7350 6210 7410
rect 6910 7350 8410 7410
rect 9110 7350 10610 7410
rect 11310 7350 12810 7410
rect 13510 7350 15010 7410
rect 15710 7350 17210 7410
rect 21310 7310 21490 7390
rect 27380 7240 27440 7330
rect 2510 7180 2690 7240
rect 3170 7180 3350 7240
rect 3830 7180 4010 7240
rect 4710 7180 4890 7240
rect 5370 7180 5550 7240
rect 6030 7180 6210 7240
rect 6910 7040 7090 7100
rect 7570 7040 7750 7100
rect 8230 7040 8410 7100
rect 9110 7040 9290 7100
rect 9770 7040 9950 7100
rect 10430 7040 10610 7100
rect 11310 7040 11490 7100
rect 11970 7040 12150 7100
rect 12630 7040 12810 7100
rect 13510 7040 13690 7100
rect 14170 7040 14350 7100
rect 14830 7040 15010 7100
rect 15710 7180 15890 7240
rect 16370 7180 16550 7240
rect 17030 7180 17210 7240
rect 17910 7180 18090 7240
rect 18570 7180 18750 7240
rect 19230 7180 19410 7240
rect 27620 7080 27680 7170
rect -70 6870 -10 6930
rect 2130 6870 2190 6930
rect 4330 6870 4390 6930
rect 6530 6870 6590 6930
rect 8730 6870 8790 6930
rect 10930 6870 10990 6930
rect 13130 6870 13190 6930
rect 15330 6870 15390 6930
rect 17530 6870 17590 6930
rect 19730 6870 19790 6930
rect 1420 6660 1480 6810
rect 6420 6760 6480 6820
rect 8840 6760 8900 6820
rect 11040 6760 11100 6820
rect 13240 6760 13300 6820
rect 15440 6760 15500 6820
rect 17420 6760 17480 6820
rect 20240 6750 20300 6900
rect 21930 6870 21990 6930
rect 27380 6925 27440 7015
rect 27620 6765 27680 6855
rect 4220 6650 4280 6710
rect 6640 6650 6700 6710
rect 8840 6650 8900 6710
rect 11040 6650 11100 6710
rect 13240 6650 13300 6710
rect 15220 6650 15280 6710
rect 430 6510 610 6590
rect 4710 6550 6210 6610
rect 6910 6550 8410 6610
rect 9110 6550 10610 6610
rect 11310 6550 12810 6610
rect 13510 6550 15010 6610
rect 15710 6550 17210 6610
rect 27380 6610 27440 6700
rect 28880 6860 28940 7080
rect 37600 8294 37718 8416
rect 35370 7800 35490 7920
rect 35350 7570 35470 7690
rect 36880 7800 37000 7920
rect 36010 7500 36130 7620
rect 31290 7090 31570 7210
rect 21310 6510 21490 6590
rect 2510 6240 2690 6300
rect 3170 6240 3350 6300
rect 3830 6240 4010 6300
rect 4710 6240 4890 6300
rect 5370 6240 5550 6300
rect 6030 6240 6210 6300
rect 6910 6380 7090 6440
rect 7570 6380 7750 6440
rect 8230 6380 8410 6440
rect 9110 6380 9290 6440
rect 9770 6380 9950 6440
rect 10430 6380 10610 6440
rect 11310 6380 11490 6440
rect 11970 6380 12150 6440
rect 12630 6380 12810 6440
rect 13510 6380 13690 6440
rect 14170 6380 14350 6440
rect 14830 6380 15010 6440
rect 15710 6240 15890 6300
rect 16370 6240 16550 6300
rect 17030 6240 17210 6300
rect 17910 6240 18090 6300
rect 18570 6240 18750 6300
rect 19230 6240 19410 6300
rect 27380 6200 27440 6290
rect -70 6070 -10 6130
rect 2130 6070 2190 6130
rect 4330 6070 4390 6130
rect 6530 6070 6590 6130
rect 8730 6070 8790 6130
rect 10930 6070 10990 6130
rect 13130 6070 13190 6130
rect 15330 6070 15390 6130
rect 17530 6070 17590 6130
rect 19730 6070 19790 6130
rect 21930 6070 21990 6130
rect 27500 6040 27560 6130
rect 4440 5960 4500 6020
rect 6640 5960 6700 6020
rect 8620 5960 8680 6020
rect 10820 5960 10880 6020
rect 13020 5960 13080 6020
rect 15220 5960 15280 6020
rect 17640 5960 17700 6020
rect 19840 5940 19900 6000
rect 2240 5850 2300 5910
rect 4440 5850 4500 5910
rect 6420 5850 6480 5910
rect 8620 5850 8680 5910
rect 10820 5850 10880 5910
rect 13020 5850 13080 5910
rect 15440 5850 15500 5910
rect 17640 5850 17700 5910
rect 27380 5885 27440 5975
rect 2510 5750 4010 5810
rect 4710 5750 6210 5810
rect 6910 5750 8410 5810
rect 9110 5750 10610 5810
rect 11310 5750 12810 5810
rect 13510 5750 15010 5810
rect 15710 5750 17210 5810
rect 17910 5750 19410 5810
rect 27500 5725 27560 5815
rect 2510 5580 2690 5640
rect 3170 5580 3350 5640
rect 3830 5580 4010 5640
rect 4710 5580 4890 5640
rect 5370 5580 5550 5640
rect 6030 5580 6210 5640
rect 6910 5440 7090 5500
rect 7570 5440 7750 5500
rect 8230 5440 8410 5500
rect 9110 5440 9290 5500
rect 9770 5440 9950 5500
rect 10430 5440 10610 5500
rect 11310 5440 11490 5500
rect 11970 5440 12150 5500
rect 12630 5440 12810 5500
rect 13510 5440 13690 5500
rect 14170 5440 14350 5500
rect 14830 5440 15010 5500
rect 15710 5580 15890 5640
rect 16370 5580 16550 5640
rect 17030 5580 17210 5640
rect 17910 5580 18090 5640
rect 18570 5580 18750 5640
rect 19230 5580 19410 5640
rect 27380 5570 27440 5660
rect 29010 5820 29070 6040
rect -70 5270 -10 5330
rect 2130 5270 2190 5330
rect 4330 5270 4390 5330
rect 6530 5270 6590 5330
rect 8730 5270 8790 5330
rect 10930 5270 10990 5330
rect 13130 5270 13190 5330
rect 15330 5270 15390 5330
rect 17530 5270 17590 5330
rect 19730 5270 19790 5330
rect 21930 5270 21990 5330
rect 4220 5160 4280 5220
rect 6420 5160 6480 5220
rect 8840 5160 8900 5220
rect 11040 5160 11100 5220
rect 13240 5160 13300 5220
rect 15440 5160 15500 5220
rect 17420 5160 17480 5220
rect 19620 5140 19680 5200
rect 27180 5110 27310 5240
rect 2020 5050 2080 5110
rect 4220 5050 4280 5110
rect 6640 5050 6700 5110
rect 8840 5050 8900 5110
rect 11040 5050 11100 5110
rect 13240 5050 13300 5110
rect 15220 5050 15280 5110
rect 17420 5050 17480 5110
rect 2510 4950 4010 5010
rect 4710 4950 6210 5010
rect 6910 4950 8410 5010
rect 9110 4950 10610 5010
rect 11310 4950 12810 5010
rect 13510 4950 15010 5010
rect 15710 4950 17210 5010
rect 17910 4950 19410 5010
rect 7800 4540 7940 4680
rect 23050 4600 23580 4970
rect 10820 4360 10880 4420
rect 13240 4360 13300 4420
rect 37494 7504 37610 7620
rect 37510 7370 37630 7490
rect 36128 6982 36810 7176
rect 8620 4250 8680 4310
rect 11040 4250 11100 4310
rect 10890 3960 11030 4100
rect 30520 4750 30640 4870
rect 30910 4750 31030 4870
rect 36230 6080 36410 6260
rect 36530 6080 36710 6260
rect 36300 5820 36390 5890
rect 37680 5820 37770 5890
rect 36300 5560 36390 5630
rect 36300 5300 36390 5370
rect 37680 5560 37770 5630
rect 37680 5300 37770 5370
rect 36300 5040 36390 5110
rect 36300 4780 36390 4850
rect 37680 5040 37770 5110
rect 37680 4780 37770 4850
rect 36300 4520 36390 4590
rect 30080 3860 30260 4040
rect 31680 3860 31860 4040
rect 32810 4010 32980 4070
rect 33130 4010 33300 4070
rect 33440 4010 33610 4070
rect 33760 4010 33930 4070
rect 34870 4010 35190 4090
rect 32850 3350 33870 3430
rect 35070 3350 35410 3430
rect 36300 4260 36390 4330
rect 37680 4520 37770 4590
rect 37680 4260 37770 4330
rect 36300 4000 36390 4070
rect 36380 3440 36520 3580
rect 37680 4000 37770 4070
rect 32466 3068 32668 3156
rect 18060 2870 18200 3010
rect 16910 2640 17130 2780
rect 17380 2640 17490 2780
rect 17740 2640 17960 2780
rect 34066 3068 34268 3156
rect 32450 2430 32690 2510
rect 34050 2430 34290 2510
rect 35666 3068 35868 3156
rect 35650 2430 35890 2510
rect 480 -4780 660 2220
rect 32450 2070 32690 2130
rect 34050 2070 34290 2130
rect 35650 2070 35890 2130
rect 2110 1310 2230 1990
rect 3710 1310 3830 1990
rect 5310 1310 5430 1990
rect 6910 1310 7030 1990
rect 8510 1310 8630 1990
rect 10110 1310 10230 1990
rect 11030 1330 11150 1950
rect 12610 1330 12730 1950
rect 13990 1330 14110 1950
rect 14910 1320 15030 1980
rect 16510 1310 16630 1990
rect 18110 1310 18230 1990
rect 19710 1310 19830 1990
rect 21310 1310 21430 1990
rect 22910 1310 23030 1990
rect 24510 1310 24630 1990
rect 26110 1310 26230 1990
rect 27710 1310 27830 1990
rect 29310 1310 29430 1990
rect 30910 1310 31030 1990
rect 32510 1310 32630 1990
rect 34110 1310 34230 1990
rect 35710 1310 35830 1990
rect 37310 1310 37430 1990
rect 1410 1030 1530 1150
rect 3010 1030 3130 1150
rect 4610 1030 4730 1150
rect 6210 1030 6330 1150
rect 7810 1030 7930 1150
rect 9410 1030 9530 1150
rect 11250 1070 11670 1230
rect 15600 1030 15700 1150
rect 17200 1030 17300 1150
rect 18800 1030 18900 1150
rect 20400 1030 20500 1150
rect 22000 1030 22100 1150
rect 23600 1030 23700 1150
rect 26800 1030 26900 1150
rect 28400 1030 28500 1150
rect 12390 750 12510 870
rect 1190 560 1310 680
rect 2790 560 2910 680
rect 4390 560 4510 680
rect 5990 560 6110 680
rect 7590 560 7710 680
rect 9190 560 9310 680
rect 15820 560 15920 680
rect 17420 560 17520 680
rect 19020 560 19120 680
rect 20620 560 20720 680
rect 22220 560 22320 680
rect 23820 560 23920 680
rect 27020 560 27120 680
rect 28620 560 28720 680
rect 31820 560 31920 680
rect 36600 550 36720 670
rect 37850 530 37970 650
rect 2110 -490 2230 190
rect 3710 -490 3830 190
rect 5310 -490 5430 190
rect 6910 -490 7030 190
rect 8510 -490 8630 190
rect 10110 -490 10230 190
rect 11710 -570 11830 190
rect 13310 -490 13430 190
rect 1410 -770 1530 -650
rect 3010 -770 3130 -650
rect 4610 -770 4730 -650
rect 6210 -770 6330 -650
rect 7810 -770 7930 -650
rect 9410 -770 9530 -650
rect 11270 -730 12270 -570
rect 14910 -570 15030 190
rect 16510 -490 16630 190
rect 18110 -490 18230 190
rect 19710 -490 19830 190
rect 21310 -490 21430 190
rect 22910 -490 23030 190
rect 24510 -490 24630 190
rect 26110 -490 26230 190
rect 27710 -490 27830 190
rect 29310 -490 29430 190
rect 30910 -490 31030 190
rect 32510 -490 32630 190
rect 34110 -490 34230 190
rect 35710 -490 35830 190
rect 12390 -810 12510 -650
rect 14470 -730 15470 -570
rect 15600 -770 15700 -650
rect 17200 -770 17300 -650
rect 18800 -770 18900 -650
rect 20400 -770 20500 -650
rect 22000 -770 22100 -650
rect 23600 -770 23700 -650
rect 26800 -770 26900 -650
rect 28400 -770 28500 -650
rect 12390 -1050 12510 -980
rect 12630 -1070 12750 -930
rect 13970 -1070 14090 -930
rect 1190 -1240 1310 -1120
rect 2790 -1240 2910 -1120
rect 4390 -1240 4510 -1120
rect 5990 -1240 6110 -1120
rect 7590 -1240 7710 -1120
rect 9190 -1240 9310 -1120
rect 12880 -1260 13240 -1110
rect 15820 -1240 15920 -1120
rect 17420 -1240 17520 -1120
rect 19020 -1240 19120 -1120
rect 20620 -1240 20720 -1120
rect 22220 -1240 22320 -1120
rect 23820 -1240 23920 -1120
rect 27020 -1240 27120 -1120
rect 28620 -1240 28720 -1120
rect 31600 -1240 31700 -1120
rect 33360 -1590 33480 -1470
rect 2110 -2290 2230 -1610
rect 3710 -2290 3830 -1610
rect 5310 -2290 5430 -1610
rect 6910 -2290 7030 -1610
rect 8510 -2290 8630 -1610
rect 10110 -2290 10230 -1610
rect 11710 -2290 11830 -1610
rect 13310 -2290 13430 -1610
rect 14910 -2290 15030 -1610
rect 16510 -2290 16630 -1610
rect 18110 -2290 18230 -1610
rect 19710 -2290 19830 -1610
rect 21310 -2290 21430 -1610
rect 22910 -2290 23030 -1610
rect 24510 -2290 24630 -1610
rect 26110 -2290 26230 -1610
rect 27710 -2290 27830 -1610
rect 29310 -2290 29430 -1610
rect 30910 -2290 31030 -1610
rect 35020 -1590 35140 -1470
rect 32510 -2290 32630 -1610
rect 34110 -2290 34230 -1610
rect 35690 -2310 35750 -1600
rect 1410 -2570 1530 -2450
rect 3010 -2570 3130 -2450
rect 4610 -2570 4730 -2450
rect 6210 -2570 6330 -2450
rect 7810 -2570 7930 -2450
rect 9410 -2570 9530 -2450
rect 15600 -2570 15700 -2450
rect 17200 -2570 17300 -2450
rect 18800 -2570 18900 -2450
rect 20400 -2570 20500 -2450
rect 22000 -2570 22100 -2450
rect 23600 -2570 23700 -2450
rect 25200 -2570 25300 -2450
rect 26800 -2570 26900 -2450
rect 28400 -2570 28500 -2450
rect 30000 -2570 30100 -2450
rect 33180 -2570 33300 -2450
rect 12390 -2850 12510 -2730
rect 1190 -3040 1310 -2920
rect 2790 -3040 2910 -2920
rect 4390 -3040 4510 -2920
rect 5990 -3040 6110 -2920
rect 7590 -3040 7710 -2920
rect 9190 -3040 9310 -2920
rect 11010 -3040 11130 -2920
rect 14210 -3040 14330 -2920
rect 14430 -3040 14550 -2920
rect 15820 -3040 15920 -2920
rect 17420 -3040 17520 -2920
rect 19020 -3040 19120 -2920
rect 20620 -3040 20720 -2920
rect 22220 -3040 22320 -2920
rect 23820 -3040 23920 -2920
rect 25420 -3040 25520 -2920
rect 27020 -3040 27120 -2920
rect 28620 -3040 28720 -2920
rect 30220 -3040 30320 -2920
rect 36400 -3030 36500 -2910
rect 12610 -3390 12730 -3290
rect 2110 -4090 2230 -3410
rect 3710 -4090 3830 -3410
rect 5310 -4090 5430 -3410
rect 6910 -4090 7030 -3410
rect 8510 -4090 8630 -3410
rect 10110 -4090 10230 -3410
rect 11710 -4090 11830 -3410
rect 13310 -4090 13430 -3410
rect 14210 -3410 14330 -3290
rect 14910 -4090 15030 -3410
rect 16510 -4090 16630 -3410
rect 18110 -4090 18230 -3410
rect 19710 -4090 19830 -3410
rect 21310 -4090 21430 -3410
rect 22910 -4090 23030 -3410
rect 24510 -4090 24630 -3410
rect 26110 -4090 26230 -3410
rect 27710 -4090 27830 -3410
rect 29310 -4090 29430 -3410
rect 30910 -4090 31030 -3410
rect 33400 -3400 33530 -3280
rect 32510 -4090 32630 -3410
rect 34110 -4090 34230 -3410
rect 35710 -4090 35830 -3410
rect 1410 -4370 1530 -4250
rect 3010 -4370 3130 -4250
rect 4610 -4370 4730 -4250
rect 6210 -4370 6330 -4250
rect 7810 -4370 7930 -4250
rect 9410 -4370 9530 -4250
rect 15600 -4370 15700 -4250
rect 17200 -4370 17300 -4250
rect 18800 -4370 18900 -4250
rect 20400 -4370 20500 -4250
rect 22000 -4370 22100 -4250
rect 23600 -4370 23700 -4250
rect 25200 -4370 25300 -4250
rect 26800 -4370 26900 -4250
rect 28400 -4370 28500 -4250
rect 30000 -4370 30100 -4250
rect 33180 -4370 33300 -4250
rect 12390 -4650 12510 -4530
rect 1190 -4840 1310 -4720
rect 2790 -4840 2910 -4720
rect 4390 -4840 4510 -4720
rect 5990 -4840 6110 -4720
rect 7590 -4840 7710 -4720
rect 9190 -4840 9310 -4720
rect 11710 -4930 11830 -4810
rect 12610 -4850 12730 -4730
rect 13630 -4910 13750 -4790
rect 14210 -4850 14330 -4730
rect 15230 -4910 15350 -4790
rect 15820 -4840 15920 -4720
rect 17420 -4840 17520 -4720
rect 19020 -4840 19120 -4720
rect 20620 -4840 20720 -4720
rect 22220 -4840 22320 -4720
rect 23820 -4840 23920 -4720
rect 25420 -4840 25520 -4720
rect 27020 -4840 27120 -4720
rect 28620 -4840 28720 -4720
rect 30220 -4840 30320 -4720
rect 36400 -4830 36500 -4710
rect 11710 -5950 11830 -5830
rect 13310 -5950 13430 -5830
rect 11710 -6170 11830 -6050
rect 13630 -6170 13750 -6050
rect 14230 -6170 14350 -6050
rect 15230 -6170 15350 -6050
rect 12630 -6390 12750 -6270
rect 16510 -6390 16630 -6270
rect 12410 -6610 12530 -6490
rect 14910 -6610 15030 -6490
rect 12950 -6990 13110 -6830
rect 7810 -7990 7930 -7870
rect 14910 -8000 15040 -7880
rect 490 -22380 670 -8090
rect 1210 -8190 1330 -8070
rect 2810 -8190 2930 -8070
rect 4410 -8190 4530 -8070
rect 6010 -8190 6130 -8070
rect 7610 -8190 7730 -8070
rect 9210 -8190 9330 -8070
rect 11710 -8230 11840 -8110
rect 15830 -8190 15950 -8070
rect 17430 -8190 17550 -8070
rect 19030 -8190 19150 -8070
rect 20630 -8190 20750 -8070
rect 22230 -8190 22350 -8070
rect 23830 -8190 23950 -8070
rect 25430 -8190 25550 -8070
rect 27030 -8190 27150 -8070
rect 28630 -8190 28750 -8070
rect 30230 -8190 30350 -8070
rect 31830 -8190 31950 -8070
rect 34810 -8190 34930 -8070
rect 10810 -8380 10930 -8260
rect 16510 -8380 16640 -8260
rect 1430 -8630 1550 -8510
rect 3030 -8630 3150 -8510
rect 4630 -8630 4750 -8510
rect 6230 -8630 6350 -8510
rect 7830 -8630 7950 -8510
rect 9430 -8630 9550 -8510
rect 2130 -9470 2230 -8810
rect 3730 -9470 3830 -8810
rect 5330 -9470 5430 -8810
rect 6930 -9470 7030 -8810
rect 8530 -9470 8630 -8810
rect 10130 -9470 10230 -8810
rect 11720 -9470 11830 -8810
rect 15610 -8640 15730 -8520
rect 17210 -8640 17330 -8520
rect 18810 -8640 18930 -8520
rect 20410 -8640 20530 -8520
rect 22010 -8640 22130 -8520
rect 23610 -8640 23730 -8520
rect 25210 -8640 25330 -8520
rect 26810 -8640 26930 -8520
rect 28410 -8640 28530 -8520
rect 30010 -8640 30130 -8520
rect 13320 -9470 13430 -8810
rect 16520 -9480 16630 -8800
rect 18120 -9480 18230 -8800
rect 19720 -9480 19830 -8800
rect 21320 -9480 21430 -8800
rect 22920 -9480 23030 -8800
rect 24520 -9480 24630 -8800
rect 26120 -9480 26230 -8800
rect 27720 -9480 27830 -8800
rect 29320 -9480 29430 -8800
rect 30920 -9480 31030 -8800
rect 32520 -9360 32630 -8800
rect 34120 -9360 34230 -8800
rect 35720 -9360 35830 -8800
rect 33410 -9630 33530 -9510
rect 1210 -9990 1330 -9870
rect 2810 -9990 2930 -9870
rect 4410 -9990 4530 -9870
rect 6010 -9990 6130 -9870
rect 7610 -9990 7730 -9870
rect 9210 -9990 9330 -9870
rect 15830 -9990 15950 -9870
rect 17430 -9990 17550 -9870
rect 19030 -9990 19150 -9870
rect 20630 -9990 20750 -9870
rect 22230 -9990 22350 -9870
rect 23830 -9990 23950 -9870
rect 25430 -9990 25550 -9870
rect 27030 -9990 27150 -9870
rect 28630 -9990 28750 -9870
rect 30230 -9990 30350 -9870
rect 31830 -9990 31950 -9870
rect 34810 -9990 34930 -9870
rect 10810 -10180 10930 -10060
rect 1430 -10430 1550 -10310
rect 3030 -10430 3150 -10310
rect 4630 -10430 4750 -10310
rect 6230 -10430 6350 -10310
rect 7830 -10430 7950 -10310
rect 9430 -10430 9550 -10310
rect 11030 -10530 11150 -10410
rect 15610 -10440 15730 -10320
rect 2130 -11270 2230 -10610
rect 3730 -11270 3830 -10610
rect 5330 -11270 5430 -10610
rect 6930 -11270 7030 -10610
rect 8530 -11270 8630 -10610
rect 10130 -11270 10230 -10610
rect 11720 -11270 11830 -10610
rect 13320 -11270 13430 -10610
rect 17210 -10440 17330 -10320
rect 18810 -10440 18930 -10320
rect 20410 -10440 20530 -10320
rect 22010 -10440 22130 -10320
rect 23610 -10440 23730 -10320
rect 25210 -10440 25330 -10320
rect 26810 -10440 26930 -10320
rect 28410 -10440 28530 -10320
rect 30010 -10440 30130 -10320
rect 31610 -10440 31730 -10320
rect 16520 -11280 16630 -10600
rect 18120 -11280 18230 -10600
rect 19720 -11280 19830 -10600
rect 21320 -11280 21430 -10600
rect 22920 -11280 23030 -10600
rect 24520 -11280 24630 -10600
rect 26120 -11280 26230 -10600
rect 27720 -11280 27830 -10600
rect 29320 -11280 29430 -10600
rect 30920 -11280 31030 -10600
rect 32520 -11110 32630 -10600
rect 34120 -11110 34230 -10600
rect 35720 -11110 35830 -10600
rect 35010 -11430 35130 -11310
rect 1210 -11790 1330 -11670
rect 2810 -11790 2930 -11670
rect 4410 -11790 4530 -11670
rect 6010 -11790 6130 -11670
rect 7610 -11790 7730 -11670
rect 9210 -11790 9330 -11670
rect 13310 -11790 13430 -11670
rect 14230 -11790 14350 -11670
rect 15830 -11790 15950 -11670
rect 17430 -11790 17550 -11670
rect 19030 -11790 19150 -11670
rect 20630 -11790 20750 -11670
rect 22230 -11790 22350 -11670
rect 23830 -11790 23950 -11670
rect 25430 -11790 25550 -11670
rect 27030 -11790 27150 -11670
rect 28630 -11790 28750 -11670
rect 30230 -11790 30350 -11670
rect 31830 -11790 31950 -11670
rect 34810 -11790 34930 -11670
rect 10810 -11980 10930 -11860
rect 1430 -12230 1550 -12110
rect 3030 -12230 3150 -12110
rect 4630 -12230 4750 -12110
rect 6230 -12230 6350 -12110
rect 7830 -12230 7950 -12110
rect 9430 -12230 9550 -12110
rect 14910 -12230 15040 -12100
rect 15610 -12240 15730 -12120
rect 17210 -12240 17330 -12120
rect 18810 -12240 18930 -12120
rect 20410 -12240 20530 -12120
rect 22010 -12240 22130 -12120
rect 23610 -12240 23730 -12120
rect 25210 -12240 25330 -12120
rect 26810 -12240 26930 -12120
rect 28410 -12240 28530 -12120
rect 30010 -12240 30130 -12120
rect 31610 -12240 31730 -12120
rect 2130 -13070 2230 -12410
rect 3730 -13070 3830 -12410
rect 5330 -13070 5430 -12410
rect 6930 -13070 7030 -12410
rect 8530 -13070 8630 -12410
rect 10130 -13070 10230 -12410
rect 11720 -13070 11830 -12410
rect 13320 -13070 13430 -12410
rect 14920 -13070 15030 -12410
rect 16520 -13080 16630 -12400
rect 18120 -13080 18230 -12400
rect 19720 -13080 19830 -12400
rect 21320 -13080 21430 -12400
rect 22920 -13080 23030 -12400
rect 24520 -13080 24630 -12400
rect 26120 -13080 26230 -12400
rect 27720 -13080 27830 -12400
rect 29320 -13080 29430 -12400
rect 30920 -13080 31030 -12400
rect 32520 -12910 32630 -12400
rect 34120 -12910 34230 -12400
rect 35720 -12910 35830 -12400
rect 11270 -13210 11650 -13150
rect 35010 -13230 35130 -13110
rect 1210 -13590 1330 -13470
rect 2810 -13590 2930 -13470
rect 4410 -13590 4530 -13470
rect 6010 -13590 6130 -13470
rect 7610 -13590 7730 -13470
rect 9210 -13590 9330 -13470
rect 14010 -13600 14130 -13480
rect 15830 -13590 15950 -13470
rect 17430 -13590 17550 -13470
rect 19030 -13590 19150 -13470
rect 20630 -13590 20750 -13470
rect 22230 -13590 22350 -13470
rect 23830 -13590 23950 -13470
rect 25430 -13590 25550 -13470
rect 27030 -13590 27150 -13470
rect 28630 -13590 28750 -13470
rect 30230 -13590 30350 -13470
rect 31830 -13590 31950 -13470
rect 34810 -13590 34930 -13470
rect 10810 -13780 10930 -13660
rect 1430 -14030 1550 -13910
rect 3030 -14030 3150 -13910
rect 4630 -14030 4750 -13910
rect 6230 -14030 6350 -13910
rect 7830 -14030 7950 -13910
rect 9430 -14030 9550 -13910
rect 11270 -14120 11650 -14060
rect 15610 -14040 15730 -13920
rect 17210 -14040 17330 -13920
rect 18810 -14040 18930 -13920
rect 20410 -14040 20530 -13920
rect 22010 -14040 22130 -13920
rect 23610 -14040 23730 -13920
rect 25210 -14040 25330 -13920
rect 26810 -14040 26930 -13920
rect 28410 -14040 28530 -13920
rect 30010 -14040 30130 -13920
rect 31610 -14040 31730 -13920
rect 2130 -14870 2230 -14210
rect 3730 -14870 3830 -14210
rect 5330 -14870 5430 -14210
rect 6930 -14870 7030 -14210
rect 8530 -14870 8630 -14210
rect 10130 -14870 10230 -14210
rect 11720 -14870 11830 -14210
rect 13320 -14870 13430 -14210
rect 14920 -14870 15030 -14210
rect 16520 -14880 16630 -14200
rect 18120 -14880 18230 -14200
rect 19720 -14880 19830 -14200
rect 21320 -14880 21430 -14200
rect 22920 -14880 23030 -14200
rect 24520 -14880 24630 -14200
rect 26120 -14880 26230 -14200
rect 27720 -14880 27830 -14200
rect 29320 -14880 29430 -14200
rect 30920 -14880 31030 -14200
rect 32520 -14710 32630 -14200
rect 34120 -14710 34230 -14200
rect 35720 -14710 35830 -14200
rect 35010 -15030 35130 -14910
rect 1210 -15390 1330 -15270
rect 2810 -15390 2930 -15270
rect 4410 -15390 4530 -15270
rect 6010 -15390 6130 -15270
rect 7610 -15390 7730 -15270
rect 9210 -15390 9330 -15270
rect 13330 -15390 13430 -15290
rect 14020 -15410 14120 -15310
rect 14930 -15390 15030 -15290
rect 15830 -15390 15950 -15270
rect 17430 -15390 17550 -15270
rect 19030 -15390 19150 -15270
rect 20630 -15390 20750 -15270
rect 22230 -15390 22350 -15270
rect 23830 -15390 23950 -15270
rect 27030 -15390 27150 -15270
rect 28630 -15390 28750 -15270
rect 31850 -15400 31970 -15280
rect 10810 -15580 10930 -15460
rect 1430 -15830 1550 -15710
rect 3030 -15830 3150 -15710
rect 4630 -15830 4750 -15710
rect 6230 -15830 6350 -15710
rect 7830 -15830 7950 -15710
rect 9430 -15830 9550 -15710
rect 2130 -16670 2230 -16010
rect 3730 -16670 3830 -16010
rect 5330 -16670 5430 -16010
rect 6930 -16670 7030 -16010
rect 8530 -16670 8630 -16010
rect 10130 -16670 10230 -16010
rect 15610 -15840 15730 -15720
rect 17210 -15840 17330 -15720
rect 18810 -15840 18930 -15720
rect 20410 -15840 20530 -15720
rect 22010 -15840 22130 -15720
rect 23610 -15840 23730 -15720
rect 26810 -15840 26930 -15720
rect 28410 -15840 28530 -15720
rect 31590 -15840 31710 -15720
rect 13320 -16670 13430 -16010
rect 14920 -16670 15030 -16010
rect 16520 -16680 16630 -16000
rect 18120 -16680 18230 -16000
rect 19720 -16680 19830 -16000
rect 21320 -16680 21430 -16000
rect 22920 -16680 23030 -16000
rect 24520 -16680 24630 -16000
rect 26120 -16680 26230 -16000
rect 27720 -16680 27830 -16000
rect 29320 -16680 29430 -16000
rect 30920 -16680 31030 -16000
rect 32520 -16680 32630 -16000
rect 34120 -16680 34230 -16000
rect 35720 -16680 35830 -16000
rect 1210 -17190 1330 -17070
rect 2810 -17190 2930 -17070
rect 4410 -17190 4530 -17070
rect 6010 -17190 6130 -17070
rect 7610 -17190 7730 -17070
rect 9210 -17190 9330 -17070
rect 12630 -17200 12750 -17080
rect 15830 -17190 15950 -17070
rect 17430 -17190 17550 -17070
rect 19030 -17190 19150 -17070
rect 20630 -17190 20750 -17070
rect 22230 -17190 22350 -17070
rect 23830 -17190 23950 -17070
rect 27030 -17190 27150 -17070
rect 28630 -17190 28750 -17070
rect 31850 -17200 31970 -17080
rect 10810 -17380 10930 -17260
rect 1430 -17630 1550 -17510
rect 3030 -17630 3150 -17510
rect 4630 -17630 4750 -17510
rect 6230 -17630 6350 -17510
rect 7830 -17630 7950 -17510
rect 9430 -17630 9550 -17510
rect 2130 -18470 2230 -17810
rect 3730 -18470 3830 -17810
rect 5330 -18470 5430 -17810
rect 6930 -18470 7030 -17810
rect 8530 -18470 8630 -17810
rect 10130 -18470 10230 -17810
rect 15610 -17640 15730 -17520
rect 17210 -17640 17330 -17520
rect 18810 -17640 18930 -17520
rect 20410 -17640 20530 -17520
rect 22010 -17640 22130 -17520
rect 23610 -17640 23730 -17520
rect 26810 -17640 26930 -17520
rect 28410 -17640 28530 -17520
rect 31590 -17640 31710 -17520
rect 13320 -18470 13430 -17810
rect 14920 -18470 15030 -17810
rect 16520 -18480 16630 -17800
rect 18120 -18480 18230 -17800
rect 19720 -18480 19830 -17800
rect 21320 -18480 21430 -17800
rect 22920 -18480 23030 -17800
rect 24520 -18480 24630 -17800
rect 26120 -18480 26230 -17800
rect 27720 -18480 27830 -17800
rect 29320 -18480 29430 -17800
rect 30920 -18480 31030 -17800
rect 32520 -18480 32630 -17800
rect 34120 -18480 34230 -17800
rect 35720 -18480 35830 -17800
rect 1210 -18990 1330 -18870
rect 2810 -18990 2930 -18870
rect 4410 -18990 4530 -18870
rect 6010 -18990 6130 -18870
rect 7610 -18990 7730 -18870
rect 9210 -18990 9330 -18870
rect 12410 -19000 12530 -18880
rect 15830 -18990 15950 -18870
rect 17430 -18990 17550 -18870
rect 19030 -18990 19150 -18870
rect 20630 -18990 20750 -18870
rect 22230 -18990 22350 -18870
rect 23830 -18990 23950 -18870
rect 27030 -18990 27150 -18870
rect 28630 -18990 28750 -18870
rect 31590 -19000 31710 -18880
rect 10810 -19180 10930 -19060
rect 1430 -19430 1550 -19310
rect 3030 -19430 3150 -19310
rect 4630 -19430 4750 -19310
rect 6230 -19430 6350 -19310
rect 7830 -19430 7950 -19310
rect 9430 -19430 9550 -19310
rect 2130 -20270 2230 -19610
rect 3730 -20270 3830 -19610
rect 5330 -20270 5430 -19610
rect 6930 -20270 7030 -19610
rect 8530 -20270 8630 -19610
rect 10130 -20270 10230 -19610
rect 15610 -19440 15730 -19320
rect 17210 -19440 17330 -19320
rect 18810 -19440 18930 -19320
rect 20410 -19440 20530 -19320
rect 22010 -19440 22130 -19320
rect 23610 -19440 23730 -19320
rect 26810 -19440 26930 -19320
rect 28410 -19440 28530 -19320
rect 31750 -19520 31810 -19240
rect 13320 -20270 13430 -19610
rect 14920 -20270 15030 -19610
rect 16520 -20280 16630 -19600
rect 18120 -20280 18230 -19600
rect 19720 -20280 19830 -19600
rect 21320 -20280 21430 -19600
rect 22920 -20280 23030 -19600
rect 24520 -20280 24630 -19600
rect 26120 -20280 26230 -19600
rect 27720 -20280 27830 -19600
rect 29320 -20280 29430 -19600
rect 30920 -20280 31030 -19600
rect 32520 -20280 32630 -19600
rect 34120 -20280 34230 -19600
rect 35720 -20280 35830 -19600
rect 33190 -20460 33310 -20340
rect 1210 -20790 1330 -20670
rect 2810 -20790 2930 -20670
rect 4410 -20790 4530 -20670
rect 6010 -20790 6130 -20670
rect 7610 -20790 7730 -20670
rect 9210 -20790 9330 -20670
rect 12410 -20800 12530 -20680
rect 15830 -20790 15950 -20670
rect 17430 -20790 17550 -20670
rect 19030 -20790 19150 -20670
rect 20630 -20790 20750 -20670
rect 22230 -20790 22350 -20670
rect 23830 -20790 23950 -20670
rect 27030 -20790 27150 -20670
rect 28630 -20790 28750 -20670
rect 31590 -20800 31710 -20680
rect 10810 -20980 10930 -20860
rect 1430 -21230 1550 -21110
rect 3030 -21230 3150 -21110
rect 4630 -21230 4750 -21110
rect 6230 -21230 6350 -21110
rect 7830 -21230 7950 -21110
rect 9430 -21230 9550 -21110
rect 15610 -21240 15730 -21120
rect 2130 -22070 2230 -21410
rect 3730 -22070 3830 -21410
rect 5330 -22070 5430 -21410
rect 6930 -22070 7030 -21410
rect 8530 -22070 8630 -21410
rect 10130 -22070 10230 -21410
rect 11710 -22080 11840 -21400
rect 17210 -21240 17330 -21120
rect 18810 -21240 18930 -21120
rect 20410 -21240 20530 -21120
rect 22010 -21240 22130 -21120
rect 23610 -21240 23730 -21120
rect 26810 -21240 26930 -21120
rect 28410 -21240 28530 -21120
rect 31750 -21320 31810 -21040
rect 16520 -22080 16630 -21400
rect 18120 -22080 18230 -21400
rect 19720 -22080 19830 -21400
rect 21320 -22080 21430 -21400
rect 22920 -22080 23030 -21400
rect 24520 -22080 24630 -21400
rect 26120 -22080 26230 -21400
rect 27720 -22080 27830 -21400
rect 29320 -22080 29430 -21400
rect 30920 -22080 31030 -21400
rect 32520 -22080 32630 -21400
rect 34120 -22080 34230 -21400
rect 35720 -22080 35830 -21400
rect 33210 -22240 33290 -22140
rect 34020 -22240 34360 -22170
rect 28150 -22870 28370 -22730
rect 28630 -22870 28740 -22740
rect 29000 -22870 29220 -22730
rect 32630 -22490 33300 -22430
rect 34040 -22490 34310 -22430
rect 32700 -23150 32910 -23070
rect 33020 -23150 33230 -23070
rect 34070 -23160 34300 -23100
rect 29750 -23590 29880 -23520
rect 33410 -23620 33910 -23560
rect 35000 -23620 37020 -23560
rect 33170 -24280 33280 -24220
rect 33410 -24280 33600 -24220
rect 33730 -24280 33920 -24220
rect 34040 -24280 34140 -24220
rect 34620 -24280 34770 -24220
rect 34990 -24280 35130 -24220
rect 35260 -24280 35450 -24220
rect 35570 -24280 35760 -24220
rect 35890 -24280 36080 -24220
rect 36200 -24280 36390 -24220
rect 36520 -24280 36710 -24220
rect 36830 -24280 37020 -24220
rect 2510 -25130 4010 -25070
rect 4710 -25130 6210 -25070
rect 6910 -25130 8410 -25070
rect 9110 -25130 10610 -25070
rect 11310 -25130 12810 -25070
rect 13510 -25130 15010 -25070
rect 15710 -25130 17210 -25070
rect 17910 -25130 19410 -25070
rect 23040 -25070 23560 -24690
rect 4440 -25230 4500 -25170
rect 6640 -25230 6700 -25170
rect 8620 -25230 8680 -25170
rect 10820 -25230 10880 -25170
rect 13020 -25230 13080 -25170
rect 15220 -25230 15280 -25170
rect 17640 -25230 17700 -25170
rect 19840 -25230 19900 -25170
rect 2240 -25320 2300 -25260
rect 4440 -25340 4500 -25280
rect 6420 -25340 6480 -25280
rect 8620 -25340 8680 -25280
rect 10820 -25340 10880 -25280
rect 13020 -25340 13080 -25280
rect 15440 -25340 15500 -25280
rect 17640 -25340 17700 -25280
rect 2510 -25760 2690 -25700
rect 3170 -25760 3350 -25700
rect 3830 -25760 4010 -25700
rect 4710 -25760 4890 -25700
rect 5370 -25760 5550 -25700
rect 6030 -25760 6210 -25700
rect 6910 -25620 7090 -25560
rect 7570 -25620 7750 -25560
rect 8230 -25620 8410 -25560
rect 9110 -25620 9290 -25560
rect 9770 -25620 9950 -25560
rect 10430 -25620 10610 -25560
rect 11310 -25620 11490 -25560
rect 11970 -25620 12150 -25560
rect 12630 -25620 12810 -25560
rect 13510 -25620 13690 -25560
rect 14170 -25620 14350 -25560
rect 14830 -25620 15010 -25560
rect 15710 -25760 15890 -25700
rect 16370 -25760 16550 -25700
rect 17030 -25760 17210 -25700
rect 17910 -25760 18090 -25700
rect 18570 -25760 18750 -25700
rect 34810 -24610 34930 -24490
rect 27260 -25600 27320 -25510
rect 19230 -25760 19410 -25700
rect 27740 -25760 27800 -25670
rect 2510 -25930 4010 -25870
rect 4710 -25930 6210 -25870
rect 6910 -25930 8410 -25870
rect 9110 -25930 10610 -25870
rect 11310 -25930 12810 -25870
rect 13510 -25930 15010 -25870
rect 15710 -25930 17210 -25870
rect 17910 -25930 19410 -25870
rect 27260 -25920 27320 -25830
rect 4220 -26030 4280 -25970
rect 6420 -26030 6480 -25970
rect 8840 -26030 8900 -25970
rect 11040 -26030 11100 -25970
rect 13240 -26030 13300 -25970
rect 15440 -26030 15500 -25970
rect 17420 -26030 17480 -25970
rect 19620 -26030 19680 -25970
rect 2020 -26120 2080 -26060
rect 27740 -26075 27800 -25985
rect 29380 -25970 29440 -25770
rect 4220 -26140 4280 -26080
rect 6640 -26140 6700 -26080
rect 8840 -26140 8900 -26080
rect 11040 -26140 11100 -26080
rect 13240 -26140 13300 -26080
rect 15220 -26140 15280 -26080
rect 17420 -26140 17480 -26080
rect 27260 -26235 27320 -26145
rect 2510 -26420 2690 -26360
rect 3170 -26420 3350 -26360
rect 3830 -26420 4010 -26360
rect 4710 -26420 4890 -26360
rect 5370 -26420 5550 -26360
rect 6030 -26420 6210 -26360
rect 6910 -26560 7090 -26500
rect 7570 -26560 7750 -26500
rect 8230 -26560 8410 -26500
rect 9110 -26560 9290 -26500
rect 9770 -26560 9950 -26500
rect 10430 -26560 10610 -26500
rect 11310 -26560 11490 -26500
rect 11970 -26560 12150 -26500
rect 12630 -26560 12810 -26500
rect 13510 -26560 13690 -26500
rect 14170 -26560 14350 -26500
rect 14830 -26560 15010 -26500
rect 15710 -26420 15890 -26360
rect 16370 -26420 16550 -26360
rect 17030 -26420 17210 -26360
rect 17910 -26420 18090 -26360
rect 18570 -26420 18750 -26360
rect 19230 -26420 19410 -26360
rect 430 -26710 610 -26630
rect 4710 -26730 6210 -26670
rect 6910 -26730 8410 -26670
rect 9110 -26730 10610 -26670
rect 11310 -26730 12810 -26670
rect 13510 -26730 15010 -26670
rect 15710 -26730 17210 -26670
rect 21310 -26710 21490 -26630
rect 27740 -26640 27800 -26550
rect 6640 -26830 6700 -26770
rect 8620 -26830 8680 -26770
rect 10820 -26830 10880 -26770
rect 13020 -26830 13080 -26770
rect 15220 -26830 15280 -26770
rect 17640 -26830 17700 -26770
rect 1420 -27020 1480 -26870
rect 4440 -26940 4500 -26880
rect 6420 -26940 6480 -26880
rect 8620 -26940 8680 -26880
rect 10820 -26940 10880 -26880
rect 13020 -26940 13080 -26880
rect 15440 -26940 15500 -26880
rect 20240 -26930 20300 -26780
rect 27380 -26800 27440 -26710
rect 27740 -26960 27800 -26870
rect 2510 -27360 2690 -27300
rect 3170 -27360 3350 -27300
rect 3830 -27360 4010 -27300
rect 4710 -27360 4890 -27300
rect 5370 -27360 5550 -27300
rect 6030 -27360 6210 -27300
rect 6910 -27220 7090 -27160
rect 7570 -27220 7750 -27160
rect 8230 -27220 8410 -27160
rect 9110 -27220 9290 -27160
rect 9770 -27220 9950 -27160
rect 10430 -27220 10610 -27160
rect 11310 -27220 11490 -27160
rect 11970 -27220 12150 -27160
rect 12630 -27220 12810 -27160
rect 13510 -27220 13690 -27160
rect 14170 -27220 14350 -27160
rect 14830 -27220 15010 -27160
rect 15710 -27360 15890 -27300
rect 16370 -27360 16550 -27300
rect 17030 -27360 17210 -27300
rect 17910 -27360 18090 -27300
rect 18570 -27360 18750 -27300
rect 27380 -27115 27440 -27025
rect 29530 -27010 29590 -26810
rect 27740 -27275 27800 -27185
rect 19230 -27360 19410 -27300
rect 34810 -25010 34900 -24940
rect 37190 -25010 37280 -24940
rect 34810 -25270 34900 -25200
rect 34810 -25530 34900 -25460
rect 37190 -25270 37280 -25200
rect 37190 -25530 37280 -25460
rect 34810 -25790 34900 -25720
rect 34810 -26050 34900 -25980
rect 37190 -25790 37280 -25720
rect 37190 -26050 37280 -25980
rect 34810 -26310 34900 -26240
rect 34810 -26570 34900 -26500
rect 37190 -26310 37280 -26240
rect 37190 -26570 37280 -26500
rect 34810 -26830 34900 -26760
rect 37190 -26830 37280 -26760
rect 36030 -27140 36410 -27010
rect 36530 -27140 36910 -27010
rect 430 -27510 610 -27430
rect 4710 -27530 6210 -27470
rect 6910 -27530 8410 -27470
rect 9110 -27530 10610 -27470
rect 11310 -27530 12810 -27470
rect 13510 -27530 15010 -27470
rect 15710 -27530 17210 -27470
rect 21310 -27510 21490 -27430
rect 6420 -27630 6480 -27570
rect 8840 -27630 8900 -27570
rect 11040 -27630 11100 -27570
rect 13240 -27630 13300 -27570
rect 15440 -27630 15500 -27570
rect 17420 -27630 17480 -27570
rect 1620 -27820 1680 -27670
rect 4220 -27740 4280 -27680
rect 6640 -27740 6700 -27680
rect 8840 -27740 8900 -27680
rect 11040 -27740 11100 -27680
rect 13240 -27740 13300 -27680
rect 15220 -27740 15280 -27680
rect 20440 -27730 20500 -27580
rect 27260 -27685 27320 -27595
rect 27500 -27840 27560 -27750
rect 2510 -28020 2690 -27960
rect 3170 -28020 3350 -27960
rect 3830 -28020 4010 -27960
rect 4710 -28020 4890 -27960
rect 5370 -28020 5550 -27960
rect 6030 -28020 6210 -27960
rect 6910 -28160 7090 -28100
rect 7570 -28160 7750 -28100
rect 8230 -28160 8410 -28100
rect 9110 -28160 9290 -28100
rect 9770 -28160 9950 -28100
rect 10430 -28160 10610 -28100
rect 11310 -28160 11490 -28100
rect 11970 -28160 12150 -28100
rect 12630 -28160 12810 -28100
rect 13510 -28160 13690 -28100
rect 14170 -28160 14350 -28100
rect 14830 -28160 15010 -28100
rect 15710 -28020 15890 -27960
rect 16370 -28020 16550 -27960
rect 17030 -28020 17210 -27960
rect 17910 -28020 18090 -27960
rect 18570 -28020 18750 -27960
rect 19230 -28020 19410 -27960
rect 27260 -28000 27320 -27910
rect 27500 -28155 27560 -28065
rect 29080 -28050 29140 -27850
rect 36920 -27900 37680 -27540
rect 430 -28310 610 -28230
rect 4710 -28330 6210 -28270
rect 6910 -28330 8410 -28270
rect 9110 -28330 10610 -28270
rect 11310 -28330 12810 -28270
rect 13510 -28330 15010 -28270
rect 15710 -28330 17210 -28270
rect 21310 -28310 21490 -28230
rect 27260 -28315 27320 -28225
rect 6420 -28430 6480 -28370
rect 8840 -28430 8900 -28370
rect 11040 -28430 11100 -28370
rect 13240 -28430 13300 -28370
rect 15440 -28430 15500 -28370
rect 17420 -28430 17480 -28370
rect 1620 -28620 1680 -28470
rect 4220 -28540 4280 -28480
rect 6640 -28540 6700 -28480
rect 8840 -28540 8900 -28480
rect 11040 -28540 11100 -28480
rect 13240 -28540 13300 -28480
rect 15220 -28540 15280 -28480
rect 20440 -28530 20500 -28380
rect 36920 -28520 37680 -28160
rect 2510 -28820 2690 -28760
rect 3170 -28820 3350 -28760
rect 3830 -28820 4010 -28760
rect 4710 -28820 4890 -28760
rect 5370 -28820 5550 -28760
rect 6030 -28820 6210 -28760
rect 6910 -28960 7090 -28900
rect 7570 -28960 7750 -28900
rect 8230 -28960 8410 -28900
rect 9110 -28960 9290 -28900
rect 9770 -28960 9950 -28900
rect 10430 -28960 10610 -28900
rect 11310 -28960 11490 -28900
rect 11970 -28960 12150 -28900
rect 12630 -28960 12810 -28900
rect 13510 -28960 13690 -28900
rect 14170 -28960 14350 -28900
rect 14830 -28960 15010 -28900
rect 15710 -28820 15890 -28760
rect 16370 -28820 16550 -28760
rect 17030 -28820 17210 -28760
rect 17910 -28820 18090 -28760
rect 18570 -28820 18750 -28760
rect 27260 -28720 27320 -28630
rect 19230 -28820 19410 -28760
rect 27620 -28880 27680 -28790
rect 430 -29110 610 -29030
rect 4710 -29130 6210 -29070
rect 6910 -29130 8410 -29070
rect 9110 -29130 10610 -29070
rect 11310 -29130 12810 -29070
rect 13510 -29130 15010 -29070
rect 15710 -29130 17210 -29070
rect 21310 -29110 21490 -29030
rect 27260 -29040 27320 -28950
rect 6640 -29230 6700 -29170
rect 8620 -29230 8680 -29170
rect 10820 -29230 10880 -29170
rect 13020 -29230 13080 -29170
rect 15220 -29230 15280 -29170
rect 17640 -29230 17700 -29170
rect 1420 -29420 1480 -29270
rect 4440 -29340 4500 -29280
rect 6420 -29340 6480 -29280
rect 8620 -29340 8680 -29280
rect 10820 -29340 10880 -29280
rect 13020 -29340 13080 -29280
rect 15440 -29340 15500 -29280
rect 20240 -29330 20300 -29180
rect 27620 -29200 27680 -29110
rect 29230 -29090 29290 -28890
rect 27260 -29350 27320 -29260
rect 2510 -29760 2690 -29700
rect 3170 -29760 3350 -29700
rect 3830 -29760 4010 -29700
rect 4710 -29760 4890 -29700
rect 5370 -29760 5550 -29700
rect 6030 -29760 6210 -29700
rect 6910 -29620 7090 -29560
rect 7570 -29620 7750 -29560
rect 8230 -29620 8410 -29560
rect 9110 -29620 9290 -29560
rect 9770 -29620 9950 -29560
rect 10430 -29620 10610 -29560
rect 11310 -29620 11490 -29560
rect 11970 -29620 12150 -29560
rect 12630 -29620 12810 -29560
rect 13510 -29620 13690 -29560
rect 14170 -29620 14350 -29560
rect 14830 -29620 15010 -29560
rect 15710 -29760 15890 -29700
rect 16370 -29760 16550 -29700
rect 17030 -29760 17210 -29700
rect 17910 -29760 18090 -29700
rect 18570 -29760 18750 -29700
rect 19230 -29760 19410 -29700
rect 27380 -29760 27440 -29670
rect 2510 -29930 4010 -29870
rect 4710 -29930 6210 -29870
rect 6910 -29930 8410 -29870
rect 9110 -29930 10610 -29870
rect 11310 -29930 12810 -29870
rect 13510 -29930 15010 -29870
rect 15710 -29930 17210 -29870
rect 17910 -29930 19410 -29870
rect 27620 -29920 27680 -29830
rect 4220 -30030 4280 -29970
rect 6420 -30030 6480 -29970
rect 8840 -30030 8900 -29970
rect 11040 -30030 11100 -29970
rect 13240 -30030 13300 -29970
rect 15440 -30030 15500 -29970
rect 17420 -30030 17480 -29970
rect 19620 -30030 19680 -29970
rect 2020 -30120 2080 -30060
rect 27380 -30075 27440 -29985
rect 4220 -30140 4280 -30080
rect 6640 -30140 6700 -30080
rect 8840 -30140 8900 -30080
rect 11040 -30140 11100 -30080
rect 13240 -30140 13300 -30080
rect 15220 -30140 15280 -30080
rect 17420 -30140 17480 -30080
rect 27620 -30235 27680 -30145
rect 29080 -30130 29140 -29930
rect 2510 -30420 2690 -30360
rect 3170 -30420 3350 -30360
rect 3830 -30420 4010 -30360
rect 4710 -30420 4890 -30360
rect 5370 -30420 5550 -30360
rect 6030 -30420 6210 -30360
rect 6910 -30560 7090 -30500
rect 7570 -30560 7750 -30500
rect 8230 -30560 8410 -30500
rect 9110 -30560 9290 -30500
rect 9770 -30560 9950 -30500
rect 10430 -30560 10610 -30500
rect 11310 -30560 11490 -30500
rect 11970 -30560 12150 -30500
rect 12630 -30560 12810 -30500
rect 13510 -30560 13690 -30500
rect 14170 -30560 14350 -30500
rect 14830 -30560 15010 -30500
rect 15710 -30420 15890 -30360
rect 16370 -30420 16550 -30360
rect 17030 -30420 17210 -30360
rect 17910 -30420 18090 -30360
rect 18570 -30420 18750 -30360
rect 19230 -30420 19410 -30360
rect 27380 -30390 27440 -30300
rect 2510 -30730 4010 -30670
rect 4710 -30730 6210 -30670
rect 6910 -30730 8410 -30670
rect 9110 -30730 10610 -30670
rect 11310 -30730 12810 -30670
rect 13510 -30730 15010 -30670
rect 15710 -30730 17210 -30670
rect 17910 -30730 19410 -30670
rect 4440 -30830 4500 -30770
rect 6640 -30830 6700 -30770
rect 8620 -30830 8680 -30770
rect 10820 -30830 10880 -30770
rect 13020 -30830 13080 -30770
rect 15220 -30830 15280 -30770
rect 17640 -30830 17700 -30770
rect 19840 -30830 19900 -30770
rect 27380 -30800 27440 -30710
rect 2240 -30920 2300 -30860
rect 4440 -30940 4500 -30880
rect 6420 -30940 6480 -30880
rect 8620 -30940 8680 -30880
rect 10820 -30940 10880 -30880
rect 13020 -30940 13080 -30880
rect 15440 -30940 15500 -30880
rect 17640 -30940 17700 -30880
rect 27500 -30960 27560 -30870
rect 2510 -31360 2690 -31300
rect 3170 -31360 3350 -31300
rect 3830 -31360 4010 -31300
rect 4710 -31360 4890 -31300
rect 5370 -31360 5550 -31300
rect 6030 -31360 6210 -31300
rect 6910 -31220 7090 -31160
rect 7570 -31220 7750 -31160
rect 8230 -31220 8410 -31160
rect 9110 -31220 9290 -31160
rect 9770 -31220 9950 -31160
rect 10430 -31220 10610 -31160
rect 11310 -31220 11490 -31160
rect 11970 -31220 12150 -31160
rect 12630 -31220 12810 -31160
rect 13510 -31220 13690 -31160
rect 14170 -31220 14350 -31160
rect 14830 -31220 15010 -31160
rect 15710 -31360 15890 -31300
rect 16370 -31360 16550 -31300
rect 17030 -31360 17210 -31300
rect 17910 -31360 18090 -31300
rect 18570 -31360 18750 -31300
rect 27380 -31115 27440 -31025
rect 29070 -31030 29290 -30960
rect 27500 -31275 27560 -31185
rect 19230 -31360 19410 -31300
rect 27380 -31430 27440 -31340
rect 25700 -31880 26220 -31510
rect 32794 -30488 32846 -30336
rect 33126 -30494 33178 -30342
rect 33794 -30488 33846 -30336
rect 34126 -30494 34178 -30342
rect 34794 -30488 34846 -30336
rect 35126 -30494 35178 -30342
rect 35794 -30488 35846 -30336
rect 36126 -30494 36178 -30342
rect 36794 -30488 36846 -30336
rect 37126 -30494 37178 -30342
rect 37794 -30488 37846 -30336
rect 38126 -30494 38178 -30342
rect 38410 -30730 38588 -30154
rect 30840 -32440 31240 -31680
rect 38406 -32314 38520 -32180
rect 38320 -32690 38520 -32314
rect 38310 -32910 38530 -32690
<< metal2 >>
rect -360 11990 -160 12000
rect -360 11610 -350 11990
rect -170 11610 -160 11990
rect 2020 11720 2080 12020
rect 2200 12010 2340 12020
rect 2200 11890 2210 12010
rect 2330 11890 2340 12010
rect 2200 11880 2340 11890
rect 1980 11710 2120 11720
rect -360 -6590 -160 11610
rect 80 11690 280 11700
rect 80 11310 90 11690
rect 270 11310 280 11690
rect 1980 11590 1990 11710
rect 2110 11590 2120 11710
rect 1980 11580 2120 11590
rect -70 10930 -10 10940
rect -70 10860 -10 10870
rect -70 10130 -10 10140
rect -70 10060 -10 10070
rect -70 9330 -10 9340
rect -70 9260 -10 9270
rect -70 8530 -10 8540
rect -70 8460 -10 8470
rect -70 7730 -10 7740
rect -70 7660 -10 7670
rect -70 6930 -10 6940
rect -70 6860 -10 6870
rect -70 6130 -10 6140
rect -70 6060 -10 6070
rect -70 5330 -10 5340
rect -70 5260 -10 5270
rect -360 -7170 -350 -6590
rect -170 -7170 -160 -6590
rect -360 -31450 -160 -7170
rect -360 -31830 -350 -31450
rect -170 -31830 -160 -31450
rect -360 -32120 -160 -31830
rect 80 -5750 280 11310
rect 2020 10830 2080 11580
rect 2130 10930 2190 10940
rect 2130 10860 2190 10870
rect 2240 10830 2300 11880
rect 4220 11720 4280 12020
rect 4400 12010 4540 12020
rect 4400 11890 4410 12010
rect 4530 11890 4540 12010
rect 4400 11880 4540 11890
rect 4180 11710 4320 11720
rect 4180 11590 4190 11710
rect 4310 11590 4320 11710
rect 4180 11580 4320 11590
rect 2500 11240 2700 11250
rect 2500 11180 2510 11240
rect 2690 11180 2700 11240
rect 2500 11170 2700 11180
rect 3160 11240 3360 11250
rect 3160 11180 3170 11240
rect 3350 11180 3360 11240
rect 3160 11170 3360 11180
rect 3820 11240 4020 11250
rect 3820 11180 3830 11240
rect 4010 11180 4020 11240
rect 3820 11170 4020 11180
rect 2500 11030 2700 11110
rect 3160 11030 3360 11110
rect 3820 11030 4020 11110
rect 4220 10830 4280 11580
rect 4330 10930 4390 10940
rect 4330 10860 4390 10870
rect 4440 10830 4500 11880
rect 6420 11720 6480 12020
rect 6600 12010 6740 12020
rect 6600 11890 6610 12010
rect 6730 11890 6740 12010
rect 6600 11880 6740 11890
rect 6380 11710 6520 11720
rect 6380 11590 6390 11710
rect 6510 11590 6520 11710
rect 6380 11580 6520 11590
rect 4700 11240 4900 11250
rect 4700 11180 4710 11240
rect 4890 11180 4900 11240
rect 4700 11170 4900 11180
rect 5360 11240 5560 11250
rect 5360 11180 5370 11240
rect 5550 11180 5560 11240
rect 5360 11170 5560 11180
rect 6020 11240 6220 11250
rect 6020 11180 6030 11240
rect 6210 11180 6220 11240
rect 6020 11170 6220 11180
rect 4700 11030 4900 11110
rect 5360 11030 5560 11110
rect 6020 11030 6220 11110
rect 6420 10830 6480 11580
rect 6530 10930 6590 10940
rect 6530 10860 6590 10870
rect 6640 10830 6700 11880
rect 8620 11720 8680 12020
rect 8800 12010 8940 12020
rect 8800 11890 8810 12010
rect 8930 11890 8940 12010
rect 8800 11880 8940 11890
rect 8580 11710 8720 11720
rect 8580 11590 8590 11710
rect 8710 11590 8720 11710
rect 8580 11580 8720 11590
rect 6900 11170 7100 11250
rect 7560 11170 7760 11250
rect 8220 11170 8420 11250
rect 6900 11100 7100 11110
rect 6900 11040 6910 11100
rect 7090 11040 7100 11100
rect 6900 11030 7100 11040
rect 7560 11100 7760 11110
rect 7560 11040 7570 11100
rect 7750 11040 7760 11100
rect 7560 11030 7760 11040
rect 8220 11100 8420 11110
rect 8220 11040 8230 11100
rect 8410 11040 8420 11100
rect 8220 11030 8420 11040
rect 8620 10830 8680 11580
rect 8730 10930 8790 10940
rect 8730 10860 8790 10870
rect 8840 10830 8900 11880
rect 10820 11720 10880 12020
rect 11000 12010 11140 12020
rect 11000 11890 11010 12010
rect 11130 11890 11140 12010
rect 11000 11880 11140 11890
rect 10780 11710 10920 11720
rect 10780 11590 10790 11710
rect 10910 11590 10920 11710
rect 10780 11580 10920 11590
rect 9100 11170 9300 11250
rect 9760 11170 9960 11250
rect 10420 11170 10620 11250
rect 9100 11100 9300 11110
rect 9100 11040 9110 11100
rect 9290 11040 9300 11100
rect 9100 11030 9300 11040
rect 9760 11100 9960 11110
rect 9760 11040 9770 11100
rect 9950 11040 9960 11100
rect 9760 11030 9960 11040
rect 10420 11100 10620 11110
rect 10420 11040 10430 11100
rect 10610 11040 10620 11100
rect 10420 11030 10620 11040
rect 10820 10830 10880 11580
rect 10930 10930 10990 10940
rect 10930 10860 10990 10870
rect 11040 10830 11100 11880
rect 13020 11720 13080 12020
rect 13200 12010 13340 12020
rect 13200 11890 13210 12010
rect 13330 11890 13340 12010
rect 13200 11880 13340 11890
rect 12980 11710 13120 11720
rect 12980 11590 12990 11710
rect 13110 11590 13120 11710
rect 12980 11580 13120 11590
rect 11300 11170 11500 11250
rect 11960 11170 12160 11250
rect 12620 11170 12820 11250
rect 11300 11100 11500 11110
rect 11300 11040 11310 11100
rect 11490 11040 11500 11100
rect 11300 11030 11500 11040
rect 11960 11100 12160 11110
rect 11960 11040 11970 11100
rect 12150 11040 12160 11100
rect 11960 11030 12160 11040
rect 12620 11100 12820 11110
rect 12620 11040 12630 11100
rect 12810 11040 12820 11100
rect 12620 11030 12820 11040
rect 13020 10830 13080 11580
rect 13130 10930 13190 10940
rect 13130 10860 13190 10870
rect 13240 10830 13300 11880
rect 15220 11720 15280 12020
rect 15400 12010 15540 12020
rect 15400 11890 15410 12010
rect 15530 11890 15540 12010
rect 15400 11880 15540 11890
rect 15180 11710 15320 11720
rect 15180 11590 15190 11710
rect 15310 11590 15320 11710
rect 15180 11580 15320 11590
rect 13500 11170 13700 11250
rect 14160 11170 14360 11250
rect 14820 11170 15020 11250
rect 13500 11100 13700 11110
rect 13500 11040 13510 11100
rect 13690 11040 13700 11100
rect 13500 11030 13700 11040
rect 14160 11100 14360 11110
rect 14160 11040 14170 11100
rect 14350 11040 14360 11100
rect 14160 11030 14360 11040
rect 14820 11100 15020 11110
rect 14820 11040 14830 11100
rect 15010 11040 15020 11100
rect 14820 11030 15020 11040
rect 15220 10830 15280 11580
rect 15330 10930 15390 10940
rect 15330 10860 15390 10870
rect 15440 10830 15500 11880
rect 17420 11720 17480 12020
rect 17600 12010 17740 12020
rect 17600 11890 17610 12010
rect 17730 11890 17740 12010
rect 17600 11880 17740 11890
rect 17380 11710 17520 11720
rect 17380 11590 17390 11710
rect 17510 11590 17520 11710
rect 17380 11580 17520 11590
rect 15700 11240 15900 11250
rect 15700 11180 15710 11240
rect 15890 11180 15900 11240
rect 15700 11170 15900 11180
rect 16360 11240 16560 11250
rect 16360 11180 16370 11240
rect 16550 11180 16560 11240
rect 16360 11170 16560 11180
rect 17020 11240 17220 11250
rect 17020 11180 17030 11240
rect 17210 11180 17220 11240
rect 17020 11170 17220 11180
rect 15700 11030 15900 11110
rect 16360 11030 16560 11110
rect 17020 11030 17220 11110
rect 17420 10830 17480 11580
rect 17530 10930 17590 10940
rect 17530 10860 17590 10870
rect 17640 10830 17700 11880
rect 19620 11720 19680 12020
rect 19800 12010 19940 12020
rect 19800 11890 19810 12010
rect 19930 11890 19940 12010
rect 31400 11959 31490 13400
rect 32200 11937 32290 13400
rect 33000 11943 33090 13400
rect 36900 12540 38300 12560
rect 36900 12280 36920 12540
rect 38280 12280 38300 12540
rect 36900 12260 38300 12280
rect 36930 12030 37080 12040
rect 19800 11880 19940 11890
rect 19580 11710 19720 11720
rect 19580 11590 19590 11710
rect 19710 11590 19720 11710
rect 19580 11580 19720 11590
rect 17900 11240 18100 11250
rect 17900 11180 17910 11240
rect 18090 11180 18100 11240
rect 17900 11170 18100 11180
rect 18560 11240 18760 11250
rect 18560 11180 18570 11240
rect 18750 11180 18760 11240
rect 18560 11170 18760 11180
rect 19220 11240 19420 11250
rect 19220 11180 19230 11240
rect 19410 11180 19420 11240
rect 19220 11170 19420 11180
rect 17900 11030 18100 11110
rect 18560 11030 18760 11110
rect 19220 11030 19420 11110
rect 2010 10710 2090 10830
rect 2010 10650 2020 10710
rect 2080 10650 2090 10710
rect 2010 10640 2090 10650
rect 2230 10640 2310 10830
rect 4210 10820 4290 10830
rect 4210 10760 4220 10820
rect 4280 10760 4290 10820
rect 4210 10710 4290 10760
rect 4210 10650 4220 10710
rect 4280 10650 4290 10710
rect 4210 10640 4290 10650
rect 4430 10640 4510 10830
rect 6410 10820 6490 10830
rect 6410 10760 6420 10820
rect 6480 10760 6490 10820
rect 6410 10640 6490 10760
rect 6630 10710 6710 10830
rect 6630 10650 6640 10710
rect 6700 10650 6710 10710
rect 6630 10640 6710 10650
rect 8610 10640 8690 10830
rect 8830 10820 8910 10830
rect 8830 10760 8840 10820
rect 8900 10760 8910 10820
rect 8830 10710 8910 10760
rect 8830 10650 8840 10710
rect 8900 10650 8910 10710
rect 8830 10640 8910 10650
rect 10810 10640 10890 10830
rect 11030 10820 11110 10830
rect 11030 10760 11040 10820
rect 11100 10760 11110 10820
rect 11030 10710 11110 10760
rect 11030 10650 11040 10710
rect 11100 10650 11110 10710
rect 11030 10640 11110 10650
rect 13010 10640 13090 10830
rect 13230 10820 13310 10830
rect 13230 10760 13240 10820
rect 13300 10760 13310 10820
rect 13230 10710 13310 10760
rect 13230 10650 13240 10710
rect 13300 10650 13310 10710
rect 13230 10640 13310 10650
rect 15210 10710 15290 10830
rect 15210 10650 15220 10710
rect 15280 10650 15290 10710
rect 15210 10640 15290 10650
rect 15430 10820 15510 10830
rect 15430 10760 15440 10820
rect 15500 10760 15510 10820
rect 15430 10640 15510 10760
rect 17410 10820 17490 10830
rect 17410 10760 17420 10820
rect 17480 10760 17490 10820
rect 17410 10710 17490 10760
rect 17410 10650 17420 10710
rect 17480 10650 17490 10710
rect 17410 10640 17490 10650
rect 17630 10640 17710 10830
rect 19620 10810 19680 11580
rect 19730 10930 19790 10940
rect 19730 10860 19790 10870
rect 19840 10810 19900 11880
rect 36930 11850 36940 12030
rect 37070 11850 37080 12030
rect 36930 11840 37080 11850
rect 37350 12030 37500 12040
rect 37350 11850 37360 12030
rect 37490 11850 37500 12030
rect 37350 11840 37500 11850
rect 37770 12030 37920 12040
rect 37770 11850 37780 12030
rect 37910 11850 37920 12030
rect 37770 11840 37920 11850
rect 25710 11780 26250 11790
rect 25710 11410 25720 11780
rect 26240 11690 26250 11780
rect 36990 11690 37050 11840
rect 37410 11690 37470 11840
rect 37830 11690 37890 11840
rect 26240 11500 27320 11690
rect 36980 11680 37060 11690
rect 26240 11490 27330 11500
rect 26240 11410 26250 11490
rect 25710 11400 26250 11410
rect 21930 10930 21990 10940
rect 21930 10860 21990 10870
rect 19610 10800 19690 10810
rect 19610 10740 19620 10800
rect 19680 10740 19690 10800
rect 19610 10640 19690 10740
rect 19830 10640 19910 10810
rect 2020 10030 2080 10640
rect 2130 10130 2190 10140
rect 2130 10060 2190 10070
rect 2240 10030 2300 10640
rect 2500 10610 4020 10620
rect 2500 10550 2510 10610
rect 4010 10550 4020 10610
rect 2500 10540 4020 10550
rect 2500 10370 2700 10450
rect 3160 10370 3360 10450
rect 3820 10370 4020 10450
rect 2500 10300 2700 10310
rect 2500 10240 2510 10300
rect 2690 10240 2700 10300
rect 2500 10230 2700 10240
rect 3160 10300 3360 10310
rect 3160 10240 3170 10300
rect 3350 10240 3360 10300
rect 3160 10230 3360 10240
rect 3820 10300 4020 10310
rect 3820 10240 3830 10300
rect 4010 10240 4020 10300
rect 3820 10230 4020 10240
rect 4220 10030 4280 10640
rect 4330 10130 4390 10140
rect 4330 10060 4390 10070
rect 4440 10030 4500 10640
rect 4700 10610 6220 10620
rect 4700 10550 4710 10610
rect 6210 10550 6220 10610
rect 4700 10540 6220 10550
rect 4700 10370 4900 10450
rect 5360 10370 5560 10450
rect 6020 10370 6220 10450
rect 4700 10300 4900 10310
rect 4700 10240 4710 10300
rect 4890 10240 4900 10300
rect 4700 10230 4900 10240
rect 5360 10300 5560 10310
rect 5360 10240 5370 10300
rect 5550 10240 5560 10300
rect 5360 10230 5560 10240
rect 6020 10300 6220 10310
rect 6020 10240 6030 10300
rect 6210 10240 6220 10300
rect 6020 10230 6220 10240
rect 6420 10030 6480 10640
rect 6530 10130 6590 10140
rect 6530 10060 6590 10070
rect 6640 10030 6700 10640
rect 6900 10610 8420 10620
rect 6900 10550 6910 10610
rect 8410 10550 8420 10610
rect 6900 10540 8420 10550
rect 6900 10440 7100 10450
rect 6900 10380 6910 10440
rect 7090 10380 7100 10440
rect 6900 10370 7100 10380
rect 7560 10440 7760 10450
rect 7560 10380 7570 10440
rect 7750 10380 7760 10440
rect 7560 10370 7760 10380
rect 8220 10440 8420 10450
rect 8220 10380 8230 10440
rect 8410 10380 8420 10440
rect 8220 10370 8420 10380
rect 6900 10230 7100 10310
rect 7560 10230 7760 10310
rect 8220 10230 8420 10310
rect 8620 10030 8680 10640
rect 8730 10130 8790 10140
rect 8730 10060 8790 10070
rect 8840 10030 8900 10640
rect 9100 10610 10620 10620
rect 9100 10550 9110 10610
rect 10610 10550 10620 10610
rect 9100 10540 10620 10550
rect 9100 10440 9300 10450
rect 9100 10380 9110 10440
rect 9290 10380 9300 10440
rect 9100 10370 9300 10380
rect 9760 10440 9960 10450
rect 9760 10380 9770 10440
rect 9950 10380 9960 10440
rect 9760 10370 9960 10380
rect 10420 10440 10620 10450
rect 10420 10380 10430 10440
rect 10610 10380 10620 10440
rect 10420 10370 10620 10380
rect 9100 10230 9300 10310
rect 9760 10230 9960 10310
rect 10420 10230 10620 10310
rect 10820 10030 10880 10640
rect 10930 10130 10990 10140
rect 10930 10060 10990 10070
rect 11040 10030 11100 10640
rect 11300 10610 12820 10620
rect 11300 10550 11310 10610
rect 12810 10550 12820 10610
rect 11300 10540 12820 10550
rect 11300 10440 11500 10450
rect 11300 10380 11310 10440
rect 11490 10380 11500 10440
rect 11300 10370 11500 10380
rect 11960 10440 12160 10450
rect 11960 10380 11970 10440
rect 12150 10380 12160 10440
rect 11960 10370 12160 10380
rect 12620 10440 12820 10450
rect 12620 10380 12630 10440
rect 12810 10380 12820 10440
rect 12620 10370 12820 10380
rect 11300 10230 11500 10310
rect 11960 10230 12160 10310
rect 12620 10230 12820 10310
rect 13020 10030 13080 10640
rect 13130 10130 13190 10140
rect 13130 10060 13190 10070
rect 13240 10030 13300 10640
rect 13500 10610 15020 10620
rect 13500 10550 13510 10610
rect 15010 10550 15020 10610
rect 13500 10540 15020 10550
rect 13500 10440 13700 10450
rect 13500 10380 13510 10440
rect 13690 10380 13700 10440
rect 13500 10370 13700 10380
rect 14160 10440 14360 10450
rect 14160 10380 14170 10440
rect 14350 10380 14360 10440
rect 14160 10370 14360 10380
rect 14820 10440 15020 10450
rect 14820 10380 14830 10440
rect 15010 10380 15020 10440
rect 14820 10370 15020 10380
rect 13500 10230 13700 10310
rect 14160 10230 14360 10310
rect 14820 10230 15020 10310
rect 15220 10030 15280 10640
rect 15330 10130 15390 10140
rect 15330 10060 15390 10070
rect 15440 10030 15500 10640
rect 15700 10610 17220 10620
rect 15700 10550 15710 10610
rect 17210 10550 17220 10610
rect 15700 10540 17220 10550
rect 15700 10370 15900 10450
rect 16360 10370 16560 10450
rect 17020 10370 17220 10450
rect 15700 10300 15900 10310
rect 15700 10240 15710 10300
rect 15890 10240 15900 10300
rect 15700 10230 15900 10240
rect 16360 10300 16560 10310
rect 16360 10240 16370 10300
rect 16550 10240 16560 10300
rect 16360 10230 16560 10240
rect 17020 10300 17220 10310
rect 17020 10240 17030 10300
rect 17210 10240 17220 10300
rect 17020 10230 17220 10240
rect 17420 10030 17480 10640
rect 17530 10130 17590 10140
rect 17530 10060 17590 10070
rect 17640 10030 17700 10640
rect 17900 10610 19420 10620
rect 17900 10550 17910 10610
rect 19410 10550 19420 10610
rect 17900 10540 19420 10550
rect 17900 10370 18100 10450
rect 18560 10370 18760 10450
rect 19220 10370 19420 10450
rect 17900 10300 18100 10310
rect 17900 10240 17910 10300
rect 18090 10240 18100 10300
rect 17900 10230 18100 10240
rect 18560 10300 18760 10310
rect 18560 10240 18570 10300
rect 18750 10240 18760 10300
rect 18560 10230 18760 10240
rect 19220 10300 19420 10310
rect 19220 10240 19230 10300
rect 19410 10240 19420 10300
rect 19220 10230 19420 10240
rect 2010 9840 2090 10030
rect 2230 9910 2310 10030
rect 2230 9850 2240 9910
rect 2300 9850 2310 9910
rect 2230 9840 2310 9850
rect 4210 9840 4290 10030
rect 4430 10020 4510 10030
rect 4430 9960 4440 10020
rect 4500 9960 4510 10020
rect 4430 9910 4510 9960
rect 4430 9850 4440 9910
rect 4500 9850 4510 9910
rect 4430 9840 4510 9850
rect 6410 9910 6490 10030
rect 6410 9850 6420 9910
rect 6480 9850 6490 9910
rect 6410 9840 6490 9850
rect 6630 10020 6710 10030
rect 6630 9960 6640 10020
rect 6700 9960 6710 10020
rect 6630 9840 6710 9960
rect 8610 10020 8690 10030
rect 8610 9960 8620 10020
rect 8680 9960 8690 10020
rect 8610 9910 8690 9960
rect 8610 9850 8620 9910
rect 8680 9850 8690 9910
rect 8610 9840 8690 9850
rect 8830 9840 8910 10030
rect 10810 10020 10890 10030
rect 10810 9960 10820 10020
rect 10880 9960 10890 10020
rect 10810 9910 10890 9960
rect 10810 9850 10820 9910
rect 10880 9850 10890 9910
rect 10810 9840 10890 9850
rect 11030 9840 11110 10030
rect 13010 10020 13090 10030
rect 13010 9960 13020 10020
rect 13080 9960 13090 10020
rect 13010 9910 13090 9960
rect 13010 9850 13020 9910
rect 13080 9850 13090 9910
rect 13010 9840 13090 9850
rect 13230 9840 13310 10030
rect 15210 10020 15290 10030
rect 15210 9960 15220 10020
rect 15280 9960 15290 10020
rect 15210 9840 15290 9960
rect 15430 9910 15510 10030
rect 15430 9850 15440 9910
rect 15500 9850 15510 9910
rect 15430 9840 15510 9850
rect 17410 9840 17490 10030
rect 17630 10020 17710 10030
rect 17630 9960 17640 10020
rect 17700 9960 17710 10020
rect 19620 10010 19680 10640
rect 19730 10130 19790 10140
rect 19730 10060 19790 10070
rect 19840 10010 19900 10640
rect 21930 10130 21990 10140
rect 21930 10060 21990 10070
rect 17630 9910 17710 9960
rect 17630 9850 17640 9910
rect 17700 9850 17710 9910
rect 17630 9840 17710 9850
rect 19610 9840 19690 10010
rect 19830 10000 19910 10010
rect 19830 9940 19840 10000
rect 19900 9940 19910 10000
rect 19830 9840 19910 9940
rect 2020 9230 2080 9840
rect 2130 9330 2190 9340
rect 2130 9260 2190 9270
rect 2240 9230 2300 9840
rect 2500 9810 4020 9820
rect 2500 9750 2510 9810
rect 4010 9750 4020 9810
rect 2500 9740 4020 9750
rect 2500 9640 2700 9650
rect 2500 9580 2510 9640
rect 2690 9580 2700 9640
rect 2500 9570 2700 9580
rect 3160 9640 3360 9650
rect 3160 9580 3170 9640
rect 3350 9580 3360 9640
rect 3160 9570 3360 9580
rect 3820 9640 4020 9650
rect 3820 9580 3830 9640
rect 4010 9580 4020 9640
rect 3820 9570 4020 9580
rect 2500 9430 2700 9510
rect 3160 9430 3360 9510
rect 3820 9430 4020 9510
rect 4220 9230 4280 9840
rect 4330 9330 4390 9340
rect 4330 9260 4390 9270
rect 4440 9230 4500 9840
rect 4700 9810 6220 9820
rect 4700 9750 4710 9810
rect 6210 9750 6220 9810
rect 4700 9740 6220 9750
rect 4700 9640 4900 9650
rect 4700 9580 4710 9640
rect 4890 9580 4900 9640
rect 4700 9570 4900 9580
rect 5360 9640 5560 9650
rect 5360 9580 5370 9640
rect 5550 9580 5560 9640
rect 5360 9570 5560 9580
rect 6020 9640 6220 9650
rect 6020 9580 6030 9640
rect 6210 9580 6220 9640
rect 6020 9570 6220 9580
rect 4700 9430 4900 9510
rect 5360 9430 5560 9510
rect 6020 9430 6220 9510
rect 6420 9230 6480 9840
rect 6530 9330 6590 9340
rect 6530 9260 6590 9270
rect 6640 9230 6700 9840
rect 6900 9810 8420 9820
rect 6900 9750 6910 9810
rect 8410 9750 8420 9810
rect 6900 9740 8420 9750
rect 6900 9570 7100 9650
rect 7560 9570 7760 9650
rect 8220 9570 8420 9650
rect 6900 9500 7100 9510
rect 6900 9440 6910 9500
rect 7090 9440 7100 9500
rect 6900 9430 7100 9440
rect 7560 9500 7760 9510
rect 7560 9440 7570 9500
rect 7750 9440 7760 9500
rect 7560 9430 7760 9440
rect 8220 9500 8420 9510
rect 8220 9440 8230 9500
rect 8410 9440 8420 9500
rect 8220 9430 8420 9440
rect 8620 9230 8680 9840
rect 8730 9330 8790 9340
rect 8730 9260 8790 9270
rect 8840 9230 8900 9840
rect 9100 9810 10620 9820
rect 9100 9750 9110 9810
rect 10610 9750 10620 9810
rect 9100 9740 10620 9750
rect 9100 9570 9300 9650
rect 9760 9570 9960 9650
rect 10420 9570 10620 9650
rect 9100 9500 9300 9510
rect 9100 9440 9110 9500
rect 9290 9440 9300 9500
rect 9100 9430 9300 9440
rect 9760 9500 9960 9510
rect 9760 9440 9770 9500
rect 9950 9440 9960 9500
rect 9760 9430 9960 9440
rect 10420 9500 10620 9510
rect 10420 9440 10430 9500
rect 10610 9440 10620 9500
rect 10420 9430 10620 9440
rect 10820 9230 10880 9840
rect 10930 9330 10990 9340
rect 10930 9260 10990 9270
rect 11040 9230 11100 9840
rect 11300 9810 12820 9820
rect 11300 9750 11310 9810
rect 12810 9750 12820 9810
rect 11300 9740 12820 9750
rect 11300 9570 11500 9650
rect 11960 9570 12160 9650
rect 12620 9570 12820 9650
rect 11300 9500 11500 9510
rect 11300 9440 11310 9500
rect 11490 9440 11500 9500
rect 11300 9430 11500 9440
rect 11960 9500 12160 9510
rect 11960 9440 11970 9500
rect 12150 9440 12160 9500
rect 11960 9430 12160 9440
rect 12620 9500 12820 9510
rect 12620 9440 12630 9500
rect 12810 9440 12820 9500
rect 12620 9430 12820 9440
rect 13020 9230 13080 9840
rect 13130 9330 13190 9340
rect 13130 9260 13190 9270
rect 13240 9230 13300 9840
rect 13500 9810 15020 9820
rect 13500 9750 13510 9810
rect 15010 9750 15020 9810
rect 13500 9740 15020 9750
rect 13500 9570 13700 9650
rect 14160 9570 14360 9650
rect 14820 9570 15020 9650
rect 13500 9500 13700 9510
rect 13500 9440 13510 9500
rect 13690 9440 13700 9500
rect 13500 9430 13700 9440
rect 14160 9500 14360 9510
rect 14160 9440 14170 9500
rect 14350 9440 14360 9500
rect 14160 9430 14360 9440
rect 14820 9500 15020 9510
rect 14820 9440 14830 9500
rect 15010 9440 15020 9500
rect 14820 9430 15020 9440
rect 15220 9230 15280 9840
rect 15330 9330 15390 9340
rect 15330 9260 15390 9270
rect 15440 9230 15500 9840
rect 15700 9810 17220 9820
rect 15700 9750 15710 9810
rect 17210 9750 17220 9810
rect 15700 9740 17220 9750
rect 15700 9640 15900 9650
rect 15700 9580 15710 9640
rect 15890 9580 15900 9640
rect 15700 9570 15900 9580
rect 16360 9640 16560 9650
rect 16360 9580 16370 9640
rect 16550 9580 16560 9640
rect 16360 9570 16560 9580
rect 17020 9640 17220 9650
rect 17020 9580 17030 9640
rect 17210 9580 17220 9640
rect 17020 9570 17220 9580
rect 15700 9430 15900 9510
rect 16360 9430 16560 9510
rect 17020 9430 17220 9510
rect 17420 9230 17480 9840
rect 17530 9330 17590 9340
rect 17530 9260 17590 9270
rect 17640 9230 17700 9840
rect 17900 9810 19420 9820
rect 17900 9750 17910 9810
rect 19410 9750 19420 9810
rect 17900 9740 19420 9750
rect 17900 9640 18100 9650
rect 17900 9580 17910 9640
rect 18090 9580 18100 9640
rect 17900 9570 18100 9580
rect 18560 9640 18760 9650
rect 18560 9580 18570 9640
rect 18750 9580 18760 9640
rect 18560 9570 18760 9580
rect 19220 9640 19420 9650
rect 19220 9580 19230 9640
rect 19410 9580 19420 9640
rect 19220 9570 19420 9580
rect 17900 9430 18100 9510
rect 18560 9430 18760 9510
rect 19220 9430 19420 9510
rect 1410 9210 1490 9220
rect 1410 9060 1420 9210
rect 1480 9060 1490 9210
rect 1410 9050 1490 9060
rect 420 8990 620 9000
rect 420 8910 430 8990
rect 610 8910 620 8990
rect 420 8900 620 8910
rect 420 8190 620 8200
rect 420 8110 430 8190
rect 610 8110 620 8190
rect 420 8100 620 8110
rect 420 7390 620 7400
rect 420 7310 430 7390
rect 610 7310 620 7390
rect 420 7300 620 7310
rect 1420 6820 1480 9050
rect 1620 8420 1680 9220
rect 2010 9040 2090 9230
rect 2230 9040 2310 9230
rect 4210 9110 4290 9230
rect 4210 9050 4220 9110
rect 4280 9050 4290 9110
rect 4210 9040 4290 9050
rect 4430 9040 4510 9230
rect 6410 9220 6490 9230
rect 6410 9160 6420 9220
rect 6480 9160 6490 9220
rect 6410 9040 6490 9160
rect 6630 9110 6710 9230
rect 6630 9050 6640 9110
rect 6700 9050 6710 9110
rect 6630 9040 6710 9050
rect 8610 9040 8690 9230
rect 8830 9220 8910 9230
rect 8830 9160 8840 9220
rect 8900 9160 8910 9220
rect 8830 9110 8910 9160
rect 8830 9050 8840 9110
rect 8900 9050 8910 9110
rect 8830 9040 8910 9050
rect 10810 9040 10890 9230
rect 11030 9220 11110 9230
rect 11030 9160 11040 9220
rect 11100 9160 11110 9220
rect 11030 9110 11110 9160
rect 11030 9050 11040 9110
rect 11100 9050 11110 9110
rect 11030 9040 11110 9050
rect 13010 9040 13090 9230
rect 13230 9220 13310 9230
rect 13230 9160 13240 9220
rect 13300 9160 13310 9220
rect 13230 9110 13310 9160
rect 13230 9050 13240 9110
rect 13300 9050 13310 9110
rect 13230 9040 13310 9050
rect 15210 9110 15290 9230
rect 15210 9050 15220 9110
rect 15280 9050 15290 9110
rect 15210 9040 15290 9050
rect 15430 9220 15510 9230
rect 15430 9160 15440 9220
rect 15500 9160 15510 9220
rect 15430 9040 15510 9160
rect 17410 9220 17490 9230
rect 17410 9160 17420 9220
rect 17480 9160 17490 9220
rect 17410 9040 17490 9160
rect 17630 9040 17710 9230
rect 19620 9210 19680 9840
rect 19730 9330 19790 9340
rect 19730 9260 19790 9270
rect 19840 9210 19900 9840
rect 21930 9330 21990 9340
rect 20230 9300 20310 9310
rect 19610 9040 19690 9210
rect 19830 9040 19910 9210
rect 20230 9150 20240 9300
rect 20300 9150 20310 9300
rect 20230 9140 20310 9150
rect 2020 8430 2080 9040
rect 2130 8530 2190 8540
rect 2130 8460 2190 8470
rect 2240 8430 2300 9040
rect 2500 8770 2700 8850
rect 3160 8770 3360 8850
rect 3820 8770 4020 8850
rect 2500 8700 2700 8710
rect 2500 8640 2510 8700
rect 2690 8640 2700 8700
rect 2500 8630 2700 8640
rect 3160 8700 3360 8710
rect 3160 8640 3170 8700
rect 3350 8640 3360 8700
rect 3160 8630 3360 8640
rect 3820 8700 4020 8710
rect 3820 8640 3830 8700
rect 4010 8640 4020 8700
rect 3820 8630 4020 8640
rect 4220 8430 4280 9040
rect 4330 8530 4390 8540
rect 4330 8460 4390 8470
rect 4440 8430 4500 9040
rect 4700 9010 6220 9020
rect 4700 8950 4710 9010
rect 6210 8950 6220 9010
rect 4700 8940 6220 8950
rect 4700 8770 4900 8850
rect 5360 8770 5560 8850
rect 6020 8770 6220 8850
rect 4700 8700 4900 8710
rect 4700 8640 4710 8700
rect 4890 8640 4900 8700
rect 4700 8630 4900 8640
rect 5360 8700 5560 8710
rect 5360 8640 5370 8700
rect 5550 8640 5560 8700
rect 5360 8630 5560 8640
rect 6020 8700 6220 8710
rect 6020 8640 6030 8700
rect 6210 8640 6220 8700
rect 6020 8630 6220 8640
rect 6420 8430 6480 9040
rect 6530 8530 6590 8540
rect 6530 8460 6590 8470
rect 6640 8430 6700 9040
rect 6900 9010 8420 9020
rect 6900 8950 6910 9010
rect 8410 8950 8420 9010
rect 6900 8940 8420 8950
rect 6900 8840 7100 8850
rect 6900 8780 6910 8840
rect 7090 8780 7100 8840
rect 6900 8770 7100 8780
rect 7560 8840 7760 8850
rect 7560 8780 7570 8840
rect 7750 8780 7760 8840
rect 7560 8770 7760 8780
rect 8220 8840 8420 8850
rect 8220 8780 8230 8840
rect 8410 8780 8420 8840
rect 8220 8770 8420 8780
rect 6900 8630 7100 8710
rect 7560 8630 7760 8710
rect 8220 8630 8420 8710
rect 8620 8430 8680 9040
rect 8730 8530 8790 8540
rect 8730 8460 8790 8470
rect 8840 8430 8900 9040
rect 9100 9010 10620 9020
rect 9100 8950 9110 9010
rect 10610 8950 10620 9010
rect 9100 8940 10620 8950
rect 9100 8840 9300 8850
rect 9100 8780 9110 8840
rect 9290 8780 9300 8840
rect 9100 8770 9300 8780
rect 9760 8840 9960 8850
rect 9760 8780 9770 8840
rect 9950 8780 9960 8840
rect 9760 8770 9960 8780
rect 10420 8840 10620 8850
rect 10420 8780 10430 8840
rect 10610 8780 10620 8840
rect 10420 8770 10620 8780
rect 9100 8630 9300 8710
rect 9760 8630 9960 8710
rect 10420 8630 10620 8710
rect 10820 8430 10880 9040
rect 10930 8530 10990 8540
rect 10930 8460 10990 8470
rect 11040 8430 11100 9040
rect 11300 9010 12820 9020
rect 11300 8950 11310 9010
rect 12810 8950 12820 9010
rect 11300 8940 12820 8950
rect 11300 8840 11500 8850
rect 11300 8780 11310 8840
rect 11490 8780 11500 8840
rect 11300 8770 11500 8780
rect 11960 8840 12160 8850
rect 11960 8780 11970 8840
rect 12150 8780 12160 8840
rect 11960 8770 12160 8780
rect 12620 8840 12820 8850
rect 12620 8780 12630 8840
rect 12810 8780 12820 8840
rect 12620 8770 12820 8780
rect 11300 8630 11500 8710
rect 11960 8630 12160 8710
rect 12620 8630 12820 8710
rect 13020 8430 13080 9040
rect 13130 8530 13190 8540
rect 13130 8460 13190 8470
rect 13240 8430 13300 9040
rect 13500 9010 15020 9020
rect 13500 8950 13510 9010
rect 15010 8950 15020 9010
rect 13500 8940 15020 8950
rect 13500 8840 13700 8850
rect 13500 8780 13510 8840
rect 13690 8780 13700 8840
rect 13500 8770 13700 8780
rect 14160 8840 14360 8850
rect 14160 8780 14170 8840
rect 14350 8780 14360 8840
rect 14160 8770 14360 8780
rect 14820 8840 15020 8850
rect 14820 8780 14830 8840
rect 15010 8780 15020 8840
rect 14820 8770 15020 8780
rect 13500 8630 13700 8710
rect 14160 8630 14360 8710
rect 14820 8630 15020 8710
rect 15220 8430 15280 9040
rect 15330 8530 15390 8540
rect 15330 8460 15390 8470
rect 15440 8430 15500 9040
rect 15700 9010 17220 9020
rect 15700 8950 15710 9010
rect 17210 8950 17220 9010
rect 15700 8940 17220 8950
rect 15700 8770 15900 8850
rect 16360 8770 16560 8850
rect 17020 8770 17220 8850
rect 15700 8700 15900 8710
rect 15700 8640 15710 8700
rect 15890 8640 15900 8700
rect 15700 8630 15900 8640
rect 16360 8700 16560 8710
rect 16360 8640 16370 8700
rect 16550 8640 16560 8700
rect 16360 8630 16560 8640
rect 17020 8700 17220 8710
rect 17020 8640 17030 8700
rect 17210 8640 17220 8700
rect 17020 8630 17220 8640
rect 17420 8430 17480 9040
rect 17530 8530 17590 8540
rect 17530 8460 17590 8470
rect 17640 8430 17700 9040
rect 17900 8770 18100 8850
rect 18560 8770 18760 8850
rect 19220 8770 19420 8850
rect 17900 8700 18100 8710
rect 17900 8640 17910 8700
rect 18090 8640 18100 8700
rect 17900 8630 18100 8640
rect 18560 8700 18760 8710
rect 18560 8640 18570 8700
rect 18750 8640 18760 8700
rect 18560 8630 18760 8640
rect 19220 8700 19420 8710
rect 19220 8640 19230 8700
rect 19410 8640 19420 8700
rect 19220 8630 19420 8640
rect 1610 8410 1690 8420
rect 1610 8260 1620 8410
rect 1680 8260 1690 8410
rect 1610 8250 1690 8260
rect 1620 7620 1680 8250
rect 2010 8240 2090 8430
rect 2230 8240 2310 8430
rect 4210 8240 4290 8430
rect 4430 8310 4510 8430
rect 4430 8250 4440 8310
rect 4500 8250 4510 8310
rect 4430 8240 4510 8250
rect 6410 8310 6490 8430
rect 6410 8250 6420 8310
rect 6480 8250 6490 8310
rect 6410 8240 6490 8250
rect 6630 8420 6710 8430
rect 6630 8360 6640 8420
rect 6700 8360 6710 8420
rect 6630 8240 6710 8360
rect 8610 8420 8690 8430
rect 8610 8360 8620 8420
rect 8680 8360 8690 8420
rect 8610 8310 8690 8360
rect 8610 8250 8620 8310
rect 8680 8250 8690 8310
rect 8610 8240 8690 8250
rect 8830 8240 8910 8430
rect 10810 8420 10890 8430
rect 10810 8360 10820 8420
rect 10880 8360 10890 8420
rect 10810 8310 10890 8360
rect 10810 8250 10820 8310
rect 10880 8250 10890 8310
rect 10810 8240 10890 8250
rect 11030 8240 11110 8430
rect 13010 8420 13090 8430
rect 13010 8360 13020 8420
rect 13080 8360 13090 8420
rect 13010 8310 13090 8360
rect 13010 8250 13020 8310
rect 13080 8250 13090 8310
rect 13010 8240 13090 8250
rect 13230 8240 13310 8430
rect 15210 8420 15290 8430
rect 15210 8360 15220 8420
rect 15280 8360 15290 8420
rect 15210 8240 15290 8360
rect 15430 8310 15510 8430
rect 15430 8250 15440 8310
rect 15500 8250 15510 8310
rect 15430 8240 15510 8250
rect 17410 8240 17490 8430
rect 17630 8420 17710 8430
rect 17630 8360 17640 8420
rect 17700 8360 17710 8420
rect 19620 8410 19680 9040
rect 19730 8530 19790 8540
rect 19730 8460 19790 8470
rect 19840 8410 19900 9040
rect 17630 8240 17710 8360
rect 19610 8240 19690 8410
rect 19830 8240 19910 8410
rect 2020 7630 2080 8240
rect 2130 7730 2190 7740
rect 2130 7660 2190 7670
rect 2240 7630 2300 8240
rect 2500 7970 2700 8050
rect 3160 7970 3360 8050
rect 3820 7970 4020 8050
rect 2500 7900 2700 7910
rect 2500 7840 2510 7900
rect 2690 7840 2700 7900
rect 2500 7830 2700 7840
rect 3160 7900 3360 7910
rect 3160 7840 3170 7900
rect 3350 7840 3360 7900
rect 3160 7830 3360 7840
rect 3820 7900 4020 7910
rect 3820 7840 3830 7900
rect 4010 7840 4020 7900
rect 3820 7830 4020 7840
rect 4220 7630 4280 8240
rect 4330 7730 4390 7740
rect 4330 7660 4390 7670
rect 4440 7630 4500 8240
rect 4700 8210 6220 8220
rect 4700 8150 4710 8210
rect 6210 8150 6220 8210
rect 4700 8140 6220 8150
rect 4700 7970 4900 8050
rect 5360 7970 5560 8050
rect 6020 7970 6220 8050
rect 4700 7900 4900 7910
rect 4700 7840 4710 7900
rect 4890 7840 4900 7900
rect 4700 7830 4900 7840
rect 5360 7900 5560 7910
rect 5360 7840 5370 7900
rect 5550 7840 5560 7900
rect 5360 7830 5560 7840
rect 6020 7900 6220 7910
rect 6020 7840 6030 7900
rect 6210 7840 6220 7900
rect 6020 7830 6220 7840
rect 6420 7630 6480 8240
rect 6530 7730 6590 7740
rect 6530 7660 6590 7670
rect 6640 7630 6700 8240
rect 6900 8210 8420 8220
rect 6900 8150 6910 8210
rect 8410 8150 8420 8210
rect 6900 8140 8420 8150
rect 6900 8040 7100 8050
rect 6900 7980 6910 8040
rect 7090 7980 7100 8040
rect 6900 7970 7100 7980
rect 7560 8040 7760 8050
rect 7560 7980 7570 8040
rect 7750 7980 7760 8040
rect 7560 7970 7760 7980
rect 8220 8040 8420 8050
rect 8220 7980 8230 8040
rect 8410 7980 8420 8040
rect 8220 7970 8420 7980
rect 6900 7830 7100 7910
rect 7560 7830 7760 7910
rect 8220 7830 8420 7910
rect 8620 7630 8680 8240
rect 8730 7730 8790 7740
rect 8730 7660 8790 7670
rect 8840 7630 8900 8240
rect 9100 8210 10620 8220
rect 9100 8150 9110 8210
rect 10610 8150 10620 8210
rect 9100 8140 10620 8150
rect 9100 8040 9300 8050
rect 9100 7980 9110 8040
rect 9290 7980 9300 8040
rect 9100 7970 9300 7980
rect 9760 8040 9960 8050
rect 9760 7980 9770 8040
rect 9950 7980 9960 8040
rect 9760 7970 9960 7980
rect 10420 8040 10620 8050
rect 10420 7980 10430 8040
rect 10610 7980 10620 8040
rect 10420 7970 10620 7980
rect 9100 7830 9300 7910
rect 9760 7830 9960 7910
rect 10420 7830 10620 7910
rect 10820 7630 10880 8240
rect 10930 7730 10990 7740
rect 10930 7660 10990 7670
rect 11040 7630 11100 8240
rect 11300 8210 12820 8220
rect 11300 8150 11310 8210
rect 12810 8150 12820 8210
rect 11300 8140 12820 8150
rect 11300 8040 11500 8050
rect 11300 7980 11310 8040
rect 11490 7980 11500 8040
rect 11300 7970 11500 7980
rect 11960 8040 12160 8050
rect 11960 7980 11970 8040
rect 12150 7980 12160 8040
rect 11960 7970 12160 7980
rect 12620 8040 12820 8050
rect 12620 7980 12630 8040
rect 12810 7980 12820 8040
rect 12620 7970 12820 7980
rect 11300 7830 11500 7910
rect 11960 7830 12160 7910
rect 12620 7830 12820 7910
rect 13020 7630 13080 8240
rect 13130 7730 13190 7740
rect 13130 7660 13190 7670
rect 13240 7630 13300 8240
rect 13500 8210 15020 8220
rect 13500 8150 13510 8210
rect 15010 8150 15020 8210
rect 13500 8140 15020 8150
rect 13500 8040 13700 8050
rect 13500 7980 13510 8040
rect 13690 7980 13700 8040
rect 13500 7970 13700 7980
rect 14160 8040 14360 8050
rect 14160 7980 14170 8040
rect 14350 7980 14360 8040
rect 14160 7970 14360 7980
rect 14820 8040 15020 8050
rect 14820 7980 14830 8040
rect 15010 7980 15020 8040
rect 14820 7970 15020 7980
rect 13500 7830 13700 7910
rect 14160 7830 14360 7910
rect 14820 7830 15020 7910
rect 15220 7630 15280 8240
rect 15330 7730 15390 7740
rect 15330 7660 15390 7670
rect 15440 7630 15500 8240
rect 15700 8210 17220 8220
rect 15700 8150 15710 8210
rect 17210 8150 17220 8210
rect 15700 8140 17220 8150
rect 15700 7970 15900 8050
rect 16360 7970 16560 8050
rect 17020 7970 17220 8050
rect 15700 7900 15900 7910
rect 15700 7840 15710 7900
rect 15890 7840 15900 7900
rect 15700 7830 15900 7840
rect 16360 7900 16560 7910
rect 16360 7840 16370 7900
rect 16550 7840 16560 7900
rect 16360 7830 16560 7840
rect 17020 7900 17220 7910
rect 17020 7840 17030 7900
rect 17210 7840 17220 7900
rect 17020 7830 17220 7840
rect 17420 7630 17480 8240
rect 17530 7730 17590 7740
rect 17530 7660 17590 7670
rect 17640 7630 17700 8240
rect 17900 7970 18100 8050
rect 18560 7970 18760 8050
rect 19220 7970 19420 8050
rect 17900 7900 18100 7910
rect 17900 7840 17910 7900
rect 18090 7840 18100 7900
rect 17900 7830 18100 7840
rect 18560 7900 18760 7910
rect 18560 7840 18570 7900
rect 18750 7840 18760 7900
rect 18560 7830 18760 7840
rect 19220 7900 19420 7910
rect 19220 7840 19230 7900
rect 19410 7840 19420 7900
rect 19220 7830 19420 7840
rect 1610 7610 1690 7620
rect 1610 7460 1620 7610
rect 1680 7460 1690 7610
rect 1610 7450 1690 7460
rect 1410 6810 1490 6820
rect 1410 6660 1420 6810
rect 1480 6660 1490 6810
rect 1410 6650 1490 6660
rect 420 6590 620 6600
rect 420 6510 430 6590
rect 610 6510 620 6590
rect 420 6500 620 6510
rect 1420 4540 1480 6650
rect 1280 4530 1480 4540
rect 1280 4350 1290 4530
rect 1470 4350 1480 4530
rect 1280 4340 1480 4350
rect 1620 4140 1680 7450
rect 2010 7440 2090 7630
rect 2230 7440 2310 7630
rect 4210 7440 4290 7630
rect 4430 7510 4510 7630
rect 4430 7450 4440 7510
rect 4500 7450 4510 7510
rect 4430 7440 4510 7450
rect 6410 7510 6490 7630
rect 6410 7450 6420 7510
rect 6480 7450 6490 7510
rect 6410 7440 6490 7450
rect 6630 7620 6710 7630
rect 6630 7560 6640 7620
rect 6700 7560 6710 7620
rect 6630 7440 6710 7560
rect 8610 7620 8690 7630
rect 8610 7560 8620 7620
rect 8680 7560 8690 7620
rect 8610 7510 8690 7560
rect 8610 7450 8620 7510
rect 8680 7450 8690 7510
rect 8610 7440 8690 7450
rect 8830 7440 8910 7630
rect 10810 7620 10890 7630
rect 10810 7560 10820 7620
rect 10880 7560 10890 7620
rect 10810 7510 10890 7560
rect 10810 7450 10820 7510
rect 10880 7450 10890 7510
rect 10810 7440 10890 7450
rect 11030 7440 11110 7630
rect 13010 7620 13090 7630
rect 13010 7560 13020 7620
rect 13080 7560 13090 7620
rect 13010 7510 13090 7560
rect 13010 7450 13020 7510
rect 13080 7450 13090 7510
rect 13010 7440 13090 7450
rect 13230 7440 13310 7630
rect 15210 7620 15290 7630
rect 15210 7560 15220 7620
rect 15280 7560 15290 7620
rect 15210 7440 15290 7560
rect 15430 7510 15510 7630
rect 15430 7450 15440 7510
rect 15500 7450 15510 7510
rect 15430 7440 15510 7450
rect 17410 7440 17490 7630
rect 17630 7620 17710 7630
rect 17630 7560 17640 7620
rect 17700 7560 17710 7620
rect 19620 7610 19680 8240
rect 19730 7730 19790 7740
rect 19730 7660 19790 7670
rect 19840 7610 19900 8240
rect 17630 7440 17710 7560
rect 19610 7440 19690 7610
rect 19830 7440 19910 7610
rect 2020 6830 2080 7440
rect 2130 6930 2190 6940
rect 2130 6860 2190 6870
rect 2240 6830 2300 7440
rect 2500 7240 2700 7250
rect 2500 7180 2510 7240
rect 2690 7180 2700 7240
rect 2500 7170 2700 7180
rect 3160 7240 3360 7250
rect 3160 7180 3170 7240
rect 3350 7180 3360 7240
rect 3160 7170 3360 7180
rect 3820 7240 4020 7250
rect 3820 7180 3830 7240
rect 4010 7180 4020 7240
rect 3820 7170 4020 7180
rect 2500 7030 2700 7110
rect 3160 7030 3360 7110
rect 3820 7030 4020 7110
rect 4220 6830 4280 7440
rect 4330 6930 4390 6940
rect 4330 6860 4390 6870
rect 4440 6830 4500 7440
rect 4700 7410 6220 7420
rect 4700 7350 4710 7410
rect 6210 7350 6220 7410
rect 4700 7340 6220 7350
rect 4700 7240 4900 7250
rect 4700 7180 4710 7240
rect 4890 7180 4900 7240
rect 4700 7170 4900 7180
rect 5360 7240 5560 7250
rect 5360 7180 5370 7240
rect 5550 7180 5560 7240
rect 5360 7170 5560 7180
rect 6020 7240 6220 7250
rect 6020 7180 6030 7240
rect 6210 7180 6220 7240
rect 6020 7170 6220 7180
rect 4700 7030 4900 7110
rect 5360 7030 5560 7110
rect 6020 7030 6220 7110
rect 6420 6830 6480 7440
rect 6530 6930 6590 6940
rect 6530 6860 6590 6870
rect 6640 6830 6700 7440
rect 6900 7410 8420 7420
rect 6900 7350 6910 7410
rect 8410 7350 8420 7410
rect 6900 7340 8420 7350
rect 6900 7170 7100 7250
rect 7560 7170 7760 7250
rect 8220 7170 8420 7250
rect 6900 7100 7100 7110
rect 6900 7040 6910 7100
rect 7090 7040 7100 7100
rect 6900 7030 7100 7040
rect 7560 7100 7760 7110
rect 7560 7040 7570 7100
rect 7750 7040 7760 7100
rect 7560 7030 7760 7040
rect 8220 7100 8420 7110
rect 8220 7040 8230 7100
rect 8410 7040 8420 7100
rect 8220 7030 8420 7040
rect 8620 6830 8680 7440
rect 8730 6930 8790 6940
rect 8730 6860 8790 6870
rect 8840 6830 8900 7440
rect 9100 7410 10620 7420
rect 9100 7350 9110 7410
rect 10610 7350 10620 7410
rect 9100 7340 10620 7350
rect 9100 7170 9300 7250
rect 9760 7170 9960 7250
rect 10420 7170 10620 7250
rect 9100 7100 9300 7110
rect 9100 7040 9110 7100
rect 9290 7040 9300 7100
rect 9100 7030 9300 7040
rect 9760 7100 9960 7110
rect 9760 7040 9770 7100
rect 9950 7040 9960 7100
rect 9760 7030 9960 7040
rect 10420 7100 10620 7110
rect 10420 7040 10430 7100
rect 10610 7040 10620 7100
rect 10420 7030 10620 7040
rect 10820 6830 10880 7440
rect 10930 6930 10990 6940
rect 10930 6860 10990 6870
rect 11040 6830 11100 7440
rect 11300 7410 12820 7420
rect 11300 7350 11310 7410
rect 12810 7350 12820 7410
rect 11300 7340 12820 7350
rect 11300 7170 11500 7250
rect 11960 7170 12160 7250
rect 12620 7170 12820 7250
rect 11300 7100 11500 7110
rect 11300 7040 11310 7100
rect 11490 7040 11500 7100
rect 11300 7030 11500 7040
rect 11960 7100 12160 7110
rect 11960 7040 11970 7100
rect 12150 7040 12160 7100
rect 11960 7030 12160 7040
rect 12620 7100 12820 7110
rect 12620 7040 12630 7100
rect 12810 7040 12820 7100
rect 12620 7030 12820 7040
rect 13020 6830 13080 7440
rect 13130 6930 13190 6940
rect 13130 6860 13190 6870
rect 13240 6830 13300 7440
rect 13500 7410 15020 7420
rect 13500 7350 13510 7410
rect 15010 7350 15020 7410
rect 13500 7340 15020 7350
rect 13500 7170 13700 7250
rect 14160 7170 14360 7250
rect 14820 7170 15020 7250
rect 13500 7100 13700 7110
rect 13500 7040 13510 7100
rect 13690 7040 13700 7100
rect 13500 7030 13700 7040
rect 14160 7100 14360 7110
rect 14160 7040 14170 7100
rect 14350 7040 14360 7100
rect 14160 7030 14360 7040
rect 14820 7100 15020 7110
rect 14820 7040 14830 7100
rect 15010 7040 15020 7100
rect 14820 7030 15020 7040
rect 15220 6830 15280 7440
rect 15330 6930 15390 6940
rect 15330 6860 15390 6870
rect 15440 6830 15500 7440
rect 15700 7410 17220 7420
rect 15700 7350 15710 7410
rect 17210 7350 17220 7410
rect 15700 7340 17220 7350
rect 15700 7240 15900 7250
rect 15700 7180 15710 7240
rect 15890 7180 15900 7240
rect 15700 7170 15900 7180
rect 16360 7240 16560 7250
rect 16360 7180 16370 7240
rect 16550 7180 16560 7240
rect 16360 7170 16560 7180
rect 17020 7240 17220 7250
rect 17020 7180 17030 7240
rect 17210 7180 17220 7240
rect 17020 7170 17220 7180
rect 15700 7030 15900 7110
rect 16360 7030 16560 7110
rect 17020 7030 17220 7110
rect 17420 6830 17480 7440
rect 17530 6930 17590 6940
rect 17530 6860 17590 6870
rect 17640 6830 17700 7440
rect 17900 7240 18100 7250
rect 17900 7180 17910 7240
rect 18090 7180 18100 7240
rect 17900 7170 18100 7180
rect 18560 7240 18760 7250
rect 18560 7180 18570 7240
rect 18750 7180 18760 7240
rect 18560 7170 18760 7180
rect 19220 7240 19420 7250
rect 19220 7180 19230 7240
rect 19410 7180 19420 7240
rect 19220 7170 19420 7180
rect 17900 7030 18100 7110
rect 18560 7030 18760 7110
rect 19220 7030 19420 7110
rect 2010 6640 2090 6830
rect 2230 6640 2310 6830
rect 4210 6710 4290 6830
rect 4210 6650 4220 6710
rect 4280 6650 4290 6710
rect 4210 6640 4290 6650
rect 4430 6640 4510 6830
rect 6410 6820 6490 6830
rect 6410 6760 6420 6820
rect 6480 6760 6490 6820
rect 6410 6640 6490 6760
rect 6630 6710 6710 6830
rect 6630 6650 6640 6710
rect 6700 6650 6710 6710
rect 6630 6640 6710 6650
rect 8610 6640 8690 6830
rect 8830 6820 8910 6830
rect 8830 6760 8840 6820
rect 8900 6760 8910 6820
rect 8830 6710 8910 6760
rect 8830 6650 8840 6710
rect 8900 6650 8910 6710
rect 8830 6640 8910 6650
rect 10810 6640 10890 6830
rect 11030 6820 11110 6830
rect 11030 6760 11040 6820
rect 11100 6760 11110 6820
rect 11030 6710 11110 6760
rect 11030 6650 11040 6710
rect 11100 6650 11110 6710
rect 11030 6640 11110 6650
rect 13010 6640 13090 6830
rect 13230 6820 13310 6830
rect 13230 6760 13240 6820
rect 13300 6760 13310 6820
rect 13230 6710 13310 6760
rect 13230 6650 13240 6710
rect 13300 6650 13310 6710
rect 13230 6640 13310 6650
rect 15210 6710 15290 6830
rect 15210 6650 15220 6710
rect 15280 6650 15290 6710
rect 15210 6640 15290 6650
rect 15430 6820 15510 6830
rect 15430 6760 15440 6820
rect 15500 6760 15510 6820
rect 15430 6640 15510 6760
rect 17410 6820 17490 6830
rect 17410 6760 17420 6820
rect 17480 6760 17490 6820
rect 17410 6640 17490 6760
rect 17630 6640 17710 6830
rect 19620 6810 19680 7440
rect 19730 6930 19790 6940
rect 19730 6860 19790 6870
rect 19840 6810 19900 7440
rect 20240 6910 20300 9140
rect 20440 8510 20500 9310
rect 21930 9260 21990 9270
rect 21300 8990 21500 9000
rect 21300 8910 21310 8990
rect 21490 8910 21500 8990
rect 21300 8900 21500 8910
rect 21930 8530 21990 8540
rect 20430 8500 20510 8510
rect 20430 8350 20440 8500
rect 20500 8350 20510 8500
rect 21930 8460 21990 8470
rect 20430 8340 20510 8350
rect 20440 7710 20500 8340
rect 21300 8190 21500 8200
rect 21300 8110 21310 8190
rect 21490 8110 21500 8190
rect 21300 8100 21500 8110
rect 21930 7730 21990 7740
rect 20430 7700 20510 7710
rect 20430 7550 20440 7700
rect 20500 7550 20510 7700
rect 21930 7660 21990 7670
rect 20430 7540 20510 7550
rect 20230 6900 20310 6910
rect 19610 6640 19690 6810
rect 19830 6640 19910 6810
rect 20230 6750 20240 6900
rect 20300 6750 20310 6900
rect 20230 6740 20310 6750
rect 2020 6030 2080 6640
rect 2130 6130 2190 6140
rect 2130 6060 2190 6070
rect 2240 6030 2300 6640
rect 2500 6370 2700 6450
rect 3160 6370 3360 6450
rect 3820 6370 4020 6450
rect 2500 6300 2700 6310
rect 2500 6240 2510 6300
rect 2690 6240 2700 6300
rect 2500 6230 2700 6240
rect 3160 6300 3360 6310
rect 3160 6240 3170 6300
rect 3350 6240 3360 6300
rect 3160 6230 3360 6240
rect 3820 6300 4020 6310
rect 3820 6240 3830 6300
rect 4010 6240 4020 6300
rect 3820 6230 4020 6240
rect 4220 6030 4280 6640
rect 4330 6130 4390 6140
rect 4330 6060 4390 6070
rect 4440 6030 4500 6640
rect 4700 6610 6220 6620
rect 4700 6550 4710 6610
rect 6210 6550 6220 6610
rect 4700 6540 6220 6550
rect 4700 6370 4900 6450
rect 5360 6370 5560 6450
rect 6020 6370 6220 6450
rect 4700 6300 4900 6310
rect 4700 6240 4710 6300
rect 4890 6240 4900 6300
rect 4700 6230 4900 6240
rect 5360 6300 5560 6310
rect 5360 6240 5370 6300
rect 5550 6240 5560 6300
rect 5360 6230 5560 6240
rect 6020 6300 6220 6310
rect 6020 6240 6030 6300
rect 6210 6240 6220 6300
rect 6020 6230 6220 6240
rect 6420 6030 6480 6640
rect 6530 6130 6590 6140
rect 6530 6060 6590 6070
rect 6640 6030 6700 6640
rect 6900 6610 8420 6620
rect 6900 6550 6910 6610
rect 8410 6550 8420 6610
rect 6900 6540 8420 6550
rect 6900 6440 7100 6450
rect 6900 6380 6910 6440
rect 7090 6380 7100 6440
rect 6900 6370 7100 6380
rect 7560 6440 7760 6450
rect 7560 6380 7570 6440
rect 7750 6380 7760 6440
rect 7560 6370 7760 6380
rect 8220 6440 8420 6450
rect 8220 6380 8230 6440
rect 8410 6380 8420 6440
rect 8220 6370 8420 6380
rect 6900 6230 7100 6310
rect 7560 6230 7760 6310
rect 8220 6230 8420 6310
rect 8620 6030 8680 6640
rect 8730 6130 8790 6140
rect 8730 6060 8790 6070
rect 8840 6030 8900 6640
rect 9100 6610 10620 6620
rect 9100 6550 9110 6610
rect 10610 6550 10620 6610
rect 9100 6540 10620 6550
rect 9100 6440 9300 6450
rect 9100 6380 9110 6440
rect 9290 6380 9300 6440
rect 9100 6370 9300 6380
rect 9760 6440 9960 6450
rect 9760 6380 9770 6440
rect 9950 6380 9960 6440
rect 9760 6370 9960 6380
rect 10420 6440 10620 6450
rect 10420 6380 10430 6440
rect 10610 6380 10620 6440
rect 10420 6370 10620 6380
rect 9100 6230 9300 6310
rect 9760 6230 9960 6310
rect 10420 6230 10620 6310
rect 10820 6030 10880 6640
rect 10930 6130 10990 6140
rect 10930 6060 10990 6070
rect 11040 6030 11100 6640
rect 11300 6610 12820 6620
rect 11300 6550 11310 6610
rect 12810 6550 12820 6610
rect 11300 6540 12820 6550
rect 11300 6440 11500 6450
rect 11300 6380 11310 6440
rect 11490 6380 11500 6440
rect 11300 6370 11500 6380
rect 11960 6440 12160 6450
rect 11960 6380 11970 6440
rect 12150 6380 12160 6440
rect 11960 6370 12160 6380
rect 12620 6440 12820 6450
rect 12620 6380 12630 6440
rect 12810 6380 12820 6440
rect 12620 6370 12820 6380
rect 11300 6230 11500 6310
rect 11960 6230 12160 6310
rect 12620 6230 12820 6310
rect 13020 6030 13080 6640
rect 13130 6130 13190 6140
rect 13130 6060 13190 6070
rect 13240 6030 13300 6640
rect 13500 6610 15020 6620
rect 13500 6550 13510 6610
rect 15010 6550 15020 6610
rect 13500 6540 15020 6550
rect 13500 6440 13700 6450
rect 13500 6380 13510 6440
rect 13690 6380 13700 6440
rect 13500 6370 13700 6380
rect 14160 6440 14360 6450
rect 14160 6380 14170 6440
rect 14350 6380 14360 6440
rect 14160 6370 14360 6380
rect 14820 6440 15020 6450
rect 14820 6380 14830 6440
rect 15010 6380 15020 6440
rect 14820 6370 15020 6380
rect 13500 6230 13700 6310
rect 14160 6230 14360 6310
rect 14820 6230 15020 6310
rect 15220 6030 15280 6640
rect 15330 6130 15390 6140
rect 15330 6060 15390 6070
rect 15440 6030 15500 6640
rect 15700 6610 17220 6620
rect 15700 6550 15710 6610
rect 17210 6550 17220 6610
rect 15700 6540 17220 6550
rect 15700 6370 15900 6450
rect 16360 6370 16560 6450
rect 17020 6370 17220 6450
rect 15700 6300 15900 6310
rect 15700 6240 15710 6300
rect 15890 6240 15900 6300
rect 15700 6230 15900 6240
rect 16360 6300 16560 6310
rect 16360 6240 16370 6300
rect 16550 6240 16560 6300
rect 16360 6230 16560 6240
rect 17020 6300 17220 6310
rect 17020 6240 17030 6300
rect 17210 6240 17220 6300
rect 17020 6230 17220 6240
rect 17420 6030 17480 6640
rect 17530 6130 17590 6140
rect 17530 6060 17590 6070
rect 17640 6030 17700 6640
rect 17900 6370 18100 6450
rect 18560 6370 18760 6450
rect 19220 6370 19420 6450
rect 17900 6300 18100 6310
rect 17900 6240 17910 6300
rect 18090 6240 18100 6300
rect 17900 6230 18100 6240
rect 18560 6300 18760 6310
rect 18560 6240 18570 6300
rect 18750 6240 18760 6300
rect 18560 6230 18760 6240
rect 19220 6300 19420 6310
rect 19220 6240 19230 6300
rect 19410 6240 19420 6300
rect 19220 6230 19420 6240
rect 2010 5840 2090 6030
rect 2230 5910 2310 6030
rect 2230 5850 2240 5910
rect 2300 5850 2310 5910
rect 2230 5840 2310 5850
rect 4210 5840 4290 6030
rect 4430 6020 4510 6030
rect 4430 5960 4440 6020
rect 4500 5960 4510 6020
rect 4430 5910 4510 5960
rect 4430 5850 4440 5910
rect 4500 5850 4510 5910
rect 4430 5840 4510 5850
rect 6410 5910 6490 6030
rect 6410 5850 6420 5910
rect 6480 5850 6490 5910
rect 6410 5840 6490 5850
rect 6630 6020 6710 6030
rect 6630 5960 6640 6020
rect 6700 5960 6710 6020
rect 6630 5840 6710 5960
rect 8610 6020 8690 6030
rect 8610 5960 8620 6020
rect 8680 5960 8690 6020
rect 8610 5910 8690 5960
rect 8610 5850 8620 5910
rect 8680 5850 8690 5910
rect 8610 5840 8690 5850
rect 8830 5840 8910 6030
rect 10810 6020 10890 6030
rect 10810 5960 10820 6020
rect 10880 5960 10890 6020
rect 10810 5910 10890 5960
rect 10810 5850 10820 5910
rect 10880 5850 10890 5910
rect 10810 5840 10890 5850
rect 11030 5840 11110 6030
rect 13010 6020 13090 6030
rect 13010 5960 13020 6020
rect 13080 5960 13090 6020
rect 13010 5910 13090 5960
rect 13010 5850 13020 5910
rect 13080 5850 13090 5910
rect 13010 5840 13090 5850
rect 13230 5840 13310 6030
rect 15210 6020 15290 6030
rect 15210 5960 15220 6020
rect 15280 5960 15290 6020
rect 15210 5840 15290 5960
rect 15430 5910 15510 6030
rect 15430 5850 15440 5910
rect 15500 5850 15510 5910
rect 15430 5840 15510 5850
rect 17410 5840 17490 6030
rect 17630 6020 17710 6030
rect 17630 5960 17640 6020
rect 17700 5960 17710 6020
rect 19620 6010 19680 6640
rect 19730 6130 19790 6140
rect 19730 6060 19790 6070
rect 19840 6010 19900 6640
rect 17630 5910 17710 5960
rect 17630 5850 17640 5910
rect 17700 5850 17710 5910
rect 17630 5840 17710 5850
rect 19610 5840 19690 6010
rect 19830 6000 19910 6010
rect 19830 5940 19840 6000
rect 19900 5940 19910 6000
rect 19830 5840 19910 5940
rect 2020 5230 2080 5840
rect 2130 5330 2190 5340
rect 2130 5260 2190 5270
rect 2240 5230 2300 5840
rect 2500 5810 4020 5820
rect 2500 5750 2510 5810
rect 4010 5750 4020 5810
rect 2500 5740 4020 5750
rect 2500 5640 2700 5650
rect 2500 5580 2510 5640
rect 2690 5580 2700 5640
rect 2500 5570 2700 5580
rect 3160 5640 3360 5650
rect 3160 5580 3170 5640
rect 3350 5580 3360 5640
rect 3160 5570 3360 5580
rect 3820 5640 4020 5650
rect 3820 5580 3830 5640
rect 4010 5580 4020 5640
rect 3820 5570 4020 5580
rect 2500 5430 2700 5510
rect 3160 5430 3360 5510
rect 3820 5430 4020 5510
rect 4220 5230 4280 5840
rect 4330 5330 4390 5340
rect 4330 5260 4390 5270
rect 4440 5230 4500 5840
rect 4700 5810 6220 5820
rect 4700 5750 4710 5810
rect 6210 5750 6220 5810
rect 4700 5740 6220 5750
rect 4700 5640 4900 5650
rect 4700 5580 4710 5640
rect 4890 5580 4900 5640
rect 4700 5570 4900 5580
rect 5360 5640 5560 5650
rect 5360 5580 5370 5640
rect 5550 5580 5560 5640
rect 5360 5570 5560 5580
rect 6020 5640 6220 5650
rect 6020 5580 6030 5640
rect 6210 5580 6220 5640
rect 6020 5570 6220 5580
rect 4700 5430 4900 5510
rect 5360 5430 5560 5510
rect 6020 5430 6220 5510
rect 6420 5230 6480 5840
rect 6530 5330 6590 5340
rect 6530 5260 6590 5270
rect 6640 5230 6700 5840
rect 6900 5810 8420 5820
rect 6900 5750 6910 5810
rect 8410 5750 8420 5810
rect 6900 5740 8420 5750
rect 6900 5570 7100 5650
rect 7560 5570 7760 5650
rect 8220 5570 8420 5650
rect 6900 5500 7100 5510
rect 6900 5440 6910 5500
rect 7090 5440 7100 5500
rect 6900 5430 7100 5440
rect 7560 5500 7760 5510
rect 7560 5440 7570 5500
rect 7750 5440 7760 5500
rect 7560 5430 7760 5440
rect 8220 5500 8420 5510
rect 8220 5440 8230 5500
rect 8410 5440 8420 5500
rect 8220 5430 8420 5440
rect 8620 5230 8680 5840
rect 8730 5330 8790 5340
rect 8730 5260 8790 5270
rect 8840 5230 8900 5840
rect 9100 5810 10620 5820
rect 9100 5750 9110 5810
rect 10610 5750 10620 5810
rect 9100 5740 10620 5750
rect 9100 5570 9300 5650
rect 9760 5570 9960 5650
rect 10420 5570 10620 5650
rect 9100 5500 9300 5510
rect 9100 5440 9110 5500
rect 9290 5440 9300 5500
rect 9100 5430 9300 5440
rect 9760 5500 9960 5510
rect 9760 5440 9770 5500
rect 9950 5440 9960 5500
rect 9760 5430 9960 5440
rect 10420 5500 10620 5510
rect 10420 5440 10430 5500
rect 10610 5440 10620 5500
rect 10420 5430 10620 5440
rect 10820 5230 10880 5840
rect 10930 5330 10990 5340
rect 10930 5260 10990 5270
rect 11040 5230 11100 5840
rect 11300 5810 12820 5820
rect 11300 5750 11310 5810
rect 12810 5750 12820 5810
rect 11300 5740 12820 5750
rect 11300 5570 11500 5650
rect 11960 5570 12160 5650
rect 12620 5570 12820 5650
rect 11300 5500 11500 5510
rect 11300 5440 11310 5500
rect 11490 5440 11500 5500
rect 11300 5430 11500 5440
rect 11960 5500 12160 5510
rect 11960 5440 11970 5500
rect 12150 5440 12160 5500
rect 11960 5430 12160 5440
rect 12620 5500 12820 5510
rect 12620 5440 12630 5500
rect 12810 5440 12820 5500
rect 12620 5430 12820 5440
rect 13020 5230 13080 5840
rect 13130 5330 13190 5340
rect 13130 5260 13190 5270
rect 13240 5230 13300 5840
rect 13500 5810 15020 5820
rect 13500 5750 13510 5810
rect 15010 5750 15020 5810
rect 13500 5740 15020 5750
rect 13500 5570 13700 5650
rect 14160 5570 14360 5650
rect 14820 5570 15020 5650
rect 13500 5500 13700 5510
rect 13500 5440 13510 5500
rect 13690 5440 13700 5500
rect 13500 5430 13700 5440
rect 14160 5500 14360 5510
rect 14160 5440 14170 5500
rect 14350 5440 14360 5500
rect 14160 5430 14360 5440
rect 14820 5500 15020 5510
rect 14820 5440 14830 5500
rect 15010 5440 15020 5500
rect 14820 5430 15020 5440
rect 15220 5230 15280 5840
rect 15330 5330 15390 5340
rect 15330 5260 15390 5270
rect 15440 5230 15500 5840
rect 15700 5810 17220 5820
rect 15700 5750 15710 5810
rect 17210 5750 17220 5810
rect 15700 5740 17220 5750
rect 15700 5640 15900 5650
rect 15700 5580 15710 5640
rect 15890 5580 15900 5640
rect 15700 5570 15900 5580
rect 16360 5640 16560 5650
rect 16360 5580 16370 5640
rect 16550 5580 16560 5640
rect 16360 5570 16560 5580
rect 17020 5640 17220 5650
rect 17020 5580 17030 5640
rect 17210 5580 17220 5640
rect 17020 5570 17220 5580
rect 15700 5430 15900 5510
rect 16360 5430 16560 5510
rect 17020 5430 17220 5510
rect 17420 5230 17480 5840
rect 17530 5330 17590 5340
rect 17530 5260 17590 5270
rect 17640 5230 17700 5840
rect 17900 5810 19420 5820
rect 17900 5750 17910 5810
rect 19410 5750 19420 5810
rect 17900 5740 19420 5750
rect 17900 5640 18100 5650
rect 17900 5580 17910 5640
rect 18090 5580 18100 5640
rect 17900 5570 18100 5580
rect 18560 5640 18760 5650
rect 18560 5580 18570 5640
rect 18750 5580 18760 5640
rect 18560 5570 18760 5580
rect 19220 5640 19420 5650
rect 19220 5580 19230 5640
rect 19410 5580 19420 5640
rect 19220 5570 19420 5580
rect 17900 5430 18100 5510
rect 18560 5430 18760 5510
rect 19220 5430 19420 5510
rect 2010 5110 2090 5230
rect 2010 5050 2020 5110
rect 2080 5050 2090 5110
rect 2010 5040 2090 5050
rect 2230 5040 2310 5230
rect 4210 5220 4290 5230
rect 4210 5160 4220 5220
rect 4280 5160 4290 5220
rect 4210 5110 4290 5160
rect 4210 5050 4220 5110
rect 4280 5050 4290 5110
rect 4210 5040 4290 5050
rect 4430 5040 4510 5230
rect 6410 5220 6490 5230
rect 6410 5160 6420 5220
rect 6480 5160 6490 5220
rect 6410 5040 6490 5160
rect 6630 5110 6710 5230
rect 6630 5050 6640 5110
rect 6700 5050 6710 5110
rect 6630 5040 6710 5050
rect 8610 5040 8690 5230
rect 8830 5220 8910 5230
rect 8830 5160 8840 5220
rect 8900 5160 8910 5220
rect 8830 5110 8910 5160
rect 8830 5050 8840 5110
rect 8900 5050 8910 5110
rect 8830 5040 8910 5050
rect 10810 5040 10890 5230
rect 11030 5220 11110 5230
rect 11030 5160 11040 5220
rect 11100 5160 11110 5220
rect 11030 5110 11110 5160
rect 11030 5050 11040 5110
rect 11100 5050 11110 5110
rect 11030 5040 11110 5050
rect 13010 5040 13090 5230
rect 13230 5220 13310 5230
rect 13230 5160 13240 5220
rect 13300 5160 13310 5220
rect 13230 5110 13310 5160
rect 13230 5050 13240 5110
rect 13300 5050 13310 5110
rect 13230 5040 13310 5050
rect 15210 5110 15290 5230
rect 15210 5050 15220 5110
rect 15280 5050 15290 5110
rect 15210 5040 15290 5050
rect 15430 5220 15510 5230
rect 15430 5160 15440 5220
rect 15500 5160 15510 5220
rect 15430 5040 15510 5160
rect 17410 5220 17490 5230
rect 17410 5160 17420 5220
rect 17480 5160 17490 5220
rect 17410 5110 17490 5160
rect 17410 5050 17420 5110
rect 17480 5050 17490 5110
rect 17410 5040 17490 5050
rect 17630 5040 17710 5230
rect 19620 5210 19680 5840
rect 19730 5330 19790 5340
rect 19730 5260 19790 5270
rect 19840 5210 19900 5840
rect 19610 5200 19690 5210
rect 19610 5140 19620 5200
rect 19680 5140 19690 5200
rect 19610 5040 19690 5140
rect 19830 5040 19910 5210
rect 2020 4830 2080 5040
rect 2240 4830 2300 5040
rect 2500 5010 4020 5020
rect 2500 4950 2510 5010
rect 4010 4950 4020 5010
rect 2500 4940 4020 4950
rect 4220 4830 4280 5040
rect 4440 4830 4500 5040
rect 4700 5010 6220 5020
rect 4700 4950 4710 5010
rect 6210 4950 6220 5010
rect 4700 4940 6220 4950
rect 6420 4830 6480 5040
rect 6640 4830 6700 5040
rect 6900 5010 8420 5020
rect 6900 4950 6910 5010
rect 8410 4950 8420 5010
rect 6900 4940 8420 4950
rect 7790 4680 7950 4690
rect 7790 4540 7800 4680
rect 7940 4540 7950 4680
rect 7790 4530 7950 4540
rect 1620 4130 1820 4140
rect 1620 3950 1630 4130
rect 1810 3950 1820 4130
rect 1620 3940 1820 3950
rect 1160 3330 1340 3340
rect 1160 3150 1170 3330
rect 1330 3150 1340 3330
rect 1160 3140 1340 3150
rect 2760 3330 2940 3340
rect 2760 3150 2770 3330
rect 2930 3150 2940 3330
rect 2760 3140 2940 3150
rect 4360 3330 4540 3340
rect 4360 3150 4370 3330
rect 4530 3150 4540 3330
rect 4360 3140 4540 3150
rect 5960 3330 6140 3340
rect 5960 3150 5970 3330
rect 6130 3150 6140 3330
rect 5960 3140 6140 3150
rect 7560 3330 7740 3340
rect 7560 3150 7570 3330
rect 7730 3150 7740 3330
rect 7560 3140 7740 3150
rect 470 2220 670 2240
rect 470 -4780 480 2220
rect 660 -4780 670 2220
rect 1200 690 1300 3140
rect 2100 2250 2240 2260
rect 2100 2090 2110 2250
rect 2230 2090 2240 2250
rect 2100 1990 2240 2090
rect 2100 1310 2110 1990
rect 2230 1310 2240 1990
rect 1420 1160 1520 1180
rect 1400 1150 1540 1160
rect 1400 1030 1410 1150
rect 1530 1030 1540 1150
rect 1400 1020 1540 1030
rect 1180 680 1320 690
rect 1180 560 1190 680
rect 1310 560 1320 680
rect 1180 550 1320 560
rect 1200 -1110 1300 550
rect 1420 -640 1520 1020
rect 2100 450 2240 1310
rect 2800 690 2900 3140
rect 3700 2250 3840 2260
rect 3700 2090 3710 2250
rect 3830 2090 3840 2250
rect 3700 1990 3840 2090
rect 3700 1310 3710 1990
rect 3830 1310 3840 1990
rect 3020 1160 3120 1180
rect 3000 1150 3140 1160
rect 3000 1030 3010 1150
rect 3130 1030 3140 1150
rect 3000 1020 3140 1030
rect 2780 680 2920 690
rect 2780 560 2790 680
rect 2910 560 2920 680
rect 2780 550 2920 560
rect 2100 290 2110 450
rect 2230 290 2240 450
rect 2100 190 2240 290
rect 2100 -490 2110 190
rect 2230 -490 2240 190
rect 1400 -650 1540 -640
rect 1400 -770 1410 -650
rect 1530 -770 1540 -650
rect 1400 -780 1540 -770
rect 1180 -1120 1320 -1110
rect 1180 -1240 1190 -1120
rect 1310 -1240 1320 -1120
rect 1180 -1250 1320 -1240
rect 1200 -2910 1300 -1250
rect 1420 -2440 1520 -780
rect 2100 -1350 2240 -490
rect 2800 -1110 2900 550
rect 3020 -640 3120 1020
rect 3700 450 3840 1310
rect 4400 690 4500 3140
rect 5300 2250 5440 2260
rect 5300 2090 5310 2250
rect 5430 2090 5440 2250
rect 5300 1990 5440 2090
rect 5300 1310 5310 1990
rect 5430 1310 5440 1990
rect 4620 1160 4720 1180
rect 4600 1150 4740 1160
rect 4600 1030 4610 1150
rect 4730 1030 4740 1150
rect 4600 1020 4740 1030
rect 4380 680 4520 690
rect 4380 560 4390 680
rect 4510 560 4520 680
rect 4380 550 4520 560
rect 3700 290 3710 450
rect 3830 290 3840 450
rect 3700 190 3840 290
rect 3700 -490 3710 190
rect 3830 -490 3840 190
rect 3000 -650 3140 -640
rect 3000 -770 3010 -650
rect 3130 -770 3140 -650
rect 3000 -780 3140 -770
rect 2780 -1120 2920 -1110
rect 2780 -1240 2790 -1120
rect 2910 -1240 2920 -1120
rect 2780 -1250 2920 -1240
rect 2100 -1510 2110 -1350
rect 2230 -1510 2240 -1350
rect 2100 -1610 2240 -1510
rect 2100 -2290 2110 -1610
rect 2230 -2290 2240 -1610
rect 1400 -2450 1540 -2440
rect 1400 -2570 1410 -2450
rect 1530 -2570 1540 -2450
rect 1400 -2580 1540 -2570
rect 1180 -2920 1320 -2910
rect 1180 -3040 1190 -2920
rect 1310 -3040 1320 -2920
rect 1180 -3050 1320 -3040
rect 1200 -4710 1300 -3050
rect 1420 -4240 1520 -2580
rect 2100 -3150 2240 -2290
rect 2800 -2910 2900 -1250
rect 3020 -2440 3120 -780
rect 3700 -1350 3840 -490
rect 4400 -1110 4500 550
rect 4620 -640 4720 1020
rect 5300 450 5440 1310
rect 6000 690 6100 3140
rect 6900 2250 7040 2260
rect 6900 2090 6910 2250
rect 7030 2090 7040 2250
rect 6900 1990 7040 2090
rect 6900 1310 6910 1990
rect 7030 1310 7040 1990
rect 6220 1160 6320 1180
rect 6200 1150 6340 1160
rect 6200 1030 6210 1150
rect 6330 1030 6340 1150
rect 6200 1020 6340 1030
rect 5980 680 6120 690
rect 5980 560 5990 680
rect 6110 560 6120 680
rect 5980 550 6120 560
rect 5300 290 5310 450
rect 5430 290 5440 450
rect 5300 190 5440 290
rect 5300 -490 5310 190
rect 5430 -490 5440 190
rect 4600 -650 4740 -640
rect 4600 -770 4610 -650
rect 4730 -770 4740 -650
rect 4600 -780 4740 -770
rect 4380 -1120 4520 -1110
rect 4380 -1240 4390 -1120
rect 4510 -1240 4520 -1120
rect 4380 -1250 4520 -1240
rect 3700 -1510 3710 -1350
rect 3830 -1510 3840 -1350
rect 3700 -1610 3840 -1510
rect 3700 -2290 3710 -1610
rect 3830 -2290 3840 -1610
rect 3000 -2450 3140 -2440
rect 3000 -2570 3010 -2450
rect 3130 -2570 3140 -2450
rect 3000 -2580 3140 -2570
rect 2780 -2920 2920 -2910
rect 2780 -3040 2790 -2920
rect 2910 -3040 2920 -2920
rect 2780 -3050 2920 -3040
rect 2100 -3310 2110 -3150
rect 2230 -3310 2240 -3150
rect 2100 -3410 2240 -3310
rect 2100 -4090 2110 -3410
rect 2230 -4090 2240 -3410
rect 2100 -4100 2240 -4090
rect 1400 -4250 1540 -4240
rect 1400 -4370 1410 -4250
rect 1530 -4370 1540 -4250
rect 1400 -4380 1540 -4370
rect 1420 -4400 1520 -4380
rect 2800 -4710 2900 -3050
rect 3020 -4240 3120 -2580
rect 3700 -3150 3840 -2290
rect 4400 -2910 4500 -1250
rect 4620 -2440 4720 -780
rect 5300 -1350 5440 -490
rect 6000 -1110 6100 550
rect 6220 -640 6320 1020
rect 6900 450 7040 1310
rect 7600 690 7700 3140
rect 7820 2940 7920 4530
rect 8620 4430 8680 5040
rect 8840 4430 8900 5040
rect 9100 5010 10620 5020
rect 9100 4950 9110 5010
rect 10610 4950 10620 5010
rect 9100 4940 10620 4950
rect 10820 4430 10880 5040
rect 11040 4430 11100 5040
rect 11300 5010 12820 5020
rect 11300 4950 11310 5010
rect 12810 4950 12820 5010
rect 11300 4940 12820 4950
rect 13020 4430 13080 5040
rect 13240 4430 13300 5040
rect 13500 5010 15020 5020
rect 13500 4950 13510 5010
rect 15010 4950 15020 5010
rect 13500 4940 15020 4950
rect 15220 4830 15280 5040
rect 15440 4830 15500 5040
rect 15700 5010 17220 5020
rect 15700 4950 15710 5010
rect 17210 4950 17220 5010
rect 15700 4940 17220 4950
rect 17420 4830 17480 5040
rect 17640 4830 17700 5040
rect 17900 5010 19420 5020
rect 17900 4950 17910 5010
rect 19410 4950 19420 5010
rect 17900 4940 19420 4950
rect 19620 4830 19680 5040
rect 19840 4830 19900 5040
rect 20240 4540 20300 6740
rect 20100 4530 20300 4540
rect 8610 4310 8690 4430
rect 8610 4250 8620 4310
rect 8680 4250 8690 4310
rect 8610 4240 8690 4250
rect 8830 4240 8910 4430
rect 10810 4420 10890 4430
rect 10810 4360 10820 4420
rect 10880 4360 10890 4420
rect 10810 4240 10890 4360
rect 11030 4310 11110 4430
rect 11030 4250 11040 4310
rect 11100 4250 11110 4310
rect 11030 4240 11110 4250
rect 13010 4240 13090 4430
rect 13230 4420 13310 4430
rect 13230 4360 13240 4420
rect 13300 4360 13310 4420
rect 13230 4240 13310 4360
rect 20100 4350 20110 4530
rect 20290 4350 20300 4530
rect 20100 4340 20300 4350
rect 8620 4230 8680 4240
rect 8840 4230 8900 4240
rect 10820 4230 10880 4240
rect 11040 4230 11100 4240
rect 13020 4230 13080 4240
rect 13240 4230 13300 4240
rect 20440 4140 20500 7540
rect 21300 7390 21500 7400
rect 21300 7310 21310 7390
rect 21490 7310 21500 7390
rect 21300 7300 21500 7310
rect 21930 6930 21990 6940
rect 21930 6860 21990 6870
rect 21300 6590 21500 6600
rect 21300 6510 21310 6590
rect 21490 6510 21500 6590
rect 21300 6500 21500 6510
rect 21930 6130 21990 6140
rect 21930 6060 21990 6070
rect 21930 5330 21990 5340
rect 21930 5260 21990 5270
rect 23040 4970 23590 4980
rect 23040 4600 23050 4970
rect 23580 4600 23590 4970
rect 23040 4590 23590 4600
rect 20440 4130 20640 4140
rect 10880 4100 11040 4110
rect 10880 3960 10890 4100
rect 11030 3960 11040 4100
rect 10880 3950 11040 3960
rect 20440 3950 20450 4130
rect 20630 3950 20640 4130
rect 9160 3330 9340 3340
rect 9160 3150 9170 3330
rect 9330 3150 9340 3330
rect 9160 3140 9340 3150
rect 7800 2930 7940 2940
rect 7800 2810 7810 2930
rect 7930 2810 7940 2930
rect 7820 2540 7920 2810
rect 8500 2250 8640 2260
rect 8500 2090 8510 2250
rect 8630 2090 8640 2250
rect 8500 1990 8640 2090
rect 8500 1310 8510 1990
rect 8630 1310 8640 1990
rect 7820 1160 7920 1180
rect 7800 1150 7940 1160
rect 7800 1030 7810 1150
rect 7930 1030 7940 1150
rect 7800 1020 7940 1030
rect 7580 680 7720 690
rect 7580 560 7590 680
rect 7710 560 7720 680
rect 7580 550 7720 560
rect 6900 290 6910 450
rect 7030 290 7040 450
rect 6900 190 7040 290
rect 6900 -490 6910 190
rect 7030 -490 7040 190
rect 6200 -650 6340 -640
rect 6200 -770 6210 -650
rect 6330 -770 6340 -650
rect 6200 -780 6340 -770
rect 5980 -1120 6120 -1110
rect 5980 -1240 5990 -1120
rect 6110 -1240 6120 -1120
rect 5980 -1250 6120 -1240
rect 5300 -1510 5310 -1350
rect 5430 -1510 5440 -1350
rect 5300 -1610 5440 -1510
rect 5300 -2290 5310 -1610
rect 5430 -2290 5440 -1610
rect 4600 -2450 4740 -2440
rect 4600 -2570 4610 -2450
rect 4730 -2570 4740 -2450
rect 4600 -2580 4740 -2570
rect 4380 -2920 4520 -2910
rect 4380 -3040 4390 -2920
rect 4510 -3040 4520 -2920
rect 4380 -3050 4520 -3040
rect 3700 -3310 3710 -3150
rect 3830 -3310 3840 -3150
rect 3700 -3410 3840 -3310
rect 3700 -4090 3710 -3410
rect 3830 -4090 3840 -3410
rect 3700 -4100 3840 -4090
rect 3000 -4250 3140 -4240
rect 3000 -4370 3010 -4250
rect 3130 -4370 3140 -4250
rect 3000 -4380 3140 -4370
rect 3020 -4400 3120 -4380
rect 4400 -4710 4500 -3050
rect 4620 -4240 4720 -2580
rect 5300 -3150 5440 -2290
rect 6000 -2910 6100 -1250
rect 6220 -2440 6320 -780
rect 6900 -1350 7040 -490
rect 7600 -1110 7700 550
rect 7820 -640 7920 1020
rect 8500 450 8640 1310
rect 9200 690 9300 3140
rect 10910 3020 11010 3950
rect 20440 3940 20640 3950
rect 23210 3090 23410 4590
rect 26590 3360 26790 11490
rect 27250 11400 27260 11490
rect 27320 11400 27330 11490
rect 27250 11390 27330 11400
rect 27260 11180 27320 11390
rect 27250 11170 27330 11180
rect 27250 11080 27260 11170
rect 27320 11080 27330 11170
rect 27250 11070 27330 11080
rect 27260 10865 27320 11070
rect 27250 10855 27330 10865
rect 27250 10765 27260 10855
rect 27320 10765 27330 10855
rect 27250 10755 27330 10765
rect 27260 9415 27320 10755
rect 27380 10300 27440 11480
rect 27370 10290 27450 10300
rect 27370 10200 27380 10290
rect 27440 10200 27450 10290
rect 27370 10190 27450 10200
rect 27380 9985 27440 10190
rect 27370 9975 27450 9985
rect 27370 9885 27380 9975
rect 27440 9885 27450 9975
rect 27370 9875 27450 9885
rect 27250 9405 27330 9415
rect 27250 9315 27260 9405
rect 27320 9315 27330 9405
rect 27250 9305 27330 9315
rect 27260 9100 27320 9305
rect 27250 9090 27330 9100
rect 27250 9000 27260 9090
rect 27320 9000 27330 9090
rect 27250 8990 27330 9000
rect 27260 8785 27320 8990
rect 27250 8775 27330 8785
rect 27250 8685 27260 8775
rect 27320 8685 27330 8775
rect 27250 8675 27330 8685
rect 27260 8380 27320 8675
rect 27250 8370 27330 8380
rect 27250 8280 27260 8370
rect 27320 8280 27330 8370
rect 27250 8270 27330 8280
rect 27260 8060 27320 8270
rect 27250 8050 27330 8060
rect 27250 7960 27260 8050
rect 27320 7960 27330 8050
rect 27250 7950 27330 7960
rect 27260 7750 27320 7950
rect 27250 7740 27330 7750
rect 27250 7650 27260 7740
rect 27320 7650 27330 7740
rect 27250 7640 27330 7650
rect 27260 5250 27320 7640
rect 27380 7340 27440 9875
rect 27500 9260 27560 11480
rect 27490 9250 27570 9260
rect 27490 9160 27500 9250
rect 27560 9160 27570 9250
rect 27490 9150 27570 9160
rect 27500 8945 27560 9150
rect 27490 8935 27570 8945
rect 27490 8845 27500 8935
rect 27560 8845 27570 8935
rect 27490 8835 27570 8845
rect 27370 7330 27450 7340
rect 27370 7240 27380 7330
rect 27440 7240 27450 7330
rect 27370 7230 27450 7240
rect 27380 7025 27440 7230
rect 27370 7015 27450 7025
rect 27370 6925 27380 7015
rect 27440 6925 27450 7015
rect 27370 6915 27450 6925
rect 27380 6710 27440 6915
rect 27370 6700 27450 6710
rect 27370 6610 27380 6700
rect 27440 6610 27450 6700
rect 27370 6600 27450 6610
rect 27380 6300 27440 6600
rect 27370 6290 27450 6300
rect 27370 6200 27380 6290
rect 27440 6200 27450 6290
rect 27370 6190 27450 6200
rect 27380 5985 27440 6190
rect 27500 6140 27560 8835
rect 27620 8220 27680 11480
rect 27740 11340 27800 11480
rect 27730 11330 27810 11340
rect 27730 11240 27740 11330
rect 27800 11240 27810 11330
rect 36980 11300 36990 11680
rect 37050 11300 37060 11680
rect 36980 11290 37060 11300
rect 37400 11680 37480 11690
rect 37400 11300 37410 11680
rect 37470 11300 37480 11680
rect 37400 11290 37480 11300
rect 37820 11680 37900 11690
rect 37820 11300 37830 11680
rect 37890 11300 37900 11680
rect 37820 11290 37900 11300
rect 27730 11230 27810 11240
rect 29260 11280 29340 11290
rect 27740 11025 27800 11230
rect 29260 11060 29270 11280
rect 29330 11060 29340 11280
rect 29260 11050 29340 11060
rect 30802 11060 31214 11082
rect 27730 11015 27810 11025
rect 27730 10925 27740 11015
rect 27800 10925 27810 11015
rect 27730 10915 27810 10925
rect 27740 10460 27800 10915
rect 29270 10800 29330 11050
rect 30802 10934 30824 11060
rect 31194 10934 31214 11060
rect 30802 10876 31214 10934
rect 29270 10790 29520 10800
rect 29270 10720 29280 10790
rect 29510 10720 29520 10790
rect 29270 10710 29520 10720
rect 28950 10640 29200 10650
rect 28950 10570 28960 10640
rect 29190 10570 29200 10640
rect 28950 10560 29200 10570
rect 28860 10480 28940 10490
rect 27730 10450 27810 10460
rect 27730 10360 27740 10450
rect 27800 10360 27810 10450
rect 27730 10350 27810 10360
rect 27740 10140 27800 10350
rect 28860 10310 28870 10480
rect 28930 10310 28940 10480
rect 28860 10300 28940 10310
rect 27730 10130 27810 10140
rect 27730 10040 27740 10130
rect 27800 10040 27810 10130
rect 27730 10030 27810 10040
rect 27740 9825 27800 10030
rect 27730 9815 27810 9825
rect 27730 9725 27740 9815
rect 27800 9725 27810 9815
rect 27730 9715 27810 9725
rect 28880 9170 28940 10300
rect 29010 10340 29090 10350
rect 29010 10170 29020 10340
rect 29080 10170 29090 10340
rect 29140 10200 29200 10560
rect 29010 10160 29090 10170
rect 29130 10190 29210 10200
rect 28870 9160 28950 9170
rect 28870 8940 28880 9160
rect 28940 8940 28950 9160
rect 28870 8930 28950 8940
rect 27610 8210 27690 8220
rect 27610 8120 27620 8210
rect 27680 8120 27690 8210
rect 27610 8110 27690 8120
rect 27620 7900 27680 8110
rect 27610 7890 27690 7900
rect 27610 7800 27620 7890
rect 27680 7800 27690 7890
rect 27610 7790 27690 7800
rect 27620 7180 27680 7790
rect 27610 7170 27690 7180
rect 27610 7080 27620 7170
rect 27680 7080 27690 7170
rect 28880 7090 28940 8930
rect 29010 8120 29070 10160
rect 29130 9970 29140 10190
rect 29200 9970 29210 10190
rect 29130 9960 29210 9970
rect 29000 8110 29080 8120
rect 29000 7890 29010 8110
rect 29070 7890 29080 8110
rect 29000 7880 29080 7890
rect 27610 7070 27690 7080
rect 28870 7080 28950 7090
rect 27620 6865 27680 7070
rect 27610 6855 27690 6865
rect 27610 6765 27620 6855
rect 27680 6765 27690 6855
rect 28870 6860 28880 7080
rect 28940 6860 28950 7080
rect 28870 6850 28950 6860
rect 27610 6755 27690 6765
rect 27490 6130 27570 6140
rect 27490 6040 27500 6130
rect 27560 6040 27570 6130
rect 27490 6030 27570 6040
rect 27370 5975 27450 5985
rect 27370 5885 27380 5975
rect 27440 5885 27450 5975
rect 27370 5875 27450 5885
rect 27380 5670 27440 5875
rect 27500 5825 27560 6030
rect 27490 5815 27570 5825
rect 27490 5725 27500 5815
rect 27560 5725 27570 5815
rect 27490 5715 27570 5725
rect 27370 5660 27450 5670
rect 27370 5570 27380 5660
rect 27440 5570 27450 5660
rect 27370 5560 27450 5570
rect 27170 5240 27320 5250
rect 27170 5110 27180 5240
rect 27310 5110 27320 5240
rect 27170 5100 27320 5110
rect 27380 5000 27440 5560
rect 27240 4930 27440 5000
rect 27240 4750 27250 4930
rect 27430 4750 27440 4930
rect 27240 4740 27440 4750
rect 27500 4600 27560 5715
rect 27360 4530 27560 4600
rect 27360 4350 27370 4530
rect 27550 4350 27560 4530
rect 27360 4340 27560 4350
rect 27620 4200 27680 6755
rect 29010 6050 29070 7880
rect 29000 6040 29080 6050
rect 29000 5820 29010 6040
rect 29070 5820 29080 6040
rect 29000 5810 29080 5820
rect 29140 4530 29200 9960
rect 29130 4520 29210 4530
rect 29130 4290 29140 4520
rect 29200 4290 29210 4520
rect 29130 4280 29210 4290
rect 29270 4270 29330 10710
rect 30802 10346 30826 10876
rect 31190 10346 31214 10876
rect 34472 11038 34876 11042
rect 34472 11022 36808 11038
rect 34472 10846 34490 11022
rect 34848 10846 36808 11022
rect 37180 11010 37350 11020
rect 37180 10860 37190 11010
rect 37340 10860 37350 11010
rect 37180 10850 37350 10860
rect 37980 10960 38130 10970
rect 34472 10824 36808 10846
rect 34472 10822 34876 10824
rect 33510 10790 33770 10800
rect 33510 10720 33520 10790
rect 33760 10720 33770 10790
rect 33510 10710 33770 10720
rect 32470 10630 32730 10640
rect 32470 10560 32480 10630
rect 32720 10560 32730 10630
rect 33540 10586 33620 10710
rect 32470 10550 32730 10560
rect 31670 10490 31930 10500
rect 31670 10420 31680 10490
rect 31920 10420 31930 10490
rect 31670 10410 31930 10420
rect 30802 10322 31214 10346
rect 31320 10350 31580 10360
rect 31320 10280 31330 10350
rect 31570 10280 31580 10350
rect 31320 10270 31580 10280
rect 31414 10262 31502 10270
rect 31414 10082 31422 10262
rect 31494 10082 31502 10262
rect 31414 10074 31502 10082
rect 31748 10262 31834 10410
rect 32554 10280 32634 10550
rect 33354 10506 33620 10586
rect 33354 10280 33434 10506
rect 31748 10082 31756 10262
rect 31828 10082 31834 10262
rect 31748 10076 31834 10082
rect 32548 10262 32634 10280
rect 32548 10082 32556 10262
rect 32628 10082 32634 10262
rect 32548 10076 32634 10082
rect 33348 10262 33434 10280
rect 33348 10082 33356 10262
rect 33428 10082 33434 10262
rect 36410 10434 36808 10824
rect 37980 10780 37990 10960
rect 38120 10780 38130 10960
rect 37980 10770 38130 10780
rect 37600 10750 37770 10760
rect 37600 10600 37610 10750
rect 37760 10600 37770 10750
rect 37600 10590 37770 10600
rect 36980 10500 37060 10510
rect 36980 10434 36990 10500
rect 36410 10320 36990 10434
rect 37050 10434 37060 10500
rect 37400 10500 37480 10510
rect 37400 10434 37410 10500
rect 37050 10320 37410 10434
rect 37470 10434 37480 10500
rect 37820 10500 37900 10510
rect 37820 10434 37830 10500
rect 37470 10320 37830 10434
rect 37890 10434 37900 10500
rect 37890 10406 39308 10434
rect 37890 10320 38298 10406
rect 36410 10160 38298 10320
rect 33348 10076 33434 10082
rect 33354 10074 33434 10076
rect 35020 10140 36340 10150
rect 35020 10070 35820 10140
rect 36010 10070 36140 10140
rect 36330 10070 36340 10140
rect 35020 10060 36340 10070
rect 30510 8290 30650 8300
rect 30510 8170 30520 8290
rect 30640 8170 30650 8290
rect 30510 8160 30650 8170
rect 30540 4880 30620 8160
rect 30900 8090 31040 8100
rect 30900 7970 30910 8090
rect 31030 7970 31040 8090
rect 30900 7960 31040 7970
rect 30930 4880 31010 7960
rect 31280 7210 31580 7220
rect 31280 7090 31290 7210
rect 31570 7180 31580 7210
rect 31570 7120 32180 7180
rect 31570 7090 31580 7120
rect 31280 7080 31580 7090
rect 30510 4870 30650 4880
rect 30510 4750 30520 4870
rect 30640 4750 30650 4870
rect 30510 4740 30650 4750
rect 30900 4870 31040 4880
rect 30900 4750 30910 4870
rect 31030 4750 31040 4870
rect 30900 4740 31040 4750
rect 29270 4260 29520 4270
rect 27620 4130 27820 4200
rect 29270 4190 29280 4260
rect 29510 4190 29520 4260
rect 29270 4180 29520 4190
rect 27620 3950 27630 4130
rect 27810 3950 27820 4130
rect 27620 3940 27820 3950
rect 30070 4040 30270 4050
rect 30070 3860 30080 4040
rect 30260 3860 30270 4040
rect 30070 3850 30270 3860
rect 31670 4040 31870 4050
rect 31670 3860 31680 4040
rect 31860 3860 31870 4040
rect 31670 3850 31870 3860
rect 32090 3750 32180 7120
rect 35020 5370 35120 10060
rect 36410 9980 36950 10160
rect 37080 9980 37370 10160
rect 37500 9980 37790 10160
rect 37920 9980 38298 10160
rect 36410 9970 38298 9980
rect 36410 9924 36560 9970
rect 35250 9664 35394 9676
rect 35250 9542 35266 9664
rect 35384 9542 35394 9664
rect 35250 9526 35394 9542
rect 35268 8426 35352 9526
rect 36410 9434 36430 9924
rect 36542 9434 36560 9924
rect 38268 9848 38298 9970
rect 39274 9970 39308 10406
rect 39274 9848 39306 9970
rect 38268 9822 39306 9848
rect 37572 9664 37716 9680
rect 37572 9542 37584 9664
rect 37702 9542 37716 9664
rect 37572 9530 37716 9542
rect 36410 9406 36560 9434
rect 37622 8428 37706 9530
rect 35238 8414 35384 8426
rect 35238 8292 35254 8414
rect 35372 8292 35384 8414
rect 35238 8280 35384 8292
rect 37586 8416 37732 8428
rect 37586 8294 37600 8416
rect 37718 8294 37732 8416
rect 37586 8282 37732 8294
rect 35360 7920 35500 7930
rect 35360 7800 35370 7920
rect 35490 7900 35500 7920
rect 36870 7920 37010 7930
rect 36870 7900 36880 7920
rect 35490 7820 36880 7900
rect 35490 7800 35500 7820
rect 35360 7790 35500 7800
rect 36870 7800 36880 7820
rect 37000 7800 37010 7920
rect 36870 7790 37010 7800
rect 35340 7690 35480 7700
rect 35340 7570 35350 7690
rect 35470 7570 35480 7690
rect 35340 7560 35480 7570
rect 36000 7620 36140 7630
rect 36000 7500 36010 7620
rect 36130 7600 36140 7620
rect 37480 7620 37620 7630
rect 37480 7600 37494 7620
rect 36130 7520 37494 7600
rect 36130 7500 36140 7520
rect 36000 7490 36140 7500
rect 37480 7504 37494 7520
rect 37610 7504 37620 7620
rect 37480 7500 37620 7504
rect 37480 7490 37640 7500
rect 37500 7370 37510 7490
rect 37630 7370 37640 7490
rect 37500 7360 37640 7370
rect 36106 7176 36838 7200
rect 36106 6982 36128 7176
rect 36810 6982 36838 7176
rect 36106 6964 36838 6982
rect 36220 6260 36420 6270
rect 36220 6080 36230 6260
rect 36410 6080 36420 6260
rect 36220 6070 36420 6080
rect 36520 6260 36720 6270
rect 36520 6080 36530 6260
rect 36710 6080 36720 6260
rect 36520 6070 36720 6080
rect 34890 5360 35120 5370
rect 34890 5280 34900 5360
rect 35110 5280 35120 5360
rect 34890 5270 35120 5280
rect 36290 5890 36400 5900
rect 36290 5820 36300 5890
rect 36390 5820 36400 5890
rect 36290 5630 36400 5820
rect 36290 5560 36300 5630
rect 36390 5560 36400 5630
rect 36290 5370 36400 5560
rect 36290 5040 36300 5370
rect 36390 5040 36400 5370
rect 36290 4850 36400 5040
rect 36290 4780 36300 4850
rect 36390 4780 36400 4850
rect 36290 4590 36400 4780
rect 36290 4520 36300 4590
rect 36390 4520 36400 4590
rect 32490 4480 32650 4490
rect 32490 4340 32500 4480
rect 32640 4340 32650 4480
rect 32490 4330 32650 4340
rect 34080 4480 34240 4490
rect 34080 4340 34090 4480
rect 34230 4340 34240 4480
rect 34080 4330 34240 4340
rect 36290 4330 36400 4520
rect 32070 3740 32220 3750
rect 31520 3730 31700 3740
rect 31520 3550 31530 3730
rect 31690 3550 31700 3730
rect 32070 3610 32080 3740
rect 32210 3610 32220 3740
rect 32070 3600 32220 3610
rect 31520 3540 31700 3550
rect 26590 3220 26620 3360
rect 26760 3220 26790 3360
rect 26590 3210 26790 3220
rect 14180 3030 14360 3040
rect 10880 3010 11040 3020
rect 10880 2870 10890 3010
rect 11030 2870 11040 3010
rect 10880 2860 11040 2870
rect 14180 2870 14190 3030
rect 14350 2870 14360 3030
rect 14180 2860 14360 2870
rect 18050 3010 18210 3020
rect 18050 2870 18060 3010
rect 18200 2870 18210 3010
rect 23210 2910 23220 3090
rect 23400 2910 23410 3090
rect 23210 2900 23410 2910
rect 18050 2860 18210 2870
rect 11690 2770 11850 2780
rect 11690 2620 11700 2770
rect 11840 2620 11850 2770
rect 11690 2610 11850 2620
rect 10990 2540 11150 2550
rect 10990 2400 11000 2540
rect 11140 2400 11150 2540
rect 10990 2390 11150 2400
rect 10100 2250 10240 2260
rect 10100 2090 10110 2250
rect 10230 2090 10240 2250
rect 10100 1990 10240 2090
rect 10100 1310 10110 1990
rect 10230 1310 10240 1990
rect 11020 1960 11120 2390
rect 11700 2250 11840 2610
rect 12590 2540 12750 2550
rect 12590 2400 12600 2540
rect 12740 2400 12750 2540
rect 12590 2390 12750 2400
rect 13970 2540 14130 2550
rect 13970 2400 13980 2540
rect 14120 2400 14130 2540
rect 13970 2390 14130 2400
rect 11700 2090 11710 2250
rect 11830 2090 11840 2250
rect 11020 1950 11160 1960
rect 11020 1330 11030 1950
rect 11150 1330 11160 1950
rect 11020 1320 11160 1330
rect 9420 1160 9520 1180
rect 9400 1150 9540 1160
rect 9400 1030 9410 1150
rect 9530 1030 9540 1150
rect 9400 1020 9540 1030
rect 9180 680 9320 690
rect 9180 560 9190 680
rect 9310 560 9320 680
rect 9180 550 9320 560
rect 8500 290 8510 450
rect 8630 290 8640 450
rect 8500 190 8640 290
rect 8500 -490 8510 190
rect 8630 -490 8640 190
rect 7800 -650 7940 -640
rect 7800 -770 7810 -650
rect 7930 -770 7940 -650
rect 7800 -780 7940 -770
rect 7580 -1120 7720 -1110
rect 7580 -1240 7590 -1120
rect 7710 -1240 7720 -1120
rect 7580 -1250 7720 -1240
rect 6900 -1510 6910 -1350
rect 7030 -1510 7040 -1350
rect 6900 -1610 7040 -1510
rect 6900 -2290 6910 -1610
rect 7030 -2290 7040 -1610
rect 6200 -2450 6340 -2440
rect 6200 -2570 6210 -2450
rect 6330 -2570 6340 -2450
rect 6200 -2580 6340 -2570
rect 5980 -2920 6120 -2910
rect 5980 -3040 5990 -2920
rect 6110 -3040 6120 -2920
rect 5980 -3050 6120 -3040
rect 5300 -3310 5310 -3150
rect 5430 -3310 5440 -3150
rect 5300 -3410 5440 -3310
rect 5300 -4090 5310 -3410
rect 5430 -4090 5440 -3410
rect 5300 -4100 5440 -4090
rect 4600 -4250 4740 -4240
rect 4600 -4370 4610 -4250
rect 4730 -4370 4740 -4250
rect 4600 -4380 4740 -4370
rect 4620 -4400 4720 -4380
rect 6000 -4710 6100 -3050
rect 6220 -4240 6320 -2580
rect 6900 -3150 7040 -2290
rect 7600 -2910 7700 -1250
rect 7820 -2440 7920 -780
rect 8500 -1350 8640 -490
rect 9200 -1110 9300 550
rect 9420 -640 9520 1020
rect 10100 450 10240 1310
rect 11700 1240 11840 2090
rect 12620 1960 12720 2390
rect 13300 2250 13440 2260
rect 13300 2090 13310 2250
rect 13430 2090 13440 2250
rect 12600 1950 12740 1960
rect 12600 1330 12610 1950
rect 12730 1330 12740 1950
rect 12600 1320 12740 1330
rect 11240 1230 11840 1240
rect 11240 1070 11250 1230
rect 11670 1070 11840 1230
rect 11240 1060 11840 1070
rect 10100 290 10110 450
rect 10230 290 10240 450
rect 10100 190 10240 290
rect 10100 -490 10110 190
rect 10230 -490 10240 190
rect 9400 -650 9540 -640
rect 9400 -770 9410 -650
rect 9530 -770 9540 -650
rect 9400 -780 9540 -770
rect 9180 -1120 9320 -1110
rect 9180 -1240 9190 -1120
rect 9310 -1240 9320 -1120
rect 9180 -1250 9320 -1240
rect 8500 -1510 8510 -1350
rect 8630 -1510 8640 -1350
rect 8500 -1610 8640 -1510
rect 8500 -2290 8510 -1610
rect 8630 -2290 8640 -1610
rect 7800 -2450 7940 -2440
rect 7800 -2570 7810 -2450
rect 7930 -2570 7940 -2450
rect 7800 -2580 7940 -2570
rect 7580 -2920 7720 -2910
rect 7580 -3040 7590 -2920
rect 7710 -3040 7720 -2920
rect 7580 -3050 7720 -3040
rect 6900 -3310 6910 -3150
rect 7030 -3310 7040 -3150
rect 6900 -3410 7040 -3310
rect 6900 -4090 6910 -3410
rect 7030 -4090 7040 -3410
rect 6900 -4100 7040 -4090
rect 6200 -4250 6340 -4240
rect 6200 -4370 6210 -4250
rect 6330 -4370 6340 -4250
rect 6200 -4380 6340 -4370
rect 6220 -4400 6320 -4380
rect 7600 -4710 7700 -3050
rect 7820 -4240 7920 -2580
rect 8500 -3150 8640 -2290
rect 9200 -2910 9300 -1250
rect 9420 -2440 9520 -780
rect 10100 -1350 10240 -490
rect 11700 450 11840 1060
rect 12380 870 12520 880
rect 12380 750 12390 870
rect 12510 750 12520 870
rect 12380 740 12520 750
rect 11700 290 11710 450
rect 11830 290 11840 450
rect 11700 190 11840 290
rect 11700 -560 11710 190
rect 11260 -570 11710 -560
rect 11830 -560 11840 190
rect 11830 -570 12280 -560
rect 11260 -730 11270 -570
rect 12270 -730 12280 -570
rect 12400 -640 12500 740
rect 11260 -740 12280 -730
rect 12380 -650 12520 -640
rect 10100 -1510 10110 -1350
rect 10230 -1510 10240 -1350
rect 10100 -1610 10240 -1510
rect 10100 -2290 10110 -1610
rect 10230 -2290 10240 -1610
rect 9400 -2450 9540 -2440
rect 9400 -2570 9410 -2450
rect 9530 -2570 9540 -2450
rect 9400 -2580 9540 -2570
rect 9180 -2920 9320 -2910
rect 9180 -3040 9190 -2920
rect 9310 -3040 9320 -2920
rect 9180 -3050 9320 -3040
rect 8500 -3310 8510 -3150
rect 8630 -3310 8640 -3150
rect 8500 -3410 8640 -3310
rect 8500 -4090 8510 -3410
rect 8630 -4090 8640 -3410
rect 8500 -4100 8640 -4090
rect 7800 -4250 7940 -4240
rect 7800 -4370 7810 -4250
rect 7930 -4370 7940 -4250
rect 7800 -4380 7940 -4370
rect 7820 -4400 7920 -4380
rect 9200 -4710 9300 -3050
rect 9420 -4240 9520 -2580
rect 10100 -3150 10240 -2290
rect 11700 -1350 11840 -740
rect 12380 -810 12390 -650
rect 12510 -810 12520 -650
rect 12380 -980 12520 -810
rect 12380 -1050 12390 -980
rect 12510 -1050 12520 -980
rect 12380 -1060 12520 -1050
rect 12620 -710 12720 1320
rect 13300 450 13440 2090
rect 14000 1960 14100 2390
rect 13980 1950 14120 1960
rect 13980 1330 13990 1950
rect 14110 1330 14120 1950
rect 13980 1320 14120 1330
rect 13300 290 13310 450
rect 13430 290 13440 450
rect 13300 190 13440 290
rect 13300 -490 13310 190
rect 13430 -490 13440 190
rect 12620 -920 12721 -710
rect 12620 -930 12760 -920
rect 11700 -1510 11710 -1350
rect 11830 -1510 11840 -1350
rect 11700 -1610 11840 -1510
rect 11700 -2290 11710 -1610
rect 11830 -2290 11840 -1610
rect 11020 -2910 11120 -2900
rect 11000 -2920 11140 -2910
rect 11000 -3040 11010 -2920
rect 11130 -3040 11140 -2920
rect 11000 -3050 11140 -3040
rect 10100 -3310 10110 -3150
rect 10230 -3310 10240 -3150
rect 10100 -3410 10240 -3310
rect 10100 -4090 10110 -3410
rect 10230 -4090 10240 -3410
rect 10100 -4100 10240 -4090
rect 9400 -4250 9540 -4240
rect 9400 -4370 9410 -4250
rect 9530 -4370 9540 -4250
rect 9400 -4380 9540 -4370
rect 9420 -4400 9520 -4380
rect 470 -4800 670 -4780
rect 1180 -4720 1320 -4710
rect 1180 -4840 1190 -4720
rect 1310 -4840 1320 -4720
rect 1180 -4850 1320 -4840
rect 2780 -4720 2920 -4710
rect 2780 -4840 2790 -4720
rect 2910 -4840 2920 -4720
rect 2780 -4850 2920 -4840
rect 4380 -4720 4520 -4710
rect 4380 -4840 4390 -4720
rect 4510 -4840 4520 -4720
rect 4380 -4850 4520 -4840
rect 5980 -4720 6120 -4710
rect 5980 -4840 5990 -4720
rect 6110 -4840 6120 -4720
rect 5980 -4850 6120 -4840
rect 7580 -4720 7720 -4710
rect 7580 -4840 7590 -4720
rect 7710 -4840 7720 -4720
rect 7580 -4850 7720 -4840
rect 9180 -4720 9320 -4710
rect 9180 -4840 9190 -4720
rect 9310 -4840 9320 -4720
rect 9180 -4850 9320 -4840
rect 11020 -4750 11120 -3050
rect 11700 -3150 11840 -2290
rect 12400 -2720 12500 -1060
rect 12620 -1070 12630 -930
rect 12750 -1070 12760 -930
rect 12620 -1100 12760 -1070
rect 12870 -1110 13250 -1100
rect 12870 -1260 12880 -1110
rect 13240 -1260 13250 -1110
rect 12870 -1270 13250 -1260
rect 13300 -1350 13440 -490
rect 14000 -920 14100 1320
rect 13960 -930 14100 -920
rect 13960 -1070 13970 -930
rect 14090 -1070 14100 -930
rect 13960 -1100 14100 -1070
rect 13300 -1510 13310 -1350
rect 13430 -1510 13440 -1350
rect 13300 -1610 13440 -1510
rect 13300 -2290 13310 -1610
rect 13430 -2290 13440 -1610
rect 12380 -2730 12520 -2720
rect 12380 -2850 12390 -2730
rect 12510 -2850 12520 -2730
rect 12380 -2860 12520 -2850
rect 11700 -3310 11710 -3150
rect 11830 -3310 11840 -3150
rect 11700 -3410 11840 -3310
rect 11700 -4090 11710 -3410
rect 11830 -4090 11840 -3410
rect 11700 -4100 11840 -4090
rect 12400 -4520 12500 -2860
rect 13300 -3150 13440 -2290
rect 14220 -2910 14320 2860
rect 16900 2780 17140 2790
rect 16900 2640 16910 2780
rect 17130 2640 17140 2780
rect 16900 2630 17140 2640
rect 17370 2780 17500 2790
rect 17370 2640 17380 2780
rect 17490 2640 17500 2780
rect 17370 2630 17500 2640
rect 17730 2780 17970 2790
rect 17730 2640 17740 2780
rect 17960 2640 17970 2780
rect 17730 2630 17970 2640
rect 16500 2250 16640 2260
rect 16500 2090 16510 2250
rect 16630 2090 16640 2250
rect 14900 1980 15040 2010
rect 14900 1320 14910 1980
rect 15030 1320 15040 1980
rect 14900 1240 15040 1320
rect 16500 1990 16640 2090
rect 16500 1310 16510 1990
rect 16630 1310 16640 1990
rect 18100 2250 18240 2260
rect 18100 2090 18110 2250
rect 18230 2090 18240 2250
rect 18100 1990 18240 2090
rect 18100 1310 18110 1990
rect 18230 1310 18240 1990
rect 19700 2250 19840 2260
rect 19700 2090 19710 2250
rect 19830 2090 19840 2250
rect 19700 1990 19840 2090
rect 19700 1310 19710 1990
rect 19830 1310 19840 1990
rect 21300 2250 21440 2260
rect 21300 2090 21310 2250
rect 21430 2090 21440 2250
rect 21300 1990 21440 2090
rect 21300 1310 21310 1990
rect 21430 1310 21440 1990
rect 22900 2250 23040 2260
rect 22900 2090 22910 2250
rect 23030 2090 23040 2250
rect 22900 1990 23040 2090
rect 22900 1310 22910 1990
rect 23030 1310 23040 1990
rect 24500 2250 24640 2260
rect 24500 2090 24510 2250
rect 24630 2090 24640 2250
rect 24500 1990 24640 2090
rect 24500 1310 24510 1990
rect 24630 1310 24640 1990
rect 26100 2250 26240 2260
rect 26100 2090 26110 2250
rect 26230 2090 26240 2250
rect 26100 1990 26240 2090
rect 26100 1310 26110 1990
rect 26230 1310 26240 1990
rect 27700 2250 27840 2260
rect 27700 2070 27710 2250
rect 27830 2070 27840 2250
rect 27700 1990 27840 2070
rect 27700 1310 27710 1990
rect 27830 1310 27840 1990
rect 29300 2250 29440 2260
rect 29300 2070 29310 2250
rect 29430 2070 29440 2250
rect 29300 1990 29440 2070
rect 29300 1310 29310 1990
rect 29430 1310 29440 1990
rect 15600 1160 15700 1310
rect 15590 1150 15710 1160
rect 15590 1030 15600 1150
rect 15700 1030 15710 1150
rect 15590 1020 15710 1030
rect 14900 190 15040 460
rect 14900 -560 14910 190
rect 14460 -570 14910 -560
rect 15030 -560 15040 190
rect 15030 -570 15480 -560
rect 14460 -730 14470 -570
rect 15470 -730 15480 -570
rect 15600 -640 15700 1020
rect 15820 690 15920 1310
rect 15810 680 15930 690
rect 15810 560 15820 680
rect 15920 560 15930 680
rect 15810 550 15930 560
rect 14460 -740 15480 -730
rect 15590 -650 15710 -640
rect 14900 -1350 15040 -1340
rect 14900 -1510 14910 -1350
rect 15030 -1510 15040 -1350
rect 14900 -1610 15040 -1510
rect 15240 -1350 15380 -740
rect 15590 -770 15600 -650
rect 15700 -770 15710 -650
rect 15590 -780 15710 -770
rect 15240 -1510 15250 -1350
rect 15370 -1510 15380 -1350
rect 15240 -1520 15380 -1510
rect 14900 -2290 14910 -1610
rect 15030 -2290 15040 -1610
rect 14200 -2920 14340 -2910
rect 14200 -3040 14210 -2920
rect 14330 -3040 14340 -2920
rect 14200 -3050 14340 -3040
rect 14420 -2920 14560 -2910
rect 14420 -3040 14430 -2920
rect 14550 -3040 14560 -2920
rect 14420 -3050 14560 -3040
rect 14440 -3110 14540 -3050
rect 12600 -3290 12740 -3280
rect 12600 -3390 12610 -3290
rect 12730 -3390 12740 -3290
rect 12600 -3400 12740 -3390
rect 13300 -3310 13310 -3150
rect 13430 -3310 13440 -3150
rect 12380 -4530 12520 -4520
rect 12380 -4650 12390 -4530
rect 12510 -4650 12520 -4530
rect 12380 -4660 12520 -4650
rect 12620 -4720 12720 -3400
rect 13300 -3410 13440 -3310
rect 13300 -4090 13310 -3410
rect 13430 -4090 13440 -3410
rect 13300 -4100 13440 -4090
rect 14000 -3220 14540 -3110
rect 14900 -3150 15040 -2290
rect 15600 -2440 15700 -780
rect 15820 -1110 15920 550
rect 16500 450 16640 1310
rect 17200 1160 17300 1310
rect 17190 1150 17310 1160
rect 17190 1030 17200 1150
rect 17300 1030 17310 1150
rect 17190 1020 17310 1030
rect 16500 290 16510 450
rect 16630 290 16640 450
rect 16500 190 16640 290
rect 16500 -490 16510 190
rect 16630 -490 16640 190
rect 15810 -1120 15930 -1110
rect 15810 -1240 15820 -1120
rect 15920 -1240 15930 -1120
rect 15810 -1250 15930 -1240
rect 15590 -2450 15710 -2440
rect 15590 -2570 15600 -2450
rect 15700 -2570 15710 -2450
rect 15590 -2580 15710 -2570
rect 12600 -4730 12740 -4720
rect 11020 -4850 11140 -4750
rect 1200 -4860 1300 -4850
rect 2800 -4880 2900 -4850
rect 4400 -4880 4500 -4850
rect 6000 -4880 6100 -4850
rect 7600 -4880 7700 -4850
rect 9200 -4880 9300 -4850
rect 80 -6330 90 -5750
rect 270 -6330 280 -5750
rect 80 -31730 280 -6330
rect 7800 -7870 7940 -7860
rect 7800 -7990 7810 -7870
rect 7930 -7990 7940 -7870
rect 7800 -8000 7940 -7990
rect 1220 -8060 1320 -8050
rect 1200 -8070 1340 -8060
rect 480 -8090 680 -8080
rect 480 -22380 490 -8090
rect 670 -22380 680 -8090
rect 1200 -8190 1210 -8070
rect 1330 -8190 1340 -8070
rect 1200 -8200 1340 -8190
rect 1220 -9860 1320 -8200
rect 1440 -8500 1540 -8050
rect 2820 -8060 2920 -8050
rect 2800 -8070 2940 -8060
rect 2800 -8190 2810 -8070
rect 2930 -8190 2940 -8070
rect 2800 -8200 2940 -8190
rect 1420 -8510 1560 -8500
rect 1420 -8630 1430 -8510
rect 1550 -8630 1560 -8510
rect 1420 -8640 1560 -8630
rect 1200 -9870 1340 -9860
rect 1200 -9990 1210 -9870
rect 1330 -9990 1340 -9870
rect 1200 -10000 1340 -9990
rect 1220 -11660 1320 -10000
rect 1440 -10300 1540 -8640
rect 2120 -8810 2240 -8780
rect 2120 -9470 2130 -8810
rect 2230 -9470 2240 -8810
rect 2120 -9590 2240 -9470
rect 2120 -9750 2130 -9590
rect 2230 -9750 2240 -9590
rect 1420 -10310 1560 -10300
rect 1420 -10430 1430 -10310
rect 1550 -10430 1560 -10310
rect 1420 -10440 1560 -10430
rect 1200 -11670 1340 -11660
rect 1200 -11790 1210 -11670
rect 1330 -11790 1340 -11670
rect 1200 -11800 1340 -11790
rect 1220 -13460 1320 -11800
rect 1440 -12100 1540 -10440
rect 2120 -10610 2240 -9750
rect 2820 -9860 2920 -8200
rect 3040 -8500 3140 -8050
rect 4420 -8060 4520 -8050
rect 4400 -8070 4540 -8060
rect 4400 -8190 4410 -8070
rect 4530 -8190 4540 -8070
rect 4400 -8200 4540 -8190
rect 3020 -8510 3160 -8500
rect 3020 -8630 3030 -8510
rect 3150 -8630 3160 -8510
rect 3020 -8640 3160 -8630
rect 2800 -9870 2940 -9860
rect 2800 -9990 2810 -9870
rect 2930 -9990 2940 -9870
rect 2800 -10000 2940 -9990
rect 2120 -11270 2130 -10610
rect 2230 -11270 2240 -10610
rect 2120 -11390 2240 -11270
rect 2120 -11550 2130 -11390
rect 2230 -11550 2240 -11390
rect 1420 -12110 1560 -12100
rect 1420 -12230 1430 -12110
rect 1550 -12230 1560 -12110
rect 1420 -12240 1560 -12230
rect 1200 -13470 1340 -13460
rect 1200 -13590 1210 -13470
rect 1330 -13590 1340 -13470
rect 1200 -13600 1340 -13590
rect 1220 -15260 1320 -13600
rect 1440 -13900 1540 -12240
rect 2120 -12410 2240 -11550
rect 2820 -11660 2920 -10000
rect 3040 -10300 3140 -8640
rect 3720 -8810 3840 -8780
rect 3720 -9470 3730 -8810
rect 3830 -9470 3840 -8810
rect 3720 -9590 3840 -9470
rect 3720 -9750 3730 -9590
rect 3830 -9750 3840 -9590
rect 3020 -10310 3160 -10300
rect 3020 -10430 3030 -10310
rect 3150 -10430 3160 -10310
rect 3020 -10440 3160 -10430
rect 2800 -11670 2940 -11660
rect 2800 -11790 2810 -11670
rect 2930 -11790 2940 -11670
rect 2800 -11800 2940 -11790
rect 2120 -13070 2130 -12410
rect 2230 -13070 2240 -12410
rect 2120 -13190 2240 -13070
rect 2120 -13350 2130 -13190
rect 2230 -13350 2240 -13190
rect 1420 -13910 1560 -13900
rect 1420 -14030 1430 -13910
rect 1550 -14030 1560 -13910
rect 1420 -14040 1560 -14030
rect 1200 -15270 1340 -15260
rect 1200 -15390 1210 -15270
rect 1330 -15390 1340 -15270
rect 1200 -15400 1340 -15390
rect 1220 -17060 1320 -15400
rect 1440 -15700 1540 -14040
rect 2120 -14210 2240 -13350
rect 2820 -13460 2920 -11800
rect 3040 -12100 3140 -10440
rect 3720 -10610 3840 -9750
rect 4420 -9860 4520 -8200
rect 4640 -8500 4740 -8050
rect 6020 -8060 6120 -8050
rect 6000 -8070 6140 -8060
rect 6000 -8190 6010 -8070
rect 6130 -8190 6140 -8070
rect 6000 -8200 6140 -8190
rect 4620 -8510 4760 -8500
rect 4620 -8630 4630 -8510
rect 4750 -8630 4760 -8510
rect 4620 -8640 4760 -8630
rect 4400 -9870 4540 -9860
rect 4400 -9990 4410 -9870
rect 4530 -9990 4540 -9870
rect 4400 -10000 4540 -9990
rect 3720 -11270 3730 -10610
rect 3830 -11270 3840 -10610
rect 3720 -11390 3840 -11270
rect 3720 -11550 3730 -11390
rect 3830 -11550 3840 -11390
rect 3020 -12110 3160 -12100
rect 3020 -12230 3030 -12110
rect 3150 -12230 3160 -12110
rect 3020 -12240 3160 -12230
rect 2800 -13470 2940 -13460
rect 2800 -13590 2810 -13470
rect 2930 -13590 2940 -13470
rect 2800 -13600 2940 -13590
rect 2120 -14870 2130 -14210
rect 2230 -14870 2240 -14210
rect 2120 -14990 2240 -14870
rect 2120 -15150 2130 -14990
rect 2230 -15150 2240 -14990
rect 1420 -15710 1560 -15700
rect 1420 -15830 1430 -15710
rect 1550 -15830 1560 -15710
rect 1420 -15840 1560 -15830
rect 1200 -17070 1340 -17060
rect 1200 -17190 1210 -17070
rect 1330 -17190 1340 -17070
rect 1200 -17200 1340 -17190
rect 1220 -18860 1320 -17200
rect 1440 -17500 1540 -15840
rect 2120 -16010 2240 -15150
rect 2820 -15260 2920 -13600
rect 3040 -13900 3140 -12240
rect 3720 -12410 3840 -11550
rect 4420 -11660 4520 -10000
rect 4640 -10300 4740 -8640
rect 5320 -8810 5440 -8780
rect 5320 -9470 5330 -8810
rect 5430 -9470 5440 -8810
rect 5320 -9590 5440 -9470
rect 5320 -9750 5330 -9590
rect 5430 -9750 5440 -9590
rect 4620 -10310 4760 -10300
rect 4620 -10430 4630 -10310
rect 4750 -10430 4760 -10310
rect 4620 -10440 4760 -10430
rect 4400 -11670 4540 -11660
rect 4400 -11790 4410 -11670
rect 4530 -11790 4540 -11670
rect 4400 -11800 4540 -11790
rect 3720 -13070 3730 -12410
rect 3830 -13070 3840 -12410
rect 3720 -13190 3840 -13070
rect 3720 -13350 3730 -13190
rect 3830 -13350 3840 -13190
rect 3020 -13910 3160 -13900
rect 3020 -14030 3030 -13910
rect 3150 -14030 3160 -13910
rect 3020 -14040 3160 -14030
rect 2800 -15270 2940 -15260
rect 2800 -15390 2810 -15270
rect 2930 -15390 2940 -15270
rect 2800 -15400 2940 -15390
rect 2120 -16670 2130 -16010
rect 2230 -16670 2240 -16010
rect 2120 -16790 2240 -16670
rect 2120 -16950 2130 -16790
rect 2230 -16950 2240 -16790
rect 1420 -17510 1560 -17500
rect 1420 -17630 1430 -17510
rect 1550 -17630 1560 -17510
rect 1420 -17640 1560 -17630
rect 1200 -18870 1340 -18860
rect 1200 -18990 1210 -18870
rect 1330 -18990 1340 -18870
rect 1200 -19000 1340 -18990
rect 1220 -20660 1320 -19000
rect 1440 -19300 1540 -17640
rect 2120 -17810 2240 -16950
rect 2820 -17060 2920 -15400
rect 3040 -15700 3140 -14040
rect 3720 -14210 3840 -13350
rect 4420 -13460 4520 -11800
rect 4640 -12100 4740 -10440
rect 5320 -10610 5440 -9750
rect 6020 -9860 6120 -8200
rect 6240 -8500 6340 -8050
rect 7620 -8060 7720 -8050
rect 9220 -8060 9320 -8050
rect 7600 -8070 7740 -8060
rect 7600 -8190 7610 -8070
rect 7730 -8190 7740 -8070
rect 7600 -8200 7740 -8190
rect 9200 -8070 9340 -8060
rect 9200 -8190 9210 -8070
rect 9330 -8190 9340 -8070
rect 9200 -8200 9340 -8190
rect 6220 -8510 6360 -8500
rect 6220 -8630 6230 -8510
rect 6350 -8630 6360 -8510
rect 6220 -8640 6360 -8630
rect 6000 -9870 6140 -9860
rect 6000 -9990 6010 -9870
rect 6130 -9990 6140 -9870
rect 6000 -10000 6140 -9990
rect 5320 -11270 5330 -10610
rect 5430 -11270 5440 -10610
rect 5320 -11390 5440 -11270
rect 5320 -11550 5330 -11390
rect 5430 -11550 5440 -11390
rect 4620 -12110 4760 -12100
rect 4620 -12230 4630 -12110
rect 4750 -12230 4760 -12110
rect 4620 -12240 4760 -12230
rect 4400 -13470 4540 -13460
rect 4400 -13590 4410 -13470
rect 4530 -13590 4540 -13470
rect 4400 -13600 4540 -13590
rect 3720 -14870 3730 -14210
rect 3830 -14870 3840 -14210
rect 3720 -14990 3840 -14870
rect 3720 -15150 3730 -14990
rect 3830 -15150 3840 -14990
rect 3020 -15710 3160 -15700
rect 3020 -15830 3030 -15710
rect 3150 -15830 3160 -15710
rect 3020 -15840 3160 -15830
rect 2800 -17070 2940 -17060
rect 2800 -17190 2810 -17070
rect 2930 -17190 2940 -17070
rect 2800 -17200 2940 -17190
rect 2120 -18470 2130 -17810
rect 2230 -18470 2240 -17810
rect 2120 -18590 2240 -18470
rect 2120 -18750 2130 -18590
rect 2230 -18750 2240 -18590
rect 1420 -19310 1560 -19300
rect 1420 -19430 1430 -19310
rect 1550 -19430 1560 -19310
rect 1420 -19440 1560 -19430
rect 1200 -20670 1340 -20660
rect 1200 -20790 1210 -20670
rect 1330 -20790 1340 -20670
rect 1200 -20800 1340 -20790
rect 480 -22400 680 -22380
rect 1220 -23260 1320 -20800
rect 1440 -21100 1540 -19440
rect 2120 -19610 2240 -18750
rect 2820 -18860 2920 -17200
rect 3040 -17500 3140 -15840
rect 3720 -16010 3840 -15150
rect 4420 -15260 4520 -13600
rect 4640 -13900 4740 -12240
rect 5320 -12410 5440 -11550
rect 6020 -11660 6120 -10000
rect 6240 -10300 6340 -8640
rect 6920 -8810 7040 -8780
rect 6920 -9470 6930 -8810
rect 7030 -9470 7040 -8810
rect 6920 -9590 7040 -9470
rect 6920 -9750 6930 -9590
rect 7030 -9750 7040 -9590
rect 6220 -10310 6360 -10300
rect 6220 -10430 6230 -10310
rect 6350 -10430 6360 -10310
rect 6220 -10440 6360 -10430
rect 6000 -11670 6140 -11660
rect 6000 -11790 6010 -11670
rect 6130 -11790 6140 -11670
rect 6000 -11800 6140 -11790
rect 5320 -13070 5330 -12410
rect 5430 -13070 5440 -12410
rect 5320 -13190 5440 -13070
rect 5320 -13350 5330 -13190
rect 5430 -13350 5440 -13190
rect 4620 -13910 4760 -13900
rect 4620 -14030 4630 -13910
rect 4750 -14030 4760 -13910
rect 4620 -14040 4760 -14030
rect 4400 -15270 4540 -15260
rect 4400 -15390 4410 -15270
rect 4530 -15390 4540 -15270
rect 4400 -15400 4540 -15390
rect 3720 -16670 3730 -16010
rect 3830 -16670 3840 -16010
rect 3720 -16790 3840 -16670
rect 3720 -16950 3730 -16790
rect 3830 -16950 3840 -16790
rect 3020 -17510 3160 -17500
rect 3020 -17630 3030 -17510
rect 3150 -17630 3160 -17510
rect 3020 -17640 3160 -17630
rect 2800 -18870 2940 -18860
rect 2800 -18990 2810 -18870
rect 2930 -18990 2940 -18870
rect 2800 -19000 2940 -18990
rect 2120 -20270 2130 -19610
rect 2230 -20270 2240 -19610
rect 2120 -20390 2240 -20270
rect 2120 -20550 2130 -20390
rect 2230 -20550 2240 -20390
rect 1420 -21110 1560 -21100
rect 1420 -21230 1430 -21110
rect 1550 -21230 1560 -21110
rect 1420 -21240 1560 -21230
rect 2120 -21410 2240 -20550
rect 2820 -20660 2920 -19000
rect 3040 -19300 3140 -17640
rect 3720 -17810 3840 -16950
rect 4420 -17060 4520 -15400
rect 4640 -15700 4740 -14040
rect 5320 -14210 5440 -13350
rect 6020 -13460 6120 -11800
rect 6240 -12100 6340 -10440
rect 6920 -10610 7040 -9750
rect 7620 -9860 7720 -8200
rect 7840 -8500 7940 -8220
rect 7820 -8510 7960 -8500
rect 7820 -8630 7830 -8510
rect 7950 -8630 7960 -8510
rect 7820 -8640 7960 -8630
rect 7600 -9870 7740 -9860
rect 7600 -9990 7610 -9870
rect 7730 -9990 7740 -9870
rect 7600 -10000 7740 -9990
rect 6920 -11270 6930 -10610
rect 7030 -11270 7040 -10610
rect 6920 -11390 7040 -11270
rect 6920 -11550 6930 -11390
rect 7030 -11550 7040 -11390
rect 6220 -12110 6360 -12100
rect 6220 -12230 6230 -12110
rect 6350 -12230 6360 -12110
rect 6220 -12240 6360 -12230
rect 6000 -13470 6140 -13460
rect 6000 -13590 6010 -13470
rect 6130 -13590 6140 -13470
rect 6000 -13600 6140 -13590
rect 5320 -14870 5330 -14210
rect 5430 -14870 5440 -14210
rect 5320 -14990 5440 -14870
rect 5320 -15150 5330 -14990
rect 5430 -15150 5440 -14990
rect 4620 -15710 4760 -15700
rect 4620 -15830 4630 -15710
rect 4750 -15830 4760 -15710
rect 4620 -15840 4760 -15830
rect 4400 -17070 4540 -17060
rect 4400 -17190 4410 -17070
rect 4530 -17190 4540 -17070
rect 4400 -17200 4540 -17190
rect 3720 -18470 3730 -17810
rect 3830 -18470 3840 -17810
rect 3720 -18590 3840 -18470
rect 3720 -18750 3730 -18590
rect 3830 -18750 3840 -18590
rect 3020 -19310 3160 -19300
rect 3020 -19430 3030 -19310
rect 3150 -19430 3160 -19310
rect 3020 -19440 3160 -19430
rect 2800 -20670 2940 -20660
rect 2800 -20790 2810 -20670
rect 2930 -20790 2940 -20670
rect 2800 -20800 2940 -20790
rect 2120 -22070 2130 -21410
rect 2230 -22070 2240 -21410
rect 2120 -22190 2240 -22070
rect 2120 -22350 2130 -22190
rect 2230 -22350 2240 -22190
rect 2120 -22360 2240 -22350
rect 2820 -23260 2920 -20800
rect 3040 -21100 3140 -19440
rect 3720 -19610 3840 -18750
rect 4420 -18860 4520 -17200
rect 4640 -17500 4740 -15840
rect 5320 -16010 5440 -15150
rect 6020 -15260 6120 -13600
rect 6240 -13900 6340 -12240
rect 6920 -12410 7040 -11550
rect 7620 -11660 7720 -10000
rect 7840 -10300 7940 -8640
rect 8520 -8810 8640 -8780
rect 8520 -9470 8530 -8810
rect 8630 -9470 8640 -8810
rect 8520 -9590 8640 -9470
rect 8520 -9750 8530 -9590
rect 8630 -9750 8640 -9590
rect 7820 -10310 7960 -10300
rect 7820 -10430 7830 -10310
rect 7950 -10430 7960 -10310
rect 7820 -10440 7960 -10430
rect 7600 -11670 7740 -11660
rect 7600 -11790 7610 -11670
rect 7730 -11790 7740 -11670
rect 7600 -11800 7740 -11790
rect 6920 -13070 6930 -12410
rect 7030 -13070 7040 -12410
rect 6920 -13190 7040 -13070
rect 6920 -13350 6930 -13190
rect 7030 -13350 7040 -13190
rect 6220 -13910 6360 -13900
rect 6220 -14030 6230 -13910
rect 6350 -14030 6360 -13910
rect 6220 -14040 6360 -14030
rect 6000 -15270 6140 -15260
rect 6000 -15390 6010 -15270
rect 6130 -15390 6140 -15270
rect 6000 -15400 6140 -15390
rect 5320 -16670 5330 -16010
rect 5430 -16670 5440 -16010
rect 5320 -16790 5440 -16670
rect 5320 -16950 5330 -16790
rect 5430 -16950 5440 -16790
rect 4620 -17510 4760 -17500
rect 4620 -17630 4630 -17510
rect 4750 -17630 4760 -17510
rect 4620 -17640 4760 -17630
rect 4400 -18870 4540 -18860
rect 4400 -18990 4410 -18870
rect 4530 -18990 4540 -18870
rect 4400 -19000 4540 -18990
rect 3720 -20270 3730 -19610
rect 3830 -20270 3840 -19610
rect 3720 -20390 3840 -20270
rect 3720 -20550 3730 -20390
rect 3830 -20550 3840 -20390
rect 3020 -21110 3160 -21100
rect 3020 -21230 3030 -21110
rect 3150 -21230 3160 -21110
rect 3020 -21240 3160 -21230
rect 3720 -21410 3840 -20550
rect 4420 -20660 4520 -19000
rect 4640 -19300 4740 -17640
rect 5320 -17810 5440 -16950
rect 6020 -17060 6120 -15400
rect 6240 -15700 6340 -14040
rect 6920 -14210 7040 -13350
rect 7620 -13460 7720 -11800
rect 7840 -12100 7940 -10440
rect 8520 -10610 8640 -9750
rect 9220 -9860 9320 -8200
rect 9440 -8500 9540 -8050
rect 10820 -8250 10920 -8030
rect 10800 -8260 10940 -8250
rect 10800 -8380 10810 -8260
rect 10930 -8380 10940 -8260
rect 10800 -8390 10940 -8380
rect 9420 -8510 9560 -8500
rect 9420 -8630 9430 -8510
rect 9550 -8630 9560 -8510
rect 9420 -8640 9560 -8630
rect 9200 -9870 9340 -9860
rect 9200 -9990 9210 -9870
rect 9330 -9990 9340 -9870
rect 9200 -10000 9340 -9990
rect 8520 -11270 8530 -10610
rect 8630 -11270 8640 -10610
rect 8520 -11390 8640 -11270
rect 8520 -11550 8530 -11390
rect 8630 -11550 8640 -11390
rect 7820 -12110 7960 -12100
rect 7820 -12230 7830 -12110
rect 7950 -12230 7960 -12110
rect 7820 -12240 7960 -12230
rect 7600 -13470 7740 -13460
rect 7600 -13590 7610 -13470
rect 7730 -13590 7740 -13470
rect 7600 -13600 7740 -13590
rect 6920 -14870 6930 -14210
rect 7030 -14870 7040 -14210
rect 6920 -14990 7040 -14870
rect 6920 -15150 6930 -14990
rect 7030 -15150 7040 -14990
rect 6220 -15710 6360 -15700
rect 6220 -15830 6230 -15710
rect 6350 -15830 6360 -15710
rect 6220 -15840 6360 -15830
rect 6000 -17070 6140 -17060
rect 6000 -17190 6010 -17070
rect 6130 -17190 6140 -17070
rect 6000 -17200 6140 -17190
rect 5320 -18470 5330 -17810
rect 5430 -18470 5440 -17810
rect 5320 -18590 5440 -18470
rect 5320 -18750 5330 -18590
rect 5430 -18750 5440 -18590
rect 4620 -19310 4760 -19300
rect 4620 -19430 4630 -19310
rect 4750 -19430 4760 -19310
rect 4620 -19440 4760 -19430
rect 4400 -20670 4540 -20660
rect 4400 -20790 4410 -20670
rect 4530 -20790 4540 -20670
rect 4400 -20800 4540 -20790
rect 3720 -22070 3730 -21410
rect 3830 -22070 3840 -21410
rect 3720 -22190 3840 -22070
rect 3720 -22350 3730 -22190
rect 3830 -22350 3840 -22190
rect 3720 -22360 3840 -22350
rect 4420 -23260 4520 -20800
rect 4640 -21100 4740 -19440
rect 5320 -19610 5440 -18750
rect 6020 -18860 6120 -17200
rect 6240 -17500 6340 -15840
rect 6920 -16010 7040 -15150
rect 7620 -15260 7720 -13600
rect 7840 -13900 7940 -12240
rect 8520 -12410 8640 -11550
rect 9220 -11660 9320 -10000
rect 9440 -10300 9540 -8640
rect 10120 -8810 10240 -8780
rect 10120 -9470 10130 -8810
rect 10230 -9470 10240 -8810
rect 10120 -9590 10240 -9470
rect 10120 -9750 10130 -9590
rect 10230 -9750 10240 -9590
rect 9420 -10310 9560 -10300
rect 9420 -10430 9430 -10310
rect 9550 -10430 9560 -10310
rect 9420 -10440 9560 -10430
rect 9200 -11670 9340 -11660
rect 9200 -11790 9210 -11670
rect 9330 -11790 9340 -11670
rect 9200 -11800 9340 -11790
rect 8520 -13070 8530 -12410
rect 8630 -13070 8640 -12410
rect 8520 -13190 8640 -13070
rect 8520 -13350 8530 -13190
rect 8630 -13350 8640 -13190
rect 7820 -13910 7960 -13900
rect 7820 -14030 7830 -13910
rect 7950 -14030 7960 -13910
rect 7820 -14040 7960 -14030
rect 7600 -15270 7740 -15260
rect 7600 -15390 7610 -15270
rect 7730 -15390 7740 -15270
rect 7600 -15400 7740 -15390
rect 6920 -16670 6930 -16010
rect 7030 -16670 7040 -16010
rect 6920 -16790 7040 -16670
rect 6920 -16950 6930 -16790
rect 7030 -16950 7040 -16790
rect 6220 -17510 6360 -17500
rect 6220 -17630 6230 -17510
rect 6350 -17630 6360 -17510
rect 6220 -17640 6360 -17630
rect 6000 -18870 6140 -18860
rect 6000 -18990 6010 -18870
rect 6130 -18990 6140 -18870
rect 6000 -19000 6140 -18990
rect 5320 -20270 5330 -19610
rect 5430 -20270 5440 -19610
rect 5320 -20390 5440 -20270
rect 5320 -20550 5330 -20390
rect 5430 -20550 5440 -20390
rect 4620 -21110 4760 -21100
rect 4620 -21230 4630 -21110
rect 4750 -21230 4760 -21110
rect 4620 -21240 4760 -21230
rect 5320 -21410 5440 -20550
rect 6020 -20660 6120 -19000
rect 6240 -19300 6340 -17640
rect 6920 -17810 7040 -16950
rect 7620 -17060 7720 -15400
rect 7840 -15700 7940 -14040
rect 8520 -14210 8640 -13350
rect 9220 -13460 9320 -11800
rect 9440 -12100 9540 -10440
rect 10120 -10610 10240 -9750
rect 10820 -10050 10920 -8390
rect 11040 -9580 11140 -4850
rect 11700 -4810 11840 -4800
rect 11700 -4930 11710 -4810
rect 11830 -4930 11840 -4810
rect 12600 -4850 12610 -4730
rect 12730 -4850 12740 -4730
rect 12600 -4860 12740 -4850
rect 13620 -4790 13760 -4780
rect 13620 -4910 13630 -4790
rect 13750 -4910 13760 -4790
rect 13620 -4920 13760 -4910
rect 11700 -4940 11840 -4930
rect 11720 -5820 11820 -4940
rect 11700 -5830 11840 -5820
rect 11700 -5950 11710 -5830
rect 11830 -5950 11840 -5830
rect 11700 -5960 11840 -5950
rect 13300 -5830 13440 -5820
rect 13300 -5950 13310 -5830
rect 13430 -5950 13440 -5830
rect 13300 -5960 13440 -5950
rect 11700 -6050 11840 -6040
rect 11700 -6170 11710 -6050
rect 11830 -6170 11840 -6050
rect 11700 -6180 11840 -6170
rect 11720 -8100 11820 -6180
rect 12620 -6270 12760 -6260
rect 12620 -6390 12630 -6270
rect 12750 -6390 12760 -6270
rect 12620 -6400 12760 -6390
rect 12400 -6490 12540 -6480
rect 12400 -6610 12410 -6490
rect 12530 -6610 12540 -6490
rect 12400 -6620 12540 -6610
rect 11700 -8110 11860 -8100
rect 11700 -8230 11710 -8110
rect 11840 -8140 11860 -8110
rect 11840 -8230 11850 -8140
rect 11700 -8240 11850 -8230
rect 11710 -8810 11840 -8240
rect 11710 -9470 11720 -8810
rect 11830 -9470 11840 -8810
rect 11710 -9480 11840 -9470
rect 11030 -9760 11150 -9580
rect 10800 -10060 10940 -10050
rect 10800 -10180 10810 -10060
rect 10930 -10180 10940 -10060
rect 10800 -10190 10940 -10180
rect 10120 -11270 10130 -10610
rect 10230 -11270 10240 -10610
rect 10120 -11390 10240 -11270
rect 10120 -11550 10130 -11390
rect 10230 -11550 10240 -11390
rect 9420 -12110 9560 -12100
rect 9420 -12230 9430 -12110
rect 9550 -12230 9560 -12110
rect 9420 -12240 9560 -12230
rect 9200 -13470 9340 -13460
rect 9200 -13590 9210 -13470
rect 9330 -13590 9340 -13470
rect 9200 -13600 9340 -13590
rect 8520 -14870 8530 -14210
rect 8630 -14870 8640 -14210
rect 8520 -14990 8640 -14870
rect 8520 -15150 8530 -14990
rect 8630 -15150 8640 -14990
rect 7820 -15710 7960 -15700
rect 7820 -15830 7830 -15710
rect 7950 -15830 7960 -15710
rect 7820 -15840 7960 -15830
rect 7600 -17070 7740 -17060
rect 7600 -17190 7610 -17070
rect 7730 -17190 7740 -17070
rect 7600 -17200 7740 -17190
rect 6920 -18470 6930 -17810
rect 7030 -18470 7040 -17810
rect 6920 -18590 7040 -18470
rect 6920 -18750 6930 -18590
rect 7030 -18750 7040 -18590
rect 6220 -19310 6360 -19300
rect 6220 -19430 6230 -19310
rect 6350 -19430 6360 -19310
rect 6220 -19440 6360 -19430
rect 6000 -20670 6140 -20660
rect 6000 -20790 6010 -20670
rect 6130 -20790 6140 -20670
rect 6000 -20800 6140 -20790
rect 5320 -22070 5330 -21410
rect 5430 -22070 5440 -21410
rect 5320 -22190 5440 -22070
rect 5320 -22350 5330 -22190
rect 5430 -22350 5440 -22190
rect 5320 -22360 5440 -22350
rect 6020 -23260 6120 -20800
rect 6240 -21100 6340 -19440
rect 6920 -19610 7040 -18750
rect 7620 -18860 7720 -17200
rect 7840 -17500 7940 -15840
rect 8520 -16010 8640 -15150
rect 9220 -15260 9320 -13600
rect 9440 -13900 9540 -12240
rect 10120 -12410 10240 -11550
rect 10820 -11850 10920 -10190
rect 11040 -10400 11140 -9760
rect 11020 -10410 11160 -10400
rect 11020 -10530 11030 -10410
rect 11150 -10530 11160 -10410
rect 11020 -10540 11160 -10530
rect 11040 -11380 11140 -10540
rect 11710 -10610 11840 -10600
rect 11710 -11270 11720 -10610
rect 11830 -11270 11840 -10610
rect 11030 -11560 11150 -11380
rect 10800 -11860 10940 -11850
rect 10800 -11980 10810 -11860
rect 10930 -11980 10940 -11860
rect 10800 -11990 10940 -11980
rect 10120 -13070 10130 -12410
rect 10230 -13070 10240 -12410
rect 10120 -13190 10240 -13070
rect 10120 -13350 10130 -13190
rect 10230 -13350 10240 -13190
rect 9420 -13910 9560 -13900
rect 9420 -14030 9430 -13910
rect 9550 -14030 9560 -13910
rect 9420 -14040 9560 -14030
rect 9200 -15270 9340 -15260
rect 9200 -15390 9210 -15270
rect 9330 -15390 9340 -15270
rect 9200 -15400 9340 -15390
rect 8520 -16670 8530 -16010
rect 8630 -16670 8640 -16010
rect 8520 -16790 8640 -16670
rect 8520 -16950 8530 -16790
rect 8630 -16950 8640 -16790
rect 7820 -17510 7960 -17500
rect 7820 -17630 7830 -17510
rect 7950 -17630 7960 -17510
rect 7820 -17640 7960 -17630
rect 7600 -18870 7740 -18860
rect 7600 -18990 7610 -18870
rect 7730 -18990 7740 -18870
rect 7600 -19000 7740 -18990
rect 6920 -20270 6930 -19610
rect 7030 -20270 7040 -19610
rect 6920 -20390 7040 -20270
rect 6920 -20550 6930 -20390
rect 7030 -20550 7040 -20390
rect 6220 -21110 6360 -21100
rect 6220 -21230 6230 -21110
rect 6350 -21230 6360 -21110
rect 6220 -21240 6360 -21230
rect 6920 -21410 7040 -20550
rect 7620 -20660 7720 -19000
rect 7840 -19300 7940 -17640
rect 8520 -17810 8640 -16950
rect 9220 -17060 9320 -15400
rect 9440 -15700 9540 -14040
rect 10120 -14210 10240 -13350
rect 10820 -13650 10920 -11990
rect 11040 -13180 11140 -11560
rect 11710 -12410 11840 -11270
rect 11710 -13070 11720 -12410
rect 11830 -13070 11840 -12410
rect 11030 -13360 11150 -13180
rect 11260 -13210 11270 -13150
rect 11650 -13210 11660 -13150
rect 10800 -13660 10940 -13650
rect 10800 -13780 10810 -13660
rect 10930 -13780 10940 -13660
rect 10800 -13790 10940 -13780
rect 10120 -14870 10130 -14210
rect 10230 -14870 10240 -14210
rect 10120 -14990 10240 -14870
rect 10120 -15150 10130 -14990
rect 10230 -15150 10240 -14990
rect 9420 -15710 9560 -15700
rect 9420 -15830 9430 -15710
rect 9550 -15830 9560 -15710
rect 9420 -15840 9560 -15830
rect 9200 -17070 9340 -17060
rect 9200 -17190 9210 -17070
rect 9330 -17190 9340 -17070
rect 9200 -17200 9340 -17190
rect 8520 -18470 8530 -17810
rect 8630 -18470 8640 -17810
rect 8520 -18590 8640 -18470
rect 8520 -18750 8530 -18590
rect 8630 -18750 8640 -18590
rect 7820 -19310 7960 -19300
rect 7820 -19430 7830 -19310
rect 7950 -19430 7960 -19310
rect 7820 -19440 7960 -19430
rect 7600 -20670 7740 -20660
rect 7600 -20790 7610 -20670
rect 7730 -20790 7740 -20670
rect 7600 -20800 7740 -20790
rect 6920 -22070 6930 -21410
rect 7030 -22070 7040 -21410
rect 6920 -22190 7040 -22070
rect 6920 -22350 6930 -22190
rect 7030 -22350 7040 -22190
rect 6920 -22360 7040 -22350
rect 7620 -23260 7720 -20800
rect 7840 -21100 7940 -19440
rect 8520 -19610 8640 -18750
rect 9220 -18860 9320 -17200
rect 9440 -17500 9540 -15840
rect 10120 -16010 10240 -15150
rect 10820 -15450 10920 -13790
rect 11040 -14980 11140 -13360
rect 11260 -14060 11660 -13210
rect 11260 -14120 11270 -14060
rect 11650 -14120 11660 -14060
rect 11260 -14130 11660 -14120
rect 11710 -14210 11840 -13070
rect 11710 -14870 11720 -14210
rect 11830 -14870 11840 -14210
rect 11710 -14880 11840 -14870
rect 11030 -15160 11150 -14980
rect 10800 -15460 10940 -15450
rect 10800 -15580 10810 -15460
rect 10930 -15580 10940 -15460
rect 10800 -15590 10940 -15580
rect 10120 -16670 10130 -16010
rect 10230 -16670 10240 -16010
rect 10120 -16790 10240 -16670
rect 10120 -16950 10130 -16790
rect 10230 -16950 10240 -16790
rect 9420 -17510 9560 -17500
rect 9420 -17630 9430 -17510
rect 9550 -17630 9560 -17510
rect 9420 -17640 9560 -17630
rect 9200 -18870 9340 -18860
rect 9200 -18990 9210 -18870
rect 9330 -18990 9340 -18870
rect 9200 -19000 9340 -18990
rect 8520 -20270 8530 -19610
rect 8630 -20270 8640 -19610
rect 8520 -20390 8640 -20270
rect 8520 -20550 8530 -20390
rect 8630 -20550 8640 -20390
rect 7820 -21110 7960 -21100
rect 7820 -21230 7830 -21110
rect 7950 -21230 7960 -21110
rect 7820 -21240 7960 -21230
rect 8520 -21410 8640 -20550
rect 9220 -20660 9320 -19000
rect 9440 -19300 9540 -17640
rect 10120 -17810 10240 -16950
rect 10820 -17250 10920 -15590
rect 11040 -16780 11140 -15160
rect 11030 -16960 11150 -16780
rect 10800 -17260 10940 -17250
rect 10800 -17380 10810 -17260
rect 10930 -17380 10940 -17260
rect 10800 -17390 10940 -17380
rect 10120 -18470 10130 -17810
rect 10230 -18470 10240 -17810
rect 10120 -18590 10240 -18470
rect 10120 -18750 10130 -18590
rect 10230 -18750 10240 -18590
rect 9420 -19310 9560 -19300
rect 9420 -19430 9430 -19310
rect 9550 -19430 9560 -19310
rect 9420 -19440 9560 -19430
rect 9200 -20670 9340 -20660
rect 9200 -20790 9210 -20670
rect 9330 -20790 9340 -20670
rect 9200 -20800 9340 -20790
rect 8520 -22070 8530 -21410
rect 8630 -22070 8640 -21410
rect 8520 -22190 8640 -22070
rect 8520 -22350 8530 -22190
rect 8630 -22350 8640 -22190
rect 8520 -22360 8640 -22350
rect 9220 -23260 9320 -20800
rect 9440 -21100 9540 -19440
rect 10120 -19610 10240 -18750
rect 10820 -19050 10920 -17390
rect 11040 -18580 11140 -16960
rect 11030 -18760 11150 -18580
rect 10800 -19060 10940 -19050
rect 10800 -19180 10810 -19060
rect 10930 -19180 10940 -19060
rect 10800 -19190 10940 -19180
rect 10120 -20270 10130 -19610
rect 10230 -20270 10240 -19610
rect 10120 -20390 10240 -20270
rect 10120 -20550 10130 -20390
rect 10230 -20550 10240 -20390
rect 9420 -21110 9560 -21100
rect 9420 -21230 9430 -21110
rect 9550 -21230 9560 -21110
rect 9420 -21240 9560 -21230
rect 10120 -21410 10240 -20550
rect 10820 -20850 10920 -19190
rect 11040 -20380 11140 -18760
rect 12420 -18870 12520 -6620
rect 12640 -17070 12740 -6400
rect 12940 -6830 13120 -6820
rect 12940 -6990 12950 -6830
rect 13110 -6990 13120 -6830
rect 12940 -7000 13120 -6990
rect 13310 -8240 13440 -5960
rect 13640 -6040 13740 -4920
rect 14000 -5070 14100 -3220
rect 14200 -3290 14340 -3280
rect 14200 -3410 14210 -3290
rect 14330 -3410 14340 -3290
rect 14200 -3420 14340 -3410
rect 14900 -3310 14910 -3150
rect 15030 -3310 15040 -3150
rect 14900 -3410 15040 -3310
rect 14220 -4720 14320 -3420
rect 14900 -4090 14910 -3410
rect 15030 -4090 15040 -3410
rect 14900 -4100 15040 -4090
rect 15600 -4240 15700 -2580
rect 15820 -2910 15920 -1250
rect 16500 -1350 16640 -490
rect 17200 -640 17300 1020
rect 17420 690 17520 1310
rect 17410 680 17530 690
rect 17410 560 17420 680
rect 17520 560 17530 680
rect 17410 550 17530 560
rect 17190 -650 17310 -640
rect 17190 -770 17200 -650
rect 17300 -770 17310 -650
rect 17190 -780 17310 -770
rect 16500 -1510 16510 -1350
rect 16630 -1510 16640 -1350
rect 16500 -1610 16640 -1510
rect 16500 -2290 16510 -1610
rect 16630 -2290 16640 -1610
rect 15810 -2920 15930 -2910
rect 15810 -3040 15820 -2920
rect 15920 -3040 15930 -2920
rect 15810 -3050 15930 -3040
rect 15590 -4250 15710 -4240
rect 15590 -4370 15600 -4250
rect 15700 -4370 15710 -4250
rect 15590 -4380 15710 -4370
rect 14200 -4730 14340 -4720
rect 14200 -4850 14210 -4730
rect 14330 -4850 14340 -4730
rect 14200 -4860 14340 -4850
rect 15220 -4790 15360 -4780
rect 15220 -4910 15230 -4790
rect 15350 -4910 15360 -4790
rect 15220 -4920 15360 -4910
rect 14000 -5200 14120 -5070
rect 13620 -6050 13760 -6040
rect 13620 -6170 13630 -6050
rect 13750 -6170 13760 -6050
rect 13620 -6180 13760 -6170
rect 13300 -8260 13450 -8240
rect 13300 -8380 13310 -8260
rect 13440 -8380 13450 -8260
rect 13300 -8390 13450 -8380
rect 13310 -8810 13440 -8390
rect 13310 -9470 13320 -8810
rect 13430 -9470 13440 -8810
rect 13310 -9480 13440 -9470
rect 13310 -10610 13440 -10600
rect 13310 -11270 13320 -10610
rect 13430 -11270 13440 -10610
rect 13310 -11280 13440 -11270
rect 13300 -11670 13440 -11660
rect 13300 -11790 13310 -11670
rect 13430 -11790 13440 -11670
rect 13300 -11800 13440 -11790
rect 13310 -12410 13440 -11800
rect 13310 -13070 13320 -12410
rect 13430 -13070 13440 -12410
rect 13310 -13160 13440 -13070
rect 13280 -13170 13470 -13160
rect 13280 -13330 13290 -13170
rect 13460 -13330 13470 -13170
rect 13280 -13340 13470 -13330
rect 13310 -14210 13440 -13340
rect 14020 -13470 14120 -5200
rect 15240 -6040 15340 -4920
rect 15600 -5160 15700 -4380
rect 15820 -4710 15920 -3050
rect 16500 -3150 16640 -2290
rect 17200 -2440 17300 -780
rect 17420 -1110 17520 550
rect 18100 450 18240 1310
rect 18800 1160 18900 1310
rect 18790 1150 18910 1160
rect 18790 1030 18800 1150
rect 18900 1030 18910 1150
rect 18790 1020 18910 1030
rect 18100 290 18110 450
rect 18230 290 18240 450
rect 18100 190 18240 290
rect 18100 -490 18110 190
rect 18230 -490 18240 190
rect 17410 -1120 17530 -1110
rect 17410 -1240 17420 -1120
rect 17520 -1240 17530 -1120
rect 17410 -1250 17530 -1240
rect 17190 -2450 17310 -2440
rect 17190 -2570 17200 -2450
rect 17300 -2570 17310 -2450
rect 17190 -2580 17310 -2570
rect 16500 -3310 16510 -3150
rect 16630 -3310 16640 -3150
rect 16500 -3410 16640 -3310
rect 16500 -4090 16510 -3410
rect 16630 -4090 16640 -3410
rect 15810 -4720 15930 -4710
rect 15810 -4840 15820 -4720
rect 15920 -4840 15930 -4720
rect 15810 -4850 15930 -4840
rect 15560 -5170 15740 -5160
rect 15560 -5350 15570 -5170
rect 15730 -5350 15740 -5170
rect 15560 -5360 15740 -5350
rect 15560 -5570 15740 -5560
rect 15560 -5750 15570 -5570
rect 15730 -5750 15740 -5570
rect 15560 -5760 15740 -5750
rect 14220 -6050 14360 -6040
rect 14220 -6170 14230 -6050
rect 14350 -6170 14360 -6050
rect 14220 -6180 14360 -6170
rect 15220 -6050 15360 -6040
rect 15220 -6170 15230 -6050
rect 15350 -6170 15360 -6050
rect 15220 -6180 15360 -6170
rect 14240 -11660 14340 -6180
rect 14900 -6490 15040 -6480
rect 14900 -6610 14910 -6490
rect 15030 -6610 15040 -6490
rect 14900 -6620 15040 -6610
rect 14900 -7880 15050 -7870
rect 14900 -8000 14910 -7880
rect 15040 -8000 15050 -7880
rect 14900 -8010 15050 -8000
rect 14220 -11670 14360 -11660
rect 14220 -11790 14230 -11670
rect 14350 -11790 14360 -11670
rect 14220 -11800 14360 -11790
rect 14000 -13480 14140 -13470
rect 14000 -13600 14010 -13480
rect 14130 -13600 14140 -13480
rect 14000 -13610 14140 -13600
rect 13310 -14870 13320 -14210
rect 13430 -14870 13440 -14210
rect 13310 -14960 13440 -14870
rect 13280 -14970 13470 -14960
rect 13280 -15130 13290 -14970
rect 13460 -15130 13470 -14970
rect 13280 -15140 13470 -15130
rect 13310 -15290 13440 -15280
rect 13310 -15390 13330 -15290
rect 13430 -15390 13440 -15290
rect 14020 -15300 14120 -13610
rect 13310 -16010 13440 -15390
rect 14010 -15310 14130 -15300
rect 14010 -15410 14020 -15310
rect 14120 -15410 14130 -15310
rect 14010 -15420 14130 -15410
rect 13310 -16670 13320 -16010
rect 13430 -16670 13440 -16010
rect 13310 -16680 13440 -16670
rect 13310 -16780 13430 -16680
rect 13290 -16790 13460 -16780
rect 13290 -16950 13300 -16790
rect 13450 -16950 13460 -16790
rect 13290 -16960 13460 -16950
rect 12620 -17080 12760 -17070
rect 12620 -17200 12630 -17080
rect 12750 -17200 12760 -17080
rect 12620 -17210 12760 -17200
rect 13310 -17800 13430 -16960
rect 13310 -17810 13440 -17800
rect 13310 -18470 13320 -17810
rect 13430 -18470 13440 -17810
rect 13310 -18580 13440 -18470
rect 13290 -18590 13460 -18580
rect 13290 -18750 13300 -18590
rect 13450 -18750 13460 -18590
rect 13290 -18760 13460 -18750
rect 12400 -18880 12540 -18870
rect 12400 -19000 12410 -18880
rect 12530 -19000 12540 -18880
rect 12400 -19010 12540 -19000
rect 14240 -19320 14340 -11800
rect 14910 -12090 15040 -8010
rect 15620 -8510 15720 -5760
rect 15820 -5960 15920 -4850
rect 15780 -5970 15960 -5960
rect 15780 -6150 15790 -5970
rect 15950 -6150 15960 -5970
rect 15780 -6160 15960 -6150
rect 15840 -8060 15940 -6160
rect 16500 -6270 16640 -4090
rect 17200 -4240 17300 -2580
rect 17420 -2910 17520 -1250
rect 18100 -1350 18240 -490
rect 18800 -640 18900 1020
rect 19020 690 19120 1310
rect 19010 680 19130 690
rect 19010 560 19020 680
rect 19120 560 19130 680
rect 19010 550 19130 560
rect 18790 -650 18910 -640
rect 18790 -770 18800 -650
rect 18900 -770 18910 -650
rect 18790 -780 18910 -770
rect 18100 -1510 18110 -1350
rect 18230 -1510 18240 -1350
rect 18100 -1610 18240 -1510
rect 18100 -2290 18110 -1610
rect 18230 -2290 18240 -1610
rect 17410 -2920 17530 -2910
rect 17410 -3040 17420 -2920
rect 17520 -3040 17530 -2920
rect 17410 -3050 17530 -3040
rect 17190 -4250 17310 -4240
rect 17190 -4370 17200 -4250
rect 17300 -4370 17310 -4250
rect 17190 -4380 17310 -4370
rect 16500 -6390 16510 -6270
rect 16630 -6390 16640 -6270
rect 16500 -6400 16640 -6390
rect 17200 -7160 17300 -4380
rect 17420 -4710 17520 -3050
rect 18100 -3150 18240 -2290
rect 18800 -2440 18900 -780
rect 19020 -1110 19120 550
rect 19700 450 19840 1310
rect 20400 1160 20500 1310
rect 20390 1150 20510 1160
rect 20390 1030 20400 1150
rect 20500 1030 20510 1150
rect 20390 1020 20510 1030
rect 19700 290 19710 450
rect 19830 290 19840 450
rect 19700 190 19840 290
rect 19700 -490 19710 190
rect 19830 -490 19840 190
rect 19010 -1120 19130 -1110
rect 19010 -1240 19020 -1120
rect 19120 -1240 19130 -1120
rect 19010 -1250 19130 -1240
rect 18790 -2450 18910 -2440
rect 18790 -2570 18800 -2450
rect 18900 -2570 18910 -2450
rect 18790 -2580 18910 -2570
rect 18100 -3310 18110 -3150
rect 18230 -3310 18240 -3150
rect 18100 -3410 18240 -3310
rect 18100 -4090 18110 -3410
rect 18230 -4090 18240 -3410
rect 18100 -4100 18240 -4090
rect 18800 -4240 18900 -2580
rect 19020 -2910 19120 -1250
rect 19700 -1350 19840 -490
rect 20400 -640 20500 1020
rect 20620 690 20720 1310
rect 20610 680 20730 690
rect 20610 560 20620 680
rect 20720 560 20730 680
rect 20610 550 20730 560
rect 20390 -650 20510 -640
rect 20390 -770 20400 -650
rect 20500 -770 20510 -650
rect 20390 -780 20510 -770
rect 19700 -1510 19710 -1350
rect 19830 -1510 19840 -1350
rect 19700 -1610 19840 -1510
rect 19700 -2290 19710 -1610
rect 19830 -2290 19840 -1610
rect 19010 -2920 19130 -2910
rect 19010 -3040 19020 -2920
rect 19120 -3040 19130 -2920
rect 19010 -3050 19130 -3040
rect 18790 -4250 18910 -4240
rect 18790 -4370 18800 -4250
rect 18900 -4370 18910 -4250
rect 18790 -4380 18910 -4370
rect 17410 -4720 17530 -4710
rect 17410 -4840 17420 -4720
rect 17520 -4840 17530 -4720
rect 17410 -4850 17530 -4840
rect 17420 -6760 17520 -4850
rect 18800 -5160 18900 -4380
rect 19020 -4710 19120 -3050
rect 19700 -3150 19840 -2290
rect 20400 -2440 20500 -780
rect 20620 -1110 20720 550
rect 21300 450 21440 1310
rect 22000 1160 22100 1310
rect 21990 1150 22110 1160
rect 21990 1030 22000 1150
rect 22100 1030 22110 1150
rect 21990 1020 22110 1030
rect 21300 290 21310 450
rect 21430 290 21440 450
rect 21300 190 21440 290
rect 21300 -490 21310 190
rect 21430 -490 21440 190
rect 20610 -1120 20730 -1110
rect 20610 -1240 20620 -1120
rect 20720 -1240 20730 -1120
rect 20610 -1250 20730 -1240
rect 20390 -2450 20510 -2440
rect 20390 -2570 20400 -2450
rect 20500 -2570 20510 -2450
rect 20390 -2580 20510 -2570
rect 19700 -3310 19710 -3150
rect 19830 -3310 19840 -3150
rect 19700 -3410 19840 -3310
rect 19700 -4090 19710 -3410
rect 19830 -4090 19840 -3410
rect 19700 -4100 19840 -4090
rect 20400 -4240 20500 -2580
rect 20620 -2910 20720 -1250
rect 21300 -1350 21440 -490
rect 22000 -640 22100 1020
rect 22220 690 22320 1310
rect 22210 680 22330 690
rect 22210 560 22220 680
rect 22320 560 22330 680
rect 22210 550 22330 560
rect 21990 -650 22110 -640
rect 21990 -770 22000 -650
rect 22100 -770 22110 -650
rect 21990 -780 22110 -770
rect 21300 -1510 21310 -1350
rect 21430 -1510 21440 -1350
rect 21300 -1610 21440 -1510
rect 21300 -2290 21310 -1610
rect 21430 -2290 21440 -1610
rect 20610 -2920 20730 -2910
rect 20610 -3040 20620 -2920
rect 20720 -3040 20730 -2920
rect 20610 -3050 20730 -3040
rect 20390 -4250 20510 -4240
rect 20390 -4370 20400 -4250
rect 20500 -4370 20510 -4250
rect 20390 -4380 20510 -4370
rect 19010 -4720 19130 -4710
rect 19010 -4840 19020 -4720
rect 19120 -4840 19130 -4720
rect 19010 -4850 19130 -4840
rect 18760 -5170 18940 -5160
rect 18760 -5350 18770 -5170
rect 18930 -5350 18940 -5170
rect 18760 -5360 18940 -5350
rect 18760 -5570 18940 -5560
rect 18760 -5750 18770 -5570
rect 18930 -5750 18940 -5570
rect 18760 -5760 18940 -5750
rect 17380 -6770 17560 -6760
rect 17380 -6950 17390 -6770
rect 17550 -6950 17560 -6770
rect 17380 -6960 17560 -6950
rect 17160 -7170 17340 -7160
rect 17160 -7350 17170 -7170
rect 17330 -7350 17340 -7170
rect 17160 -7360 17340 -7350
rect 17160 -7570 17340 -7560
rect 17160 -7750 17170 -7570
rect 17330 -7750 17340 -7570
rect 17160 -7760 17340 -7750
rect 15820 -8070 15960 -8060
rect 15820 -8190 15830 -8070
rect 15950 -8190 15960 -8070
rect 15820 -8200 15960 -8190
rect 15600 -8520 15740 -8510
rect 15600 -8640 15610 -8520
rect 15730 -8640 15740 -8520
rect 15600 -8650 15740 -8640
rect 15620 -10310 15720 -8650
rect 15840 -9860 15940 -8200
rect 16500 -8260 16650 -8250
rect 16500 -8380 16510 -8260
rect 16640 -8380 16650 -8260
rect 16500 -8390 16650 -8380
rect 17220 -8510 17320 -7760
rect 17440 -8060 17540 -6960
rect 17420 -8070 17560 -8060
rect 17420 -8190 17430 -8070
rect 17550 -8190 17560 -8070
rect 17420 -8200 17560 -8190
rect 17200 -8520 17340 -8510
rect 17200 -8640 17210 -8520
rect 17330 -8640 17340 -8520
rect 17200 -8650 17340 -8640
rect 16510 -8800 16640 -8790
rect 16510 -9480 16520 -8800
rect 16630 -9480 16640 -8800
rect 16510 -9560 16640 -9480
rect 16500 -9570 16650 -9560
rect 16500 -9730 16510 -9570
rect 16640 -9730 16650 -9570
rect 16500 -9740 16650 -9730
rect 15820 -9870 15960 -9860
rect 15820 -9990 15830 -9870
rect 15950 -9990 15960 -9870
rect 15820 -10000 15960 -9990
rect 15600 -10320 15740 -10310
rect 15600 -10440 15610 -10320
rect 15730 -10440 15740 -10320
rect 15600 -10450 15740 -10440
rect 14900 -12100 15050 -12090
rect 14900 -12230 14910 -12100
rect 15040 -12230 15050 -12100
rect 15620 -12110 15720 -10450
rect 15840 -11660 15940 -10000
rect 16510 -10600 16640 -9740
rect 17220 -10310 17320 -8650
rect 17440 -9860 17540 -8200
rect 18820 -8510 18920 -5760
rect 19020 -5960 19120 -4850
rect 18980 -5970 19160 -5960
rect 18980 -6150 18990 -5970
rect 19150 -6150 19160 -5970
rect 18980 -6160 19160 -6150
rect 19040 -8060 19140 -6160
rect 20400 -7160 20500 -4380
rect 20620 -4710 20720 -3050
rect 21300 -3150 21440 -2290
rect 22000 -2440 22100 -780
rect 22220 -1110 22320 550
rect 22900 450 23040 1310
rect 23600 1160 23700 1310
rect 23590 1150 23710 1160
rect 23590 1030 23600 1150
rect 23700 1030 23710 1150
rect 23590 1020 23710 1030
rect 22900 290 22910 450
rect 23030 290 23040 450
rect 22900 190 23040 290
rect 22900 -490 22910 190
rect 23030 -490 23040 190
rect 22210 -1120 22330 -1110
rect 22210 -1240 22220 -1120
rect 22320 -1240 22330 -1120
rect 22210 -1250 22330 -1240
rect 21990 -2450 22110 -2440
rect 21990 -2570 22000 -2450
rect 22100 -2570 22110 -2450
rect 21990 -2580 22110 -2570
rect 21300 -3310 21310 -3150
rect 21430 -3310 21440 -3150
rect 21300 -3410 21440 -3310
rect 21300 -4090 21310 -3410
rect 21430 -4090 21440 -3410
rect 21300 -4100 21440 -4090
rect 22000 -4240 22100 -2580
rect 22220 -2910 22320 -1250
rect 22900 -1350 23040 -490
rect 23600 -640 23700 1020
rect 23820 690 23920 1310
rect 23810 680 23930 690
rect 23810 560 23820 680
rect 23920 560 23930 680
rect 23810 550 23930 560
rect 23590 -650 23710 -640
rect 23590 -770 23600 -650
rect 23700 -770 23710 -650
rect 23590 -780 23710 -770
rect 22900 -1510 22910 -1350
rect 23030 -1510 23040 -1350
rect 22900 -1610 23040 -1510
rect 22900 -2290 22910 -1610
rect 23030 -2290 23040 -1610
rect 22210 -2920 22330 -2910
rect 22210 -3040 22220 -2920
rect 22320 -3040 22330 -2920
rect 22210 -3050 22330 -3040
rect 21990 -4250 22110 -4240
rect 21990 -4370 22000 -4250
rect 22100 -4370 22110 -4250
rect 21990 -4380 22110 -4370
rect 20610 -4720 20730 -4710
rect 20610 -4840 20620 -4720
rect 20720 -4840 20730 -4720
rect 20610 -4850 20730 -4840
rect 20620 -6760 20720 -4850
rect 22000 -5160 22100 -4380
rect 22220 -4710 22320 -3050
rect 22900 -3150 23040 -2290
rect 23600 -2440 23700 -780
rect 23820 -1110 23920 550
rect 24500 450 24640 1310
rect 24500 290 24510 450
rect 24630 290 24640 450
rect 24500 190 24640 290
rect 24500 -490 24510 190
rect 24630 -490 24640 190
rect 23810 -1120 23930 -1110
rect 23810 -1240 23820 -1120
rect 23920 -1240 23930 -1120
rect 23810 -1250 23930 -1240
rect 23590 -2450 23710 -2440
rect 23590 -2570 23600 -2450
rect 23700 -2570 23710 -2450
rect 23590 -2580 23710 -2570
rect 22900 -3310 22910 -3150
rect 23030 -3310 23040 -3150
rect 22900 -3410 23040 -3310
rect 22900 -4090 22910 -3410
rect 23030 -4090 23040 -3410
rect 22900 -4100 23040 -4090
rect 23600 -4240 23700 -2580
rect 23820 -2910 23920 -1250
rect 24500 -1350 24640 -490
rect 24500 -1510 24510 -1350
rect 24630 -1510 24640 -1350
rect 24500 -1610 24640 -1510
rect 24500 -2290 24510 -1610
rect 24630 -2290 24640 -1610
rect 23810 -2920 23930 -2910
rect 23810 -3040 23820 -2920
rect 23920 -3040 23930 -2920
rect 23810 -3050 23930 -3040
rect 23590 -4250 23710 -4240
rect 23590 -4370 23600 -4250
rect 23700 -4370 23710 -4250
rect 23590 -4380 23710 -4370
rect 22210 -4720 22330 -4710
rect 22210 -4840 22220 -4720
rect 22320 -4840 22330 -4720
rect 22210 -4850 22330 -4840
rect 21960 -5170 22140 -5160
rect 21960 -5350 21970 -5170
rect 22130 -5350 22140 -5170
rect 21960 -5360 22140 -5350
rect 21960 -5570 22140 -5560
rect 21960 -5750 21970 -5570
rect 22130 -5750 22140 -5570
rect 21960 -5760 22140 -5750
rect 20580 -6770 20760 -6760
rect 20580 -6950 20590 -6770
rect 20750 -6950 20760 -6770
rect 20580 -6960 20760 -6950
rect 20360 -7170 20540 -7160
rect 20360 -7350 20370 -7170
rect 20530 -7350 20540 -7170
rect 20360 -7360 20540 -7350
rect 20360 -7570 20540 -7560
rect 20360 -7750 20370 -7570
rect 20530 -7750 20540 -7570
rect 20360 -7760 20540 -7750
rect 19020 -8070 19160 -8060
rect 19020 -8190 19030 -8070
rect 19150 -8190 19160 -8070
rect 19020 -8200 19160 -8190
rect 18800 -8520 18940 -8510
rect 18800 -8640 18810 -8520
rect 18930 -8640 18940 -8520
rect 18800 -8650 18940 -8640
rect 18110 -8800 18240 -8790
rect 18110 -9480 18120 -8800
rect 18230 -9480 18240 -8800
rect 18110 -9560 18240 -9480
rect 18100 -9570 18250 -9560
rect 18100 -9730 18110 -9570
rect 18240 -9730 18250 -9570
rect 18100 -9740 18250 -9730
rect 17420 -9870 17560 -9860
rect 17420 -9990 17430 -9870
rect 17550 -9990 17560 -9870
rect 17420 -10000 17560 -9990
rect 17200 -10320 17340 -10310
rect 17200 -10440 17210 -10320
rect 17330 -10440 17340 -10320
rect 17200 -10450 17340 -10440
rect 16510 -11280 16520 -10600
rect 16630 -11280 16640 -10600
rect 16510 -11360 16640 -11280
rect 16500 -11370 16650 -11360
rect 16500 -11530 16510 -11370
rect 16640 -11530 16650 -11370
rect 16500 -11540 16650 -11530
rect 15820 -11670 15960 -11660
rect 15820 -11790 15830 -11670
rect 15950 -11790 15960 -11670
rect 15820 -11800 15960 -11790
rect 14900 -12240 15050 -12230
rect 15600 -12120 15740 -12110
rect 15600 -12240 15610 -12120
rect 15730 -12240 15740 -12120
rect 15600 -12250 15740 -12240
rect 14910 -12410 15040 -12400
rect 14910 -13070 14920 -12410
rect 15030 -13070 15040 -12410
rect 14910 -13160 15040 -13070
rect 14880 -13170 15070 -13160
rect 14880 -13330 14890 -13170
rect 15060 -13330 15070 -13170
rect 14880 -13340 15070 -13330
rect 14910 -14210 15040 -13340
rect 15620 -13910 15720 -12250
rect 15840 -13460 15940 -11800
rect 16510 -12400 16640 -11540
rect 17220 -12110 17320 -10450
rect 17440 -11660 17540 -10000
rect 18110 -10600 18240 -9740
rect 18820 -10310 18920 -8650
rect 19040 -9860 19140 -8200
rect 20420 -8510 20520 -7760
rect 20640 -8060 20740 -6960
rect 20620 -8070 20760 -8060
rect 20620 -8190 20630 -8070
rect 20750 -8190 20760 -8070
rect 20620 -8200 20760 -8190
rect 20400 -8520 20540 -8510
rect 20400 -8640 20410 -8520
rect 20530 -8640 20540 -8520
rect 20400 -8650 20540 -8640
rect 19710 -8800 19840 -8790
rect 19710 -9480 19720 -8800
rect 19830 -9480 19840 -8800
rect 19710 -9560 19840 -9480
rect 19700 -9570 19850 -9560
rect 19700 -9730 19710 -9570
rect 19840 -9730 19850 -9570
rect 19700 -9740 19850 -9730
rect 19020 -9870 19160 -9860
rect 19020 -9990 19030 -9870
rect 19150 -9990 19160 -9870
rect 19020 -10000 19160 -9990
rect 18800 -10320 18940 -10310
rect 18800 -10440 18810 -10320
rect 18930 -10440 18940 -10320
rect 18800 -10450 18940 -10440
rect 18110 -11280 18120 -10600
rect 18230 -11280 18240 -10600
rect 18110 -11360 18240 -11280
rect 18100 -11370 18250 -11360
rect 18100 -11530 18110 -11370
rect 18240 -11530 18250 -11370
rect 18100 -11540 18250 -11530
rect 17420 -11670 17560 -11660
rect 17420 -11790 17430 -11670
rect 17550 -11790 17560 -11670
rect 17420 -11800 17560 -11790
rect 17200 -12120 17340 -12110
rect 17200 -12240 17210 -12120
rect 17330 -12240 17340 -12120
rect 17200 -12250 17340 -12240
rect 16510 -13080 16520 -12400
rect 16630 -13080 16640 -12400
rect 16510 -13160 16640 -13080
rect 16500 -13170 16650 -13160
rect 16500 -13330 16510 -13170
rect 16640 -13330 16650 -13170
rect 16500 -13340 16650 -13330
rect 15820 -13470 15960 -13460
rect 15820 -13590 15830 -13470
rect 15950 -13590 15960 -13470
rect 15820 -13600 15960 -13590
rect 15600 -13920 15740 -13910
rect 15600 -14040 15610 -13920
rect 15730 -14040 15740 -13920
rect 15600 -14050 15740 -14040
rect 14910 -14870 14920 -14210
rect 15030 -14870 15040 -14210
rect 14910 -14960 15040 -14870
rect 14880 -14970 15070 -14960
rect 14880 -15130 14890 -14970
rect 15060 -15130 15070 -14970
rect 14880 -15140 15070 -15130
rect 14910 -15290 15040 -15280
rect 14910 -15390 14930 -15290
rect 15030 -15390 15040 -15290
rect 14910 -16010 15040 -15390
rect 15620 -15710 15720 -14050
rect 15840 -15260 15940 -13600
rect 16510 -14200 16640 -13340
rect 17220 -13910 17320 -12250
rect 17440 -13460 17540 -11800
rect 18110 -12400 18240 -11540
rect 18820 -12110 18920 -10450
rect 19040 -11660 19140 -10000
rect 19710 -10600 19840 -9740
rect 20420 -10310 20520 -8650
rect 20640 -9860 20740 -8200
rect 22020 -8510 22120 -5760
rect 22220 -5960 22320 -4850
rect 22180 -5970 22360 -5960
rect 22180 -6150 22190 -5970
rect 22350 -6150 22360 -5970
rect 22180 -6160 22360 -6150
rect 22240 -8060 22340 -6160
rect 23600 -7160 23700 -4380
rect 23820 -4710 23920 -3050
rect 24500 -3150 24640 -2290
rect 25200 -2440 25300 1310
rect 25190 -2450 25310 -2440
rect 25190 -2570 25200 -2450
rect 25300 -2570 25310 -2450
rect 25190 -2580 25310 -2570
rect 24500 -3310 24510 -3150
rect 24630 -3310 24640 -3150
rect 24500 -3410 24640 -3310
rect 24500 -4090 24510 -3410
rect 24630 -4090 24640 -3410
rect 24500 -4100 24640 -4090
rect 25200 -4240 25300 -2580
rect 25420 -2910 25520 1310
rect 26100 450 26240 1310
rect 26800 1160 26900 1310
rect 26790 1150 26910 1160
rect 26790 1030 26800 1150
rect 26900 1030 26910 1150
rect 26790 1020 26910 1030
rect 26100 290 26110 450
rect 26230 290 26240 450
rect 26100 190 26240 290
rect 26100 -490 26110 190
rect 26230 -490 26240 190
rect 26100 -1350 26240 -490
rect 26800 -640 26900 1020
rect 27020 690 27120 1310
rect 27010 680 27130 690
rect 27010 560 27020 680
rect 27120 560 27130 680
rect 27010 550 27130 560
rect 26790 -650 26910 -640
rect 26790 -770 26800 -650
rect 26900 -770 26910 -650
rect 26790 -780 26910 -770
rect 26100 -1510 26110 -1350
rect 26230 -1510 26240 -1350
rect 26100 -1610 26240 -1510
rect 26100 -2290 26110 -1610
rect 26230 -2290 26240 -1610
rect 25410 -2920 25530 -2910
rect 25410 -3040 25420 -2920
rect 25520 -3040 25530 -2920
rect 25410 -3050 25530 -3040
rect 25190 -4250 25310 -4240
rect 25190 -4370 25200 -4250
rect 25300 -4370 25310 -4250
rect 25190 -4380 25310 -4370
rect 23810 -4720 23930 -4710
rect 23810 -4840 23820 -4720
rect 23920 -4840 23930 -4720
rect 23810 -4850 23930 -4840
rect 23820 -6760 23920 -4850
rect 25200 -5160 25300 -4380
rect 25420 -4710 25520 -3050
rect 26100 -3150 26240 -2290
rect 26800 -2440 26900 -780
rect 27020 -1110 27120 550
rect 27700 450 27840 1310
rect 28400 1160 28500 1310
rect 28391 1150 28510 1160
rect 28391 1030 28400 1150
rect 28500 1030 28510 1150
rect 28391 1020 28510 1030
rect 27700 270 27710 450
rect 27830 270 27840 450
rect 27700 190 27840 270
rect 27700 -490 27710 190
rect 27830 -490 27840 190
rect 27010 -1120 27130 -1110
rect 27010 -1240 27020 -1120
rect 27120 -1240 27130 -1120
rect 27010 -1250 27130 -1240
rect 26791 -2450 26910 -2440
rect 26791 -2570 26800 -2450
rect 26900 -2570 26910 -2450
rect 26791 -2580 26910 -2570
rect 26100 -3310 26110 -3150
rect 26230 -3310 26240 -3150
rect 26100 -3410 26240 -3310
rect 26100 -4090 26110 -3410
rect 26230 -4090 26240 -3410
rect 26100 -4100 26240 -4090
rect 26800 -4240 26900 -2580
rect 27020 -2910 27120 -1250
rect 27700 -1350 27840 -490
rect 28400 -640 28500 1020
rect 28620 690 28720 1310
rect 28611 680 28730 690
rect 28611 560 28620 680
rect 28720 560 28730 680
rect 28611 550 28730 560
rect 28391 -650 28510 -640
rect 28391 -770 28400 -650
rect 28500 -770 28510 -650
rect 28391 -780 28510 -770
rect 27700 -1530 27710 -1350
rect 27830 -1530 27840 -1350
rect 27700 -1610 27840 -1530
rect 27700 -2290 27710 -1610
rect 27830 -2290 27840 -1610
rect 27011 -2920 27130 -2910
rect 27011 -3040 27020 -2920
rect 27120 -3040 27130 -2920
rect 27011 -3050 27130 -3040
rect 26791 -4250 26910 -4240
rect 26791 -4370 26800 -4250
rect 26900 -4370 26910 -4250
rect 26791 -4380 26910 -4370
rect 25410 -4720 25530 -4710
rect 25410 -4840 25420 -4720
rect 25520 -4840 25530 -4720
rect 25410 -4850 25530 -4840
rect 25160 -5170 25340 -5160
rect 25160 -5350 25170 -5170
rect 25330 -5350 25340 -5170
rect 25160 -5360 25340 -5350
rect 25160 -5570 25340 -5560
rect 25160 -5750 25170 -5570
rect 25330 -5750 25340 -5570
rect 25160 -5760 25340 -5750
rect 23780 -6770 23960 -6760
rect 23780 -6950 23790 -6770
rect 23950 -6950 23960 -6770
rect 23780 -6960 23960 -6950
rect 23560 -7170 23740 -7160
rect 23560 -7350 23570 -7170
rect 23730 -7350 23740 -7170
rect 23560 -7360 23740 -7350
rect 23560 -7570 23740 -7560
rect 23560 -7750 23570 -7570
rect 23730 -7750 23740 -7570
rect 23560 -7760 23740 -7750
rect 22220 -8070 22360 -8060
rect 22220 -8190 22230 -8070
rect 22350 -8190 22360 -8070
rect 22220 -8200 22360 -8190
rect 22000 -8520 22140 -8510
rect 22000 -8640 22010 -8520
rect 22130 -8640 22140 -8520
rect 22000 -8650 22140 -8640
rect 21310 -8800 21440 -8790
rect 21310 -9480 21320 -8800
rect 21430 -9480 21440 -8800
rect 21310 -9560 21440 -9480
rect 21300 -9570 21450 -9560
rect 21300 -9730 21310 -9570
rect 21440 -9730 21450 -9570
rect 21300 -9740 21450 -9730
rect 20620 -9870 20760 -9860
rect 20620 -9990 20630 -9870
rect 20750 -9990 20760 -9870
rect 20620 -10000 20760 -9990
rect 20400 -10320 20540 -10310
rect 20400 -10440 20410 -10320
rect 20530 -10440 20540 -10320
rect 20400 -10450 20540 -10440
rect 19710 -11280 19720 -10600
rect 19830 -11280 19840 -10600
rect 19710 -11360 19840 -11280
rect 19700 -11370 19850 -11360
rect 19700 -11530 19710 -11370
rect 19840 -11530 19850 -11370
rect 19700 -11540 19850 -11530
rect 19020 -11670 19160 -11660
rect 19020 -11790 19030 -11670
rect 19150 -11790 19160 -11670
rect 19020 -11800 19160 -11790
rect 18800 -12120 18940 -12110
rect 18800 -12240 18810 -12120
rect 18930 -12240 18940 -12120
rect 18800 -12250 18940 -12240
rect 18110 -13080 18120 -12400
rect 18230 -13080 18240 -12400
rect 18110 -13160 18240 -13080
rect 18100 -13170 18250 -13160
rect 18100 -13330 18110 -13170
rect 18240 -13330 18250 -13170
rect 18100 -13340 18250 -13330
rect 17420 -13470 17560 -13460
rect 17420 -13590 17430 -13470
rect 17550 -13590 17560 -13470
rect 17420 -13600 17560 -13590
rect 17200 -13920 17340 -13910
rect 17200 -14040 17210 -13920
rect 17330 -14040 17340 -13920
rect 17200 -14050 17340 -14040
rect 16510 -14880 16520 -14200
rect 16630 -14880 16640 -14200
rect 16510 -14960 16640 -14880
rect 16500 -14970 16650 -14960
rect 16500 -15130 16510 -14970
rect 16640 -15130 16650 -14970
rect 16500 -15140 16650 -15130
rect 15820 -15270 15960 -15260
rect 15820 -15390 15830 -15270
rect 15950 -15390 15960 -15270
rect 15820 -15400 15960 -15390
rect 15600 -15720 15740 -15710
rect 15600 -15840 15610 -15720
rect 15730 -15840 15740 -15720
rect 15600 -15850 15740 -15840
rect 14910 -16670 14920 -16010
rect 15030 -16670 15040 -16010
rect 14910 -16680 15040 -16670
rect 14910 -16780 15030 -16680
rect 14890 -16790 15060 -16780
rect 14890 -16950 14900 -16790
rect 15050 -16950 15060 -16790
rect 14890 -16960 15060 -16950
rect 14910 -17800 15030 -16960
rect 15620 -17510 15720 -15850
rect 15840 -17060 15940 -15400
rect 16510 -16000 16640 -15140
rect 17220 -15710 17320 -14050
rect 17440 -15260 17540 -13600
rect 18110 -14200 18240 -13340
rect 18820 -13910 18920 -12250
rect 19040 -13460 19140 -11800
rect 19710 -12400 19840 -11540
rect 20420 -12110 20520 -10450
rect 20640 -11660 20740 -10000
rect 21310 -10600 21440 -9740
rect 22020 -10310 22120 -8650
rect 22240 -9860 22340 -8200
rect 23620 -8510 23720 -7760
rect 23840 -8060 23940 -6960
rect 23820 -8070 23960 -8060
rect 23820 -8190 23830 -8070
rect 23950 -8190 23960 -8070
rect 23820 -8200 23960 -8190
rect 23600 -8520 23740 -8510
rect 23600 -8640 23610 -8520
rect 23730 -8640 23740 -8520
rect 23600 -8650 23740 -8640
rect 22910 -8800 23040 -8790
rect 22910 -9480 22920 -8800
rect 23030 -9480 23040 -8800
rect 22910 -9560 23040 -9480
rect 22900 -9570 23050 -9560
rect 22900 -9730 22910 -9570
rect 23040 -9730 23050 -9570
rect 22900 -9740 23050 -9730
rect 22220 -9870 22360 -9860
rect 22220 -9990 22230 -9870
rect 22350 -9990 22360 -9870
rect 22220 -10000 22360 -9990
rect 22000 -10320 22140 -10310
rect 22000 -10440 22010 -10320
rect 22130 -10440 22140 -10320
rect 22000 -10450 22140 -10440
rect 21310 -11280 21320 -10600
rect 21430 -11280 21440 -10600
rect 21310 -11360 21440 -11280
rect 21300 -11370 21450 -11360
rect 21300 -11530 21310 -11370
rect 21440 -11530 21450 -11370
rect 21300 -11540 21450 -11530
rect 20620 -11670 20760 -11660
rect 20620 -11790 20630 -11670
rect 20750 -11790 20760 -11670
rect 20620 -11800 20760 -11790
rect 20400 -12120 20540 -12110
rect 20400 -12240 20410 -12120
rect 20530 -12240 20540 -12120
rect 20400 -12250 20540 -12240
rect 19710 -13080 19720 -12400
rect 19830 -13080 19840 -12400
rect 19710 -13160 19840 -13080
rect 19700 -13170 19850 -13160
rect 19700 -13330 19710 -13170
rect 19840 -13330 19850 -13170
rect 19700 -13340 19850 -13330
rect 19020 -13470 19160 -13460
rect 19020 -13590 19030 -13470
rect 19150 -13590 19160 -13470
rect 19020 -13600 19160 -13590
rect 18800 -13920 18940 -13910
rect 18800 -14040 18810 -13920
rect 18930 -14040 18940 -13920
rect 18800 -14050 18940 -14040
rect 18110 -14880 18120 -14200
rect 18230 -14880 18240 -14200
rect 18110 -14960 18240 -14880
rect 18100 -14970 18250 -14960
rect 18100 -15130 18110 -14970
rect 18240 -15130 18250 -14970
rect 18100 -15140 18250 -15130
rect 17420 -15270 17560 -15260
rect 17420 -15390 17430 -15270
rect 17550 -15390 17560 -15270
rect 17420 -15400 17560 -15390
rect 17200 -15720 17340 -15710
rect 17200 -15840 17210 -15720
rect 17330 -15840 17340 -15720
rect 17200 -15850 17340 -15840
rect 16510 -16680 16520 -16000
rect 16630 -16680 16640 -16000
rect 16510 -16760 16640 -16680
rect 16500 -16770 16650 -16760
rect 16500 -16930 16510 -16770
rect 16640 -16930 16650 -16770
rect 16500 -16940 16650 -16930
rect 15820 -17070 15960 -17060
rect 15820 -17190 15830 -17070
rect 15950 -17190 15960 -17070
rect 15820 -17200 15960 -17190
rect 15600 -17520 15740 -17510
rect 15600 -17640 15610 -17520
rect 15730 -17640 15740 -17520
rect 15600 -17650 15740 -17640
rect 14910 -17810 15040 -17800
rect 14910 -18470 14920 -17810
rect 15030 -18470 15040 -17810
rect 14910 -18580 15040 -18470
rect 14890 -18590 15060 -18580
rect 14890 -18750 14900 -18590
rect 15050 -18750 15060 -18590
rect 14890 -18760 15060 -18750
rect 15620 -19310 15720 -17650
rect 15840 -18860 15940 -17200
rect 16510 -17800 16640 -16940
rect 17220 -17510 17320 -15850
rect 17440 -17060 17540 -15400
rect 18110 -16000 18240 -15140
rect 18820 -15710 18920 -14050
rect 19040 -15260 19140 -13600
rect 19710 -14200 19840 -13340
rect 20420 -13910 20520 -12250
rect 20640 -13460 20740 -11800
rect 21310 -12400 21440 -11540
rect 22020 -12110 22120 -10450
rect 22240 -11660 22340 -10000
rect 22910 -10600 23040 -9740
rect 23620 -10310 23720 -8650
rect 23840 -9860 23940 -8200
rect 25220 -8510 25320 -5760
rect 25420 -5960 25520 -4850
rect 25380 -5970 25560 -5960
rect 25380 -6150 25390 -5970
rect 25550 -6150 25560 -5970
rect 25380 -6160 25560 -6150
rect 25440 -8060 25540 -6160
rect 26800 -7160 26900 -4380
rect 27020 -4710 27120 -3050
rect 27700 -3150 27840 -2290
rect 28400 -2440 28500 -780
rect 28620 -1110 28720 550
rect 29300 450 29440 1310
rect 29300 270 29310 450
rect 29430 270 29440 450
rect 29300 190 29440 270
rect 29300 -490 29310 190
rect 29430 -490 29440 190
rect 28611 -1120 28730 -1110
rect 28611 -1240 28620 -1120
rect 28720 -1240 28730 -1120
rect 28611 -1250 28730 -1240
rect 28390 -2450 28510 -2440
rect 28390 -2570 28400 -2450
rect 28500 -2570 28510 -2450
rect 28390 -2580 28510 -2570
rect 27700 -3330 27710 -3150
rect 27830 -3330 27840 -3150
rect 27700 -3410 27840 -3330
rect 27700 -4090 27710 -3410
rect 27830 -4090 27840 -3410
rect 27011 -4720 27130 -4710
rect 27011 -4840 27020 -4720
rect 27120 -4840 27130 -4720
rect 27011 -4850 27130 -4840
rect 27020 -6760 27120 -4850
rect 27700 -5960 27840 -4090
rect 28400 -4240 28500 -2580
rect 28620 -2910 28720 -1250
rect 29300 -1350 29440 -490
rect 29300 -1530 29310 -1350
rect 29430 -1530 29440 -1350
rect 29300 -1610 29440 -1530
rect 29300 -2290 29310 -1610
rect 29430 -2290 29440 -1610
rect 28610 -2920 28730 -2910
rect 28610 -3040 28620 -2920
rect 28720 -3040 28730 -2920
rect 28610 -3050 28730 -3040
rect 28390 -4250 28510 -4240
rect 28390 -4370 28400 -4250
rect 28500 -4370 28510 -4250
rect 28390 -4380 28510 -4370
rect 28400 -5160 28500 -4380
rect 28620 -4710 28720 -3050
rect 29300 -3150 29440 -2290
rect 30900 2250 31040 2260
rect 30900 2070 30910 2250
rect 31030 2070 31040 2250
rect 30900 1990 31040 2070
rect 30900 1310 30910 1990
rect 31030 1310 31040 1990
rect 30900 450 31040 1310
rect 30900 270 30910 450
rect 31030 270 31040 450
rect 30900 190 31040 270
rect 30900 -490 30910 190
rect 31030 -490 31040 190
rect 30900 -1350 31040 -490
rect 31600 -1110 31700 3540
rect 32530 3162 32620 4330
rect 33120 4110 33300 4120
rect 33120 4080 33130 4110
rect 32800 4070 33130 4080
rect 33290 4080 33300 4110
rect 33290 4070 33940 4080
rect 32800 4010 32810 4070
rect 32980 4010 33130 4070
rect 33300 4010 33440 4070
rect 33610 4010 33760 4070
rect 33930 4010 33940 4070
rect 32800 4000 33940 4010
rect 32840 3430 33880 3440
rect 32840 3350 32850 3430
rect 33870 3350 33880 3430
rect 32840 3340 33880 3350
rect 32460 3156 32674 3162
rect 31820 3090 32000 3100
rect 31820 2910 31830 3090
rect 31990 2910 32000 3090
rect 32460 3068 32466 3156
rect 32668 3068 32674 3156
rect 32460 3062 32674 3068
rect 31820 2900 32000 2910
rect 31820 690 31920 2900
rect 33170 2550 33340 2560
rect 32440 2510 32700 2520
rect 32440 2430 32450 2510
rect 32690 2430 32700 2510
rect 32440 2130 32700 2430
rect 33170 2390 33180 2550
rect 33330 2390 33340 2550
rect 33170 2380 33340 2390
rect 32440 2070 32450 2130
rect 32690 2070 32700 2130
rect 32440 2060 32700 2070
rect 32500 1990 32640 2000
rect 32500 1310 32510 1990
rect 32630 1310 32640 1990
rect 32500 1150 32640 1310
rect 32500 1030 32510 1150
rect 32630 1030 32640 1150
rect 32500 1020 32640 1030
rect 31810 680 31930 690
rect 31810 560 31820 680
rect 31920 560 31930 680
rect 31810 550 31930 560
rect 33190 450 33320 2380
rect 33170 440 33340 450
rect 33170 280 33180 440
rect 33330 280 33340 440
rect 33170 270 33340 280
rect 32500 190 32640 200
rect 32500 -490 32510 190
rect 32630 -490 32640 190
rect 32500 -500 32640 -490
rect 31590 -1120 31710 -1110
rect 31590 -1240 31600 -1120
rect 31700 -1240 31710 -1120
rect 31590 -1250 31710 -1240
rect 30900 -1530 30910 -1350
rect 31030 -1530 31040 -1350
rect 33440 -1460 33560 3340
rect 34120 3162 34210 4330
rect 35690 4290 35850 4300
rect 35690 4150 35700 4290
rect 35840 4150 35850 4290
rect 35690 4140 35850 4150
rect 36290 4260 36300 4330
rect 36390 4260 36400 4330
rect 34860 4090 35200 4100
rect 34860 4010 34870 4090
rect 35190 4010 35200 4090
rect 34860 4000 35200 4010
rect 35040 3430 35420 3440
rect 35040 3350 35070 3430
rect 35410 3350 35420 3430
rect 35040 3340 35420 3350
rect 34060 3156 34274 3162
rect 34060 3068 34066 3156
rect 34268 3068 34274 3156
rect 34060 3062 34274 3068
rect 34770 2780 34940 2790
rect 34770 2620 34780 2780
rect 34930 2620 34940 2780
rect 34770 2610 34940 2620
rect 34040 2510 34300 2520
rect 34040 2430 34050 2510
rect 34290 2430 34300 2510
rect 34040 2130 34300 2430
rect 34040 2070 34050 2130
rect 34290 2070 34300 2130
rect 34040 2060 34300 2070
rect 34100 1990 34240 2000
rect 34100 1310 34110 1990
rect 34230 1310 34240 1990
rect 34100 1150 34240 1310
rect 34790 1160 34920 2610
rect 34100 1030 34110 1150
rect 34230 1030 34240 1150
rect 34100 1020 34240 1030
rect 34780 1150 34930 1160
rect 34780 1030 34790 1150
rect 34920 1030 34930 1150
rect 34780 1020 34930 1030
rect 34100 190 34240 200
rect 34100 -490 34110 190
rect 34230 -490 34240 190
rect 34100 -500 34240 -490
rect 30900 -1610 31040 -1530
rect 33350 -1470 33560 -1460
rect 33350 -1590 33360 -1470
rect 33480 -1590 33560 -1470
rect 33350 -1600 33560 -1590
rect 30900 -2290 30910 -1610
rect 31030 -2290 31040 -1610
rect 29990 -2450 30110 -2440
rect 29990 -2570 30000 -2450
rect 30100 -2570 30110 -2450
rect 29990 -2580 30110 -2570
rect 29300 -3330 29310 -3150
rect 29430 -3330 29440 -3150
rect 29300 -3410 29440 -3330
rect 29300 -4090 29310 -3410
rect 29430 -4090 29440 -3410
rect 28610 -4720 28730 -4710
rect 28610 -4840 28620 -4720
rect 28720 -4840 28730 -4720
rect 28610 -4850 28730 -4840
rect 28360 -5170 28540 -5160
rect 28360 -5350 28370 -5170
rect 28530 -5350 28540 -5170
rect 28360 -5360 28540 -5350
rect 28360 -5570 28540 -5560
rect 28360 -5750 28370 -5570
rect 28530 -5750 28540 -5570
rect 28360 -5760 28540 -5750
rect 27680 -5970 27860 -5960
rect 27680 -6150 27690 -5970
rect 27850 -6150 27860 -5970
rect 27680 -6160 27860 -6150
rect 26980 -6770 27160 -6760
rect 26980 -6950 26990 -6770
rect 27150 -6950 27160 -6770
rect 26980 -6960 27160 -6950
rect 26760 -7170 26940 -7160
rect 26760 -7350 26770 -7170
rect 26930 -7350 26940 -7170
rect 26760 -7360 26940 -7350
rect 26760 -7570 26940 -7560
rect 26760 -7750 26770 -7570
rect 26930 -7750 26940 -7570
rect 26760 -7760 26940 -7750
rect 25420 -8070 25560 -8060
rect 25420 -8190 25430 -8070
rect 25550 -8190 25560 -8070
rect 25420 -8200 25560 -8190
rect 25200 -8520 25340 -8510
rect 25200 -8640 25210 -8520
rect 25330 -8640 25340 -8520
rect 25200 -8650 25340 -8640
rect 24510 -8800 24640 -8790
rect 24510 -9480 24520 -8800
rect 24630 -9480 24640 -8800
rect 24510 -9560 24640 -9480
rect 24500 -9570 24650 -9560
rect 24500 -9730 24510 -9570
rect 24640 -9730 24650 -9570
rect 24500 -9740 24650 -9730
rect 23820 -9870 23960 -9860
rect 23820 -9990 23830 -9870
rect 23950 -9990 23960 -9870
rect 23820 -10000 23960 -9990
rect 23600 -10320 23740 -10310
rect 23600 -10440 23610 -10320
rect 23730 -10440 23740 -10320
rect 23600 -10450 23740 -10440
rect 22910 -11280 22920 -10600
rect 23030 -11280 23040 -10600
rect 22910 -11360 23040 -11280
rect 22900 -11370 23050 -11360
rect 22900 -11530 22910 -11370
rect 23040 -11530 23050 -11370
rect 22900 -11540 23050 -11530
rect 22220 -11670 22360 -11660
rect 22220 -11790 22230 -11670
rect 22350 -11790 22360 -11670
rect 22220 -11800 22360 -11790
rect 22000 -12120 22140 -12110
rect 22000 -12240 22010 -12120
rect 22130 -12240 22140 -12120
rect 22000 -12250 22140 -12240
rect 21310 -13080 21320 -12400
rect 21430 -13080 21440 -12400
rect 21310 -13160 21440 -13080
rect 21300 -13170 21450 -13160
rect 21300 -13330 21310 -13170
rect 21440 -13330 21450 -13170
rect 21300 -13340 21450 -13330
rect 20620 -13470 20760 -13460
rect 20620 -13590 20630 -13470
rect 20750 -13590 20760 -13470
rect 20620 -13600 20760 -13590
rect 20400 -13920 20540 -13910
rect 20400 -14040 20410 -13920
rect 20530 -14040 20540 -13920
rect 20400 -14050 20540 -14040
rect 19710 -14880 19720 -14200
rect 19830 -14880 19840 -14200
rect 19710 -14960 19840 -14880
rect 19700 -14970 19850 -14960
rect 19700 -15130 19710 -14970
rect 19840 -15130 19850 -14970
rect 19700 -15140 19850 -15130
rect 19020 -15270 19160 -15260
rect 19020 -15390 19030 -15270
rect 19150 -15390 19160 -15270
rect 19020 -15400 19160 -15390
rect 18800 -15720 18940 -15710
rect 18800 -15840 18810 -15720
rect 18930 -15840 18940 -15720
rect 18800 -15850 18940 -15840
rect 18110 -16680 18120 -16000
rect 18230 -16680 18240 -16000
rect 18110 -16760 18240 -16680
rect 18100 -16770 18250 -16760
rect 18100 -16930 18110 -16770
rect 18240 -16930 18250 -16770
rect 18100 -16940 18250 -16930
rect 17420 -17070 17560 -17060
rect 17420 -17190 17430 -17070
rect 17550 -17190 17560 -17070
rect 17420 -17200 17560 -17190
rect 17200 -17520 17340 -17510
rect 17200 -17640 17210 -17520
rect 17330 -17640 17340 -17520
rect 17200 -17650 17340 -17640
rect 16510 -18480 16520 -17800
rect 16630 -18480 16640 -17800
rect 16510 -18560 16640 -18480
rect 16500 -18570 16650 -18560
rect 16500 -18730 16510 -18570
rect 16640 -18730 16650 -18570
rect 16500 -18740 16650 -18730
rect 15820 -18870 15960 -18860
rect 15820 -18990 15830 -18870
rect 15950 -18990 15960 -18870
rect 15820 -19000 15960 -18990
rect 15600 -19320 15740 -19310
rect 13310 -19440 15040 -19320
rect 13310 -19610 13440 -19440
rect 13310 -20270 13320 -19610
rect 13430 -20270 13440 -19610
rect 13310 -20280 13440 -20270
rect 14910 -19610 15040 -19440
rect 15600 -19440 15610 -19320
rect 15730 -19440 15740 -19320
rect 15600 -19450 15740 -19440
rect 14910 -20270 14920 -19610
rect 15030 -20270 15040 -19610
rect 14910 -20280 15040 -20270
rect 11030 -20560 11150 -20380
rect 10800 -20860 10940 -20850
rect 10800 -20980 10810 -20860
rect 10930 -20980 10940 -20860
rect 10800 -20990 10940 -20980
rect 10120 -22070 10130 -21410
rect 10230 -22070 10240 -21410
rect 10120 -22190 10240 -22070
rect 10820 -22190 10920 -20990
rect 11040 -22180 11140 -20560
rect 12400 -20680 12540 -20670
rect 12400 -20800 12410 -20680
rect 12530 -20800 12540 -20680
rect 12400 -20810 12540 -20800
rect 11700 -21400 11850 -21390
rect 11700 -22080 11710 -21400
rect 11840 -22080 11850 -21400
rect 11700 -22090 11850 -22080
rect 10120 -22350 10130 -22190
rect 10230 -22350 10240 -22190
rect 10120 -22440 10240 -22350
rect 11030 -22360 11150 -22180
rect 10100 -22450 10260 -22440
rect 10100 -22590 10110 -22450
rect 10250 -22590 10260 -22450
rect 10100 -22600 10260 -22590
rect 11040 -22730 11150 -22360
rect 11720 -22730 11830 -22090
rect 11040 -22740 11160 -22730
rect 11040 -22850 11050 -22740
rect 11150 -22850 11160 -22740
rect 11040 -22860 11160 -22850
rect 11710 -22740 11830 -22730
rect 11710 -22850 11720 -22740
rect 11820 -22850 11830 -22740
rect 11710 -22860 11830 -22850
rect 12420 -22970 12520 -20810
rect 15620 -21110 15720 -19450
rect 15840 -20660 15940 -19000
rect 16510 -19600 16640 -18740
rect 17220 -19310 17320 -17650
rect 17440 -18860 17540 -17200
rect 18110 -17800 18240 -16940
rect 18820 -17510 18920 -15850
rect 19040 -17060 19140 -15400
rect 19710 -16000 19840 -15140
rect 20420 -15710 20520 -14050
rect 20640 -15260 20740 -13600
rect 21310 -14200 21440 -13340
rect 22020 -13910 22120 -12250
rect 22240 -13460 22340 -11800
rect 22910 -12400 23040 -11540
rect 23620 -12110 23720 -10450
rect 23840 -11660 23940 -10000
rect 24510 -10600 24640 -9740
rect 25220 -10310 25320 -8650
rect 25440 -9860 25540 -8200
rect 26820 -8510 26920 -7760
rect 27040 -8060 27140 -6960
rect 27020 -8070 27160 -8060
rect 27020 -8190 27030 -8070
rect 27150 -8190 27160 -8070
rect 27020 -8200 27160 -8190
rect 26800 -8520 26940 -8510
rect 26800 -8640 26810 -8520
rect 26930 -8640 26940 -8520
rect 26800 -8650 26940 -8640
rect 26110 -8800 26240 -8790
rect 26110 -9480 26120 -8800
rect 26230 -9480 26240 -8800
rect 26110 -9560 26240 -9480
rect 26100 -9570 26250 -9560
rect 26100 -9730 26110 -9570
rect 26240 -9730 26250 -9570
rect 26100 -9740 26250 -9730
rect 25420 -9870 25560 -9860
rect 25420 -9990 25430 -9870
rect 25550 -9990 25560 -9870
rect 25420 -10000 25560 -9990
rect 25200 -10320 25340 -10310
rect 25200 -10440 25210 -10320
rect 25330 -10440 25340 -10320
rect 25200 -10450 25340 -10440
rect 24510 -11280 24520 -10600
rect 24630 -11280 24640 -10600
rect 24510 -11360 24640 -11280
rect 24500 -11370 24650 -11360
rect 24500 -11530 24510 -11370
rect 24640 -11530 24650 -11370
rect 24500 -11540 24650 -11530
rect 23820 -11670 23960 -11660
rect 23820 -11790 23830 -11670
rect 23950 -11790 23960 -11670
rect 23820 -11800 23960 -11790
rect 23600 -12120 23740 -12110
rect 23600 -12240 23610 -12120
rect 23730 -12240 23740 -12120
rect 23600 -12250 23740 -12240
rect 22910 -13080 22920 -12400
rect 23030 -13080 23040 -12400
rect 22910 -13160 23040 -13080
rect 22900 -13170 23050 -13160
rect 22900 -13330 22910 -13170
rect 23040 -13330 23050 -13170
rect 22900 -13340 23050 -13330
rect 22220 -13470 22360 -13460
rect 22220 -13590 22230 -13470
rect 22350 -13590 22360 -13470
rect 22220 -13600 22360 -13590
rect 22000 -13920 22140 -13910
rect 22000 -14040 22010 -13920
rect 22130 -14040 22140 -13920
rect 22000 -14050 22140 -14040
rect 21310 -14880 21320 -14200
rect 21430 -14880 21440 -14200
rect 21310 -14960 21440 -14880
rect 21300 -14970 21450 -14960
rect 21300 -15130 21310 -14970
rect 21440 -15130 21450 -14970
rect 21300 -15140 21450 -15130
rect 20620 -15270 20760 -15260
rect 20620 -15390 20630 -15270
rect 20750 -15390 20760 -15270
rect 20620 -15400 20760 -15390
rect 20400 -15720 20540 -15710
rect 20400 -15840 20410 -15720
rect 20530 -15840 20540 -15720
rect 20400 -15850 20540 -15840
rect 19710 -16680 19720 -16000
rect 19830 -16680 19840 -16000
rect 19710 -16760 19840 -16680
rect 19700 -16770 19850 -16760
rect 19700 -16930 19710 -16770
rect 19840 -16930 19850 -16770
rect 19700 -16940 19850 -16930
rect 19020 -17070 19160 -17060
rect 19020 -17190 19030 -17070
rect 19150 -17190 19160 -17070
rect 19020 -17200 19160 -17190
rect 18800 -17520 18940 -17510
rect 18800 -17640 18810 -17520
rect 18930 -17640 18940 -17520
rect 18800 -17650 18940 -17640
rect 18110 -18480 18120 -17800
rect 18230 -18480 18240 -17800
rect 18110 -18560 18240 -18480
rect 18100 -18570 18250 -18560
rect 18100 -18730 18110 -18570
rect 18240 -18730 18250 -18570
rect 18100 -18740 18250 -18730
rect 17420 -18870 17560 -18860
rect 17420 -18990 17430 -18870
rect 17550 -18990 17560 -18870
rect 17420 -19000 17560 -18990
rect 17200 -19320 17340 -19310
rect 17200 -19440 17210 -19320
rect 17330 -19440 17340 -19320
rect 17200 -19450 17340 -19440
rect 16510 -20280 16520 -19600
rect 16630 -20280 16640 -19600
rect 16510 -20360 16640 -20280
rect 16500 -20370 16650 -20360
rect 16500 -20530 16510 -20370
rect 16640 -20530 16650 -20370
rect 16500 -20540 16650 -20530
rect 15820 -20670 15960 -20660
rect 15820 -20790 15830 -20670
rect 15950 -20790 15960 -20670
rect 15820 -20800 15960 -20790
rect 15600 -21120 15740 -21110
rect 15600 -21240 15610 -21120
rect 15730 -21240 15740 -21120
rect 15600 -21250 15740 -21240
rect 15620 -21370 15720 -21250
rect 15840 -21370 15940 -20800
rect 16510 -21400 16640 -20540
rect 17220 -21110 17320 -19450
rect 17440 -20660 17540 -19000
rect 18110 -19600 18240 -18740
rect 18820 -19310 18920 -17650
rect 19040 -18860 19140 -17200
rect 19710 -17800 19840 -16940
rect 20420 -17510 20520 -15850
rect 20640 -17060 20740 -15400
rect 21310 -16000 21440 -15140
rect 22020 -15710 22120 -14050
rect 22240 -15260 22340 -13600
rect 22910 -14200 23040 -13340
rect 23620 -13910 23720 -12250
rect 23840 -13460 23940 -11800
rect 24510 -12400 24640 -11540
rect 25220 -12110 25320 -10450
rect 25440 -11660 25540 -10000
rect 26110 -10600 26240 -9740
rect 26820 -10310 26920 -8650
rect 27040 -9860 27140 -8200
rect 28420 -8510 28520 -5760
rect 28620 -5960 28720 -4850
rect 29300 -5960 29440 -4090
rect 30000 -4240 30100 -2580
rect 30210 -2920 30330 -2910
rect 30210 -3040 30220 -2920
rect 30320 -3040 30330 -2920
rect 30210 -3050 30330 -3040
rect 29990 -4250 30110 -4240
rect 29990 -4370 30000 -4250
rect 30100 -4370 30110 -4250
rect 29990 -4380 30110 -4370
rect 28580 -5970 28760 -5960
rect 28580 -6150 28590 -5970
rect 28750 -6150 28760 -5970
rect 28580 -6160 28760 -6150
rect 29280 -5970 29460 -5960
rect 29280 -6150 29290 -5970
rect 29450 -6150 29460 -5970
rect 29280 -6160 29460 -6150
rect 28640 -8060 28740 -6160
rect 30000 -7160 30100 -4380
rect 30220 -4710 30320 -3050
rect 30900 -3150 31040 -2290
rect 30900 -3330 30910 -3150
rect 31030 -3330 31040 -3150
rect 30900 -3410 31040 -3330
rect 30900 -4090 30910 -3410
rect 31030 -4090 31040 -3410
rect 30210 -4720 30330 -4710
rect 30210 -4840 30220 -4720
rect 30320 -4840 30330 -4720
rect 30210 -4850 30330 -4840
rect 30220 -6760 30320 -4850
rect 30900 -5960 31040 -4090
rect 32500 -1610 32640 -1600
rect 32500 -2290 32510 -1610
rect 32630 -2290 32640 -1610
rect 32500 -2450 32640 -2290
rect 32500 -2570 32510 -2450
rect 32630 -2570 32640 -2450
rect 32500 -3410 32640 -2570
rect 32500 -4090 32510 -3410
rect 32630 -4090 32640 -3410
rect 32500 -4100 32640 -4090
rect 33170 -2450 33310 -2440
rect 33170 -2570 33180 -2450
rect 33300 -2570 33310 -2450
rect 33170 -4250 33310 -2570
rect 33440 -3270 33560 -1600
rect 33390 -3280 33560 -3270
rect 33390 -3400 33400 -3280
rect 33530 -3400 33560 -3280
rect 33390 -3410 33560 -3400
rect 33440 -3660 33560 -3410
rect 34100 -1610 34240 -1600
rect 34100 -2290 34110 -1610
rect 34230 -2290 34240 -1610
rect 34100 -2450 34240 -2290
rect 34790 -2440 34920 1020
rect 35040 -1460 35160 3340
rect 35720 3162 35810 4140
rect 36290 4070 36400 4260
rect 36290 4000 36300 4070
rect 36390 4000 36400 4070
rect 36290 3990 36400 4000
rect 37670 5890 37780 5900
rect 37670 5820 37680 5890
rect 37770 5820 37780 5890
rect 37670 5630 37780 5820
rect 37670 5560 37680 5630
rect 37770 5560 37780 5630
rect 37670 5370 37780 5560
rect 37670 5040 37680 5370
rect 37770 5040 37780 5370
rect 37670 4850 37780 5040
rect 37670 4780 37680 4850
rect 37770 4780 37780 4850
rect 37670 4590 37780 4780
rect 37670 4520 37680 4590
rect 37770 4520 37780 4590
rect 37670 4330 37780 4520
rect 37670 4260 37680 4330
rect 37770 4260 37780 4330
rect 37670 4070 37780 4260
rect 37670 4000 37680 4070
rect 37770 4000 37780 4070
rect 37670 3990 37780 4000
rect 37870 3710 38020 3720
rect 36370 3580 36530 3590
rect 36370 3440 36380 3580
rect 36520 3440 36530 3580
rect 37870 3580 37880 3710
rect 38010 3580 38020 3710
rect 37870 3570 38020 3580
rect 36370 3430 36530 3440
rect 35660 3156 35874 3162
rect 35660 3068 35666 3156
rect 35868 3068 35874 3156
rect 35660 3062 35874 3068
rect 35640 2510 35900 2520
rect 35640 2430 35650 2510
rect 35890 2430 35900 2510
rect 35640 2130 35900 2430
rect 35640 2070 35650 2130
rect 35890 2070 35900 2130
rect 35640 2060 35900 2070
rect 35700 1990 35840 2000
rect 35700 1310 35710 1990
rect 35830 1310 35840 1990
rect 35700 1150 35840 1310
rect 35700 1030 35710 1150
rect 35830 1030 35840 1150
rect 35700 1020 35840 1030
rect 35700 190 35840 200
rect 35700 -490 35710 190
rect 35830 -490 35840 190
rect 35700 -500 35840 -490
rect 35010 -1470 35160 -1460
rect 35010 -1590 35020 -1470
rect 35140 -1570 35160 -1470
rect 35140 -1590 35150 -1570
rect 35010 -1600 35150 -1590
rect 35680 -1600 35760 -1590
rect 35680 -2310 35690 -1600
rect 35750 -2310 35760 -1600
rect 35680 -2350 35760 -2310
rect 35700 -2360 35760 -2350
rect 34100 -2570 34110 -2450
rect 34230 -2570 34240 -2450
rect 34100 -3410 34240 -2570
rect 34780 -2450 34930 -2440
rect 34780 -2570 34790 -2450
rect 34920 -2570 34930 -2450
rect 34780 -2580 34930 -2570
rect 35700 -2450 35840 -2360
rect 35700 -2570 35710 -2450
rect 35830 -2570 35840 -2450
rect 34100 -4090 34110 -3410
rect 34230 -4090 34240 -3410
rect 34100 -4100 34240 -4090
rect 35700 -3410 35840 -2570
rect 36400 -2900 36500 3430
rect 36580 3360 36740 3370
rect 36580 3220 36590 3360
rect 36730 3220 36740 3360
rect 36580 3210 36740 3220
rect 36600 680 36720 3210
rect 37300 1990 37440 2000
rect 37300 1310 37310 1990
rect 37430 1310 37440 1990
rect 37300 1150 37440 1310
rect 37300 1030 37310 1150
rect 37430 1030 37440 1150
rect 37300 1020 37440 1030
rect 36590 670 36730 680
rect 36590 550 36600 670
rect 36720 550 36730 670
rect 37900 660 38020 3570
rect 36590 540 36730 550
rect 37840 650 38020 660
rect 37840 530 37850 650
rect 37970 530 38020 650
rect 37840 520 38020 530
rect 36390 -2910 36510 -2900
rect 36390 -3030 36400 -2910
rect 36500 -3030 36510 -2910
rect 36390 -3040 36510 -3030
rect 35700 -4090 35710 -3410
rect 35830 -4090 35840 -3410
rect 35700 -4100 35840 -4090
rect 33170 -4370 33180 -4250
rect 33300 -4370 33310 -4250
rect 33170 -4380 33310 -4370
rect 36400 -4700 36500 -3040
rect 36390 -4710 36510 -4700
rect 36390 -4830 36400 -4710
rect 36500 -4830 36510 -4710
rect 36390 -4840 36510 -4830
rect 30880 -5970 31060 -5960
rect 30880 -6150 30890 -5970
rect 31050 -6150 31060 -5970
rect 30880 -6160 31060 -6150
rect 30180 -6770 30360 -6760
rect 30180 -6950 30190 -6770
rect 30350 -6950 30360 -6770
rect 30180 -6960 30360 -6950
rect 29960 -7170 30140 -7160
rect 29960 -7350 29970 -7170
rect 30130 -7350 30140 -7170
rect 29960 -7360 30140 -7350
rect 29960 -7570 30140 -7560
rect 29960 -7750 29970 -7570
rect 30130 -7750 30140 -7570
rect 29960 -7760 30140 -7750
rect 28620 -8070 28760 -8060
rect 28620 -8190 28630 -8070
rect 28750 -8190 28760 -8070
rect 28620 -8200 28760 -8190
rect 28400 -8520 28540 -8510
rect 28400 -8640 28410 -8520
rect 28530 -8640 28540 -8520
rect 28400 -8650 28540 -8640
rect 27710 -8800 27840 -8790
rect 27710 -9480 27720 -8800
rect 27830 -9480 27840 -8800
rect 27710 -9560 27840 -9480
rect 27700 -9570 27850 -9560
rect 27700 -9730 27710 -9570
rect 27840 -9730 27850 -9570
rect 27700 -9740 27850 -9730
rect 27020 -9870 27160 -9860
rect 27020 -9990 27030 -9870
rect 27150 -9990 27160 -9870
rect 27020 -10000 27160 -9990
rect 26800 -10320 26940 -10310
rect 26800 -10440 26810 -10320
rect 26930 -10440 26940 -10320
rect 26800 -10450 26940 -10440
rect 26110 -11280 26120 -10600
rect 26230 -11280 26240 -10600
rect 26110 -11360 26240 -11280
rect 26100 -11370 26250 -11360
rect 26100 -11530 26110 -11370
rect 26240 -11530 26250 -11370
rect 26100 -11540 26250 -11530
rect 25420 -11670 25560 -11660
rect 25420 -11790 25430 -11670
rect 25550 -11790 25560 -11670
rect 25420 -11800 25560 -11790
rect 25200 -12120 25340 -12110
rect 25200 -12240 25210 -12120
rect 25330 -12240 25340 -12120
rect 25200 -12250 25340 -12240
rect 24510 -13080 24520 -12400
rect 24630 -13080 24640 -12400
rect 24510 -13160 24640 -13080
rect 24500 -13170 24650 -13160
rect 24500 -13330 24510 -13170
rect 24640 -13330 24650 -13170
rect 24500 -13340 24650 -13330
rect 23820 -13470 23960 -13460
rect 23820 -13590 23830 -13470
rect 23950 -13590 23960 -13470
rect 23820 -13600 23960 -13590
rect 23600 -13920 23740 -13910
rect 23600 -14040 23610 -13920
rect 23730 -14040 23740 -13920
rect 23600 -14050 23740 -14040
rect 22910 -14880 22920 -14200
rect 23030 -14880 23040 -14200
rect 22910 -14960 23040 -14880
rect 22900 -14970 23050 -14960
rect 22900 -15130 22910 -14970
rect 23040 -15130 23050 -14970
rect 22900 -15140 23050 -15130
rect 22220 -15270 22360 -15260
rect 22220 -15390 22230 -15270
rect 22350 -15390 22360 -15270
rect 22220 -15400 22360 -15390
rect 22000 -15720 22140 -15710
rect 22000 -15840 22010 -15720
rect 22130 -15840 22140 -15720
rect 22000 -15850 22140 -15840
rect 21310 -16680 21320 -16000
rect 21430 -16680 21440 -16000
rect 21310 -16760 21440 -16680
rect 21300 -16770 21450 -16760
rect 21300 -16930 21310 -16770
rect 21440 -16930 21450 -16770
rect 21300 -16940 21450 -16930
rect 20620 -17070 20760 -17060
rect 20620 -17190 20630 -17070
rect 20750 -17190 20760 -17070
rect 20620 -17200 20760 -17190
rect 20400 -17520 20540 -17510
rect 20400 -17640 20410 -17520
rect 20530 -17640 20540 -17520
rect 20400 -17650 20540 -17640
rect 19710 -18480 19720 -17800
rect 19830 -18480 19840 -17800
rect 19710 -18560 19840 -18480
rect 19700 -18570 19850 -18560
rect 19700 -18730 19710 -18570
rect 19840 -18730 19850 -18570
rect 19700 -18740 19850 -18730
rect 19020 -18870 19160 -18860
rect 19020 -18990 19030 -18870
rect 19150 -18990 19160 -18870
rect 19020 -19000 19160 -18990
rect 18800 -19320 18940 -19310
rect 18800 -19440 18810 -19320
rect 18930 -19440 18940 -19320
rect 18800 -19450 18940 -19440
rect 18110 -20280 18120 -19600
rect 18230 -20280 18240 -19600
rect 18110 -20360 18240 -20280
rect 18100 -20370 18250 -20360
rect 18100 -20530 18110 -20370
rect 18240 -20530 18250 -20370
rect 18100 -20540 18250 -20530
rect 17420 -20670 17560 -20660
rect 17420 -20790 17430 -20670
rect 17550 -20790 17560 -20670
rect 17420 -20800 17560 -20790
rect 17200 -21120 17340 -21110
rect 17200 -21240 17210 -21120
rect 17330 -21240 17340 -21120
rect 17200 -21250 17340 -21240
rect 17220 -21370 17320 -21250
rect 17440 -21370 17540 -20800
rect 16510 -22080 16520 -21400
rect 16630 -22080 16640 -21400
rect 16510 -22160 16640 -22080
rect 18110 -21400 18240 -20540
rect 18820 -21110 18920 -19450
rect 19040 -20660 19140 -19000
rect 19710 -19600 19840 -18740
rect 20420 -19310 20520 -17650
rect 20640 -18860 20740 -17200
rect 21310 -17800 21440 -16940
rect 22020 -17510 22120 -15850
rect 22240 -17060 22340 -15400
rect 22910 -16000 23040 -15140
rect 23620 -15710 23720 -14050
rect 23840 -15260 23940 -13600
rect 24510 -14200 24640 -13340
rect 25220 -13910 25320 -12250
rect 25440 -13460 25540 -11800
rect 26110 -12400 26240 -11540
rect 26820 -12110 26920 -10450
rect 27040 -11660 27140 -10000
rect 27710 -10600 27840 -9740
rect 28420 -10310 28520 -8650
rect 28640 -9860 28740 -8200
rect 30020 -8510 30120 -7760
rect 30240 -8060 30340 -6960
rect 30220 -8070 30360 -8060
rect 30220 -8190 30230 -8070
rect 30350 -8190 30360 -8070
rect 30220 -8200 30360 -8190
rect 30000 -8520 30140 -8510
rect 30000 -8640 30010 -8520
rect 30130 -8640 30140 -8520
rect 30000 -8650 30140 -8640
rect 29310 -8800 29440 -8790
rect 29310 -9480 29320 -8800
rect 29430 -9480 29440 -8800
rect 29310 -9560 29440 -9480
rect 29300 -9570 29450 -9560
rect 29300 -9730 29310 -9570
rect 29440 -9730 29450 -9570
rect 29300 -9740 29450 -9730
rect 28620 -9870 28760 -9860
rect 28620 -9990 28630 -9870
rect 28750 -9990 28760 -9870
rect 28620 -10000 28760 -9990
rect 28400 -10320 28540 -10310
rect 28400 -10440 28410 -10320
rect 28530 -10440 28540 -10320
rect 28400 -10450 28540 -10440
rect 27710 -11280 27720 -10600
rect 27830 -11280 27840 -10600
rect 27710 -11360 27840 -11280
rect 27700 -11370 27850 -11360
rect 27700 -11530 27710 -11370
rect 27840 -11530 27850 -11370
rect 27700 -11540 27850 -11530
rect 27020 -11670 27160 -11660
rect 27020 -11790 27030 -11670
rect 27150 -11790 27160 -11670
rect 27020 -11800 27160 -11790
rect 26800 -12120 26940 -12110
rect 26800 -12240 26810 -12120
rect 26930 -12240 26940 -12120
rect 26800 -12250 26940 -12240
rect 26110 -13080 26120 -12400
rect 26230 -13080 26240 -12400
rect 26110 -13160 26240 -13080
rect 26100 -13170 26250 -13160
rect 26100 -13330 26110 -13170
rect 26240 -13330 26250 -13170
rect 26100 -13340 26250 -13330
rect 25420 -13470 25560 -13460
rect 25420 -13590 25430 -13470
rect 25550 -13590 25560 -13470
rect 25420 -13600 25560 -13590
rect 25200 -13920 25340 -13910
rect 25200 -14040 25210 -13920
rect 25330 -14040 25340 -13920
rect 25200 -14050 25340 -14040
rect 24510 -14880 24520 -14200
rect 24630 -14880 24640 -14200
rect 24510 -14960 24640 -14880
rect 24500 -14970 24650 -14960
rect 24500 -15130 24510 -14970
rect 24640 -15130 24650 -14970
rect 24500 -15140 24650 -15130
rect 23820 -15270 23960 -15260
rect 23820 -15390 23830 -15270
rect 23950 -15390 23960 -15270
rect 23820 -15400 23960 -15390
rect 23600 -15720 23740 -15710
rect 23600 -15840 23610 -15720
rect 23730 -15840 23740 -15720
rect 23600 -15850 23740 -15840
rect 22910 -16680 22920 -16000
rect 23030 -16680 23040 -16000
rect 22910 -16760 23040 -16680
rect 22900 -16770 23050 -16760
rect 22900 -16930 22910 -16770
rect 23040 -16930 23050 -16770
rect 22900 -16940 23050 -16930
rect 22220 -17070 22360 -17060
rect 22220 -17190 22230 -17070
rect 22350 -17190 22360 -17070
rect 22220 -17200 22360 -17190
rect 22000 -17520 22140 -17510
rect 22000 -17640 22010 -17520
rect 22130 -17640 22140 -17520
rect 22000 -17650 22140 -17640
rect 21310 -18480 21320 -17800
rect 21430 -18480 21440 -17800
rect 21310 -18560 21440 -18480
rect 21300 -18570 21450 -18560
rect 21300 -18730 21310 -18570
rect 21440 -18730 21450 -18570
rect 21300 -18740 21450 -18730
rect 20620 -18870 20760 -18860
rect 20620 -18990 20630 -18870
rect 20750 -18990 20760 -18870
rect 20620 -19000 20760 -18990
rect 20400 -19320 20540 -19310
rect 20400 -19440 20410 -19320
rect 20530 -19440 20540 -19320
rect 20400 -19450 20540 -19440
rect 19710 -20280 19720 -19600
rect 19830 -20280 19840 -19600
rect 19710 -20360 19840 -20280
rect 19700 -20370 19850 -20360
rect 19700 -20530 19710 -20370
rect 19840 -20530 19850 -20370
rect 19700 -20540 19850 -20530
rect 19020 -20670 19160 -20660
rect 19020 -20790 19030 -20670
rect 19150 -20790 19160 -20670
rect 19020 -20800 19160 -20790
rect 18800 -21120 18940 -21110
rect 18800 -21240 18810 -21120
rect 18930 -21240 18940 -21120
rect 18800 -21250 18940 -21240
rect 18820 -21370 18920 -21250
rect 19040 -21370 19140 -20800
rect 18110 -22080 18120 -21400
rect 18230 -22080 18240 -21400
rect 18110 -22160 18240 -22080
rect 19710 -21400 19840 -20540
rect 20420 -21110 20520 -19450
rect 20640 -20660 20740 -19000
rect 21310 -19600 21440 -18740
rect 22020 -19310 22120 -17650
rect 22240 -18860 22340 -17200
rect 22910 -17800 23040 -16940
rect 23620 -17510 23720 -15850
rect 23840 -17060 23940 -15400
rect 24510 -16000 24640 -15140
rect 25220 -15220 25320 -14050
rect 25440 -15220 25540 -13600
rect 26110 -14200 26240 -13340
rect 26820 -13910 26920 -12250
rect 27040 -13460 27140 -11800
rect 27710 -12400 27840 -11540
rect 28420 -12110 28520 -10450
rect 28640 -11660 28740 -10000
rect 29310 -10600 29440 -9740
rect 30020 -10310 30120 -8650
rect 30240 -9860 30340 -8200
rect 30910 -8650 31040 -8030
rect 34820 -8060 34920 -8030
rect 31820 -8070 31960 -8060
rect 31820 -8190 31830 -8070
rect 31950 -8190 31960 -8070
rect 31820 -8200 31960 -8190
rect 34800 -8070 34940 -8060
rect 34800 -8190 34810 -8070
rect 34930 -8190 34940 -8070
rect 34800 -8200 34940 -8190
rect 30910 -8800 31040 -8790
rect 30910 -9480 30920 -8800
rect 31030 -9480 31040 -8800
rect 30910 -9560 31040 -9480
rect 30900 -9570 31050 -9560
rect 30900 -9730 30910 -9570
rect 31040 -9730 31050 -9570
rect 30900 -9740 31050 -9730
rect 30220 -9870 30360 -9860
rect 30220 -9990 30230 -9870
rect 30350 -9990 30360 -9870
rect 30220 -10000 30360 -9990
rect 30000 -10320 30140 -10310
rect 30000 -10440 30010 -10320
rect 30130 -10440 30140 -10320
rect 30000 -10450 30140 -10440
rect 29310 -11280 29320 -10600
rect 29430 -11280 29440 -10600
rect 29310 -11360 29440 -11280
rect 29300 -11370 29450 -11360
rect 29300 -11530 29310 -11370
rect 29440 -11530 29450 -11370
rect 29300 -11540 29450 -11530
rect 28620 -11670 28760 -11660
rect 28620 -11790 28630 -11670
rect 28750 -11790 28760 -11670
rect 28620 -11800 28760 -11790
rect 28400 -12120 28540 -12110
rect 28400 -12240 28410 -12120
rect 28530 -12240 28540 -12120
rect 28400 -12250 28540 -12240
rect 27710 -13080 27720 -12400
rect 27830 -13080 27840 -12400
rect 27710 -13160 27840 -13080
rect 27700 -13170 27850 -13160
rect 27700 -13330 27710 -13170
rect 27840 -13330 27850 -13170
rect 27700 -13340 27850 -13330
rect 27020 -13470 27160 -13460
rect 27020 -13590 27030 -13470
rect 27150 -13590 27160 -13470
rect 27020 -13600 27160 -13590
rect 26800 -13920 26940 -13910
rect 26800 -14040 26810 -13920
rect 26930 -14040 26940 -13920
rect 26800 -14050 26940 -14040
rect 26110 -14880 26120 -14200
rect 26230 -14880 26240 -14200
rect 26110 -14960 26240 -14880
rect 26100 -14970 26250 -14960
rect 26100 -15130 26110 -14970
rect 26240 -15130 26250 -14970
rect 26100 -15140 26250 -15130
rect 24510 -16680 24520 -16000
rect 24630 -16680 24640 -16000
rect 24510 -16760 24640 -16680
rect 26110 -16000 26240 -15140
rect 26820 -15710 26920 -14050
rect 27040 -15260 27140 -13600
rect 27710 -14200 27840 -13340
rect 28420 -13910 28520 -12250
rect 28640 -13460 28740 -11800
rect 29310 -12400 29440 -11540
rect 30020 -12110 30120 -10450
rect 30240 -11660 30340 -10000
rect 30910 -10600 31040 -9740
rect 31840 -9860 31940 -8200
rect 32510 -8800 32640 -8790
rect 32510 -9360 32520 -8800
rect 32630 -9360 32640 -8800
rect 32510 -9560 32640 -9360
rect 34110 -8800 34240 -8790
rect 34110 -9360 34120 -8800
rect 34230 -9360 34240 -8800
rect 33400 -9510 33540 -9500
rect 32500 -9570 32650 -9560
rect 32500 -9730 32510 -9570
rect 32640 -9730 32650 -9570
rect 33400 -9630 33410 -9510
rect 33530 -9630 33540 -9510
rect 34110 -9560 34240 -9360
rect 33400 -9640 33540 -9630
rect 32500 -9740 32650 -9730
rect 31820 -9870 31960 -9860
rect 31820 -9990 31830 -9870
rect 31950 -9990 31960 -9870
rect 31820 -10000 31960 -9990
rect 31600 -10320 31740 -10310
rect 31600 -10440 31610 -10320
rect 31730 -10440 31740 -10320
rect 31600 -10450 31740 -10440
rect 30910 -11280 30920 -10600
rect 31030 -11280 31040 -10600
rect 30910 -11360 31040 -11280
rect 30900 -11370 31050 -11360
rect 30900 -11530 30910 -11370
rect 31040 -11530 31050 -11370
rect 30900 -11540 31050 -11530
rect 30220 -11670 30360 -11660
rect 30220 -11790 30230 -11670
rect 30350 -11790 30360 -11670
rect 30220 -11800 30360 -11790
rect 30000 -12120 30140 -12110
rect 30000 -12240 30010 -12120
rect 30130 -12240 30140 -12120
rect 30000 -12250 30140 -12240
rect 29310 -13080 29320 -12400
rect 29430 -13080 29440 -12400
rect 29310 -13160 29440 -13080
rect 29300 -13170 29450 -13160
rect 29300 -13330 29310 -13170
rect 29440 -13330 29450 -13170
rect 29300 -13340 29450 -13330
rect 28620 -13470 28760 -13460
rect 28620 -13590 28630 -13470
rect 28750 -13590 28760 -13470
rect 28620 -13600 28760 -13590
rect 28400 -13920 28540 -13910
rect 28400 -14040 28410 -13920
rect 28530 -14040 28540 -13920
rect 28400 -14050 28540 -14040
rect 27710 -14880 27720 -14200
rect 27830 -14880 27840 -14200
rect 27710 -14960 27840 -14880
rect 27700 -14970 27850 -14960
rect 27700 -15130 27710 -14970
rect 27840 -15130 27850 -14970
rect 27700 -15140 27850 -15130
rect 27020 -15270 27160 -15260
rect 27020 -15390 27030 -15270
rect 27150 -15390 27160 -15270
rect 27020 -15400 27160 -15390
rect 26800 -15720 26940 -15710
rect 26800 -15840 26810 -15720
rect 26930 -15840 26940 -15720
rect 26800 -15850 26940 -15840
rect 26110 -16680 26120 -16000
rect 26230 -16680 26240 -16000
rect 26110 -16760 26240 -16680
rect 24500 -16770 24650 -16760
rect 24500 -16930 24510 -16770
rect 24640 -16930 24650 -16770
rect 24500 -16940 24650 -16930
rect 26100 -16770 26250 -16760
rect 26100 -16930 26110 -16770
rect 26240 -16930 26250 -16770
rect 26100 -16940 26250 -16930
rect 23820 -17070 23960 -17060
rect 23820 -17190 23830 -17070
rect 23950 -17190 23960 -17070
rect 23820 -17200 23960 -17190
rect 23600 -17520 23740 -17510
rect 23600 -17640 23610 -17520
rect 23730 -17640 23740 -17520
rect 23600 -17650 23740 -17640
rect 22910 -18480 22920 -17800
rect 23030 -18480 23040 -17800
rect 22910 -18560 23040 -18480
rect 22900 -18570 23050 -18560
rect 22900 -18730 22910 -18570
rect 23040 -18730 23050 -18570
rect 22900 -18740 23050 -18730
rect 22220 -18870 22360 -18860
rect 22220 -18990 22230 -18870
rect 22350 -18990 22360 -18870
rect 22220 -19000 22360 -18990
rect 22000 -19320 22140 -19310
rect 22000 -19440 22010 -19320
rect 22130 -19440 22140 -19320
rect 22000 -19450 22140 -19440
rect 21310 -20280 21320 -19600
rect 21430 -20280 21440 -19600
rect 21310 -20360 21440 -20280
rect 21300 -20370 21450 -20360
rect 21300 -20530 21310 -20370
rect 21440 -20530 21450 -20370
rect 21300 -20540 21450 -20530
rect 20620 -20670 20760 -20660
rect 20620 -20790 20630 -20670
rect 20750 -20790 20760 -20670
rect 20620 -20800 20760 -20790
rect 20400 -21120 20540 -21110
rect 20400 -21240 20410 -21120
rect 20530 -21240 20540 -21120
rect 20400 -21250 20540 -21240
rect 20420 -21370 20520 -21250
rect 20640 -21370 20740 -20800
rect 19710 -22080 19720 -21400
rect 19830 -22080 19840 -21400
rect 19710 -22160 19840 -22080
rect 21310 -21400 21440 -20540
rect 22020 -21110 22120 -19450
rect 22240 -20660 22340 -19000
rect 22910 -19600 23040 -18740
rect 23620 -19310 23720 -17650
rect 23840 -18860 23940 -17200
rect 24510 -17800 24640 -16940
rect 24510 -18480 24520 -17800
rect 24630 -18480 24640 -17800
rect 24510 -18560 24640 -18480
rect 26110 -17800 26240 -16940
rect 26820 -17510 26920 -15850
rect 27040 -17060 27140 -15400
rect 27710 -16000 27840 -15140
rect 28420 -15710 28520 -14050
rect 28640 -15260 28740 -13600
rect 29310 -14200 29440 -13340
rect 30020 -13910 30120 -12250
rect 30240 -13460 30340 -11800
rect 30910 -12400 31040 -11540
rect 31620 -12110 31720 -10450
rect 31840 -11660 31940 -10000
rect 32510 -10600 32640 -9740
rect 32510 -11110 32520 -10600
rect 32630 -11110 32640 -10600
rect 32510 -11360 32640 -11110
rect 32500 -11370 32650 -11360
rect 32500 -11530 32510 -11370
rect 32640 -11530 32650 -11370
rect 32500 -11540 32650 -11530
rect 31820 -11670 31960 -11660
rect 31820 -11790 31830 -11670
rect 31950 -11790 31960 -11670
rect 31820 -11800 31960 -11790
rect 31600 -12120 31740 -12110
rect 31600 -12240 31610 -12120
rect 31730 -12240 31740 -12120
rect 31600 -12250 31740 -12240
rect 30910 -13080 30920 -12400
rect 31030 -13080 31040 -12400
rect 30910 -13160 31040 -13080
rect 30900 -13170 31050 -13160
rect 30900 -13330 30910 -13170
rect 31040 -13330 31050 -13170
rect 30900 -13340 31050 -13330
rect 30220 -13470 30360 -13460
rect 30220 -13590 30230 -13470
rect 30350 -13590 30360 -13470
rect 30220 -13600 30360 -13590
rect 30000 -13920 30140 -13910
rect 30000 -14040 30010 -13920
rect 30130 -14040 30140 -13920
rect 30000 -14050 30140 -14040
rect 29310 -14880 29320 -14200
rect 29430 -14880 29440 -14200
rect 29310 -14960 29440 -14880
rect 29300 -14970 29450 -14960
rect 29300 -15130 29310 -14970
rect 29440 -15130 29450 -14970
rect 29300 -15140 29450 -15130
rect 28620 -15270 28760 -15260
rect 28620 -15390 28630 -15270
rect 28750 -15390 28760 -15270
rect 28620 -15400 28760 -15390
rect 28400 -15720 28540 -15710
rect 28400 -15840 28410 -15720
rect 28530 -15840 28540 -15720
rect 28400 -15850 28540 -15840
rect 27710 -16680 27720 -16000
rect 27830 -16680 27840 -16000
rect 27710 -16760 27840 -16680
rect 27700 -16770 27850 -16760
rect 27700 -16930 27710 -16770
rect 27840 -16930 27850 -16770
rect 27700 -16940 27850 -16930
rect 27020 -17070 27160 -17060
rect 27020 -17190 27030 -17070
rect 27150 -17190 27160 -17070
rect 27020 -17200 27160 -17190
rect 26800 -17520 26940 -17510
rect 26800 -17640 26810 -17520
rect 26930 -17640 26940 -17520
rect 26800 -17650 26940 -17640
rect 26110 -18480 26120 -17800
rect 26230 -18480 26240 -17800
rect 26110 -18560 26240 -18480
rect 24500 -18570 24650 -18560
rect 24500 -18730 24510 -18570
rect 24640 -18730 24650 -18570
rect 24500 -18740 24650 -18730
rect 26100 -18570 26250 -18560
rect 26100 -18730 26110 -18570
rect 26240 -18730 26250 -18570
rect 26100 -18740 26250 -18730
rect 23820 -18870 23960 -18860
rect 23820 -18990 23830 -18870
rect 23950 -18990 23960 -18870
rect 23820 -19000 23960 -18990
rect 23600 -19320 23740 -19310
rect 23600 -19440 23610 -19320
rect 23730 -19440 23740 -19320
rect 23600 -19450 23740 -19440
rect 22910 -20280 22920 -19600
rect 23030 -20280 23040 -19600
rect 22910 -20360 23040 -20280
rect 22900 -20370 23050 -20360
rect 22900 -20530 22910 -20370
rect 23040 -20530 23050 -20370
rect 22900 -20540 23050 -20530
rect 22220 -20670 22360 -20660
rect 22220 -20790 22230 -20670
rect 22350 -20790 22360 -20670
rect 22220 -20800 22360 -20790
rect 22000 -21120 22140 -21110
rect 22000 -21240 22010 -21120
rect 22130 -21240 22140 -21120
rect 22000 -21250 22140 -21240
rect 22020 -21370 22120 -21250
rect 22240 -21370 22340 -20800
rect 21310 -22080 21320 -21400
rect 21430 -22080 21440 -21400
rect 21310 -22160 21440 -22080
rect 22910 -21400 23040 -20540
rect 23620 -21110 23720 -19450
rect 23840 -20660 23940 -19000
rect 24510 -19600 24640 -18740
rect 24510 -20280 24520 -19600
rect 24630 -20280 24640 -19600
rect 24510 -20360 24640 -20280
rect 26110 -19600 26240 -18740
rect 26820 -19310 26920 -17650
rect 27040 -18860 27140 -17200
rect 27710 -17800 27840 -16940
rect 28420 -17510 28520 -15850
rect 28640 -17060 28740 -15400
rect 29310 -16000 29440 -15140
rect 29310 -16680 29320 -16000
rect 29430 -16680 29440 -16000
rect 29310 -16760 29440 -16680
rect 29300 -16770 29450 -16760
rect 29300 -16930 29310 -16770
rect 29440 -16930 29450 -16770
rect 29300 -16940 29450 -16930
rect 28620 -17070 28760 -17060
rect 28620 -17190 28630 -17070
rect 28750 -17190 28760 -17070
rect 28620 -17200 28760 -17190
rect 28400 -17520 28540 -17510
rect 28400 -17640 28410 -17520
rect 28530 -17640 28540 -17520
rect 28400 -17650 28540 -17640
rect 27710 -18480 27720 -17800
rect 27830 -18480 27840 -17800
rect 27710 -18560 27840 -18480
rect 27700 -18570 27850 -18560
rect 27700 -18730 27710 -18570
rect 27840 -18730 27850 -18570
rect 27700 -18740 27850 -18730
rect 27020 -18870 27160 -18860
rect 27020 -18990 27030 -18870
rect 27150 -18990 27160 -18870
rect 27020 -19000 27160 -18990
rect 26800 -19320 26940 -19310
rect 26800 -19440 26810 -19320
rect 26930 -19440 26940 -19320
rect 26800 -19450 26940 -19440
rect 26110 -20280 26120 -19600
rect 26230 -20280 26240 -19600
rect 26110 -20360 26240 -20280
rect 24500 -20370 24650 -20360
rect 24500 -20530 24510 -20370
rect 24640 -20530 24650 -20370
rect 24500 -20540 24650 -20530
rect 26100 -20370 26250 -20360
rect 26100 -20530 26110 -20370
rect 26240 -20530 26250 -20370
rect 26100 -20540 26250 -20530
rect 23820 -20670 23960 -20660
rect 23820 -20790 23830 -20670
rect 23950 -20790 23960 -20670
rect 23820 -20800 23960 -20790
rect 23600 -21120 23740 -21110
rect 23600 -21240 23610 -21120
rect 23730 -21240 23740 -21120
rect 23600 -21250 23740 -21240
rect 23620 -21370 23720 -21250
rect 23840 -21370 23940 -20800
rect 22910 -22080 22920 -21400
rect 23030 -22080 23040 -21400
rect 22910 -22160 23040 -22080
rect 24510 -21400 24640 -20540
rect 24510 -22080 24520 -21400
rect 24630 -22080 24640 -21400
rect 24510 -22160 24640 -22080
rect 26110 -21400 26240 -20540
rect 26820 -21110 26920 -19450
rect 27040 -20660 27140 -19000
rect 27710 -19600 27840 -18740
rect 28420 -19310 28520 -17650
rect 28640 -18860 28740 -17200
rect 29310 -17800 29440 -16940
rect 29310 -18480 29320 -17800
rect 29430 -18480 29440 -17800
rect 29310 -18560 29440 -18480
rect 29300 -18570 29450 -18560
rect 29300 -18730 29310 -18570
rect 29440 -18730 29450 -18570
rect 29300 -18740 29450 -18730
rect 28620 -18870 28760 -18860
rect 28620 -18990 28630 -18870
rect 28750 -18990 28760 -18870
rect 28620 -19000 28760 -18990
rect 28400 -19320 28540 -19310
rect 28400 -19440 28410 -19320
rect 28530 -19440 28540 -19320
rect 28400 -19450 28540 -19440
rect 27710 -20280 27720 -19600
rect 27830 -20280 27840 -19600
rect 27710 -20360 27840 -20280
rect 27700 -20370 27850 -20360
rect 27700 -20530 27710 -20370
rect 27840 -20530 27850 -20370
rect 27700 -20540 27850 -20530
rect 27020 -20670 27160 -20660
rect 27020 -20790 27030 -20670
rect 27150 -20790 27160 -20670
rect 27020 -20800 27160 -20790
rect 26800 -21120 26940 -21110
rect 26800 -21240 26810 -21120
rect 26930 -21240 26940 -21120
rect 26800 -21250 26940 -21240
rect 26820 -21370 26920 -21250
rect 27040 -21370 27140 -20800
rect 26110 -22080 26120 -21400
rect 26230 -22080 26240 -21400
rect 26110 -22160 26240 -22080
rect 27710 -21400 27840 -20540
rect 28420 -21110 28520 -19450
rect 28640 -20660 28740 -19000
rect 29310 -19600 29440 -18740
rect 29310 -20280 29320 -19600
rect 29430 -20280 29440 -19600
rect 29310 -20360 29440 -20280
rect 29300 -20370 29450 -20360
rect 29300 -20530 29310 -20370
rect 29440 -20530 29450 -20370
rect 29300 -20540 29450 -20530
rect 28620 -20670 28760 -20660
rect 28620 -20790 28630 -20670
rect 28750 -20790 28760 -20670
rect 28620 -20800 28760 -20790
rect 28400 -21120 28540 -21110
rect 28400 -21240 28410 -21120
rect 28530 -21240 28540 -21120
rect 28400 -21250 28540 -21240
rect 28420 -21370 28520 -21250
rect 28640 -21370 28740 -20800
rect 27710 -22080 27720 -21400
rect 27830 -22080 27840 -21400
rect 27710 -22160 27840 -22080
rect 29310 -21400 29440 -20540
rect 30020 -21370 30120 -14050
rect 30240 -21370 30340 -13600
rect 30910 -14200 31040 -13340
rect 31620 -13910 31720 -12250
rect 31840 -13460 31940 -11800
rect 32510 -12400 32640 -11540
rect 32510 -12910 32520 -12400
rect 32630 -12910 32640 -12400
rect 32510 -13160 32640 -12910
rect 32500 -13170 32650 -13160
rect 32500 -13330 32510 -13170
rect 32640 -13330 32650 -13170
rect 32500 -13340 32650 -13330
rect 31820 -13470 31960 -13460
rect 31820 -13590 31830 -13470
rect 31950 -13590 31960 -13470
rect 31820 -13600 31960 -13590
rect 31600 -13920 31740 -13910
rect 31600 -14040 31610 -13920
rect 31730 -14040 31740 -13920
rect 31600 -14050 31740 -14040
rect 30910 -14880 30920 -14200
rect 31030 -14880 31040 -14200
rect 30910 -14960 31040 -14880
rect 32510 -14200 32640 -13340
rect 32510 -14710 32520 -14200
rect 32630 -14710 32640 -14200
rect 32510 -14890 32640 -14710
rect 30900 -14970 31050 -14960
rect 30900 -15130 30910 -14970
rect 31040 -15130 31050 -14970
rect 30900 -15140 31050 -15130
rect 30910 -16000 31040 -15140
rect 31840 -15280 31980 -15270
rect 31840 -15400 31850 -15280
rect 31970 -15400 31980 -15280
rect 31840 -15410 31980 -15400
rect 31580 -15720 31720 -15710
rect 31580 -15840 31590 -15720
rect 31710 -15840 31720 -15720
rect 31580 -15850 31720 -15840
rect 30910 -16680 30920 -16000
rect 31030 -16680 31040 -16000
rect 30910 -16760 31040 -16680
rect 30900 -16770 31050 -16760
rect 30900 -16930 30910 -16770
rect 31040 -16930 31050 -16770
rect 30900 -16940 31050 -16930
rect 30910 -17800 31040 -16940
rect 31600 -17510 31700 -15850
rect 31860 -17070 31960 -15410
rect 32510 -16000 32640 -15990
rect 32510 -16680 32520 -16000
rect 32630 -16680 32640 -16000
rect 32510 -16770 32640 -16680
rect 32510 -16920 32520 -16770
rect 32630 -16920 32640 -16770
rect 31840 -17080 31980 -17070
rect 31840 -17200 31850 -17080
rect 31970 -17200 31980 -17080
rect 31840 -17210 31980 -17200
rect 31580 -17520 31720 -17510
rect 31580 -17640 31590 -17520
rect 31710 -17640 31720 -17520
rect 31580 -17650 31720 -17640
rect 30910 -18480 30920 -17800
rect 31030 -18480 31040 -17800
rect 30910 -18560 31040 -18480
rect 30900 -18570 31050 -18560
rect 30900 -18730 30910 -18570
rect 31040 -18730 31050 -18570
rect 30900 -18740 31050 -18730
rect 30910 -19600 31040 -18740
rect 31580 -18880 31720 -18870
rect 31580 -19000 31590 -18880
rect 31710 -19000 31720 -18880
rect 31580 -19010 31720 -19000
rect 30910 -20280 30920 -19600
rect 31030 -20280 31040 -19600
rect 30910 -20360 31040 -20280
rect 30900 -20370 31050 -20360
rect 30900 -20530 30910 -20370
rect 31040 -20530 31050 -20370
rect 30900 -20540 31050 -20530
rect 29310 -22080 29320 -21400
rect 29430 -22080 29440 -21400
rect 29310 -22160 29440 -22080
rect 30910 -21400 31040 -20540
rect 31600 -20670 31700 -19010
rect 31740 -19240 31820 -19230
rect 31740 -19520 31750 -19240
rect 31810 -19520 31820 -19240
rect 31740 -19530 31820 -19520
rect 31580 -20680 31720 -20670
rect 31580 -20800 31590 -20680
rect 31710 -20800 31720 -20680
rect 31580 -20810 31720 -20800
rect 30910 -22080 30920 -21400
rect 31030 -22080 31040 -21400
rect 30910 -22160 31040 -22080
rect 16500 -22170 16650 -22160
rect 16500 -22330 16510 -22170
rect 16640 -22330 16650 -22170
rect 16500 -22340 16650 -22330
rect 18100 -22170 18250 -22160
rect 18100 -22330 18110 -22170
rect 18240 -22330 18250 -22170
rect 18100 -22340 18250 -22330
rect 19700 -22170 19850 -22160
rect 19700 -22330 19710 -22170
rect 19840 -22330 19850 -22170
rect 19700 -22340 19850 -22330
rect 21300 -22170 21450 -22160
rect 21300 -22330 21310 -22170
rect 21440 -22330 21450 -22170
rect 21300 -22340 21450 -22330
rect 22900 -22170 23050 -22160
rect 22900 -22330 22910 -22170
rect 23040 -22330 23050 -22170
rect 22900 -22340 23050 -22330
rect 24500 -22170 24650 -22160
rect 24500 -22330 24510 -22170
rect 24640 -22330 24650 -22170
rect 24500 -22340 24650 -22330
rect 26100 -22170 26250 -22160
rect 26100 -22330 26110 -22170
rect 26240 -22330 26250 -22170
rect 26100 -22340 26250 -22330
rect 27700 -22170 27850 -22160
rect 27700 -22330 27710 -22170
rect 27840 -22330 27850 -22170
rect 27700 -22340 27850 -22330
rect 29300 -22170 29450 -22160
rect 29300 -22330 29310 -22170
rect 29440 -22330 29450 -22170
rect 29300 -22340 29450 -22330
rect 30900 -22170 31050 -22160
rect 30900 -22330 30910 -22170
rect 31040 -22330 31050 -22170
rect 30900 -22340 31050 -22330
rect 27710 -22740 27840 -22340
rect 27710 -22850 27720 -22740
rect 27830 -22850 27840 -22740
rect 27710 -22860 27840 -22850
rect 28140 -22730 28380 -22720
rect 28990 -22730 29230 -22720
rect 28140 -22870 28150 -22730
rect 28370 -22870 28380 -22730
rect 28140 -22880 28380 -22870
rect 28620 -22740 28750 -22730
rect 28620 -22870 28630 -22740
rect 28740 -22870 28750 -22740
rect 28620 -22880 28750 -22870
rect 28990 -22870 29000 -22730
rect 29220 -22870 29230 -22730
rect 29310 -22740 29440 -22340
rect 29310 -22850 29320 -22740
rect 29430 -22850 29440 -22740
rect 29310 -22860 29440 -22850
rect 30910 -22740 31040 -22340
rect 30910 -22850 30920 -22740
rect 31030 -22850 31040 -22740
rect 30910 -22860 31040 -22850
rect 28990 -22880 29230 -22870
rect 12410 -22980 12530 -22970
rect 12410 -23090 12420 -22980
rect 12520 -23090 12530 -22980
rect 12410 -23100 12530 -23090
rect 26520 -22980 26720 -22970
rect 26520 -23160 26530 -22980
rect 26710 -23160 26720 -22980
rect 1180 -23270 1360 -23260
rect 1180 -23450 1190 -23270
rect 1350 -23450 1360 -23270
rect 1180 -23460 1360 -23450
rect 2780 -23270 2960 -23260
rect 2780 -23450 2790 -23270
rect 2950 -23450 2960 -23270
rect 2780 -23460 2960 -23450
rect 4380 -23270 4560 -23260
rect 4380 -23450 4390 -23270
rect 4550 -23450 4560 -23270
rect 4380 -23460 4560 -23450
rect 5980 -23270 6160 -23260
rect 5980 -23450 5990 -23270
rect 6150 -23450 6160 -23270
rect 5980 -23460 6160 -23450
rect 7580 -23270 7760 -23260
rect 7580 -23450 7590 -23270
rect 7750 -23450 7760 -23270
rect 7580 -23460 7760 -23450
rect 9180 -23270 9360 -23260
rect 9180 -23450 9190 -23270
rect 9350 -23450 9360 -23270
rect 9180 -23460 9360 -23450
rect 23200 -23300 23400 -23290
rect 23200 -23480 23210 -23300
rect 23390 -23480 23400 -23300
rect 1620 -24070 1820 -24060
rect 1620 -24250 1630 -24070
rect 1810 -24250 1820 -24070
rect 1620 -24260 1820 -24250
rect 1280 -24470 1480 -24460
rect 1280 -24650 1290 -24470
rect 1470 -24650 1480 -24470
rect 1280 -24660 1480 -24650
rect 420 -26630 620 -26620
rect 420 -26710 430 -26630
rect 610 -26710 620 -26630
rect 420 -26720 620 -26710
rect 1420 -26860 1480 -24660
rect 1410 -26870 1490 -26860
rect 1410 -27020 1420 -26870
rect 1480 -27020 1490 -26870
rect 1410 -27030 1490 -27020
rect 420 -27430 620 -27420
rect 420 -27510 430 -27430
rect 610 -27510 620 -27430
rect 420 -27520 620 -27510
rect 420 -28230 620 -28220
rect 420 -28310 430 -28230
rect 610 -28310 620 -28230
rect 420 -28320 620 -28310
rect 420 -29030 620 -29020
rect 420 -29110 430 -29030
rect 610 -29110 620 -29030
rect 420 -29120 620 -29110
rect 1420 -29260 1480 -27030
rect 1620 -27660 1680 -24260
rect 2020 -25160 2080 -23820
rect 2240 -25160 2300 -23820
rect 2500 -25070 4020 -25060
rect 2500 -25130 2510 -25070
rect 4010 -25130 4020 -25070
rect 2500 -25140 4020 -25130
rect 4220 -25160 4280 -23820
rect 4440 -25160 4500 -23820
rect 4700 -25070 6220 -25060
rect 4700 -25130 4710 -25070
rect 6210 -25130 6220 -25070
rect 4700 -25140 6220 -25130
rect 6420 -25160 6480 -23820
rect 6640 -25160 6700 -23820
rect 6900 -25070 8420 -25060
rect 6900 -25130 6910 -25070
rect 8410 -25130 8420 -25070
rect 6900 -25140 8420 -25130
rect 8620 -25160 8680 -23820
rect 8840 -25160 8900 -23820
rect 9100 -25070 10620 -25060
rect 9100 -25130 9110 -25070
rect 10610 -25130 10620 -25070
rect 9100 -25140 10620 -25130
rect 10820 -25160 10880 -23820
rect 11040 -25160 11100 -23820
rect 11300 -25070 12820 -25060
rect 11300 -25130 11310 -25070
rect 12810 -25130 12820 -25070
rect 11300 -25140 12820 -25130
rect 13020 -25160 13080 -23820
rect 13240 -25160 13300 -23820
rect 13500 -25070 15020 -25060
rect 13500 -25130 13510 -25070
rect 15010 -25130 15020 -25070
rect 13500 -25140 15020 -25130
rect 15220 -25160 15280 -23820
rect 15440 -25160 15500 -23820
rect 15700 -25070 17220 -25060
rect 15700 -25130 15710 -25070
rect 17210 -25130 17220 -25070
rect 15700 -25140 17220 -25130
rect 17420 -25160 17480 -23820
rect 17640 -25160 17700 -23820
rect 17900 -25070 19420 -25060
rect 17900 -25130 17910 -25070
rect 19410 -25130 19420 -25070
rect 17900 -25140 19420 -25130
rect 19620 -25160 19680 -23820
rect 19840 -25160 19900 -23820
rect 20440 -24070 20640 -24060
rect 20440 -24250 20450 -24070
rect 20630 -24250 20640 -24070
rect 20440 -24260 20640 -24250
rect 20100 -24470 20300 -24460
rect 20100 -24650 20110 -24470
rect 20290 -24650 20300 -24470
rect 20100 -24660 20300 -24650
rect 2010 -25330 2090 -25160
rect 2230 -25260 2310 -25160
rect 2230 -25320 2240 -25260
rect 2300 -25320 2310 -25260
rect 2230 -25330 2310 -25320
rect 2020 -25960 2080 -25330
rect 2240 -25960 2300 -25330
rect 4210 -25350 4290 -25160
rect 4430 -25170 4510 -25160
rect 4430 -25230 4440 -25170
rect 4500 -25230 4510 -25170
rect 4430 -25280 4510 -25230
rect 4430 -25340 4440 -25280
rect 4500 -25340 4510 -25280
rect 4430 -25350 4510 -25340
rect 6410 -25280 6490 -25160
rect 6410 -25340 6420 -25280
rect 6480 -25340 6490 -25280
rect 6410 -25350 6490 -25340
rect 6630 -25170 6710 -25160
rect 6630 -25230 6640 -25170
rect 6700 -25230 6710 -25170
rect 6630 -25350 6710 -25230
rect 8610 -25170 8690 -25160
rect 8610 -25230 8620 -25170
rect 8680 -25230 8690 -25170
rect 8610 -25280 8690 -25230
rect 8610 -25340 8620 -25280
rect 8680 -25340 8690 -25280
rect 8610 -25350 8690 -25340
rect 8830 -25350 8910 -25160
rect 10810 -25170 10890 -25160
rect 10810 -25230 10820 -25170
rect 10880 -25230 10890 -25170
rect 10810 -25280 10890 -25230
rect 10810 -25340 10820 -25280
rect 10880 -25340 10890 -25280
rect 10810 -25350 10890 -25340
rect 11030 -25350 11110 -25160
rect 13010 -25170 13090 -25160
rect 13010 -25230 13020 -25170
rect 13080 -25230 13090 -25170
rect 13010 -25280 13090 -25230
rect 13010 -25340 13020 -25280
rect 13080 -25340 13090 -25280
rect 13010 -25350 13090 -25340
rect 13230 -25350 13310 -25160
rect 15210 -25170 15290 -25160
rect 15210 -25230 15220 -25170
rect 15280 -25230 15290 -25170
rect 15210 -25350 15290 -25230
rect 15430 -25280 15510 -25160
rect 15430 -25340 15440 -25280
rect 15500 -25340 15510 -25280
rect 15430 -25350 15510 -25340
rect 17410 -25350 17490 -25160
rect 17630 -25170 17710 -25160
rect 17630 -25230 17640 -25170
rect 17700 -25230 17710 -25170
rect 17630 -25280 17710 -25230
rect 17630 -25340 17640 -25280
rect 17700 -25340 17710 -25280
rect 17630 -25350 17710 -25340
rect 19610 -25350 19690 -25160
rect 19830 -25170 19910 -25160
rect 19830 -25230 19840 -25170
rect 19900 -25230 19910 -25170
rect 19830 -25350 19910 -25230
rect 2500 -25630 2700 -25550
rect 3160 -25630 3360 -25550
rect 3820 -25630 4020 -25550
rect 2500 -25700 2700 -25690
rect 2500 -25760 2510 -25700
rect 2690 -25760 2700 -25700
rect 2500 -25770 2700 -25760
rect 3160 -25700 3360 -25690
rect 3160 -25760 3170 -25700
rect 3350 -25760 3360 -25700
rect 3160 -25770 3360 -25760
rect 3820 -25700 4020 -25690
rect 3820 -25760 3830 -25700
rect 4010 -25760 4020 -25700
rect 3820 -25770 4020 -25760
rect 2500 -25870 4020 -25860
rect 2500 -25930 2510 -25870
rect 4010 -25930 4020 -25870
rect 2500 -25940 4020 -25930
rect 4220 -25960 4280 -25350
rect 4440 -25960 4500 -25350
rect 4700 -25630 4900 -25550
rect 5360 -25630 5560 -25550
rect 6020 -25630 6220 -25550
rect 4700 -25700 4900 -25690
rect 4700 -25760 4710 -25700
rect 4890 -25760 4900 -25700
rect 4700 -25770 4900 -25760
rect 5360 -25700 5560 -25690
rect 5360 -25760 5370 -25700
rect 5550 -25760 5560 -25700
rect 5360 -25770 5560 -25760
rect 6020 -25700 6220 -25690
rect 6020 -25760 6030 -25700
rect 6210 -25760 6220 -25700
rect 6020 -25770 6220 -25760
rect 4700 -25870 6220 -25860
rect 4700 -25930 4710 -25870
rect 6210 -25930 6220 -25870
rect 4700 -25940 6220 -25930
rect 6420 -25960 6480 -25350
rect 6640 -25960 6700 -25350
rect 6900 -25560 7100 -25550
rect 6900 -25620 6910 -25560
rect 7090 -25620 7100 -25560
rect 6900 -25630 7100 -25620
rect 7560 -25560 7760 -25550
rect 7560 -25620 7570 -25560
rect 7750 -25620 7760 -25560
rect 7560 -25630 7760 -25620
rect 8220 -25560 8420 -25550
rect 8220 -25620 8230 -25560
rect 8410 -25620 8420 -25560
rect 8220 -25630 8420 -25620
rect 6900 -25770 7100 -25690
rect 7560 -25770 7760 -25690
rect 8220 -25770 8420 -25690
rect 6900 -25870 8420 -25860
rect 6900 -25930 6910 -25870
rect 8410 -25930 8420 -25870
rect 6900 -25940 8420 -25930
rect 8620 -25960 8680 -25350
rect 8840 -25960 8900 -25350
rect 9100 -25560 9300 -25550
rect 9100 -25620 9110 -25560
rect 9290 -25620 9300 -25560
rect 9100 -25630 9300 -25620
rect 9760 -25560 9960 -25550
rect 9760 -25620 9770 -25560
rect 9950 -25620 9960 -25560
rect 9760 -25630 9960 -25620
rect 10420 -25560 10620 -25550
rect 10420 -25620 10430 -25560
rect 10610 -25620 10620 -25560
rect 10420 -25630 10620 -25620
rect 9100 -25770 9300 -25690
rect 9760 -25770 9960 -25690
rect 10420 -25770 10620 -25690
rect 9100 -25870 10620 -25860
rect 9100 -25930 9110 -25870
rect 10610 -25930 10620 -25870
rect 9100 -25940 10620 -25930
rect 10820 -25960 10880 -25350
rect 11040 -25960 11100 -25350
rect 11300 -25560 11500 -25550
rect 11300 -25620 11310 -25560
rect 11490 -25620 11500 -25560
rect 11300 -25630 11500 -25620
rect 11960 -25560 12160 -25550
rect 11960 -25620 11970 -25560
rect 12150 -25620 12160 -25560
rect 11960 -25630 12160 -25620
rect 12620 -25560 12820 -25550
rect 12620 -25620 12630 -25560
rect 12810 -25620 12820 -25560
rect 12620 -25630 12820 -25620
rect 11300 -25770 11500 -25690
rect 11960 -25770 12160 -25690
rect 12620 -25770 12820 -25690
rect 11300 -25870 12820 -25860
rect 11300 -25930 11310 -25870
rect 12810 -25930 12820 -25870
rect 11300 -25940 12820 -25930
rect 13020 -25960 13080 -25350
rect 13240 -25960 13300 -25350
rect 13500 -25560 13700 -25550
rect 13500 -25620 13510 -25560
rect 13690 -25620 13700 -25560
rect 13500 -25630 13700 -25620
rect 14160 -25560 14360 -25550
rect 14160 -25620 14170 -25560
rect 14350 -25620 14360 -25560
rect 14160 -25630 14360 -25620
rect 14820 -25560 15020 -25550
rect 14820 -25620 14830 -25560
rect 15010 -25620 15020 -25560
rect 14820 -25630 15020 -25620
rect 13500 -25770 13700 -25690
rect 14160 -25770 14360 -25690
rect 14820 -25770 15020 -25690
rect 13500 -25870 15020 -25860
rect 13500 -25930 13510 -25870
rect 15010 -25930 15020 -25870
rect 13500 -25940 15020 -25930
rect 15220 -25960 15280 -25350
rect 15440 -25960 15500 -25350
rect 15700 -25630 15900 -25550
rect 16360 -25630 16560 -25550
rect 17020 -25630 17220 -25550
rect 15700 -25700 15900 -25690
rect 15700 -25760 15710 -25700
rect 15890 -25760 15900 -25700
rect 15700 -25770 15900 -25760
rect 16360 -25700 16560 -25690
rect 16360 -25760 16370 -25700
rect 16550 -25760 16560 -25700
rect 16360 -25770 16560 -25760
rect 17020 -25700 17220 -25690
rect 17020 -25760 17030 -25700
rect 17210 -25760 17220 -25700
rect 17020 -25770 17220 -25760
rect 15700 -25870 17220 -25860
rect 15700 -25930 15710 -25870
rect 17210 -25930 17220 -25870
rect 15700 -25940 17220 -25930
rect 17420 -25960 17480 -25350
rect 17640 -25960 17700 -25350
rect 17900 -25630 18100 -25550
rect 18560 -25630 18760 -25550
rect 19220 -25630 19420 -25550
rect 17900 -25700 18100 -25690
rect 17900 -25760 17910 -25700
rect 18090 -25760 18100 -25700
rect 17900 -25770 18100 -25760
rect 18560 -25700 18760 -25690
rect 18560 -25760 18570 -25700
rect 18750 -25760 18760 -25700
rect 18560 -25770 18760 -25760
rect 19220 -25700 19420 -25690
rect 19220 -25760 19230 -25700
rect 19410 -25760 19420 -25700
rect 19220 -25770 19420 -25760
rect 17900 -25870 19420 -25860
rect 17900 -25930 17910 -25870
rect 19410 -25930 19420 -25870
rect 17900 -25940 19420 -25930
rect 19620 -25960 19680 -25350
rect 19840 -25960 19900 -25350
rect 2010 -26060 2090 -25960
rect 2010 -26120 2020 -26060
rect 2080 -26120 2090 -26060
rect 2010 -26130 2090 -26120
rect 2230 -26130 2310 -25960
rect 4210 -25970 4290 -25960
rect 4210 -26030 4220 -25970
rect 4280 -26030 4290 -25970
rect 4210 -26080 4290 -26030
rect 2020 -26760 2080 -26130
rect 2240 -26760 2300 -26130
rect 4210 -26140 4220 -26080
rect 4280 -26140 4290 -26080
rect 4210 -26150 4290 -26140
rect 4430 -26150 4510 -25960
rect 6410 -25970 6490 -25960
rect 6410 -26030 6420 -25970
rect 6480 -26030 6490 -25970
rect 6410 -26150 6490 -26030
rect 6630 -26080 6710 -25960
rect 6630 -26140 6640 -26080
rect 6700 -26140 6710 -26080
rect 6630 -26150 6710 -26140
rect 8610 -26150 8690 -25960
rect 8830 -25970 8910 -25960
rect 8830 -26030 8840 -25970
rect 8900 -26030 8910 -25970
rect 8830 -26080 8910 -26030
rect 8830 -26140 8840 -26080
rect 8900 -26140 8910 -26080
rect 8830 -26150 8910 -26140
rect 10810 -26150 10890 -25960
rect 11030 -25970 11110 -25960
rect 11030 -26030 11040 -25970
rect 11100 -26030 11110 -25970
rect 11030 -26080 11110 -26030
rect 11030 -26140 11040 -26080
rect 11100 -26140 11110 -26080
rect 11030 -26150 11110 -26140
rect 13010 -26150 13090 -25960
rect 13230 -25970 13310 -25960
rect 13230 -26030 13240 -25970
rect 13300 -26030 13310 -25970
rect 13230 -26080 13310 -26030
rect 13230 -26140 13240 -26080
rect 13300 -26140 13310 -26080
rect 13230 -26150 13310 -26140
rect 15210 -26080 15290 -25960
rect 15210 -26140 15220 -26080
rect 15280 -26140 15290 -26080
rect 15210 -26150 15290 -26140
rect 15430 -25970 15510 -25960
rect 15430 -26030 15440 -25970
rect 15500 -26030 15510 -25970
rect 15430 -26150 15510 -26030
rect 17410 -25970 17490 -25960
rect 17410 -26030 17420 -25970
rect 17480 -26030 17490 -25970
rect 17410 -26080 17490 -26030
rect 17410 -26140 17420 -26080
rect 17480 -26140 17490 -26080
rect 17410 -26150 17490 -26140
rect 17630 -26150 17710 -25960
rect 19610 -25970 19690 -25960
rect 19610 -26030 19620 -25970
rect 19680 -26030 19690 -25970
rect 19610 -26150 19690 -26030
rect 19830 -26150 19910 -25960
rect 2500 -26360 2700 -26350
rect 2500 -26420 2510 -26360
rect 2690 -26420 2700 -26360
rect 2500 -26430 2700 -26420
rect 3160 -26360 3360 -26350
rect 3160 -26420 3170 -26360
rect 3350 -26420 3360 -26360
rect 3160 -26430 3360 -26420
rect 3820 -26360 4020 -26350
rect 3820 -26420 3830 -26360
rect 4010 -26420 4020 -26360
rect 3820 -26430 4020 -26420
rect 2500 -26570 2700 -26490
rect 3160 -26570 3360 -26490
rect 3820 -26570 4020 -26490
rect 4220 -26760 4280 -26150
rect 4440 -26760 4500 -26150
rect 4700 -26360 4900 -26350
rect 4700 -26420 4710 -26360
rect 4890 -26420 4900 -26360
rect 4700 -26430 4900 -26420
rect 5360 -26360 5560 -26350
rect 5360 -26420 5370 -26360
rect 5550 -26420 5560 -26360
rect 5360 -26430 5560 -26420
rect 6020 -26360 6220 -26350
rect 6020 -26420 6030 -26360
rect 6210 -26420 6220 -26360
rect 6020 -26430 6220 -26420
rect 4700 -26570 4900 -26490
rect 5360 -26570 5560 -26490
rect 6020 -26570 6220 -26490
rect 4700 -26670 6220 -26660
rect 4700 -26730 4710 -26670
rect 6210 -26730 6220 -26670
rect 4700 -26740 6220 -26730
rect 6420 -26760 6480 -26150
rect 6640 -26760 6700 -26150
rect 6900 -26430 7100 -26350
rect 7560 -26430 7760 -26350
rect 8220 -26430 8420 -26350
rect 6900 -26500 7100 -26490
rect 6900 -26560 6910 -26500
rect 7090 -26560 7100 -26500
rect 6900 -26570 7100 -26560
rect 7560 -26500 7760 -26490
rect 7560 -26560 7570 -26500
rect 7750 -26560 7760 -26500
rect 7560 -26570 7760 -26560
rect 8220 -26500 8420 -26490
rect 8220 -26560 8230 -26500
rect 8410 -26560 8420 -26500
rect 8220 -26570 8420 -26560
rect 6900 -26670 8420 -26660
rect 6900 -26730 6910 -26670
rect 8410 -26730 8420 -26670
rect 6900 -26740 8420 -26730
rect 8620 -26760 8680 -26150
rect 8840 -26760 8900 -26150
rect 9100 -26430 9300 -26350
rect 9760 -26430 9960 -26350
rect 10420 -26430 10620 -26350
rect 9100 -26500 9300 -26490
rect 9100 -26560 9110 -26500
rect 9290 -26560 9300 -26500
rect 9100 -26570 9300 -26560
rect 9760 -26500 9960 -26490
rect 9760 -26560 9770 -26500
rect 9950 -26560 9960 -26500
rect 9760 -26570 9960 -26560
rect 10420 -26500 10620 -26490
rect 10420 -26560 10430 -26500
rect 10610 -26560 10620 -26500
rect 10420 -26570 10620 -26560
rect 9100 -26670 10620 -26660
rect 9100 -26730 9110 -26670
rect 10610 -26730 10620 -26670
rect 9100 -26740 10620 -26730
rect 10820 -26760 10880 -26150
rect 11040 -26760 11100 -26150
rect 11300 -26430 11500 -26350
rect 11960 -26430 12160 -26350
rect 12620 -26430 12820 -26350
rect 11300 -26500 11500 -26490
rect 11300 -26560 11310 -26500
rect 11490 -26560 11500 -26500
rect 11300 -26570 11500 -26560
rect 11960 -26500 12160 -26490
rect 11960 -26560 11970 -26500
rect 12150 -26560 12160 -26500
rect 11960 -26570 12160 -26560
rect 12620 -26500 12820 -26490
rect 12620 -26560 12630 -26500
rect 12810 -26560 12820 -26500
rect 12620 -26570 12820 -26560
rect 11300 -26670 12820 -26660
rect 11300 -26730 11310 -26670
rect 12810 -26730 12820 -26670
rect 11300 -26740 12820 -26730
rect 13020 -26760 13080 -26150
rect 13240 -26760 13300 -26150
rect 13500 -26430 13700 -26350
rect 14160 -26430 14360 -26350
rect 14820 -26430 15020 -26350
rect 13500 -26500 13700 -26490
rect 13500 -26560 13510 -26500
rect 13690 -26560 13700 -26500
rect 13500 -26570 13700 -26560
rect 14160 -26500 14360 -26490
rect 14160 -26560 14170 -26500
rect 14350 -26560 14360 -26500
rect 14160 -26570 14360 -26560
rect 14820 -26500 15020 -26490
rect 14820 -26560 14830 -26500
rect 15010 -26560 15020 -26500
rect 14820 -26570 15020 -26560
rect 13500 -26670 15020 -26660
rect 13500 -26730 13510 -26670
rect 15010 -26730 15020 -26670
rect 13500 -26740 15020 -26730
rect 15220 -26760 15280 -26150
rect 15440 -26760 15500 -26150
rect 15700 -26360 15900 -26350
rect 15700 -26420 15710 -26360
rect 15890 -26420 15900 -26360
rect 15700 -26430 15900 -26420
rect 16360 -26360 16560 -26350
rect 16360 -26420 16370 -26360
rect 16550 -26420 16560 -26360
rect 16360 -26430 16560 -26420
rect 17020 -26360 17220 -26350
rect 17020 -26420 17030 -26360
rect 17210 -26420 17220 -26360
rect 17020 -26430 17220 -26420
rect 15700 -26570 15900 -26490
rect 16360 -26570 16560 -26490
rect 17020 -26570 17220 -26490
rect 15700 -26670 17220 -26660
rect 15700 -26730 15710 -26670
rect 17210 -26730 17220 -26670
rect 15700 -26740 17220 -26730
rect 17420 -26760 17480 -26150
rect 17640 -26760 17700 -26150
rect 17900 -26360 18100 -26350
rect 17900 -26420 17910 -26360
rect 18090 -26420 18100 -26360
rect 17900 -26430 18100 -26420
rect 18560 -26360 18760 -26350
rect 18560 -26420 18570 -26360
rect 18750 -26420 18760 -26360
rect 18560 -26430 18760 -26420
rect 19220 -26360 19420 -26350
rect 19220 -26420 19230 -26360
rect 19410 -26420 19420 -26360
rect 19220 -26430 19420 -26420
rect 17900 -26570 18100 -26490
rect 18560 -26570 18760 -26490
rect 19220 -26570 19420 -26490
rect 19620 -26760 19680 -26150
rect 19840 -26760 19900 -26150
rect 2010 -26930 2090 -26760
rect 2230 -26930 2310 -26760
rect 2020 -27560 2080 -26930
rect 2240 -27560 2300 -26930
rect 4210 -26950 4290 -26760
rect 4430 -26880 4510 -26760
rect 4430 -26940 4440 -26880
rect 4500 -26940 4510 -26880
rect 4430 -26950 4510 -26940
rect 6410 -26880 6490 -26760
rect 6410 -26940 6420 -26880
rect 6480 -26940 6490 -26880
rect 6410 -26950 6490 -26940
rect 6630 -26770 6710 -26760
rect 6630 -26830 6640 -26770
rect 6700 -26830 6710 -26770
rect 6630 -26950 6710 -26830
rect 8610 -26770 8690 -26760
rect 8610 -26830 8620 -26770
rect 8680 -26830 8690 -26770
rect 8610 -26880 8690 -26830
rect 8610 -26940 8620 -26880
rect 8680 -26940 8690 -26880
rect 8610 -26950 8690 -26940
rect 8830 -26950 8910 -26760
rect 10810 -26770 10890 -26760
rect 10810 -26830 10820 -26770
rect 10880 -26830 10890 -26770
rect 10810 -26880 10890 -26830
rect 10810 -26940 10820 -26880
rect 10880 -26940 10890 -26880
rect 10810 -26950 10890 -26940
rect 11030 -26950 11110 -26760
rect 13010 -26770 13090 -26760
rect 13010 -26830 13020 -26770
rect 13080 -26830 13090 -26770
rect 13010 -26880 13090 -26830
rect 13010 -26940 13020 -26880
rect 13080 -26940 13090 -26880
rect 13010 -26950 13090 -26940
rect 13230 -26950 13310 -26760
rect 15210 -26770 15290 -26760
rect 15210 -26830 15220 -26770
rect 15280 -26830 15290 -26770
rect 15210 -26950 15290 -26830
rect 15430 -26880 15510 -26760
rect 15430 -26940 15440 -26880
rect 15500 -26940 15510 -26880
rect 15430 -26950 15510 -26940
rect 17410 -26950 17490 -26760
rect 17630 -26770 17710 -26760
rect 17630 -26830 17640 -26770
rect 17700 -26830 17710 -26770
rect 17630 -26950 17710 -26830
rect 19610 -26950 19690 -26760
rect 19830 -26950 19910 -26760
rect 20240 -26770 20300 -24660
rect 20230 -26780 20310 -26770
rect 20230 -26930 20240 -26780
rect 20300 -26930 20310 -26780
rect 20230 -26940 20310 -26930
rect 2500 -27230 2700 -27150
rect 3160 -27230 3360 -27150
rect 3820 -27230 4020 -27150
rect 2500 -27300 2700 -27290
rect 2500 -27360 2510 -27300
rect 2690 -27360 2700 -27300
rect 2500 -27370 2700 -27360
rect 3160 -27300 3360 -27290
rect 3160 -27360 3170 -27300
rect 3350 -27360 3360 -27300
rect 3160 -27370 3360 -27360
rect 3820 -27300 4020 -27290
rect 3820 -27360 3830 -27300
rect 4010 -27360 4020 -27300
rect 3820 -27370 4020 -27360
rect 4220 -27560 4280 -26950
rect 4440 -27560 4500 -26950
rect 4700 -27230 4900 -27150
rect 5360 -27230 5560 -27150
rect 6020 -27230 6220 -27150
rect 4700 -27300 4900 -27290
rect 4700 -27360 4710 -27300
rect 4890 -27360 4900 -27300
rect 4700 -27370 4900 -27360
rect 5360 -27300 5560 -27290
rect 5360 -27360 5370 -27300
rect 5550 -27360 5560 -27300
rect 5360 -27370 5560 -27360
rect 6020 -27300 6220 -27290
rect 6020 -27360 6030 -27300
rect 6210 -27360 6220 -27300
rect 6020 -27370 6220 -27360
rect 4700 -27470 6220 -27460
rect 4700 -27530 4710 -27470
rect 6210 -27530 6220 -27470
rect 4700 -27540 6220 -27530
rect 6420 -27560 6480 -26950
rect 6640 -27560 6700 -26950
rect 6900 -27160 7100 -27150
rect 6900 -27220 6910 -27160
rect 7090 -27220 7100 -27160
rect 6900 -27230 7100 -27220
rect 7560 -27160 7760 -27150
rect 7560 -27220 7570 -27160
rect 7750 -27220 7760 -27160
rect 7560 -27230 7760 -27220
rect 8220 -27160 8420 -27150
rect 8220 -27220 8230 -27160
rect 8410 -27220 8420 -27160
rect 8220 -27230 8420 -27220
rect 6900 -27370 7100 -27290
rect 7560 -27370 7760 -27290
rect 8220 -27370 8420 -27290
rect 6900 -27470 8420 -27460
rect 6900 -27530 6910 -27470
rect 8410 -27530 8420 -27470
rect 6900 -27540 8420 -27530
rect 8620 -27560 8680 -26950
rect 8840 -27560 8900 -26950
rect 9100 -27160 9300 -27150
rect 9100 -27220 9110 -27160
rect 9290 -27220 9300 -27160
rect 9100 -27230 9300 -27220
rect 9760 -27160 9960 -27150
rect 9760 -27220 9770 -27160
rect 9950 -27220 9960 -27160
rect 9760 -27230 9960 -27220
rect 10420 -27160 10620 -27150
rect 10420 -27220 10430 -27160
rect 10610 -27220 10620 -27160
rect 10420 -27230 10620 -27220
rect 9100 -27370 9300 -27290
rect 9760 -27370 9960 -27290
rect 10420 -27370 10620 -27290
rect 9100 -27470 10620 -27460
rect 9100 -27530 9110 -27470
rect 10610 -27530 10620 -27470
rect 9100 -27540 10620 -27530
rect 10820 -27560 10880 -26950
rect 11040 -27560 11100 -26950
rect 11300 -27160 11500 -27150
rect 11300 -27220 11310 -27160
rect 11490 -27220 11500 -27160
rect 11300 -27230 11500 -27220
rect 11960 -27160 12160 -27150
rect 11960 -27220 11970 -27160
rect 12150 -27220 12160 -27160
rect 11960 -27230 12160 -27220
rect 12620 -27160 12820 -27150
rect 12620 -27220 12630 -27160
rect 12810 -27220 12820 -27160
rect 12620 -27230 12820 -27220
rect 11300 -27370 11500 -27290
rect 11960 -27370 12160 -27290
rect 12620 -27370 12820 -27290
rect 11300 -27470 12820 -27460
rect 11300 -27530 11310 -27470
rect 12810 -27530 12820 -27470
rect 11300 -27540 12820 -27530
rect 13020 -27560 13080 -26950
rect 13240 -27560 13300 -26950
rect 13500 -27160 13700 -27150
rect 13500 -27220 13510 -27160
rect 13690 -27220 13700 -27160
rect 13500 -27230 13700 -27220
rect 14160 -27160 14360 -27150
rect 14160 -27220 14170 -27160
rect 14350 -27220 14360 -27160
rect 14160 -27230 14360 -27220
rect 14820 -27160 15020 -27150
rect 14820 -27220 14830 -27160
rect 15010 -27220 15020 -27160
rect 14820 -27230 15020 -27220
rect 13500 -27370 13700 -27290
rect 14160 -27370 14360 -27290
rect 14820 -27370 15020 -27290
rect 13500 -27470 15020 -27460
rect 13500 -27530 13510 -27470
rect 15010 -27530 15020 -27470
rect 13500 -27540 15020 -27530
rect 15220 -27560 15280 -26950
rect 15440 -27560 15500 -26950
rect 15700 -27230 15900 -27150
rect 16360 -27230 16560 -27150
rect 17020 -27230 17220 -27150
rect 15700 -27300 15900 -27290
rect 15700 -27360 15710 -27300
rect 15890 -27360 15900 -27300
rect 15700 -27370 15900 -27360
rect 16360 -27300 16560 -27290
rect 16360 -27360 16370 -27300
rect 16550 -27360 16560 -27300
rect 16360 -27370 16560 -27360
rect 17020 -27300 17220 -27290
rect 17020 -27360 17030 -27300
rect 17210 -27360 17220 -27300
rect 17020 -27370 17220 -27360
rect 15700 -27470 17220 -27460
rect 15700 -27530 15710 -27470
rect 17210 -27530 17220 -27470
rect 15700 -27540 17220 -27530
rect 17420 -27560 17480 -26950
rect 17640 -27560 17700 -26950
rect 17900 -27230 18100 -27150
rect 18560 -27230 18760 -27150
rect 19220 -27230 19420 -27150
rect 17900 -27300 18100 -27290
rect 17900 -27360 17910 -27300
rect 18090 -27360 18100 -27300
rect 17900 -27370 18100 -27360
rect 18560 -27300 18760 -27290
rect 18560 -27360 18570 -27300
rect 18750 -27360 18760 -27300
rect 18560 -27370 18760 -27360
rect 19220 -27300 19420 -27290
rect 19220 -27360 19230 -27300
rect 19410 -27360 19420 -27300
rect 19220 -27370 19420 -27360
rect 19620 -27560 19680 -26950
rect 19840 -27560 19900 -26950
rect 1610 -27670 1690 -27660
rect 1610 -27820 1620 -27670
rect 1680 -27820 1690 -27670
rect 2010 -27730 2090 -27560
rect 2230 -27730 2310 -27560
rect 4210 -27680 4290 -27560
rect 1610 -27830 1690 -27820
rect 1620 -28460 1680 -27830
rect 2020 -28360 2080 -27730
rect 2240 -28360 2300 -27730
rect 4210 -27740 4220 -27680
rect 4280 -27740 4290 -27680
rect 4210 -27750 4290 -27740
rect 4430 -27750 4510 -27560
rect 6410 -27570 6490 -27560
rect 6410 -27630 6420 -27570
rect 6480 -27630 6490 -27570
rect 6410 -27750 6490 -27630
rect 6630 -27680 6710 -27560
rect 6630 -27740 6640 -27680
rect 6700 -27740 6710 -27680
rect 6630 -27750 6710 -27740
rect 8610 -27750 8690 -27560
rect 8830 -27570 8910 -27560
rect 8830 -27630 8840 -27570
rect 8900 -27630 8910 -27570
rect 8830 -27680 8910 -27630
rect 8830 -27740 8840 -27680
rect 8900 -27740 8910 -27680
rect 8830 -27750 8910 -27740
rect 10810 -27750 10890 -27560
rect 11030 -27570 11110 -27560
rect 11030 -27630 11040 -27570
rect 11100 -27630 11110 -27570
rect 11030 -27680 11110 -27630
rect 11030 -27740 11040 -27680
rect 11100 -27740 11110 -27680
rect 11030 -27750 11110 -27740
rect 13010 -27750 13090 -27560
rect 13230 -27570 13310 -27560
rect 13230 -27630 13240 -27570
rect 13300 -27630 13310 -27570
rect 13230 -27680 13310 -27630
rect 13230 -27740 13240 -27680
rect 13300 -27740 13310 -27680
rect 13230 -27750 13310 -27740
rect 15210 -27680 15290 -27560
rect 15210 -27740 15220 -27680
rect 15280 -27740 15290 -27680
rect 15210 -27750 15290 -27740
rect 15430 -27570 15510 -27560
rect 15430 -27630 15440 -27570
rect 15500 -27630 15510 -27570
rect 15430 -27750 15510 -27630
rect 17410 -27570 17490 -27560
rect 17410 -27630 17420 -27570
rect 17480 -27630 17490 -27570
rect 17410 -27750 17490 -27630
rect 17630 -27750 17710 -27560
rect 19610 -27750 19690 -27560
rect 19830 -27750 19910 -27560
rect 2500 -27960 2700 -27950
rect 2500 -28020 2510 -27960
rect 2690 -28020 2700 -27960
rect 2500 -28030 2700 -28020
rect 3160 -27960 3360 -27950
rect 3160 -28020 3170 -27960
rect 3350 -28020 3360 -27960
rect 3160 -28030 3360 -28020
rect 3820 -27960 4020 -27950
rect 3820 -28020 3830 -27960
rect 4010 -28020 4020 -27960
rect 3820 -28030 4020 -28020
rect 2500 -28170 2700 -28090
rect 3160 -28170 3360 -28090
rect 3820 -28170 4020 -28090
rect 4220 -28360 4280 -27750
rect 4440 -28360 4500 -27750
rect 4700 -27960 4900 -27950
rect 4700 -28020 4710 -27960
rect 4890 -28020 4900 -27960
rect 4700 -28030 4900 -28020
rect 5360 -27960 5560 -27950
rect 5360 -28020 5370 -27960
rect 5550 -28020 5560 -27960
rect 5360 -28030 5560 -28020
rect 6020 -27960 6220 -27950
rect 6020 -28020 6030 -27960
rect 6210 -28020 6220 -27960
rect 6020 -28030 6220 -28020
rect 4700 -28170 4900 -28090
rect 5360 -28170 5560 -28090
rect 6020 -28170 6220 -28090
rect 4700 -28270 6220 -28260
rect 4700 -28330 4710 -28270
rect 6210 -28330 6220 -28270
rect 4700 -28340 6220 -28330
rect 6420 -28360 6480 -27750
rect 6640 -28360 6700 -27750
rect 6900 -28030 7100 -27950
rect 7560 -28030 7760 -27950
rect 8220 -28030 8420 -27950
rect 6900 -28100 7100 -28090
rect 6900 -28160 6910 -28100
rect 7090 -28160 7100 -28100
rect 6900 -28170 7100 -28160
rect 7560 -28100 7760 -28090
rect 7560 -28160 7570 -28100
rect 7750 -28160 7760 -28100
rect 7560 -28170 7760 -28160
rect 8220 -28100 8420 -28090
rect 8220 -28160 8230 -28100
rect 8410 -28160 8420 -28100
rect 8220 -28170 8420 -28160
rect 6900 -28270 8420 -28260
rect 6900 -28330 6910 -28270
rect 8410 -28330 8420 -28270
rect 6900 -28340 8420 -28330
rect 8620 -28360 8680 -27750
rect 8840 -28360 8900 -27750
rect 9100 -28030 9300 -27950
rect 9760 -28030 9960 -27950
rect 10420 -28030 10620 -27950
rect 9100 -28100 9300 -28090
rect 9100 -28160 9110 -28100
rect 9290 -28160 9300 -28100
rect 9100 -28170 9300 -28160
rect 9760 -28100 9960 -28090
rect 9760 -28160 9770 -28100
rect 9950 -28160 9960 -28100
rect 9760 -28170 9960 -28160
rect 10420 -28100 10620 -28090
rect 10420 -28160 10430 -28100
rect 10610 -28160 10620 -28100
rect 10420 -28170 10620 -28160
rect 9100 -28270 10620 -28260
rect 9100 -28330 9110 -28270
rect 10610 -28330 10620 -28270
rect 9100 -28340 10620 -28330
rect 10820 -28360 10880 -27750
rect 11040 -28360 11100 -27750
rect 11300 -28030 11500 -27950
rect 11960 -28030 12160 -27950
rect 12620 -28030 12820 -27950
rect 11300 -28100 11500 -28090
rect 11300 -28160 11310 -28100
rect 11490 -28160 11500 -28100
rect 11300 -28170 11500 -28160
rect 11960 -28100 12160 -28090
rect 11960 -28160 11970 -28100
rect 12150 -28160 12160 -28100
rect 11960 -28170 12160 -28160
rect 12620 -28100 12820 -28090
rect 12620 -28160 12630 -28100
rect 12810 -28160 12820 -28100
rect 12620 -28170 12820 -28160
rect 11300 -28270 12820 -28260
rect 11300 -28330 11310 -28270
rect 12810 -28330 12820 -28270
rect 11300 -28340 12820 -28330
rect 13020 -28360 13080 -27750
rect 13240 -28360 13300 -27750
rect 13500 -28030 13700 -27950
rect 14160 -28030 14360 -27950
rect 14820 -28030 15020 -27950
rect 13500 -28100 13700 -28090
rect 13500 -28160 13510 -28100
rect 13690 -28160 13700 -28100
rect 13500 -28170 13700 -28160
rect 14160 -28100 14360 -28090
rect 14160 -28160 14170 -28100
rect 14350 -28160 14360 -28100
rect 14160 -28170 14360 -28160
rect 14820 -28100 15020 -28090
rect 14820 -28160 14830 -28100
rect 15010 -28160 15020 -28100
rect 14820 -28170 15020 -28160
rect 13500 -28270 15020 -28260
rect 13500 -28330 13510 -28270
rect 15010 -28330 15020 -28270
rect 13500 -28340 15020 -28330
rect 15220 -28360 15280 -27750
rect 15440 -28360 15500 -27750
rect 15700 -27960 15900 -27950
rect 15700 -28020 15710 -27960
rect 15890 -28020 15900 -27960
rect 15700 -28030 15900 -28020
rect 16360 -27960 16560 -27950
rect 16360 -28020 16370 -27960
rect 16550 -28020 16560 -27960
rect 16360 -28030 16560 -28020
rect 17020 -27960 17220 -27950
rect 17020 -28020 17030 -27960
rect 17210 -28020 17220 -27960
rect 17020 -28030 17220 -28020
rect 15700 -28170 15900 -28090
rect 16360 -28170 16560 -28090
rect 17020 -28170 17220 -28090
rect 15700 -28270 17220 -28260
rect 15700 -28330 15710 -28270
rect 17210 -28330 17220 -28270
rect 15700 -28340 17220 -28330
rect 17420 -28360 17480 -27750
rect 17640 -28360 17700 -27750
rect 17900 -27960 18100 -27950
rect 17900 -28020 17910 -27960
rect 18090 -28020 18100 -27960
rect 17900 -28030 18100 -28020
rect 18560 -27960 18760 -27950
rect 18560 -28020 18570 -27960
rect 18750 -28020 18760 -27960
rect 18560 -28030 18760 -28020
rect 19220 -27960 19420 -27950
rect 19220 -28020 19230 -27960
rect 19410 -28020 19420 -27960
rect 19220 -28030 19420 -28020
rect 17900 -28170 18100 -28090
rect 18560 -28170 18760 -28090
rect 19220 -28170 19420 -28090
rect 19620 -28360 19680 -27750
rect 19840 -28360 19900 -27750
rect 1610 -28470 1690 -28460
rect 1610 -28620 1620 -28470
rect 1680 -28620 1690 -28470
rect 2010 -28530 2090 -28360
rect 2230 -28530 2310 -28360
rect 4210 -28480 4290 -28360
rect 1610 -28630 1690 -28620
rect 1410 -29270 1490 -29260
rect 1410 -29420 1420 -29270
rect 1480 -29420 1490 -29270
rect 1410 -29430 1490 -29420
rect 1620 -29430 1680 -28630
rect 2020 -29160 2080 -28530
rect 2240 -29160 2300 -28530
rect 4210 -28540 4220 -28480
rect 4280 -28540 4290 -28480
rect 4210 -28550 4290 -28540
rect 4430 -28550 4510 -28360
rect 6410 -28370 6490 -28360
rect 6410 -28430 6420 -28370
rect 6480 -28430 6490 -28370
rect 6410 -28550 6490 -28430
rect 6630 -28480 6710 -28360
rect 6630 -28540 6640 -28480
rect 6700 -28540 6710 -28480
rect 6630 -28550 6710 -28540
rect 8610 -28550 8690 -28360
rect 8830 -28370 8910 -28360
rect 8830 -28430 8840 -28370
rect 8900 -28430 8910 -28370
rect 8830 -28480 8910 -28430
rect 8830 -28540 8840 -28480
rect 8900 -28540 8910 -28480
rect 8830 -28550 8910 -28540
rect 10810 -28550 10890 -28360
rect 11030 -28370 11110 -28360
rect 11030 -28430 11040 -28370
rect 11100 -28430 11110 -28370
rect 11030 -28480 11110 -28430
rect 11030 -28540 11040 -28480
rect 11100 -28540 11110 -28480
rect 11030 -28550 11110 -28540
rect 13010 -28550 13090 -28360
rect 13230 -28370 13310 -28360
rect 13230 -28430 13240 -28370
rect 13300 -28430 13310 -28370
rect 13230 -28480 13310 -28430
rect 13230 -28540 13240 -28480
rect 13300 -28540 13310 -28480
rect 13230 -28550 13310 -28540
rect 15210 -28480 15290 -28360
rect 15210 -28540 15220 -28480
rect 15280 -28540 15290 -28480
rect 15210 -28550 15290 -28540
rect 15430 -28370 15510 -28360
rect 15430 -28430 15440 -28370
rect 15500 -28430 15510 -28370
rect 15430 -28550 15510 -28430
rect 17410 -28370 17490 -28360
rect 17410 -28430 17420 -28370
rect 17480 -28430 17490 -28370
rect 17410 -28550 17490 -28430
rect 17630 -28550 17710 -28360
rect 19610 -28550 19690 -28360
rect 19830 -28550 19910 -28360
rect 2500 -28760 2700 -28750
rect 2500 -28820 2510 -28760
rect 2690 -28820 2700 -28760
rect 2500 -28830 2700 -28820
rect 3160 -28760 3360 -28750
rect 3160 -28820 3170 -28760
rect 3350 -28820 3360 -28760
rect 3160 -28830 3360 -28820
rect 3820 -28760 4020 -28750
rect 3820 -28820 3830 -28760
rect 4010 -28820 4020 -28760
rect 3820 -28830 4020 -28820
rect 2500 -28970 2700 -28890
rect 3160 -28970 3360 -28890
rect 3820 -28970 4020 -28890
rect 4220 -29160 4280 -28550
rect 4440 -29160 4500 -28550
rect 4700 -28760 4900 -28750
rect 4700 -28820 4710 -28760
rect 4890 -28820 4900 -28760
rect 4700 -28830 4900 -28820
rect 5360 -28760 5560 -28750
rect 5360 -28820 5370 -28760
rect 5550 -28820 5560 -28760
rect 5360 -28830 5560 -28820
rect 6020 -28760 6220 -28750
rect 6020 -28820 6030 -28760
rect 6210 -28820 6220 -28760
rect 6020 -28830 6220 -28820
rect 4700 -28970 4900 -28890
rect 5360 -28970 5560 -28890
rect 6020 -28970 6220 -28890
rect 4700 -29070 6220 -29060
rect 4700 -29130 4710 -29070
rect 6210 -29130 6220 -29070
rect 4700 -29140 6220 -29130
rect 6420 -29160 6480 -28550
rect 6640 -29160 6700 -28550
rect 6900 -28830 7100 -28750
rect 7560 -28830 7760 -28750
rect 8220 -28830 8420 -28750
rect 6900 -28900 7100 -28890
rect 6900 -28960 6910 -28900
rect 7090 -28960 7100 -28900
rect 6900 -28970 7100 -28960
rect 7560 -28900 7760 -28890
rect 7560 -28960 7570 -28900
rect 7750 -28960 7760 -28900
rect 7560 -28970 7760 -28960
rect 8220 -28900 8420 -28890
rect 8220 -28960 8230 -28900
rect 8410 -28960 8420 -28900
rect 8220 -28970 8420 -28960
rect 6900 -29070 8420 -29060
rect 6900 -29130 6910 -29070
rect 8410 -29130 8420 -29070
rect 6900 -29140 8420 -29130
rect 8620 -29160 8680 -28550
rect 8840 -29160 8900 -28550
rect 9100 -28830 9300 -28750
rect 9760 -28830 9960 -28750
rect 10420 -28830 10620 -28750
rect 9100 -28900 9300 -28890
rect 9100 -28960 9110 -28900
rect 9290 -28960 9300 -28900
rect 9100 -28970 9300 -28960
rect 9760 -28900 9960 -28890
rect 9760 -28960 9770 -28900
rect 9950 -28960 9960 -28900
rect 9760 -28970 9960 -28960
rect 10420 -28900 10620 -28890
rect 10420 -28960 10430 -28900
rect 10610 -28960 10620 -28900
rect 10420 -28970 10620 -28960
rect 9100 -29070 10620 -29060
rect 9100 -29130 9110 -29070
rect 10610 -29130 10620 -29070
rect 9100 -29140 10620 -29130
rect 10820 -29160 10880 -28550
rect 11040 -29160 11100 -28550
rect 11300 -28830 11500 -28750
rect 11960 -28830 12160 -28750
rect 12620 -28830 12820 -28750
rect 11300 -28900 11500 -28890
rect 11300 -28960 11310 -28900
rect 11490 -28960 11500 -28900
rect 11300 -28970 11500 -28960
rect 11960 -28900 12160 -28890
rect 11960 -28960 11970 -28900
rect 12150 -28960 12160 -28900
rect 11960 -28970 12160 -28960
rect 12620 -28900 12820 -28890
rect 12620 -28960 12630 -28900
rect 12810 -28960 12820 -28900
rect 12620 -28970 12820 -28960
rect 11300 -29070 12820 -29060
rect 11300 -29130 11310 -29070
rect 12810 -29130 12820 -29070
rect 11300 -29140 12820 -29130
rect 13020 -29160 13080 -28550
rect 13240 -29160 13300 -28550
rect 13500 -28830 13700 -28750
rect 14160 -28830 14360 -28750
rect 14820 -28830 15020 -28750
rect 13500 -28900 13700 -28890
rect 13500 -28960 13510 -28900
rect 13690 -28960 13700 -28900
rect 13500 -28970 13700 -28960
rect 14160 -28900 14360 -28890
rect 14160 -28960 14170 -28900
rect 14350 -28960 14360 -28900
rect 14160 -28970 14360 -28960
rect 14820 -28900 15020 -28890
rect 14820 -28960 14830 -28900
rect 15010 -28960 15020 -28900
rect 14820 -28970 15020 -28960
rect 13500 -29070 15020 -29060
rect 13500 -29130 13510 -29070
rect 15010 -29130 15020 -29070
rect 13500 -29140 15020 -29130
rect 15220 -29160 15280 -28550
rect 15440 -29160 15500 -28550
rect 15700 -28760 15900 -28750
rect 15700 -28820 15710 -28760
rect 15890 -28820 15900 -28760
rect 15700 -28830 15900 -28820
rect 16360 -28760 16560 -28750
rect 16360 -28820 16370 -28760
rect 16550 -28820 16560 -28760
rect 16360 -28830 16560 -28820
rect 17020 -28760 17220 -28750
rect 17020 -28820 17030 -28760
rect 17210 -28820 17220 -28760
rect 17020 -28830 17220 -28820
rect 15700 -28970 15900 -28890
rect 16360 -28970 16560 -28890
rect 17020 -28970 17220 -28890
rect 15700 -29070 17220 -29060
rect 15700 -29130 15710 -29070
rect 17210 -29130 17220 -29070
rect 15700 -29140 17220 -29130
rect 17420 -29160 17480 -28550
rect 17640 -29160 17700 -28550
rect 17900 -28760 18100 -28750
rect 17900 -28820 17910 -28760
rect 18090 -28820 18100 -28760
rect 17900 -28830 18100 -28820
rect 18560 -28760 18760 -28750
rect 18560 -28820 18570 -28760
rect 18750 -28820 18760 -28760
rect 18560 -28830 18760 -28820
rect 19220 -28760 19420 -28750
rect 19220 -28820 19230 -28760
rect 19410 -28820 19420 -28760
rect 19220 -28830 19420 -28820
rect 17900 -28970 18100 -28890
rect 18560 -28970 18760 -28890
rect 19220 -28970 19420 -28890
rect 19620 -29160 19680 -28550
rect 19840 -29160 19900 -28550
rect 2010 -29330 2090 -29160
rect 2230 -29330 2310 -29160
rect 2020 -29960 2080 -29330
rect 2240 -29960 2300 -29330
rect 4210 -29350 4290 -29160
rect 4430 -29280 4510 -29160
rect 4430 -29340 4440 -29280
rect 4500 -29340 4510 -29280
rect 4430 -29350 4510 -29340
rect 6410 -29280 6490 -29160
rect 6410 -29340 6420 -29280
rect 6480 -29340 6490 -29280
rect 6410 -29350 6490 -29340
rect 6630 -29170 6710 -29160
rect 6630 -29230 6640 -29170
rect 6700 -29230 6710 -29170
rect 6630 -29350 6710 -29230
rect 8610 -29170 8690 -29160
rect 8610 -29230 8620 -29170
rect 8680 -29230 8690 -29170
rect 8610 -29280 8690 -29230
rect 8610 -29340 8620 -29280
rect 8680 -29340 8690 -29280
rect 8610 -29350 8690 -29340
rect 8830 -29350 8910 -29160
rect 10810 -29170 10890 -29160
rect 10810 -29230 10820 -29170
rect 10880 -29230 10890 -29170
rect 10810 -29280 10890 -29230
rect 10810 -29340 10820 -29280
rect 10880 -29340 10890 -29280
rect 10810 -29350 10890 -29340
rect 11030 -29350 11110 -29160
rect 13010 -29170 13090 -29160
rect 13010 -29230 13020 -29170
rect 13080 -29230 13090 -29170
rect 13010 -29280 13090 -29230
rect 13010 -29340 13020 -29280
rect 13080 -29340 13090 -29280
rect 13010 -29350 13090 -29340
rect 13230 -29350 13310 -29160
rect 15210 -29170 15290 -29160
rect 15210 -29230 15220 -29170
rect 15280 -29230 15290 -29170
rect 15210 -29350 15290 -29230
rect 15430 -29280 15510 -29160
rect 15430 -29340 15440 -29280
rect 15500 -29340 15510 -29280
rect 15430 -29350 15510 -29340
rect 17410 -29350 17490 -29160
rect 17630 -29170 17710 -29160
rect 17630 -29230 17640 -29170
rect 17700 -29230 17710 -29170
rect 17630 -29350 17710 -29230
rect 19610 -29350 19690 -29160
rect 19830 -29350 19910 -29160
rect 20240 -29170 20300 -26940
rect 20440 -27570 20500 -24260
rect 23200 -24680 23400 -23480
rect 23030 -24690 23570 -24680
rect 23030 -25070 23040 -24690
rect 23560 -25070 23570 -24690
rect 23030 -25080 23570 -25070
rect 26520 -25500 26720 -23160
rect 31600 -23290 31700 -20810
rect 31750 -21030 31810 -19530
rect 31740 -21040 31820 -21030
rect 31740 -21320 31750 -21040
rect 31810 -21320 31820 -21040
rect 31740 -21330 31820 -21320
rect 31550 -23300 31750 -23290
rect 31550 -23480 31560 -23300
rect 31740 -23480 31750 -23300
rect 31550 -23490 31750 -23480
rect 29740 -23520 29890 -23510
rect 29740 -23590 29750 -23520
rect 29880 -23590 29890 -23520
rect 29740 -23600 29890 -23590
rect 28490 -24040 28670 -24030
rect 27620 -24070 27820 -24060
rect 27620 -24250 27630 -24070
rect 27810 -24250 27820 -24070
rect 28490 -24200 28500 -24040
rect 28660 -24050 28670 -24040
rect 28660 -24110 29740 -24050
rect 28660 -24200 28670 -24110
rect 28490 -24210 28670 -24200
rect 27620 -24260 27820 -24250
rect 27390 -24470 27590 -24460
rect 27390 -24650 27400 -24470
rect 27580 -24650 27590 -24470
rect 27390 -24660 27590 -24650
rect 27240 -24890 27440 -24880
rect 27240 -25070 27250 -24890
rect 27430 -25070 27440 -24890
rect 27240 -25080 27440 -25070
rect 26520 -25510 27330 -25500
rect 26520 -25600 27260 -25510
rect 27320 -25600 27330 -25510
rect 26520 -25610 27330 -25600
rect 26520 -25630 27320 -25610
rect 21300 -26630 21500 -26620
rect 21300 -26710 21310 -26630
rect 21490 -26710 21500 -26630
rect 21300 -26720 21500 -26710
rect 21300 -27430 21500 -27420
rect 21300 -27510 21310 -27430
rect 21490 -27510 21500 -27430
rect 21300 -27520 21500 -27510
rect 20430 -27580 20510 -27570
rect 20430 -27730 20440 -27580
rect 20500 -27730 20510 -27580
rect 20430 -27740 20510 -27730
rect 20440 -28370 20500 -27740
rect 21300 -28230 21500 -28220
rect 21300 -28310 21310 -28230
rect 21490 -28310 21500 -28230
rect 21300 -28320 21500 -28310
rect 20430 -28380 20510 -28370
rect 20430 -28530 20440 -28380
rect 20500 -28530 20510 -28380
rect 20430 -28540 20510 -28530
rect 20230 -29180 20310 -29170
rect 20230 -29330 20240 -29180
rect 20300 -29330 20310 -29180
rect 20230 -29340 20310 -29330
rect 20440 -29340 20500 -28540
rect 21300 -29030 21500 -29020
rect 21300 -29110 21310 -29030
rect 21490 -29110 21500 -29030
rect 21300 -29120 21500 -29110
rect 2500 -29630 2700 -29550
rect 3160 -29630 3360 -29550
rect 3820 -29630 4020 -29550
rect 2500 -29700 2700 -29690
rect 2500 -29760 2510 -29700
rect 2690 -29760 2700 -29700
rect 2500 -29770 2700 -29760
rect 3160 -29700 3360 -29690
rect 3160 -29760 3170 -29700
rect 3350 -29760 3360 -29700
rect 3160 -29770 3360 -29760
rect 3820 -29700 4020 -29690
rect 3820 -29760 3830 -29700
rect 4010 -29760 4020 -29700
rect 3820 -29770 4020 -29760
rect 2500 -29870 4020 -29860
rect 2500 -29930 2510 -29870
rect 4010 -29930 4020 -29870
rect 2500 -29940 4020 -29930
rect 4220 -29960 4280 -29350
rect 4440 -29960 4500 -29350
rect 4700 -29630 4900 -29550
rect 5360 -29630 5560 -29550
rect 6020 -29630 6220 -29550
rect 4700 -29700 4900 -29690
rect 4700 -29760 4710 -29700
rect 4890 -29760 4900 -29700
rect 4700 -29770 4900 -29760
rect 5360 -29700 5560 -29690
rect 5360 -29760 5370 -29700
rect 5550 -29760 5560 -29700
rect 5360 -29770 5560 -29760
rect 6020 -29700 6220 -29690
rect 6020 -29760 6030 -29700
rect 6210 -29760 6220 -29700
rect 6020 -29770 6220 -29760
rect 4700 -29870 6220 -29860
rect 4700 -29930 4710 -29870
rect 6210 -29930 6220 -29870
rect 4700 -29940 6220 -29930
rect 6420 -29960 6480 -29350
rect 6640 -29960 6700 -29350
rect 6900 -29560 7100 -29550
rect 6900 -29620 6910 -29560
rect 7090 -29620 7100 -29560
rect 6900 -29630 7100 -29620
rect 7560 -29560 7760 -29550
rect 7560 -29620 7570 -29560
rect 7750 -29620 7760 -29560
rect 7560 -29630 7760 -29620
rect 8220 -29560 8420 -29550
rect 8220 -29620 8230 -29560
rect 8410 -29620 8420 -29560
rect 8220 -29630 8420 -29620
rect 6900 -29770 7100 -29690
rect 7560 -29770 7760 -29690
rect 8220 -29770 8420 -29690
rect 6900 -29870 8420 -29860
rect 6900 -29930 6910 -29870
rect 8410 -29930 8420 -29870
rect 6900 -29940 8420 -29930
rect 8620 -29960 8680 -29350
rect 8840 -29960 8900 -29350
rect 9100 -29560 9300 -29550
rect 9100 -29620 9110 -29560
rect 9290 -29620 9300 -29560
rect 9100 -29630 9300 -29620
rect 9760 -29560 9960 -29550
rect 9760 -29620 9770 -29560
rect 9950 -29620 9960 -29560
rect 9760 -29630 9960 -29620
rect 10420 -29560 10620 -29550
rect 10420 -29620 10430 -29560
rect 10610 -29620 10620 -29560
rect 10420 -29630 10620 -29620
rect 9100 -29770 9300 -29690
rect 9760 -29770 9960 -29690
rect 10420 -29770 10620 -29690
rect 9100 -29870 10620 -29860
rect 9100 -29930 9110 -29870
rect 10610 -29930 10620 -29870
rect 9100 -29940 10620 -29930
rect 10820 -29960 10880 -29350
rect 11040 -29960 11100 -29350
rect 11300 -29560 11500 -29550
rect 11300 -29620 11310 -29560
rect 11490 -29620 11500 -29560
rect 11300 -29630 11500 -29620
rect 11960 -29560 12160 -29550
rect 11960 -29620 11970 -29560
rect 12150 -29620 12160 -29560
rect 11960 -29630 12160 -29620
rect 12620 -29560 12820 -29550
rect 12620 -29620 12630 -29560
rect 12810 -29620 12820 -29560
rect 12620 -29630 12820 -29620
rect 11300 -29770 11500 -29690
rect 11960 -29770 12160 -29690
rect 12620 -29770 12820 -29690
rect 11300 -29870 12820 -29860
rect 11300 -29930 11310 -29870
rect 12810 -29930 12820 -29870
rect 11300 -29940 12820 -29930
rect 13020 -29960 13080 -29350
rect 13240 -29960 13300 -29350
rect 13500 -29560 13700 -29550
rect 13500 -29620 13510 -29560
rect 13690 -29620 13700 -29560
rect 13500 -29630 13700 -29620
rect 14160 -29560 14360 -29550
rect 14160 -29620 14170 -29560
rect 14350 -29620 14360 -29560
rect 14160 -29630 14360 -29620
rect 14820 -29560 15020 -29550
rect 14820 -29620 14830 -29560
rect 15010 -29620 15020 -29560
rect 14820 -29630 15020 -29620
rect 13500 -29770 13700 -29690
rect 14160 -29770 14360 -29690
rect 14820 -29770 15020 -29690
rect 13500 -29870 15020 -29860
rect 13500 -29930 13510 -29870
rect 15010 -29930 15020 -29870
rect 13500 -29940 15020 -29930
rect 15220 -29960 15280 -29350
rect 15440 -29960 15500 -29350
rect 15700 -29630 15900 -29550
rect 16360 -29630 16560 -29550
rect 17020 -29630 17220 -29550
rect 15700 -29700 15900 -29690
rect 15700 -29760 15710 -29700
rect 15890 -29760 15900 -29700
rect 15700 -29770 15900 -29760
rect 16360 -29700 16560 -29690
rect 16360 -29760 16370 -29700
rect 16550 -29760 16560 -29700
rect 16360 -29770 16560 -29760
rect 17020 -29700 17220 -29690
rect 17020 -29760 17030 -29700
rect 17210 -29760 17220 -29700
rect 17020 -29770 17220 -29760
rect 15700 -29870 17220 -29860
rect 15700 -29930 15710 -29870
rect 17210 -29930 17220 -29870
rect 15700 -29940 17220 -29930
rect 17420 -29960 17480 -29350
rect 17640 -29960 17700 -29350
rect 17900 -29630 18100 -29550
rect 18560 -29630 18760 -29550
rect 19220 -29630 19420 -29550
rect 17900 -29700 18100 -29690
rect 17900 -29760 17910 -29700
rect 18090 -29760 18100 -29700
rect 17900 -29770 18100 -29760
rect 18560 -29700 18760 -29690
rect 18560 -29760 18570 -29700
rect 18750 -29760 18760 -29700
rect 18560 -29770 18760 -29760
rect 19220 -29700 19420 -29690
rect 19220 -29760 19230 -29700
rect 19410 -29760 19420 -29700
rect 19220 -29770 19420 -29760
rect 17900 -29870 19420 -29860
rect 17900 -29930 17910 -29870
rect 19410 -29930 19420 -29870
rect 17900 -29940 19420 -29930
rect 19620 -29960 19680 -29350
rect 19840 -29960 19900 -29350
rect 2010 -30060 2090 -29960
rect 2010 -30120 2020 -30060
rect 2080 -30120 2090 -30060
rect 2010 -30130 2090 -30120
rect 2230 -30130 2310 -29960
rect 4210 -29970 4290 -29960
rect 4210 -30030 4220 -29970
rect 4280 -30030 4290 -29970
rect 4210 -30080 4290 -30030
rect 2020 -30760 2080 -30130
rect 2240 -30760 2300 -30130
rect 4210 -30140 4220 -30080
rect 4280 -30140 4290 -30080
rect 4210 -30150 4290 -30140
rect 4430 -30150 4510 -29960
rect 6410 -29970 6490 -29960
rect 6410 -30030 6420 -29970
rect 6480 -30030 6490 -29970
rect 6410 -30150 6490 -30030
rect 6630 -30080 6710 -29960
rect 6630 -30140 6640 -30080
rect 6700 -30140 6710 -30080
rect 6630 -30150 6710 -30140
rect 8610 -30150 8690 -29960
rect 8830 -29970 8910 -29960
rect 8830 -30030 8840 -29970
rect 8900 -30030 8910 -29970
rect 8830 -30080 8910 -30030
rect 8830 -30140 8840 -30080
rect 8900 -30140 8910 -30080
rect 8830 -30150 8910 -30140
rect 10810 -30150 10890 -29960
rect 11030 -29970 11110 -29960
rect 11030 -30030 11040 -29970
rect 11100 -30030 11110 -29970
rect 11030 -30080 11110 -30030
rect 11030 -30140 11040 -30080
rect 11100 -30140 11110 -30080
rect 11030 -30150 11110 -30140
rect 13010 -30150 13090 -29960
rect 13230 -29970 13310 -29960
rect 13230 -30030 13240 -29970
rect 13300 -30030 13310 -29970
rect 13230 -30080 13310 -30030
rect 13230 -30140 13240 -30080
rect 13300 -30140 13310 -30080
rect 13230 -30150 13310 -30140
rect 15210 -30080 15290 -29960
rect 15210 -30140 15220 -30080
rect 15280 -30140 15290 -30080
rect 15210 -30150 15290 -30140
rect 15430 -29970 15510 -29960
rect 15430 -30030 15440 -29970
rect 15500 -30030 15510 -29970
rect 15430 -30150 15510 -30030
rect 17410 -29970 17490 -29960
rect 17410 -30030 17420 -29970
rect 17480 -30030 17490 -29970
rect 17410 -30080 17490 -30030
rect 17410 -30140 17420 -30080
rect 17480 -30140 17490 -30080
rect 17410 -30150 17490 -30140
rect 17630 -30150 17710 -29960
rect 19610 -29970 19690 -29960
rect 19610 -30030 19620 -29970
rect 19680 -30030 19690 -29970
rect 19610 -30150 19690 -30030
rect 19830 -30150 19910 -29960
rect 2500 -30360 2700 -30350
rect 2500 -30420 2510 -30360
rect 2690 -30420 2700 -30360
rect 2500 -30430 2700 -30420
rect 3160 -30360 3360 -30350
rect 3160 -30420 3170 -30360
rect 3350 -30420 3360 -30360
rect 3160 -30430 3360 -30420
rect 3820 -30360 4020 -30350
rect 3820 -30420 3830 -30360
rect 4010 -30420 4020 -30360
rect 3820 -30430 4020 -30420
rect 2500 -30570 2700 -30490
rect 3160 -30570 3360 -30490
rect 3820 -30570 4020 -30490
rect 2500 -30670 4020 -30660
rect 2500 -30730 2510 -30670
rect 4010 -30730 4020 -30670
rect 2500 -30740 4020 -30730
rect 4220 -30760 4280 -30150
rect 4440 -30760 4500 -30150
rect 4700 -30360 4900 -30350
rect 4700 -30420 4710 -30360
rect 4890 -30420 4900 -30360
rect 4700 -30430 4900 -30420
rect 5360 -30360 5560 -30350
rect 5360 -30420 5370 -30360
rect 5550 -30420 5560 -30360
rect 5360 -30430 5560 -30420
rect 6020 -30360 6220 -30350
rect 6020 -30420 6030 -30360
rect 6210 -30420 6220 -30360
rect 6020 -30430 6220 -30420
rect 4700 -30570 4900 -30490
rect 5360 -30570 5560 -30490
rect 6020 -30570 6220 -30490
rect 4700 -30670 6220 -30660
rect 4700 -30730 4710 -30670
rect 6210 -30730 6220 -30670
rect 4700 -30740 6220 -30730
rect 6420 -30760 6480 -30150
rect 6640 -30760 6700 -30150
rect 6900 -30430 7100 -30350
rect 7560 -30430 7760 -30350
rect 8220 -30430 8420 -30350
rect 6900 -30500 7100 -30490
rect 6900 -30560 6910 -30500
rect 7090 -30560 7100 -30500
rect 6900 -30570 7100 -30560
rect 7560 -30500 7760 -30490
rect 7560 -30560 7570 -30500
rect 7750 -30560 7760 -30500
rect 7560 -30570 7760 -30560
rect 8220 -30500 8420 -30490
rect 8220 -30560 8230 -30500
rect 8410 -30560 8420 -30500
rect 8220 -30570 8420 -30560
rect 6900 -30670 8420 -30660
rect 6900 -30730 6910 -30670
rect 8410 -30730 8420 -30670
rect 6900 -30740 8420 -30730
rect 8620 -30760 8680 -30150
rect 8840 -30760 8900 -30150
rect 9100 -30430 9300 -30350
rect 9760 -30430 9960 -30350
rect 10420 -30430 10620 -30350
rect 9100 -30500 9300 -30490
rect 9100 -30560 9110 -30500
rect 9290 -30560 9300 -30500
rect 9100 -30570 9300 -30560
rect 9760 -30500 9960 -30490
rect 9760 -30560 9770 -30500
rect 9950 -30560 9960 -30500
rect 9760 -30570 9960 -30560
rect 10420 -30500 10620 -30490
rect 10420 -30560 10430 -30500
rect 10610 -30560 10620 -30500
rect 10420 -30570 10620 -30560
rect 9100 -30670 10620 -30660
rect 9100 -30730 9110 -30670
rect 10610 -30730 10620 -30670
rect 9100 -30740 10620 -30730
rect 10820 -30760 10880 -30150
rect 11040 -30760 11100 -30150
rect 11300 -30430 11500 -30350
rect 11960 -30430 12160 -30350
rect 12620 -30430 12820 -30350
rect 11300 -30500 11500 -30490
rect 11300 -30560 11310 -30500
rect 11490 -30560 11500 -30500
rect 11300 -30570 11500 -30560
rect 11960 -30500 12160 -30490
rect 11960 -30560 11970 -30500
rect 12150 -30560 12160 -30500
rect 11960 -30570 12160 -30560
rect 12620 -30500 12820 -30490
rect 12620 -30560 12630 -30500
rect 12810 -30560 12820 -30500
rect 12620 -30570 12820 -30560
rect 11300 -30670 12820 -30660
rect 11300 -30730 11310 -30670
rect 12810 -30730 12820 -30670
rect 11300 -30740 12820 -30730
rect 13020 -30760 13080 -30150
rect 13240 -30760 13300 -30150
rect 13500 -30430 13700 -30350
rect 14160 -30430 14360 -30350
rect 14820 -30430 15020 -30350
rect 13500 -30500 13700 -30490
rect 13500 -30560 13510 -30500
rect 13690 -30560 13700 -30500
rect 13500 -30570 13700 -30560
rect 14160 -30500 14360 -30490
rect 14160 -30560 14170 -30500
rect 14350 -30560 14360 -30500
rect 14160 -30570 14360 -30560
rect 14820 -30500 15020 -30490
rect 14820 -30560 14830 -30500
rect 15010 -30560 15020 -30500
rect 14820 -30570 15020 -30560
rect 13500 -30670 15020 -30660
rect 13500 -30730 13510 -30670
rect 15010 -30730 15020 -30670
rect 13500 -30740 15020 -30730
rect 15220 -30760 15280 -30150
rect 15440 -30760 15500 -30150
rect 15700 -30360 15900 -30350
rect 15700 -30420 15710 -30360
rect 15890 -30420 15900 -30360
rect 15700 -30430 15900 -30420
rect 16360 -30360 16560 -30350
rect 16360 -30420 16370 -30360
rect 16550 -30420 16560 -30360
rect 16360 -30430 16560 -30420
rect 17020 -30360 17220 -30350
rect 17020 -30420 17030 -30360
rect 17210 -30420 17220 -30360
rect 17020 -30430 17220 -30420
rect 15700 -30570 15900 -30490
rect 16360 -30570 16560 -30490
rect 17020 -30570 17220 -30490
rect 15700 -30670 17220 -30660
rect 15700 -30730 15710 -30670
rect 17210 -30730 17220 -30670
rect 15700 -30740 17220 -30730
rect 17420 -30760 17480 -30150
rect 17640 -30760 17700 -30150
rect 17900 -30360 18100 -30350
rect 17900 -30420 17910 -30360
rect 18090 -30420 18100 -30360
rect 17900 -30430 18100 -30420
rect 18560 -30360 18760 -30350
rect 18560 -30420 18570 -30360
rect 18750 -30420 18760 -30360
rect 18560 -30430 18760 -30420
rect 19220 -30360 19420 -30350
rect 19220 -30420 19230 -30360
rect 19410 -30420 19420 -30360
rect 19220 -30430 19420 -30420
rect 17900 -30570 18100 -30490
rect 18560 -30570 18760 -30490
rect 19220 -30570 19420 -30490
rect 17900 -30670 19420 -30660
rect 17900 -30730 17910 -30670
rect 19410 -30730 19420 -30670
rect 17900 -30740 19420 -30730
rect 19620 -30760 19680 -30150
rect 19840 -30760 19900 -30150
rect 2010 -30930 2090 -30760
rect 2230 -30860 2310 -30760
rect 2230 -30920 2240 -30860
rect 2300 -30920 2310 -30860
rect 2230 -30930 2310 -30920
rect 2020 -31700 2080 -30930
rect 80 -32110 90 -31730
rect 270 -32110 280 -31730
rect 1980 -31710 2120 -31700
rect 1980 -31830 1990 -31710
rect 2110 -31830 2120 -31710
rect 1980 -31840 2120 -31830
rect 80 -32120 280 -32110
rect 2020 -32140 2080 -31840
rect 2240 -32000 2300 -30930
rect 4210 -30950 4290 -30760
rect 4430 -30770 4510 -30760
rect 4430 -30830 4440 -30770
rect 4500 -30830 4510 -30770
rect 4430 -30880 4510 -30830
rect 4430 -30940 4440 -30880
rect 4500 -30940 4510 -30880
rect 4430 -30950 4510 -30940
rect 6410 -30880 6490 -30760
rect 6410 -30940 6420 -30880
rect 6480 -30940 6490 -30880
rect 6410 -30950 6490 -30940
rect 6630 -30770 6710 -30760
rect 6630 -30830 6640 -30770
rect 6700 -30830 6710 -30770
rect 6630 -30950 6710 -30830
rect 8610 -30770 8690 -30760
rect 8610 -30830 8620 -30770
rect 8680 -30830 8690 -30770
rect 8610 -30880 8690 -30830
rect 8610 -30940 8620 -30880
rect 8680 -30940 8690 -30880
rect 8610 -30950 8690 -30940
rect 8830 -30950 8910 -30760
rect 10810 -30770 10890 -30760
rect 10810 -30830 10820 -30770
rect 10880 -30830 10890 -30770
rect 10810 -30880 10890 -30830
rect 10810 -30940 10820 -30880
rect 10880 -30940 10890 -30880
rect 10810 -30950 10890 -30940
rect 11030 -30950 11110 -30760
rect 13010 -30770 13090 -30760
rect 13010 -30830 13020 -30770
rect 13080 -30830 13090 -30770
rect 13010 -30880 13090 -30830
rect 13010 -30940 13020 -30880
rect 13080 -30940 13090 -30880
rect 13010 -30950 13090 -30940
rect 13230 -30950 13310 -30760
rect 15210 -30770 15290 -30760
rect 15210 -30830 15220 -30770
rect 15280 -30830 15290 -30770
rect 15210 -30950 15290 -30830
rect 15430 -30880 15510 -30760
rect 15430 -30940 15440 -30880
rect 15500 -30940 15510 -30880
rect 15430 -30950 15510 -30940
rect 17410 -30950 17490 -30760
rect 17630 -30770 17710 -30760
rect 17630 -30830 17640 -30770
rect 17700 -30830 17710 -30770
rect 17630 -30880 17710 -30830
rect 17630 -30940 17640 -30880
rect 17700 -30940 17710 -30880
rect 17630 -30950 17710 -30940
rect 19610 -30950 19690 -30760
rect 19830 -30770 19910 -30760
rect 19830 -30830 19840 -30770
rect 19900 -30830 19910 -30770
rect 19830 -30950 19910 -30830
rect 2500 -31230 2700 -31150
rect 3160 -31230 3360 -31150
rect 3820 -31230 4020 -31150
rect 2500 -31300 2700 -31290
rect 2500 -31360 2510 -31300
rect 2690 -31360 2700 -31300
rect 2500 -31370 2700 -31360
rect 3160 -31300 3360 -31290
rect 3160 -31360 3170 -31300
rect 3350 -31360 3360 -31300
rect 3160 -31370 3360 -31360
rect 3820 -31300 4020 -31290
rect 3820 -31360 3830 -31300
rect 4010 -31360 4020 -31300
rect 3820 -31370 4020 -31360
rect 4220 -31700 4280 -30950
rect 4180 -31710 4320 -31700
rect 4180 -31830 4190 -31710
rect 4310 -31830 4320 -31710
rect 4180 -31840 4320 -31830
rect 2200 -32010 2340 -32000
rect 2200 -32130 2210 -32010
rect 2330 -32130 2340 -32010
rect 2200 -32140 2340 -32130
rect 4220 -32140 4280 -31840
rect 4440 -32000 4500 -30950
rect 4700 -31230 4900 -31150
rect 5360 -31230 5560 -31150
rect 6020 -31230 6220 -31150
rect 4700 -31300 4900 -31290
rect 4700 -31360 4710 -31300
rect 4890 -31360 4900 -31300
rect 4700 -31370 4900 -31360
rect 5360 -31300 5560 -31290
rect 5360 -31360 5370 -31300
rect 5550 -31360 5560 -31300
rect 5360 -31370 5560 -31360
rect 6020 -31300 6220 -31290
rect 6020 -31360 6030 -31300
rect 6210 -31360 6220 -31300
rect 6020 -31370 6220 -31360
rect 6420 -31700 6480 -30950
rect 6380 -31710 6520 -31700
rect 6380 -31830 6390 -31710
rect 6510 -31830 6520 -31710
rect 6380 -31840 6520 -31830
rect 4400 -32010 4540 -32000
rect 4400 -32130 4410 -32010
rect 4530 -32130 4540 -32010
rect 4400 -32140 4540 -32130
rect 6420 -32140 6480 -31840
rect 6640 -32000 6700 -30950
rect 6900 -31160 7100 -31150
rect 6900 -31220 6910 -31160
rect 7090 -31220 7100 -31160
rect 6900 -31230 7100 -31220
rect 7560 -31160 7760 -31150
rect 7560 -31220 7570 -31160
rect 7750 -31220 7760 -31160
rect 7560 -31230 7760 -31220
rect 8220 -31160 8420 -31150
rect 8220 -31220 8230 -31160
rect 8410 -31220 8420 -31160
rect 8220 -31230 8420 -31220
rect 6900 -31370 7100 -31290
rect 7560 -31370 7760 -31290
rect 8220 -31370 8420 -31290
rect 8620 -31700 8680 -30950
rect 8580 -31710 8720 -31700
rect 8580 -31830 8590 -31710
rect 8710 -31830 8720 -31710
rect 8580 -31840 8720 -31830
rect 6600 -32010 6740 -32000
rect 6600 -32130 6610 -32010
rect 6730 -32130 6740 -32010
rect 6600 -32140 6740 -32130
rect 8620 -32140 8680 -31840
rect 8840 -32000 8900 -30950
rect 9100 -31160 9300 -31150
rect 9100 -31220 9110 -31160
rect 9290 -31220 9300 -31160
rect 9100 -31230 9300 -31220
rect 9760 -31160 9960 -31150
rect 9760 -31220 9770 -31160
rect 9950 -31220 9960 -31160
rect 9760 -31230 9960 -31220
rect 10420 -31160 10620 -31150
rect 10420 -31220 10430 -31160
rect 10610 -31220 10620 -31160
rect 10420 -31230 10620 -31220
rect 9100 -31370 9300 -31290
rect 9760 -31370 9960 -31290
rect 10420 -31370 10620 -31290
rect 10820 -31700 10880 -30950
rect 10780 -31710 10920 -31700
rect 10780 -31830 10790 -31710
rect 10910 -31830 10920 -31710
rect 10780 -31840 10920 -31830
rect 8800 -32010 8940 -32000
rect 8800 -32130 8810 -32010
rect 8930 -32130 8940 -32010
rect 8800 -32140 8940 -32130
rect 10820 -32140 10880 -31840
rect 11040 -32000 11100 -30950
rect 11300 -31160 11500 -31150
rect 11300 -31220 11310 -31160
rect 11490 -31220 11500 -31160
rect 11300 -31230 11500 -31220
rect 11960 -31160 12160 -31150
rect 11960 -31220 11970 -31160
rect 12150 -31220 12160 -31160
rect 11960 -31230 12160 -31220
rect 12620 -31160 12820 -31150
rect 12620 -31220 12630 -31160
rect 12810 -31220 12820 -31160
rect 12620 -31230 12820 -31220
rect 11300 -31370 11500 -31290
rect 11960 -31370 12160 -31290
rect 12620 -31370 12820 -31290
rect 13020 -31700 13080 -30950
rect 12980 -31710 13120 -31700
rect 12980 -31830 12990 -31710
rect 13110 -31830 13120 -31710
rect 12980 -31840 13120 -31830
rect 11000 -32010 11140 -32000
rect 11000 -32130 11010 -32010
rect 11130 -32130 11140 -32010
rect 11000 -32140 11140 -32130
rect 13020 -32140 13080 -31840
rect 13240 -32000 13300 -30950
rect 13500 -31160 13700 -31150
rect 13500 -31220 13510 -31160
rect 13690 -31220 13700 -31160
rect 13500 -31230 13700 -31220
rect 14160 -31160 14360 -31150
rect 14160 -31220 14170 -31160
rect 14350 -31220 14360 -31160
rect 14160 -31230 14360 -31220
rect 14820 -31160 15020 -31150
rect 14820 -31220 14830 -31160
rect 15010 -31220 15020 -31160
rect 14820 -31230 15020 -31220
rect 13500 -31370 13700 -31290
rect 14160 -31370 14360 -31290
rect 14820 -31370 15020 -31290
rect 15220 -31700 15280 -30950
rect 15180 -31710 15320 -31700
rect 15180 -31830 15190 -31710
rect 15310 -31830 15320 -31710
rect 15180 -31840 15320 -31830
rect 13200 -32010 13340 -32000
rect 13200 -32130 13210 -32010
rect 13330 -32130 13340 -32010
rect 13200 -32140 13340 -32130
rect 15220 -32140 15280 -31840
rect 15440 -32000 15500 -30950
rect 15700 -31230 15900 -31150
rect 16360 -31230 16560 -31150
rect 17020 -31230 17220 -31150
rect 15700 -31300 15900 -31290
rect 15700 -31360 15710 -31300
rect 15890 -31360 15900 -31300
rect 15700 -31370 15900 -31360
rect 16360 -31300 16560 -31290
rect 16360 -31360 16370 -31300
rect 16550 -31360 16560 -31300
rect 16360 -31370 16560 -31360
rect 17020 -31300 17220 -31290
rect 17020 -31360 17030 -31300
rect 17210 -31360 17220 -31300
rect 17020 -31370 17220 -31360
rect 17420 -31700 17480 -30950
rect 17380 -31710 17520 -31700
rect 17380 -31830 17390 -31710
rect 17510 -31830 17520 -31710
rect 17380 -31840 17520 -31830
rect 15400 -32010 15540 -32000
rect 15400 -32130 15410 -32010
rect 15530 -32130 15540 -32010
rect 15400 -32140 15540 -32130
rect 17420 -32140 17480 -31840
rect 17640 -32000 17700 -30950
rect 17900 -31230 18100 -31150
rect 18560 -31230 18760 -31150
rect 19220 -31230 19420 -31150
rect 17900 -31300 18100 -31290
rect 17900 -31360 17910 -31300
rect 18090 -31360 18100 -31300
rect 17900 -31370 18100 -31360
rect 18560 -31300 18760 -31290
rect 18560 -31360 18570 -31300
rect 18750 -31360 18760 -31300
rect 18560 -31370 18760 -31360
rect 19220 -31300 19420 -31290
rect 19220 -31360 19230 -31300
rect 19410 -31360 19420 -31300
rect 19220 -31370 19420 -31360
rect 19620 -31700 19680 -30950
rect 19580 -31710 19720 -31700
rect 19580 -31830 19590 -31710
rect 19710 -31830 19720 -31710
rect 19580 -31840 19720 -31830
rect 17600 -32010 17740 -32000
rect 17600 -32130 17610 -32010
rect 17730 -32130 17740 -32010
rect 17600 -32140 17740 -32130
rect 19620 -32140 19680 -31840
rect 19840 -32000 19900 -30950
rect 25690 -31510 26230 -31500
rect 25690 -31880 25700 -31510
rect 26220 -31600 26230 -31510
rect 26520 -31600 26720 -25630
rect 27260 -25820 27320 -25630
rect 27250 -25830 27330 -25820
rect 27250 -25920 27260 -25830
rect 27320 -25920 27330 -25830
rect 27250 -25930 27330 -25920
rect 27260 -26135 27320 -25930
rect 27250 -26145 27330 -26135
rect 27250 -26235 27260 -26145
rect 27320 -26235 27330 -26145
rect 27250 -26245 27330 -26235
rect 27260 -27585 27320 -26245
rect 27380 -26700 27440 -25080
rect 27370 -26710 27450 -26700
rect 27370 -26800 27380 -26710
rect 27440 -26800 27450 -26710
rect 27370 -26810 27450 -26800
rect 27380 -27015 27440 -26810
rect 27370 -27025 27450 -27015
rect 27370 -27115 27380 -27025
rect 27440 -27115 27450 -27025
rect 27370 -27125 27450 -27115
rect 27250 -27595 27330 -27585
rect 27250 -27685 27260 -27595
rect 27320 -27685 27330 -27595
rect 27250 -27695 27330 -27685
rect 27260 -27900 27320 -27695
rect 27250 -27910 27330 -27900
rect 27250 -28000 27260 -27910
rect 27320 -28000 27330 -27910
rect 27250 -28010 27330 -28000
rect 27260 -28215 27320 -28010
rect 27250 -28225 27330 -28215
rect 27250 -28315 27260 -28225
rect 27320 -28315 27330 -28225
rect 27250 -28325 27330 -28315
rect 27260 -28620 27320 -28325
rect 27250 -28630 27330 -28620
rect 27250 -28720 27260 -28630
rect 27320 -28720 27330 -28630
rect 27250 -28730 27330 -28720
rect 27260 -28940 27320 -28730
rect 27250 -28950 27330 -28940
rect 27250 -29040 27260 -28950
rect 27320 -29040 27330 -28950
rect 27250 -29050 27330 -29040
rect 27260 -29250 27320 -29050
rect 27250 -29260 27330 -29250
rect 27250 -29350 27260 -29260
rect 27320 -29350 27330 -29260
rect 27250 -29360 27330 -29350
rect 27260 -31600 27320 -29360
rect 27380 -29660 27440 -27125
rect 27500 -27740 27560 -24660
rect 27490 -27750 27570 -27740
rect 27490 -27840 27500 -27750
rect 27560 -27840 27570 -27750
rect 27490 -27850 27570 -27840
rect 27500 -28055 27560 -27850
rect 27490 -28065 27570 -28055
rect 27490 -28155 27500 -28065
rect 27560 -28155 27570 -28065
rect 27490 -28165 27570 -28155
rect 27370 -29670 27450 -29660
rect 27370 -29760 27380 -29670
rect 27440 -29760 27450 -29670
rect 27370 -29770 27450 -29760
rect 27380 -29975 27440 -29770
rect 27370 -29985 27450 -29975
rect 27370 -30075 27380 -29985
rect 27440 -30075 27450 -29985
rect 27370 -30085 27450 -30075
rect 27380 -30290 27440 -30085
rect 27370 -30300 27450 -30290
rect 27370 -30390 27380 -30300
rect 27440 -30390 27450 -30300
rect 27370 -30400 27450 -30390
rect 27380 -30700 27440 -30400
rect 27370 -30710 27450 -30700
rect 27370 -30800 27380 -30710
rect 27440 -30800 27450 -30710
rect 27370 -30810 27450 -30800
rect 27380 -31015 27440 -30810
rect 27500 -30860 27560 -28165
rect 27620 -28780 27680 -24260
rect 29370 -24490 29450 -24480
rect 29370 -24720 29380 -24490
rect 29440 -24720 29450 -24490
rect 29370 -24730 29450 -24720
rect 29520 -24640 29600 -24630
rect 27730 -25670 27810 -25660
rect 27730 -25760 27740 -25670
rect 27800 -25760 27810 -25670
rect 29380 -25760 29440 -24730
rect 29520 -24870 29530 -24640
rect 29590 -24870 29600 -24640
rect 29520 -24880 29600 -24870
rect 27730 -25770 27810 -25760
rect 29370 -25770 29450 -25760
rect 27740 -25975 27800 -25770
rect 29370 -25970 29380 -25770
rect 29440 -25970 29450 -25770
rect 27730 -25985 27810 -25975
rect 29370 -25980 29450 -25970
rect 27730 -26075 27740 -25985
rect 27800 -26075 27810 -25985
rect 27730 -26085 27810 -26075
rect 27740 -26540 27800 -26085
rect 27730 -26550 27810 -26540
rect 27730 -26640 27740 -26550
rect 27800 -26640 27810 -26550
rect 27730 -26650 27810 -26640
rect 27740 -26860 27800 -26650
rect 27730 -26870 27810 -26860
rect 27730 -26960 27740 -26870
rect 27800 -26960 27810 -26870
rect 27730 -26970 27810 -26960
rect 27740 -27175 27800 -26970
rect 27730 -27185 27810 -27175
rect 27730 -27275 27740 -27185
rect 27800 -27275 27810 -27185
rect 27730 -27285 27810 -27275
rect 29070 -27850 29150 -27840
rect 29070 -28050 29080 -27850
rect 29140 -28050 29150 -27850
rect 29070 -28060 29150 -28050
rect 27610 -28790 27690 -28780
rect 27610 -28880 27620 -28790
rect 27680 -28880 27690 -28790
rect 27610 -28890 27690 -28880
rect 27620 -29100 27680 -28890
rect 27610 -29110 27690 -29100
rect 27610 -29200 27620 -29110
rect 27680 -29200 27690 -29110
rect 27610 -29210 27690 -29200
rect 27620 -29820 27680 -29210
rect 27610 -29830 27690 -29820
rect 27610 -29920 27620 -29830
rect 27680 -29920 27690 -29830
rect 29080 -29920 29140 -28060
rect 29220 -28890 29300 -28880
rect 29220 -29090 29230 -28890
rect 29290 -29090 29300 -28890
rect 29220 -29100 29300 -29090
rect 27610 -29930 27690 -29920
rect 29070 -29930 29150 -29920
rect 27620 -30135 27680 -29930
rect 29070 -30130 29080 -29930
rect 29140 -30130 29150 -29930
rect 27610 -30145 27690 -30135
rect 29070 -30140 29150 -30130
rect 27610 -30235 27620 -30145
rect 27680 -30235 27690 -30145
rect 27610 -30245 27690 -30235
rect 27490 -30870 27570 -30860
rect 27490 -30960 27500 -30870
rect 27560 -30960 27570 -30870
rect 27490 -30970 27570 -30960
rect 27370 -31025 27450 -31015
rect 27370 -31115 27380 -31025
rect 27440 -31115 27450 -31025
rect 27370 -31125 27450 -31115
rect 27380 -31330 27440 -31125
rect 27500 -31175 27560 -30970
rect 27490 -31185 27570 -31175
rect 27490 -31275 27500 -31185
rect 27560 -31275 27570 -31185
rect 27490 -31285 27570 -31275
rect 27370 -31340 27450 -31330
rect 27370 -31430 27380 -31340
rect 27440 -31430 27450 -31340
rect 27370 -31440 27450 -31430
rect 27380 -31600 27440 -31440
rect 27500 -31600 27560 -31285
rect 27620 -31600 27680 -30245
rect 29080 -30400 29140 -30140
rect 28930 -30410 29170 -30400
rect 28930 -30480 28940 -30410
rect 29160 -30480 29170 -30410
rect 28930 -30490 29170 -30480
rect 29230 -30550 29290 -29100
rect 29060 -30560 29300 -30550
rect 29060 -30630 29070 -30560
rect 29290 -30630 29300 -30560
rect 29060 -30640 29300 -30630
rect 29060 -30950 29150 -30640
rect 29380 -30700 29440 -25980
rect 29530 -26800 29590 -24880
rect 29520 -26810 29600 -26800
rect 29520 -27010 29530 -26810
rect 29590 -27010 29600 -26810
rect 29520 -27020 29600 -27010
rect 29210 -30710 29450 -30700
rect 29210 -30780 29220 -30710
rect 29440 -30780 29450 -30710
rect 29210 -30790 29450 -30780
rect 29530 -30850 29590 -27020
rect 29680 -28710 29740 -24110
rect 29670 -28720 29750 -28710
rect 29670 -28940 29680 -28720
rect 29740 -28940 29750 -28720
rect 29830 -28860 29890 -23600
rect 31860 -23660 31960 -17210
rect 32510 -17800 32640 -16920
rect 32510 -18480 32520 -17800
rect 32630 -18480 32640 -17800
rect 32510 -18490 32640 -18480
rect 32510 -19600 32640 -19590
rect 32510 -20280 32520 -19600
rect 32630 -20280 32640 -19600
rect 32510 -20360 32640 -20280
rect 33180 -20340 33320 -20330
rect 32500 -20370 32650 -20360
rect 32500 -20530 32510 -20370
rect 32640 -20530 32650 -20370
rect 33180 -20460 33190 -20340
rect 33310 -20460 33320 -20340
rect 33180 -20470 33320 -20460
rect 32500 -20540 32650 -20530
rect 32510 -21400 32640 -20540
rect 32510 -22080 32520 -21400
rect 32630 -22080 32640 -21400
rect 32510 -22090 32640 -22080
rect 33200 -22140 33300 -20470
rect 33200 -22240 33210 -22140
rect 33290 -22240 33300 -22140
rect 33200 -22420 33300 -22240
rect 32620 -22430 33310 -22420
rect 32620 -22490 32630 -22430
rect 33300 -22490 33310 -22430
rect 32620 -22500 33310 -22490
rect 32690 -23070 33240 -23060
rect 32690 -23150 32700 -23070
rect 32910 -23150 33020 -23070
rect 33230 -23150 33240 -23070
rect 32690 -23160 33240 -23150
rect 31810 -23670 32010 -23660
rect 31810 -23850 31820 -23670
rect 32000 -23850 32010 -23670
rect 31810 -23860 32010 -23850
rect 29970 -24140 30050 -24130
rect 29970 -24370 29980 -24140
rect 30040 -24370 30050 -24140
rect 29970 -24380 30050 -24370
rect 29670 -28950 29750 -28940
rect 29820 -28870 29900 -28860
rect 29820 -29090 29830 -28870
rect 29890 -29090 29900 -28870
rect 29980 -29010 30040 -24380
rect 32880 -24470 32940 -23160
rect 33440 -23550 33540 -9640
rect 34100 -9570 34250 -9560
rect 34100 -9730 34110 -9570
rect 34240 -9730 34250 -9570
rect 34100 -9740 34250 -9730
rect 34110 -10600 34240 -9740
rect 34820 -9860 34920 -8200
rect 35710 -8800 35840 -8790
rect 35710 -9360 35720 -8800
rect 35830 -9360 35840 -8800
rect 35710 -9560 35840 -9360
rect 35700 -9570 35850 -9560
rect 35700 -9730 35710 -9570
rect 35840 -9730 35850 -9570
rect 35700 -9740 35850 -9730
rect 34800 -9870 34940 -9860
rect 34800 -9990 34810 -9870
rect 34930 -9990 34940 -9870
rect 34800 -10000 34940 -9990
rect 34110 -11110 34120 -10600
rect 34230 -11110 34240 -10600
rect 34110 -11360 34240 -11110
rect 34100 -11370 34250 -11360
rect 34100 -11530 34110 -11370
rect 34240 -11530 34250 -11370
rect 34100 -11540 34250 -11530
rect 34110 -12400 34240 -11540
rect 34820 -11660 34920 -10000
rect 35710 -10600 35840 -9740
rect 35710 -11110 35720 -10600
rect 35830 -11110 35840 -10600
rect 35000 -11310 35140 -11300
rect 35000 -11430 35010 -11310
rect 35130 -11430 35140 -11310
rect 35710 -11360 35840 -11110
rect 35000 -11440 35140 -11430
rect 34800 -11670 34940 -11660
rect 34800 -11790 34810 -11670
rect 34930 -11790 34940 -11670
rect 34800 -11800 34940 -11790
rect 34110 -12910 34120 -12400
rect 34230 -12910 34240 -12400
rect 34110 -13160 34240 -12910
rect 34100 -13170 34250 -13160
rect 34100 -13330 34110 -13170
rect 34240 -13330 34250 -13170
rect 34100 -13340 34250 -13330
rect 34110 -14200 34240 -13340
rect 34820 -13460 34920 -11800
rect 35040 -13100 35140 -11440
rect 35700 -11370 35850 -11360
rect 35700 -11530 35710 -11370
rect 35840 -11530 35850 -11370
rect 35700 -11540 35850 -11530
rect 35000 -13110 35140 -13100
rect 35000 -13230 35010 -13110
rect 35130 -13230 35140 -13110
rect 35710 -12400 35840 -11540
rect 35710 -12910 35720 -12400
rect 35830 -12910 35840 -12400
rect 35710 -13160 35840 -12910
rect 35000 -13240 35140 -13230
rect 34800 -13470 34940 -13460
rect 34800 -13590 34810 -13470
rect 34930 -13590 34940 -13470
rect 34800 -13600 34940 -13590
rect 34110 -14710 34120 -14200
rect 34230 -14710 34240 -14200
rect 34110 -14890 34240 -14710
rect 34110 -16000 34240 -15990
rect 34110 -16680 34120 -16000
rect 34230 -16680 34240 -16000
rect 34110 -16770 34240 -16680
rect 34110 -16920 34120 -16770
rect 34230 -16920 34240 -16770
rect 34110 -17800 34240 -16920
rect 34110 -18480 34120 -17800
rect 34230 -18480 34240 -17800
rect 34110 -18490 34240 -18480
rect 34110 -19600 34240 -19590
rect 34110 -20280 34120 -19600
rect 34230 -20280 34240 -19600
rect 34110 -20360 34240 -20280
rect 34100 -20370 34250 -20360
rect 34100 -20530 34110 -20370
rect 34240 -20530 34250 -20370
rect 34100 -20540 34250 -20530
rect 34110 -21400 34240 -20540
rect 34110 -22080 34120 -21400
rect 34230 -22080 34240 -21400
rect 34110 -22090 34240 -22080
rect 34010 -22170 34370 -22160
rect 34010 -22240 34020 -22170
rect 34360 -22240 34370 -22170
rect 34010 -22250 34370 -22240
rect 34030 -22430 34320 -22250
rect 34030 -22490 34040 -22430
rect 34310 -22490 34320 -22430
rect 34030 -22500 34320 -22490
rect 34060 -23100 34310 -23090
rect 34060 -23160 34070 -23100
rect 34300 -23160 34310 -23100
rect 34060 -23170 34310 -23160
rect 33400 -23560 33920 -23550
rect 33400 -23620 33410 -23560
rect 33910 -23620 33920 -23560
rect 33400 -23630 33920 -23620
rect 33160 -24220 34150 -24210
rect 33160 -24280 33170 -24220
rect 33280 -24280 33410 -24220
rect 33600 -24280 33730 -24220
rect 33920 -24280 34040 -24220
rect 34140 -24280 34150 -24220
rect 33160 -24290 34150 -24280
rect 32790 -24480 33040 -24470
rect 32790 -24550 32800 -24480
rect 33030 -24550 33040 -24480
rect 32790 -24560 33040 -24550
rect 33640 -24770 33700 -24290
rect 34200 -24620 34260 -23170
rect 34820 -23460 34920 -13600
rect 35040 -14900 35140 -13240
rect 35700 -13170 35850 -13160
rect 35700 -13330 35710 -13170
rect 35840 -13330 35850 -13170
rect 35700 -13340 35850 -13330
rect 35710 -14200 35840 -13340
rect 35710 -14710 35720 -14200
rect 35830 -14710 35840 -14200
rect 35710 -14890 35840 -14710
rect 35000 -14910 35140 -14900
rect 35000 -15030 35010 -14910
rect 35130 -15030 35140 -14910
rect 35000 -15040 35140 -15030
rect 34610 -24220 34780 -24210
rect 34610 -24280 34620 -24220
rect 34770 -24280 34780 -24220
rect 34610 -24290 34780 -24280
rect 34840 -24480 34900 -23460
rect 35040 -23550 35140 -15040
rect 35710 -16000 35840 -15990
rect 35710 -16680 35720 -16000
rect 35830 -16680 35840 -16000
rect 35710 -16770 35840 -16680
rect 35710 -16920 35720 -16770
rect 35830 -16920 35840 -16770
rect 35710 -17800 35840 -16920
rect 35710 -18480 35720 -17800
rect 35830 -18480 35840 -17800
rect 35710 -18490 35840 -18480
rect 35710 -19600 35840 -19590
rect 35710 -20280 35720 -19600
rect 35830 -20280 35840 -19600
rect 35710 -20360 35840 -20280
rect 35700 -20370 35850 -20360
rect 35700 -20530 35710 -20370
rect 35840 -20530 35850 -20370
rect 35700 -20540 35850 -20530
rect 35710 -21400 35840 -20540
rect 35710 -22080 35720 -21400
rect 35830 -22080 35840 -21400
rect 35710 -22090 35840 -22080
rect 35000 -23560 37030 -23550
rect 37020 -23620 37030 -23560
rect 35000 -23630 37030 -23620
rect 34980 -24220 37030 -24210
rect 34980 -24280 34990 -24220
rect 37020 -24280 37030 -24220
rect 34980 -24290 37030 -24280
rect 34800 -24490 34940 -24480
rect 34800 -24610 34810 -24490
rect 34930 -24610 34940 -24490
rect 34800 -24620 34940 -24610
rect 34110 -24630 34360 -24620
rect 34110 -24700 34120 -24630
rect 34350 -24700 34360 -24630
rect 37120 -24640 37290 -24630
rect 34110 -24710 34360 -24700
rect 34800 -24660 34910 -24650
rect 30280 -24780 30520 -24770
rect 30280 -24850 30290 -24780
rect 30510 -24850 30520 -24780
rect 30280 -24860 30520 -24850
rect 33550 -24780 33800 -24770
rect 33550 -24850 33560 -24780
rect 33790 -24850 33800 -24780
rect 33550 -24860 33800 -24850
rect 34800 -24860 34810 -24660
rect 34900 -24860 34910 -24660
rect 37120 -24780 37130 -24640
rect 37270 -24780 37290 -24640
rect 37120 -24790 37290 -24780
rect 30120 -24940 30200 -24930
rect 30120 -25170 30130 -24940
rect 30190 -25170 30200 -24940
rect 30120 -25180 30200 -25170
rect 29820 -29100 29900 -29090
rect 29970 -29020 30050 -29010
rect 29970 -29240 29980 -29020
rect 30040 -29240 30050 -29020
rect 30130 -29160 30190 -25180
rect 29970 -29250 30050 -29240
rect 30120 -29170 30200 -29160
rect 30120 -29390 30130 -29170
rect 30190 -29390 30200 -29170
rect 30280 -29310 30340 -24860
rect 34800 -24940 34910 -24860
rect 34800 -25010 34810 -24940
rect 34900 -25010 34910 -24940
rect 30420 -25090 30500 -25080
rect 30420 -25320 30430 -25090
rect 30490 -25320 30500 -25090
rect 30420 -25330 30500 -25320
rect 34800 -25200 34910 -25010
rect 34800 -25270 34810 -25200
rect 34900 -25270 34910 -25200
rect 30120 -29400 30200 -29390
rect 30270 -29320 30350 -29310
rect 30270 -29540 30280 -29320
rect 30340 -29540 30350 -29320
rect 30430 -29460 30490 -25330
rect 34800 -25460 34910 -25270
rect 34800 -25530 34810 -25460
rect 34900 -25530 34910 -25460
rect 34800 -25720 34910 -25530
rect 34800 -25790 34810 -25720
rect 34900 -25790 34910 -25720
rect 34800 -25980 34910 -25790
rect 34800 -26050 34810 -25980
rect 34900 -26050 34910 -25980
rect 34800 -26240 34910 -26050
rect 34800 -26310 34810 -26240
rect 34900 -26310 34910 -26240
rect 34800 -26500 34910 -26310
rect 34800 -26570 34810 -26500
rect 34900 -26570 34910 -26500
rect 34800 -26760 34910 -26570
rect 34800 -26830 34810 -26760
rect 34900 -26830 34910 -26760
rect 34800 -26840 34910 -26830
rect 37180 -24940 37290 -24790
rect 37180 -25010 37190 -24940
rect 37280 -25010 37290 -24940
rect 37180 -25200 37290 -25010
rect 37180 -25270 37190 -25200
rect 37280 -25270 37290 -25200
rect 37180 -25460 37290 -25270
rect 37180 -25530 37190 -25460
rect 37280 -25530 37290 -25460
rect 37180 -25720 37290 -25530
rect 37180 -25790 37190 -25720
rect 37280 -25790 37290 -25720
rect 37180 -25980 37290 -25790
rect 37180 -26050 37190 -25980
rect 37280 -26050 37290 -25980
rect 37180 -26240 37290 -26050
rect 37180 -26310 37190 -26240
rect 37280 -26310 37290 -26240
rect 37180 -26500 37290 -26310
rect 37180 -26570 37190 -26500
rect 37280 -26570 37290 -26500
rect 37180 -26760 37290 -26570
rect 37180 -26830 37190 -26760
rect 37280 -26830 37290 -26760
rect 37180 -26840 37290 -26830
rect 36020 -27010 36420 -27000
rect 36020 -27140 36030 -27010
rect 36410 -27140 36420 -27010
rect 36020 -27150 36420 -27140
rect 36520 -27010 36920 -27000
rect 36520 -27140 36530 -27010
rect 36910 -27140 36920 -27010
rect 36520 -27150 36920 -27140
rect 36900 -27540 38600 -27520
rect 36900 -27900 36920 -27540
rect 37680 -27900 38600 -27540
rect 36900 -27920 38600 -27900
rect 36900 -28160 37700 -28140
rect 36900 -28520 36920 -28160
rect 37680 -28520 37700 -28160
rect 36900 -28540 37700 -28520
rect 35780 -28850 35860 -28670
rect 36110 -28700 36190 -28670
rect 36020 -28710 36280 -28700
rect 36020 -28780 36030 -28710
rect 36270 -28780 36280 -28710
rect 36020 -28790 36280 -28780
rect 35680 -28860 35940 -28850
rect 35680 -28930 35690 -28860
rect 35930 -28930 35940 -28860
rect 35680 -28940 35940 -28930
rect 30270 -29550 30350 -29540
rect 30420 -29470 30500 -29460
rect 30420 -29690 30430 -29470
rect 30490 -29690 30500 -29470
rect 30420 -29700 30500 -29690
rect 32780 -30336 32860 -30320
rect 32780 -30400 32794 -30336
rect 32600 -30410 32794 -30400
rect 32846 -30410 32860 -30336
rect 32600 -30480 32610 -30410
rect 32850 -30480 32860 -30410
rect 32600 -30488 32794 -30480
rect 32846 -30488 32860 -30480
rect 32600 -30490 32860 -30488
rect 32780 -30504 32860 -30490
rect 33110 -30342 33190 -30320
rect 33110 -30494 33126 -30342
rect 33178 -30424 33190 -30342
rect 33780 -30336 33860 -30320
rect 33178 -30494 33398 -30424
rect 33110 -30504 33398 -30494
rect 33780 -30488 33794 -30336
rect 33846 -30488 33860 -30336
rect 33780 -30504 33860 -30488
rect 34110 -30342 34190 -30320
rect 34110 -30494 34126 -30342
rect 34178 -30424 34190 -30342
rect 34780 -30336 34860 -30320
rect 34178 -30494 34450 -30424
rect 34110 -30504 34450 -30494
rect 34780 -30488 34794 -30336
rect 34846 -30488 34860 -30336
rect 34780 -30504 34860 -30488
rect 35110 -30342 35190 -30320
rect 35110 -30494 35126 -30342
rect 35178 -30424 35190 -30342
rect 35780 -30336 35860 -28940
rect 35178 -30494 35436 -30424
rect 35110 -30504 35436 -30494
rect 35780 -30488 35794 -30336
rect 35846 -30488 35860 -30336
rect 35780 -30504 35860 -30488
rect 36110 -30342 36190 -28790
rect 36780 -29150 36860 -28670
rect 37110 -29000 37190 -28670
rect 37020 -29010 37280 -29000
rect 37020 -29080 37030 -29010
rect 37270 -29080 37280 -29010
rect 37020 -29090 37280 -29080
rect 36690 -29160 36950 -29150
rect 36690 -29230 36700 -29160
rect 36940 -29230 36950 -29160
rect 36690 -29240 36950 -29230
rect 36110 -30494 36126 -30342
rect 36178 -30494 36190 -30342
rect 36110 -30504 36190 -30494
rect 36780 -30336 36860 -29240
rect 36780 -30488 36794 -30336
rect 36846 -30488 36860 -30336
rect 36780 -30504 36860 -30488
rect 37110 -30342 37190 -29090
rect 37780 -29450 37860 -28670
rect 38110 -29300 38190 -28670
rect 38020 -29310 38280 -29300
rect 38020 -29380 38030 -29310
rect 38270 -29380 38280 -29310
rect 38020 -29390 38280 -29380
rect 37690 -29460 37950 -29450
rect 37690 -29530 37700 -29460
rect 37940 -29530 37950 -29460
rect 37690 -29540 37950 -29530
rect 37110 -30494 37126 -30342
rect 37178 -30494 37190 -30342
rect 37110 -30504 37190 -30494
rect 37780 -30336 37860 -29540
rect 37780 -30488 37794 -30336
rect 37846 -30488 37860 -30336
rect 37780 -30504 37860 -30488
rect 38110 -30342 38190 -29390
rect 38110 -30494 38126 -30342
rect 38178 -30494 38190 -30342
rect 38110 -30504 38190 -30494
rect 38400 -30154 38600 -27920
rect 33318 -30550 33398 -30504
rect 33310 -30560 33570 -30550
rect 33310 -30630 33320 -30560
rect 33560 -30630 33570 -30560
rect 33310 -30640 33570 -30630
rect 34370 -30700 34450 -30504
rect 34310 -30712 34570 -30700
rect 34310 -30782 34320 -30712
rect 34560 -30782 34570 -30712
rect 34310 -30790 34570 -30782
rect 35356 -30850 35436 -30504
rect 38400 -30730 38410 -30154
rect 38588 -30730 38600 -30154
rect 38400 -30750 38600 -30730
rect 29360 -30860 29600 -30850
rect 29360 -30930 29370 -30860
rect 29590 -30930 29600 -30860
rect 29360 -30940 29600 -30930
rect 35310 -30860 35570 -30850
rect 35310 -30930 35320 -30860
rect 35560 -30930 35570 -30860
rect 35310 -30940 35570 -30930
rect 29060 -30960 29300 -30950
rect 29060 -31030 29070 -30960
rect 29290 -31030 29300 -30960
rect 29060 -31040 29300 -31030
rect 26220 -31800 27320 -31600
rect 30820 -31680 31260 -31660
rect 26220 -31880 26230 -31800
rect 25690 -31890 26230 -31880
rect 19800 -32010 19940 -32000
rect 19800 -32130 19810 -32010
rect 19930 -32130 19940 -32010
rect 19800 -32140 19940 -32130
rect 30820 -32440 30840 -31680
rect 31240 -32440 31260 -31680
rect 30820 -32460 31260 -32440
rect 33120 -33520 33220 -31814
rect 34120 -33520 34220 -31876
rect 35120 -33520 35220 -31842
rect 36120 -33520 36220 -31820
rect 37120 -33520 37220 -31894
rect 38120 -33520 38220 -31894
rect 38406 -32180 38540 -32160
rect 38300 -32690 38320 -32314
rect 38520 -32690 38540 -32180
rect 38300 -32910 38310 -32690
rect 38530 -32910 38540 -32690
rect 38300 -32920 38540 -32910
<< via2 >>
rect -350 11610 -170 11990
rect 2210 11890 2330 12010
rect 90 11310 270 11690
rect 1990 11590 2110 11710
rect -70 10870 -10 10930
rect -70 10070 -10 10130
rect -70 9270 -10 9330
rect -70 8470 -10 8530
rect -70 7670 -10 7730
rect -70 6870 -10 6930
rect -70 6070 -10 6130
rect -70 5270 -10 5330
rect -350 -7170 -170 -6590
rect -350 -31830 -170 -31450
rect 2130 10870 2190 10930
rect 4410 11890 4530 12010
rect 4190 11590 4310 11710
rect 2510 11180 2690 11240
rect 3170 11180 3350 11240
rect 3830 11180 4010 11240
rect 4330 10870 4390 10930
rect 6610 11890 6730 12010
rect 6390 11590 6510 11710
rect 4710 11180 4890 11240
rect 5370 11180 5550 11240
rect 6030 11180 6210 11240
rect 6530 10870 6590 10930
rect 8810 11890 8930 12010
rect 8590 11590 8710 11710
rect 6910 11040 7090 11100
rect 7570 11040 7750 11100
rect 8230 11040 8410 11100
rect 8730 10870 8790 10930
rect 11010 11890 11130 12010
rect 10790 11590 10910 11710
rect 9110 11040 9290 11100
rect 9770 11040 9950 11100
rect 10430 11040 10610 11100
rect 10930 10870 10990 10930
rect 13210 11890 13330 12010
rect 12990 11590 13110 11710
rect 11310 11040 11490 11100
rect 11970 11040 12150 11100
rect 12630 11040 12810 11100
rect 13130 10870 13190 10930
rect 15410 11890 15530 12010
rect 15190 11590 15310 11710
rect 13510 11040 13690 11100
rect 14170 11040 14350 11100
rect 14830 11040 15010 11100
rect 15330 10870 15390 10930
rect 17610 11890 17730 12010
rect 17390 11590 17510 11710
rect 15710 11180 15890 11240
rect 16370 11180 16550 11240
rect 17030 11180 17210 11240
rect 17530 10870 17590 10930
rect 19810 11890 19930 12010
rect 36920 12280 38280 12540
rect 19590 11590 19710 11710
rect 17910 11180 18090 11240
rect 18570 11180 18750 11240
rect 19230 11180 19410 11240
rect 19730 10870 19790 10930
rect 21930 10870 21990 10930
rect 2130 10070 2190 10130
rect 2510 10550 4010 10610
rect 2510 10240 2690 10300
rect 3170 10240 3350 10300
rect 3830 10240 4010 10300
rect 4330 10070 4390 10130
rect 4710 10550 6210 10610
rect 4710 10240 4890 10300
rect 5370 10240 5550 10300
rect 6030 10240 6210 10300
rect 6530 10070 6590 10130
rect 6910 10550 8410 10610
rect 6910 10380 7090 10440
rect 7570 10380 7750 10440
rect 8230 10380 8410 10440
rect 8730 10070 8790 10130
rect 9110 10550 10610 10610
rect 9110 10380 9290 10440
rect 9770 10380 9950 10440
rect 10430 10380 10610 10440
rect 10930 10070 10990 10130
rect 11310 10550 12810 10610
rect 11310 10380 11490 10440
rect 11970 10380 12150 10440
rect 12630 10380 12810 10440
rect 13130 10070 13190 10130
rect 13510 10550 15010 10610
rect 13510 10380 13690 10440
rect 14170 10380 14350 10440
rect 14830 10380 15010 10440
rect 15330 10070 15390 10130
rect 15710 10550 17210 10610
rect 15710 10240 15890 10300
rect 16370 10240 16550 10300
rect 17030 10240 17210 10300
rect 17530 10070 17590 10130
rect 17910 10550 19410 10610
rect 17910 10240 18090 10300
rect 18570 10240 18750 10300
rect 19230 10240 19410 10300
rect 19730 10070 19790 10130
rect 21930 10070 21990 10130
rect 2130 9270 2190 9330
rect 2510 9750 4010 9810
rect 2510 9580 2690 9640
rect 3170 9580 3350 9640
rect 3830 9580 4010 9640
rect 4330 9270 4390 9330
rect 4710 9750 6210 9810
rect 4710 9580 4890 9640
rect 5370 9580 5550 9640
rect 6030 9580 6210 9640
rect 6530 9270 6590 9330
rect 6910 9750 8410 9810
rect 6910 9440 7090 9500
rect 7570 9440 7750 9500
rect 8230 9440 8410 9500
rect 8730 9270 8790 9330
rect 9110 9750 10610 9810
rect 9110 9440 9290 9500
rect 9770 9440 9950 9500
rect 10430 9440 10610 9500
rect 10930 9270 10990 9330
rect 11310 9750 12810 9810
rect 11310 9440 11490 9500
rect 11970 9440 12150 9500
rect 12630 9440 12810 9500
rect 13130 9270 13190 9330
rect 13510 9750 15010 9810
rect 13510 9440 13690 9500
rect 14170 9440 14350 9500
rect 14830 9440 15010 9500
rect 15330 9270 15390 9330
rect 15710 9750 17210 9810
rect 15710 9580 15890 9640
rect 16370 9580 16550 9640
rect 17030 9580 17210 9640
rect 17530 9270 17590 9330
rect 17910 9750 19410 9810
rect 17910 9580 18090 9640
rect 18570 9580 18750 9640
rect 19230 9580 19410 9640
rect 430 8910 610 8990
rect 430 8110 610 8190
rect 430 7310 610 7390
rect 19730 9270 19790 9330
rect 2130 8470 2190 8530
rect 2510 8640 2690 8700
rect 3170 8640 3350 8700
rect 3830 8640 4010 8700
rect 4330 8470 4390 8530
rect 4710 8950 6210 9010
rect 4710 8640 4890 8700
rect 5370 8640 5550 8700
rect 6030 8640 6210 8700
rect 6530 8470 6590 8530
rect 6910 8950 8410 9010
rect 6910 8780 7090 8840
rect 7570 8780 7750 8840
rect 8230 8780 8410 8840
rect 8730 8470 8790 8530
rect 9110 8950 10610 9010
rect 9110 8780 9290 8840
rect 9770 8780 9950 8840
rect 10430 8780 10610 8840
rect 10930 8470 10990 8530
rect 11310 8950 12810 9010
rect 11310 8780 11490 8840
rect 11970 8780 12150 8840
rect 12630 8780 12810 8840
rect 13130 8470 13190 8530
rect 13510 8950 15010 9010
rect 13510 8780 13690 8840
rect 14170 8780 14350 8840
rect 14830 8780 15010 8840
rect 15330 8470 15390 8530
rect 15710 8950 17210 9010
rect 15710 8640 15890 8700
rect 16370 8640 16550 8700
rect 17030 8640 17210 8700
rect 17530 8470 17590 8530
rect 17910 8640 18090 8700
rect 18570 8640 18750 8700
rect 19230 8640 19410 8700
rect 19730 8470 19790 8530
rect 2130 7670 2190 7730
rect 2510 7840 2690 7900
rect 3170 7840 3350 7900
rect 3830 7840 4010 7900
rect 4330 7670 4390 7730
rect 4710 8150 6210 8210
rect 4710 7840 4890 7900
rect 5370 7840 5550 7900
rect 6030 7840 6210 7900
rect 6530 7670 6590 7730
rect 6910 8150 8410 8210
rect 6910 7980 7090 8040
rect 7570 7980 7750 8040
rect 8230 7980 8410 8040
rect 8730 7670 8790 7730
rect 9110 8150 10610 8210
rect 9110 7980 9290 8040
rect 9770 7980 9950 8040
rect 10430 7980 10610 8040
rect 10930 7670 10990 7730
rect 11310 8150 12810 8210
rect 11310 7980 11490 8040
rect 11970 7980 12150 8040
rect 12630 7980 12810 8040
rect 13130 7670 13190 7730
rect 13510 8150 15010 8210
rect 13510 7980 13690 8040
rect 14170 7980 14350 8040
rect 14830 7980 15010 8040
rect 15330 7670 15390 7730
rect 15710 8150 17210 8210
rect 15710 7840 15890 7900
rect 16370 7840 16550 7900
rect 17030 7840 17210 7900
rect 17530 7670 17590 7730
rect 17910 7840 18090 7900
rect 18570 7840 18750 7900
rect 19230 7840 19410 7900
rect 430 6510 610 6590
rect 1290 4350 1470 4530
rect 19730 7670 19790 7730
rect 2130 6870 2190 6930
rect 2510 7180 2690 7240
rect 3170 7180 3350 7240
rect 3830 7180 4010 7240
rect 4330 6870 4390 6930
rect 4710 7350 6210 7410
rect 4710 7180 4890 7240
rect 5370 7180 5550 7240
rect 6030 7180 6210 7240
rect 6530 6870 6590 6930
rect 6910 7350 8410 7410
rect 6910 7040 7090 7100
rect 7570 7040 7750 7100
rect 8230 7040 8410 7100
rect 8730 6870 8790 6930
rect 9110 7350 10610 7410
rect 9110 7040 9290 7100
rect 9770 7040 9950 7100
rect 10430 7040 10610 7100
rect 10930 6870 10990 6930
rect 11310 7350 12810 7410
rect 11310 7040 11490 7100
rect 11970 7040 12150 7100
rect 12630 7040 12810 7100
rect 13130 6870 13190 6930
rect 13510 7350 15010 7410
rect 13510 7040 13690 7100
rect 14170 7040 14350 7100
rect 14830 7040 15010 7100
rect 15330 6870 15390 6930
rect 15710 7350 17210 7410
rect 15710 7180 15890 7240
rect 16370 7180 16550 7240
rect 17030 7180 17210 7240
rect 17530 6870 17590 6930
rect 17910 7180 18090 7240
rect 18570 7180 18750 7240
rect 19230 7180 19410 7240
rect 19730 6870 19790 6930
rect 21930 9270 21990 9330
rect 21310 8910 21490 8990
rect 21930 8470 21990 8530
rect 21310 8110 21490 8190
rect 21930 7670 21990 7730
rect 2130 6070 2190 6130
rect 2510 6240 2690 6300
rect 3170 6240 3350 6300
rect 3830 6240 4010 6300
rect 4330 6070 4390 6130
rect 4710 6550 6210 6610
rect 4710 6240 4890 6300
rect 5370 6240 5550 6300
rect 6030 6240 6210 6300
rect 6530 6070 6590 6130
rect 6910 6550 8410 6610
rect 6910 6380 7090 6440
rect 7570 6380 7750 6440
rect 8230 6380 8410 6440
rect 8730 6070 8790 6130
rect 9110 6550 10610 6610
rect 9110 6380 9290 6440
rect 9770 6380 9950 6440
rect 10430 6380 10610 6440
rect 10930 6070 10990 6130
rect 11310 6550 12810 6610
rect 11310 6380 11490 6440
rect 11970 6380 12150 6440
rect 12630 6380 12810 6440
rect 13130 6070 13190 6130
rect 13510 6550 15010 6610
rect 13510 6380 13690 6440
rect 14170 6380 14350 6440
rect 14830 6380 15010 6440
rect 15330 6070 15390 6130
rect 15710 6550 17210 6610
rect 15710 6240 15890 6300
rect 16370 6240 16550 6300
rect 17030 6240 17210 6300
rect 17530 6070 17590 6130
rect 17910 6240 18090 6300
rect 18570 6240 18750 6300
rect 19230 6240 19410 6300
rect 19730 6070 19790 6130
rect 2130 5270 2190 5330
rect 2510 5750 4010 5810
rect 2510 5580 2690 5640
rect 3170 5580 3350 5640
rect 3830 5580 4010 5640
rect 4330 5270 4390 5330
rect 4710 5750 6210 5810
rect 4710 5580 4890 5640
rect 5370 5580 5550 5640
rect 6030 5580 6210 5640
rect 6530 5270 6590 5330
rect 6910 5750 8410 5810
rect 6910 5440 7090 5500
rect 7570 5440 7750 5500
rect 8230 5440 8410 5500
rect 8730 5270 8790 5330
rect 9110 5750 10610 5810
rect 9110 5440 9290 5500
rect 9770 5440 9950 5500
rect 10430 5440 10610 5500
rect 10930 5270 10990 5330
rect 11310 5750 12810 5810
rect 11310 5440 11490 5500
rect 11970 5440 12150 5500
rect 12630 5440 12810 5500
rect 13130 5270 13190 5330
rect 13510 5750 15010 5810
rect 13510 5440 13690 5500
rect 14170 5440 14350 5500
rect 14830 5440 15010 5500
rect 15330 5270 15390 5330
rect 15710 5750 17210 5810
rect 15710 5580 15890 5640
rect 16370 5580 16550 5640
rect 17030 5580 17210 5640
rect 17530 5270 17590 5330
rect 17910 5750 19410 5810
rect 17910 5580 18090 5640
rect 18570 5580 18750 5640
rect 19230 5580 19410 5640
rect 19730 5270 19790 5330
rect 2510 4950 4010 5010
rect 4710 4950 6210 5010
rect 6910 4950 8410 5010
rect 1630 3950 1810 4130
rect 1170 3150 1330 3330
rect 2770 3150 2930 3330
rect 4370 3150 4530 3330
rect 5970 3150 6130 3330
rect 7570 3150 7730 3330
rect 480 -4780 660 2220
rect 2110 2090 2230 2250
rect 3710 2090 3830 2250
rect 2110 290 2230 450
rect 5310 2090 5430 2250
rect 3710 290 3830 450
rect 2110 -1510 2230 -1350
rect 6910 2090 7030 2250
rect 5310 290 5430 450
rect 3710 -1510 3830 -1350
rect 2110 -3310 2230 -3150
rect 9110 4950 10610 5010
rect 11310 4950 12810 5010
rect 13510 4950 15010 5010
rect 15710 4950 17210 5010
rect 17910 4950 19410 5010
rect 20110 4350 20290 4530
rect 21310 7310 21490 7390
rect 21930 6870 21990 6930
rect 21310 6510 21490 6590
rect 21930 6070 21990 6130
rect 21930 5270 21990 5330
rect 23050 4710 23580 4970
rect 20450 3950 20630 4130
rect 9170 3150 9330 3330
rect 7810 2810 7930 2930
rect 8510 2090 8630 2250
rect 6910 290 7030 450
rect 5310 -1510 5430 -1350
rect 3710 -3310 3830 -3150
rect 30824 10934 31194 11060
rect 29280 10720 29510 10790
rect 28960 10570 29190 10640
rect 28870 10310 28930 10480
rect 29020 10170 29080 10340
rect 27250 4750 27430 4930
rect 27370 4350 27550 4530
rect 29140 4290 29200 4520
rect 37190 10860 37340 11010
rect 33520 10720 33760 10790
rect 32480 10560 32720 10630
rect 31680 10420 31920 10490
rect 31330 10280 31570 10350
rect 37990 10780 38120 10960
rect 37610 10600 37760 10750
rect 30520 8170 30640 8290
rect 30910 7970 31030 8090
rect 29280 4190 29510 4260
rect 27630 3950 27810 4130
rect 30080 3860 30260 4040
rect 31680 3860 31860 4040
rect 35350 7570 35470 7690
rect 37510 7370 37630 7490
rect 36128 6982 36810 7176
rect 36230 6080 36410 6260
rect 36530 6080 36710 6260
rect 34900 5280 35110 5360
rect 36300 5300 36390 5370
rect 36300 5110 36390 5300
rect 36300 5040 36390 5110
rect 32500 4340 32640 4480
rect 34090 4340 34230 4480
rect 31530 3550 31690 3730
rect 32080 3610 32210 3740
rect 26620 3220 26760 3360
rect 10890 2870 11030 3010
rect 14190 2870 14350 3030
rect 18060 2870 18200 3010
rect 23220 2910 23400 3090
rect 11700 2620 11840 2770
rect 11000 2400 11140 2540
rect 10110 2090 10230 2250
rect 12600 2400 12740 2540
rect 13980 2400 14120 2540
rect 11710 2090 11830 2250
rect 8510 290 8630 450
rect 6910 -1510 7030 -1350
rect 5310 -3310 5430 -3150
rect 13310 2090 13430 2250
rect 10110 290 10230 450
rect 8510 -1510 8630 -1350
rect 6910 -3310 7030 -3150
rect 11710 290 11830 450
rect 10110 -1510 10230 -1350
rect 8510 -3310 8630 -3150
rect 13310 290 13430 450
rect 11710 -1510 11830 -1350
rect 10110 -3310 10230 -3150
rect 12880 -1260 13240 -1110
rect 13310 -1510 13430 -1350
rect 11710 -3310 11830 -3150
rect 16910 2640 17130 2780
rect 17380 2640 17490 2780
rect 17740 2640 17960 2780
rect 16510 2090 16630 2250
rect 14910 1320 15030 1980
rect 18110 2090 18230 2250
rect 19710 2090 19830 2250
rect 21310 2090 21430 2250
rect 22910 2090 23030 2250
rect 24510 2090 24630 2250
rect 26110 2090 26230 2250
rect 27710 2070 27830 2250
rect 29310 2070 29430 2250
rect 14910 -1510 15030 -1350
rect 15250 -1510 15370 -1350
rect 13310 -3310 13430 -3150
rect 16510 290 16630 450
rect 90 -6330 270 -5750
rect 7810 -7990 7930 -7870
rect 490 -22380 670 -8090
rect 2130 -9750 2230 -9590
rect 2130 -11550 2230 -11390
rect 3730 -9750 3830 -9590
rect 2130 -13350 2230 -13190
rect 3730 -11550 3830 -11390
rect 2130 -15150 2230 -14990
rect 5330 -9750 5430 -9590
rect 3730 -13350 3830 -13190
rect 2130 -16950 2230 -16790
rect 5330 -11550 5430 -11390
rect 3730 -15150 3830 -14990
rect 2130 -18750 2230 -18590
rect 6930 -9750 7030 -9590
rect 5330 -13350 5430 -13190
rect 3730 -16950 3830 -16790
rect 2130 -20550 2230 -20390
rect 6930 -11550 7030 -11390
rect 5330 -15150 5430 -14990
rect 3730 -18750 3830 -18590
rect 2130 -22350 2230 -22190
rect 8530 -9750 8630 -9590
rect 6930 -13350 7030 -13190
rect 5330 -16950 5430 -16790
rect 3730 -20550 3830 -20390
rect 10810 -8380 10930 -8260
rect 8530 -11550 8630 -11390
rect 6930 -15150 7030 -14990
rect 5330 -18750 5430 -18590
rect 3730 -22350 3830 -22190
rect 10130 -9750 10230 -9590
rect 8530 -13350 8630 -13190
rect 6930 -16950 7030 -16790
rect 5330 -20550 5430 -20390
rect 10130 -11550 10230 -11390
rect 8530 -15150 8630 -14990
rect 6930 -18750 7030 -18590
rect 5330 -22350 5430 -22190
rect 10130 -13350 10230 -13190
rect 8530 -16950 8630 -16790
rect 6930 -20550 7030 -20390
rect 10130 -15150 10230 -14990
rect 8530 -18750 8630 -18590
rect 6930 -22350 7030 -22190
rect 10130 -16950 10230 -16790
rect 8530 -20550 8630 -20390
rect 10130 -18750 10230 -18590
rect 8530 -22350 8630 -22190
rect 10130 -20550 10230 -20390
rect 12950 -6990 13110 -6830
rect 14910 -3310 15030 -3150
rect 16510 -1510 16630 -1350
rect 13310 -8380 13440 -8260
rect 13290 -13330 13460 -13170
rect 18110 290 18230 450
rect 16510 -3310 16630 -3150
rect 15570 -5350 15730 -5170
rect 15570 -5750 15730 -5570
rect 14910 -6610 15030 -6490
rect 13290 -15130 13460 -14970
rect 13300 -16950 13450 -16790
rect 13300 -18750 13450 -18590
rect 15790 -6150 15950 -5970
rect 18110 -1510 18230 -1350
rect 19710 290 19830 450
rect 18110 -3310 18230 -3150
rect 19710 -1510 19830 -1350
rect 21310 290 21430 450
rect 19710 -3310 19830 -3150
rect 21310 -1510 21430 -1350
rect 18770 -5350 18930 -5170
rect 18770 -5750 18930 -5570
rect 17390 -6950 17550 -6770
rect 17170 -7350 17330 -7170
rect 17170 -7750 17330 -7570
rect 16510 -8380 16640 -8260
rect 16510 -9730 16640 -9570
rect 18990 -6150 19150 -5970
rect 22910 290 23030 450
rect 21310 -3310 21430 -3150
rect 22910 -1510 23030 -1350
rect 24510 290 24630 450
rect 22910 -3310 23030 -3150
rect 24510 -1510 24630 -1350
rect 21970 -5350 22130 -5170
rect 21970 -5750 22130 -5570
rect 20590 -6950 20750 -6770
rect 20370 -7350 20530 -7170
rect 20370 -7750 20530 -7570
rect 18110 -9730 18240 -9570
rect 16510 -11530 16640 -11370
rect 14890 -13330 15060 -13170
rect 19710 -9730 19840 -9570
rect 18110 -11530 18240 -11370
rect 16510 -13330 16640 -13170
rect 14890 -15130 15060 -14970
rect 22190 -6150 22350 -5970
rect 24510 -3310 24630 -3150
rect 26110 290 26230 450
rect 26110 -1510 26230 -1350
rect 27710 270 27830 450
rect 26110 -3310 26230 -3150
rect 27710 -1530 27830 -1350
rect 25170 -5350 25330 -5170
rect 25170 -5750 25330 -5570
rect 23790 -6950 23950 -6770
rect 23570 -7350 23730 -7170
rect 23570 -7750 23730 -7570
rect 21310 -9730 21440 -9570
rect 19710 -11530 19840 -11370
rect 18110 -13330 18240 -13170
rect 16510 -15130 16640 -14970
rect 14900 -16950 15050 -16790
rect 22910 -9730 23040 -9570
rect 21310 -11530 21440 -11370
rect 19710 -13330 19840 -13170
rect 18110 -15130 18240 -14970
rect 16510 -16930 16640 -16770
rect 14900 -18750 15050 -18590
rect 25390 -6150 25550 -5970
rect 29310 270 29430 450
rect 27710 -3330 27830 -3150
rect 29310 -1530 29430 -1350
rect 30910 2070 31030 2250
rect 30910 270 31030 450
rect 33130 4070 33290 4110
rect 33130 4010 33290 4070
rect 31830 2910 31990 3090
rect 33180 2390 33330 2550
rect 32510 1030 32630 1150
rect 33180 280 33330 440
rect 32510 -490 32630 190
rect 30910 -1530 31030 -1350
rect 35700 4150 35840 4290
rect 34870 4010 35190 4090
rect 34780 2620 34930 2780
rect 34110 1030 34230 1150
rect 34790 1030 34920 1150
rect 34110 -490 34230 190
rect 29310 -3330 29430 -3150
rect 28370 -5350 28530 -5170
rect 28370 -5750 28530 -5570
rect 27690 -6150 27850 -5970
rect 26990 -6950 27150 -6770
rect 26770 -7350 26930 -7170
rect 26770 -7750 26930 -7570
rect 24510 -9730 24640 -9570
rect 22910 -11530 23040 -11370
rect 21310 -13330 21440 -13170
rect 19710 -15130 19840 -14970
rect 18110 -16930 18240 -16770
rect 16510 -18730 16640 -18570
rect 10130 -22350 10230 -22190
rect 10110 -22590 10250 -22450
rect 11050 -22850 11150 -22740
rect 11720 -22850 11820 -22740
rect 26110 -9730 26240 -9570
rect 24510 -11530 24640 -11370
rect 22910 -13330 23040 -13170
rect 21310 -15130 21440 -14970
rect 19710 -16930 19840 -16770
rect 18110 -18730 18240 -18570
rect 16510 -20530 16640 -20370
rect 28590 -6150 28750 -5970
rect 29290 -6150 29450 -5970
rect 30910 -3330 31030 -3150
rect 32510 -2570 32630 -2450
rect 37680 5300 37770 5370
rect 37680 5110 37770 5300
rect 37680 5040 37770 5110
rect 37880 3580 38010 3710
rect 35710 1030 35830 1150
rect 35710 -490 35830 190
rect 34110 -2570 34230 -2450
rect 34790 -2570 34920 -2450
rect 35710 -2570 35830 -2450
rect 36590 3220 36730 3360
rect 37310 1030 37430 1150
rect 30890 -6150 31050 -5970
rect 30190 -6950 30350 -6770
rect 29970 -7350 30130 -7170
rect 29970 -7750 30130 -7570
rect 27710 -9730 27840 -9570
rect 26110 -11530 26240 -11370
rect 24510 -13330 24640 -13170
rect 22910 -15130 23040 -14970
rect 21310 -16930 21440 -16770
rect 19710 -18730 19840 -18570
rect 18110 -20530 18240 -20370
rect 29310 -9730 29440 -9570
rect 27710 -11530 27840 -11370
rect 26110 -13330 26240 -13170
rect 24510 -15130 24640 -14970
rect 22910 -16930 23040 -16770
rect 21310 -18730 21440 -18570
rect 19710 -20530 19840 -20370
rect 30910 -9730 31040 -9570
rect 29310 -11530 29440 -11370
rect 27710 -13330 27840 -13170
rect 26110 -15130 26240 -14970
rect 32510 -9730 32640 -9570
rect 30910 -11530 31040 -11370
rect 29310 -13330 29440 -13170
rect 27710 -15130 27840 -14970
rect 24510 -16930 24640 -16770
rect 26110 -16930 26240 -16770
rect 22910 -18730 23040 -18570
rect 21310 -20530 21440 -20370
rect 32510 -11530 32640 -11370
rect 30910 -13330 31040 -13170
rect 29310 -15130 29440 -14970
rect 27710 -16930 27840 -16770
rect 24510 -18730 24640 -18570
rect 26110 -18730 26240 -18570
rect 22910 -20530 23040 -20370
rect 29310 -16930 29440 -16770
rect 27710 -18730 27840 -18570
rect 24510 -20530 24640 -20370
rect 26110 -20530 26240 -20370
rect 29310 -18730 29440 -18570
rect 27710 -20530 27840 -20370
rect 29310 -20530 29440 -20370
rect 32510 -13330 32640 -13170
rect 30910 -15130 31040 -14970
rect 30910 -16930 31040 -16770
rect 32520 -16920 32630 -16770
rect 30910 -18730 31040 -18570
rect 30910 -20530 31040 -20370
rect 16510 -22330 16640 -22170
rect 18110 -22330 18240 -22170
rect 19710 -22330 19840 -22170
rect 21310 -22330 21440 -22170
rect 22910 -22330 23040 -22170
rect 24510 -22330 24640 -22170
rect 26110 -22330 26240 -22170
rect 27710 -22330 27840 -22170
rect 29310 -22330 29440 -22170
rect 30910 -22330 31040 -22170
rect 27720 -22850 27830 -22740
rect 28150 -22870 28370 -22730
rect 28630 -22870 28740 -22740
rect 29000 -22870 29220 -22730
rect 29320 -22850 29430 -22740
rect 30920 -22850 31030 -22740
rect 12420 -23090 12520 -22980
rect 26530 -23160 26710 -22980
rect 1190 -23450 1350 -23270
rect 2790 -23450 2950 -23270
rect 4390 -23450 4550 -23270
rect 5990 -23450 6150 -23270
rect 7590 -23450 7750 -23270
rect 9190 -23450 9350 -23270
rect 23210 -23480 23390 -23300
rect 1630 -24250 1810 -24070
rect 1290 -24650 1470 -24470
rect 430 -26710 610 -26630
rect 430 -27510 610 -27430
rect 430 -28310 610 -28230
rect 430 -29110 610 -29030
rect 2510 -25130 4010 -25070
rect 4710 -25130 6210 -25070
rect 6910 -25130 8410 -25070
rect 9110 -25130 10610 -25070
rect 11310 -25130 12810 -25070
rect 13510 -25130 15010 -25070
rect 15710 -25130 17210 -25070
rect 17910 -25130 19410 -25070
rect 20450 -24250 20630 -24070
rect 20110 -24650 20290 -24470
rect 2510 -25760 2690 -25700
rect 3170 -25760 3350 -25700
rect 3830 -25760 4010 -25700
rect 2510 -25930 4010 -25870
rect 4710 -25760 4890 -25700
rect 5370 -25760 5550 -25700
rect 6030 -25760 6210 -25700
rect 4710 -25930 6210 -25870
rect 6910 -25620 7090 -25560
rect 7570 -25620 7750 -25560
rect 8230 -25620 8410 -25560
rect 6910 -25930 8410 -25870
rect 9110 -25620 9290 -25560
rect 9770 -25620 9950 -25560
rect 10430 -25620 10610 -25560
rect 9110 -25930 10610 -25870
rect 11310 -25620 11490 -25560
rect 11970 -25620 12150 -25560
rect 12630 -25620 12810 -25560
rect 11310 -25930 12810 -25870
rect 13510 -25620 13690 -25560
rect 14170 -25620 14350 -25560
rect 14830 -25620 15010 -25560
rect 13510 -25930 15010 -25870
rect 15710 -25760 15890 -25700
rect 16370 -25760 16550 -25700
rect 17030 -25760 17210 -25700
rect 15710 -25930 17210 -25870
rect 17910 -25760 18090 -25700
rect 18570 -25760 18750 -25700
rect 19230 -25760 19410 -25700
rect 17910 -25930 19410 -25870
rect 2510 -26420 2690 -26360
rect 3170 -26420 3350 -26360
rect 3830 -26420 4010 -26360
rect 4710 -26420 4890 -26360
rect 5370 -26420 5550 -26360
rect 6030 -26420 6210 -26360
rect 4710 -26730 6210 -26670
rect 6910 -26560 7090 -26500
rect 7570 -26560 7750 -26500
rect 8230 -26560 8410 -26500
rect 6910 -26730 8410 -26670
rect 9110 -26560 9290 -26500
rect 9770 -26560 9950 -26500
rect 10430 -26560 10610 -26500
rect 9110 -26730 10610 -26670
rect 11310 -26560 11490 -26500
rect 11970 -26560 12150 -26500
rect 12630 -26560 12810 -26500
rect 11310 -26730 12810 -26670
rect 13510 -26560 13690 -26500
rect 14170 -26560 14350 -26500
rect 14830 -26560 15010 -26500
rect 13510 -26730 15010 -26670
rect 15710 -26420 15890 -26360
rect 16370 -26420 16550 -26360
rect 17030 -26420 17210 -26360
rect 15710 -26730 17210 -26670
rect 17910 -26420 18090 -26360
rect 18570 -26420 18750 -26360
rect 19230 -26420 19410 -26360
rect 2510 -27360 2690 -27300
rect 3170 -27360 3350 -27300
rect 3830 -27360 4010 -27300
rect 4710 -27360 4890 -27300
rect 5370 -27360 5550 -27300
rect 6030 -27360 6210 -27300
rect 4710 -27530 6210 -27470
rect 6910 -27220 7090 -27160
rect 7570 -27220 7750 -27160
rect 8230 -27220 8410 -27160
rect 6910 -27530 8410 -27470
rect 9110 -27220 9290 -27160
rect 9770 -27220 9950 -27160
rect 10430 -27220 10610 -27160
rect 9110 -27530 10610 -27470
rect 11310 -27220 11490 -27160
rect 11970 -27220 12150 -27160
rect 12630 -27220 12810 -27160
rect 11310 -27530 12810 -27470
rect 13510 -27220 13690 -27160
rect 14170 -27220 14350 -27160
rect 14830 -27220 15010 -27160
rect 13510 -27530 15010 -27470
rect 15710 -27360 15890 -27300
rect 16370 -27360 16550 -27300
rect 17030 -27360 17210 -27300
rect 15710 -27530 17210 -27470
rect 17910 -27360 18090 -27300
rect 18570 -27360 18750 -27300
rect 19230 -27360 19410 -27300
rect 2510 -28020 2690 -27960
rect 3170 -28020 3350 -27960
rect 3830 -28020 4010 -27960
rect 4710 -28020 4890 -27960
rect 5370 -28020 5550 -27960
rect 6030 -28020 6210 -27960
rect 4710 -28330 6210 -28270
rect 6910 -28160 7090 -28100
rect 7570 -28160 7750 -28100
rect 8230 -28160 8410 -28100
rect 6910 -28330 8410 -28270
rect 9110 -28160 9290 -28100
rect 9770 -28160 9950 -28100
rect 10430 -28160 10610 -28100
rect 9110 -28330 10610 -28270
rect 11310 -28160 11490 -28100
rect 11970 -28160 12150 -28100
rect 12630 -28160 12810 -28100
rect 11310 -28330 12810 -28270
rect 13510 -28160 13690 -28100
rect 14170 -28160 14350 -28100
rect 14830 -28160 15010 -28100
rect 13510 -28330 15010 -28270
rect 15710 -28020 15890 -27960
rect 16370 -28020 16550 -27960
rect 17030 -28020 17210 -27960
rect 15710 -28330 17210 -28270
rect 17910 -28020 18090 -27960
rect 18570 -28020 18750 -27960
rect 19230 -28020 19410 -27960
rect 2510 -28820 2690 -28760
rect 3170 -28820 3350 -28760
rect 3830 -28820 4010 -28760
rect 4710 -28820 4890 -28760
rect 5370 -28820 5550 -28760
rect 6030 -28820 6210 -28760
rect 4710 -29130 6210 -29070
rect 6910 -28960 7090 -28900
rect 7570 -28960 7750 -28900
rect 8230 -28960 8410 -28900
rect 6910 -29130 8410 -29070
rect 9110 -28960 9290 -28900
rect 9770 -28960 9950 -28900
rect 10430 -28960 10610 -28900
rect 9110 -29130 10610 -29070
rect 11310 -28960 11490 -28900
rect 11970 -28960 12150 -28900
rect 12630 -28960 12810 -28900
rect 11310 -29130 12810 -29070
rect 13510 -28960 13690 -28900
rect 14170 -28960 14350 -28900
rect 14830 -28960 15010 -28900
rect 13510 -29130 15010 -29070
rect 15710 -28820 15890 -28760
rect 16370 -28820 16550 -28760
rect 17030 -28820 17210 -28760
rect 15710 -29130 17210 -29070
rect 17910 -28820 18090 -28760
rect 18570 -28820 18750 -28760
rect 19230 -28820 19410 -28760
rect 23040 -25070 23560 -24820
rect 31560 -23480 31740 -23300
rect 27630 -24250 27810 -24070
rect 28500 -24200 28660 -24040
rect 27400 -24650 27580 -24470
rect 27250 -25070 27430 -24890
rect 21310 -26710 21490 -26630
rect 21310 -27510 21490 -27430
rect 21310 -28310 21490 -28230
rect 21310 -29110 21490 -29030
rect 2510 -29760 2690 -29700
rect 3170 -29760 3350 -29700
rect 3830 -29760 4010 -29700
rect 2510 -29930 4010 -29870
rect 4710 -29760 4890 -29700
rect 5370 -29760 5550 -29700
rect 6030 -29760 6210 -29700
rect 4710 -29930 6210 -29870
rect 6910 -29620 7090 -29560
rect 7570 -29620 7750 -29560
rect 8230 -29620 8410 -29560
rect 6910 -29930 8410 -29870
rect 9110 -29620 9290 -29560
rect 9770 -29620 9950 -29560
rect 10430 -29620 10610 -29560
rect 9110 -29930 10610 -29870
rect 11310 -29620 11490 -29560
rect 11970 -29620 12150 -29560
rect 12630 -29620 12810 -29560
rect 11310 -29930 12810 -29870
rect 13510 -29620 13690 -29560
rect 14170 -29620 14350 -29560
rect 14830 -29620 15010 -29560
rect 13510 -29930 15010 -29870
rect 15710 -29760 15890 -29700
rect 16370 -29760 16550 -29700
rect 17030 -29760 17210 -29700
rect 15710 -29930 17210 -29870
rect 17910 -29760 18090 -29700
rect 18570 -29760 18750 -29700
rect 19230 -29760 19410 -29700
rect 17910 -29930 19410 -29870
rect 2510 -30420 2690 -30360
rect 3170 -30420 3350 -30360
rect 3830 -30420 4010 -30360
rect 2510 -30730 4010 -30670
rect 4710 -30420 4890 -30360
rect 5370 -30420 5550 -30360
rect 6030 -30420 6210 -30360
rect 4710 -30730 6210 -30670
rect 6910 -30560 7090 -30500
rect 7570 -30560 7750 -30500
rect 8230 -30560 8410 -30500
rect 6910 -30730 8410 -30670
rect 9110 -30560 9290 -30500
rect 9770 -30560 9950 -30500
rect 10430 -30560 10610 -30500
rect 9110 -30730 10610 -30670
rect 11310 -30560 11490 -30500
rect 11970 -30560 12150 -30500
rect 12630 -30560 12810 -30500
rect 11310 -30730 12810 -30670
rect 13510 -30560 13690 -30500
rect 14170 -30560 14350 -30500
rect 14830 -30560 15010 -30500
rect 13510 -30730 15010 -30670
rect 15710 -30420 15890 -30360
rect 16370 -30420 16550 -30360
rect 17030 -30420 17210 -30360
rect 15710 -30730 17210 -30670
rect 17910 -30420 18090 -30360
rect 18570 -30420 18750 -30360
rect 19230 -30420 19410 -30360
rect 17910 -30730 19410 -30670
rect 90 -32110 270 -31730
rect 1990 -31830 2110 -31710
rect 2510 -31360 2690 -31300
rect 3170 -31360 3350 -31300
rect 3830 -31360 4010 -31300
rect 4190 -31830 4310 -31710
rect 2210 -32130 2330 -32010
rect 4710 -31360 4890 -31300
rect 5370 -31360 5550 -31300
rect 6030 -31360 6210 -31300
rect 6390 -31830 6510 -31710
rect 4410 -32130 4530 -32010
rect 6910 -31220 7090 -31160
rect 7570 -31220 7750 -31160
rect 8230 -31220 8410 -31160
rect 8590 -31830 8710 -31710
rect 6610 -32130 6730 -32010
rect 9110 -31220 9290 -31160
rect 9770 -31220 9950 -31160
rect 10430 -31220 10610 -31160
rect 10790 -31830 10910 -31710
rect 8810 -32130 8930 -32010
rect 11310 -31220 11490 -31160
rect 11970 -31220 12150 -31160
rect 12630 -31220 12810 -31160
rect 12990 -31830 13110 -31710
rect 11010 -32130 11130 -32010
rect 13510 -31220 13690 -31160
rect 14170 -31220 14350 -31160
rect 14830 -31220 15010 -31160
rect 15190 -31830 15310 -31710
rect 13210 -32130 13330 -32010
rect 15710 -31360 15890 -31300
rect 16370 -31360 16550 -31300
rect 17030 -31360 17210 -31300
rect 17390 -31830 17510 -31710
rect 15410 -32130 15530 -32010
rect 17910 -31360 18090 -31300
rect 18570 -31360 18750 -31300
rect 19230 -31360 19410 -31300
rect 19590 -31830 19710 -31710
rect 17610 -32130 17730 -32010
rect 29380 -24720 29440 -24490
rect 29530 -24870 29590 -24640
rect 28940 -30480 29160 -30410
rect 29070 -30630 29290 -30560
rect 29220 -30780 29440 -30710
rect 29680 -28940 29740 -28720
rect 32510 -20530 32640 -20370
rect 31820 -23850 32000 -23670
rect 29980 -24370 30040 -24140
rect 29830 -29090 29890 -28870
rect 34110 -9730 34240 -9570
rect 35710 -9730 35840 -9570
rect 34110 -11530 34240 -11370
rect 34110 -13330 34240 -13170
rect 35710 -11530 35840 -11370
rect 34120 -16920 34230 -16770
rect 34110 -20530 34240 -20370
rect 32800 -24550 33030 -24480
rect 35710 -13330 35840 -13170
rect 34620 -24280 34770 -24220
rect 35720 -16920 35830 -16770
rect 35710 -20530 35840 -20370
rect 34990 -24280 35130 -24220
rect 35130 -24280 35260 -24220
rect 35260 -24280 35450 -24220
rect 35450 -24280 35570 -24220
rect 35570 -24280 35760 -24220
rect 35760 -24280 35890 -24220
rect 35890 -24280 36080 -24220
rect 36080 -24280 36200 -24220
rect 36200 -24280 36390 -24220
rect 36390 -24280 36520 -24220
rect 36520 -24280 36710 -24220
rect 36710 -24280 36830 -24220
rect 36830 -24280 37020 -24220
rect 34120 -24700 34350 -24630
rect 30290 -24850 30510 -24780
rect 33560 -24850 33790 -24780
rect 34810 -24860 34900 -24660
rect 37130 -24780 37270 -24640
rect 30130 -25170 30190 -24940
rect 29980 -29240 30040 -29020
rect 30130 -29390 30190 -29170
rect 30430 -25320 30490 -25090
rect 30280 -29540 30340 -29320
rect 36030 -27140 36410 -27010
rect 36530 -27140 36910 -27010
rect 36920 -27900 37680 -27540
rect 36920 -28520 37680 -28160
rect 36030 -28780 36270 -28710
rect 35690 -28930 35930 -28860
rect 30430 -29690 30490 -29470
rect 32610 -30480 32794 -30410
rect 32794 -30480 32846 -30410
rect 32846 -30480 32850 -30410
rect 37030 -29080 37270 -29010
rect 36700 -29230 36940 -29160
rect 38030 -29380 38270 -29310
rect 37700 -29530 37940 -29460
rect 33320 -30630 33560 -30560
rect 34320 -30782 34560 -30712
rect 29370 -30930 29590 -30860
rect 35320 -30930 35560 -30860
rect 19810 -32130 19930 -32010
rect 30840 -32440 31240 -31680
rect 38406 -32314 38520 -32180
rect 38320 -32690 38520 -32314
rect 38310 -32910 38530 -32690
<< metal3 >>
rect 36900 12540 38300 12560
rect 36900 12280 36920 12540
rect 38280 12280 38300 12540
rect 36900 12260 38300 12280
rect 2200 12010 2340 12020
rect 2200 12000 2210 12010
rect -360 11990 2210 12000
rect -360 11610 -350 11990
rect -170 11900 2210 11990
rect -170 11610 -160 11900
rect 2200 11890 2210 11900
rect 2330 12000 2340 12010
rect 4400 12010 4540 12020
rect 4400 12000 4410 12010
rect 2330 11900 4410 12000
rect 2330 11890 2340 11900
rect 2200 11880 2340 11890
rect 4400 11890 4410 11900
rect 4530 12000 4540 12010
rect 6600 12010 6740 12020
rect 6600 12000 6610 12010
rect 4530 11900 6610 12000
rect 4530 11890 4540 11900
rect 4400 11880 4540 11890
rect 6600 11890 6610 11900
rect 6730 12000 6740 12010
rect 8800 12010 8940 12020
rect 8800 12000 8810 12010
rect 6730 11900 8810 12000
rect 6730 11890 6740 11900
rect 6600 11880 6740 11890
rect 8800 11890 8810 11900
rect 8930 12000 8940 12010
rect 11000 12010 11140 12020
rect 11000 12000 11010 12010
rect 8930 11900 11010 12000
rect 8930 11890 8940 11900
rect 8800 11880 8940 11890
rect 11000 11890 11010 11900
rect 11130 12000 11140 12010
rect 13200 12010 13340 12020
rect 13200 12000 13210 12010
rect 11130 11900 13210 12000
rect 11130 11890 11140 11900
rect 11000 11880 11140 11890
rect 13200 11890 13210 11900
rect 13330 12000 13340 12010
rect 15400 12010 15540 12020
rect 15400 12000 15410 12010
rect 13330 11900 15410 12000
rect 13330 11890 13340 11900
rect 13200 11880 13340 11890
rect 15400 11890 15410 11900
rect 15530 12000 15540 12010
rect 17600 12010 17740 12020
rect 17600 12000 17610 12010
rect 15530 11900 17610 12000
rect 15530 11890 15540 11900
rect 15400 11880 15540 11890
rect 17600 11890 17610 11900
rect 17730 12000 17740 12010
rect 19800 12010 19940 12020
rect 19800 12000 19810 12010
rect 17730 11900 19810 12000
rect 17730 11890 17740 11900
rect 17600 11880 17740 11890
rect 19800 11890 19810 11900
rect 19930 12000 19940 12010
rect 19930 11900 22160 12000
rect 19930 11890 19940 11900
rect 19800 11880 19940 11890
rect 1980 11710 2120 11720
rect 1980 11700 1990 11710
rect -360 11600 -160 11610
rect 80 11690 1990 11700
rect 80 11310 90 11690
rect 270 11600 1990 11690
rect 270 11310 280 11600
rect 1980 11590 1990 11600
rect 2110 11700 2120 11710
rect 4180 11710 4320 11720
rect 4180 11700 4190 11710
rect 2110 11600 4190 11700
rect 2110 11590 2120 11600
rect 1980 11580 2120 11590
rect 4180 11590 4190 11600
rect 4310 11700 4320 11710
rect 6380 11710 6520 11720
rect 6380 11700 6390 11710
rect 4310 11600 6390 11700
rect 4310 11590 4320 11600
rect 4180 11580 4320 11590
rect 6380 11590 6390 11600
rect 6510 11700 6520 11710
rect 8580 11710 8720 11720
rect 8580 11700 8590 11710
rect 6510 11600 8590 11700
rect 6510 11590 6520 11600
rect 6380 11580 6520 11590
rect 8580 11590 8590 11600
rect 8710 11700 8720 11710
rect 10780 11710 10920 11720
rect 10780 11700 10790 11710
rect 8710 11600 10790 11700
rect 8710 11590 8720 11600
rect 8580 11580 8720 11590
rect 10780 11590 10790 11600
rect 10910 11700 10920 11710
rect 12980 11710 13120 11720
rect 12980 11700 12990 11710
rect 10910 11600 12990 11700
rect 10910 11590 10920 11600
rect 10780 11580 10920 11590
rect 12980 11590 12990 11600
rect 13110 11700 13120 11710
rect 15180 11710 15320 11720
rect 15180 11700 15190 11710
rect 13110 11600 15190 11700
rect 13110 11590 13120 11600
rect 12980 11580 13120 11590
rect 15180 11590 15190 11600
rect 15310 11700 15320 11710
rect 17380 11710 17520 11720
rect 17380 11700 17390 11710
rect 15310 11600 17390 11700
rect 15310 11590 15320 11600
rect 15180 11580 15320 11590
rect 17380 11590 17390 11600
rect 17510 11700 17520 11710
rect 19580 11710 19720 11720
rect 19580 11700 19590 11710
rect 17510 11600 19590 11700
rect 17510 11590 17520 11600
rect 17380 11580 17520 11590
rect 19580 11590 19590 11600
rect 19710 11700 19720 11710
rect 19710 11600 22160 11700
rect 19710 11590 19720 11600
rect 19580 11580 19720 11590
rect 80 11300 280 11310
rect 820 11250 1020 11260
rect 20500 11250 20700 11260
rect 820 11240 830 11250
rect -220 11180 830 11240
rect 820 11170 830 11180
rect 1010 11240 1020 11250
rect 2500 11240 2700 11250
rect 3160 11240 3360 11250
rect 3820 11240 4020 11250
rect 4700 11240 4900 11250
rect 5360 11240 5560 11250
rect 6020 11240 6220 11250
rect 6900 11240 7100 11250
rect 7560 11240 7760 11250
rect 8220 11240 8420 11250
rect 9100 11240 9300 11250
rect 9760 11240 9960 11250
rect 10420 11240 10620 11250
rect 11300 11240 11500 11250
rect 11960 11240 12160 11250
rect 12620 11240 12820 11250
rect 13500 11240 13700 11250
rect 14160 11240 14360 11250
rect 14820 11240 15020 11250
rect 15700 11240 15900 11250
rect 16360 11240 16560 11250
rect 17020 11240 17220 11250
rect 17900 11240 18100 11250
rect 18560 11240 18760 11250
rect 19220 11240 19420 11250
rect 20500 11240 20510 11250
rect 1010 11180 2510 11240
rect 2690 11180 3170 11240
rect 3350 11180 3830 11240
rect 4010 11180 4710 11240
rect 4890 11180 5370 11240
rect 5550 11180 6030 11240
rect 6210 11180 15710 11240
rect 15890 11180 16370 11240
rect 16550 11180 17030 11240
rect 17210 11180 17910 11240
rect 18090 11180 18570 11240
rect 18750 11180 19230 11240
rect 19410 11180 20510 11240
rect 1010 11170 1020 11180
rect 2500 11170 2700 11180
rect 3160 11170 3360 11180
rect 3820 11170 4020 11180
rect 4700 11170 4900 11180
rect 5360 11170 5560 11180
rect 6020 11170 6220 11180
rect 6900 11170 7100 11180
rect 7560 11170 7760 11180
rect 8220 11170 8420 11180
rect 9100 11170 9300 11180
rect 9760 11170 9960 11180
rect 10420 11170 10620 11180
rect 11300 11170 11500 11180
rect 11960 11170 12160 11180
rect 12620 11170 12820 11180
rect 13500 11170 13700 11180
rect 14160 11170 14360 11180
rect 14820 11170 15020 11180
rect 15700 11170 15900 11180
rect 16360 11170 16560 11180
rect 17020 11170 17220 11180
rect 17900 11170 18100 11180
rect 18560 11170 18760 11180
rect 19220 11170 19420 11180
rect 20500 11170 20510 11180
rect 20690 11240 20700 11250
rect 20690 11180 22180 11240
rect 20690 11170 20700 11180
rect 820 11160 1020 11170
rect 20500 11160 20700 11170
rect 1220 11110 1420 11120
rect 20900 11110 21100 11120
rect 1220 11100 1230 11110
rect -220 11040 1230 11100
rect 1220 11030 1230 11040
rect 1410 11100 1420 11110
rect 2500 11100 2700 11110
rect 3160 11100 3360 11110
rect 3820 11100 4020 11110
rect 4700 11100 4900 11110
rect 5360 11100 5560 11110
rect 6020 11100 6220 11110
rect 6900 11100 7100 11110
rect 7560 11100 7760 11110
rect 8220 11100 8420 11110
rect 9100 11100 9300 11110
rect 9760 11100 9960 11110
rect 10420 11100 10620 11110
rect 11300 11100 11500 11110
rect 11960 11100 12160 11110
rect 12620 11100 12820 11110
rect 13500 11100 13700 11110
rect 14160 11100 14360 11110
rect 14820 11100 15020 11110
rect 15700 11100 15900 11110
rect 16360 11100 16560 11110
rect 17020 11100 17220 11110
rect 17900 11100 18100 11110
rect 18560 11100 18760 11110
rect 19220 11100 19420 11110
rect 20900 11100 20910 11110
rect 1410 11040 6910 11100
rect 7090 11040 7570 11100
rect 7750 11040 8230 11100
rect 8410 11040 9110 11100
rect 9290 11040 9770 11100
rect 9950 11040 10430 11100
rect 10610 11040 11310 11100
rect 11490 11040 11970 11100
rect 12150 11040 12630 11100
rect 12810 11040 13510 11100
rect 13690 11040 14170 11100
rect 14350 11040 14830 11100
rect 15010 11040 20910 11100
rect 1410 11030 1420 11040
rect 2500 11030 2700 11040
rect 3160 11030 3360 11040
rect 3820 11030 4020 11040
rect 4700 11030 4900 11040
rect 5360 11030 5560 11040
rect 6020 11030 6220 11040
rect 6900 11030 7100 11040
rect 7560 11030 7760 11040
rect 8220 11030 8420 11040
rect 9100 11030 9300 11040
rect 9760 11030 9960 11040
rect 10420 11030 10620 11040
rect 11300 11030 11500 11040
rect 11960 11030 12160 11040
rect 12620 11030 12820 11040
rect 13500 11030 13700 11040
rect 14160 11030 14360 11040
rect 14820 11030 15020 11040
rect 15700 11030 15900 11040
rect 16360 11030 16560 11040
rect 17020 11030 17220 11040
rect 17900 11030 18100 11040
rect 18560 11030 18760 11040
rect 19220 11030 19420 11040
rect 20900 11030 20910 11040
rect 21090 11100 21100 11110
rect 21090 11040 22180 11100
rect 30302 11060 31214 11082
rect 21090 11030 21100 11040
rect 1220 11020 1420 11030
rect 20900 11020 21100 11030
rect -110 10940 30 10960
rect -110 10690 -80 10940
rect 0 10690 30 10940
rect -110 10660 30 10690
rect 2090 10940 2230 10960
rect 2090 10690 2120 10940
rect 2200 10690 2230 10940
rect 2090 10660 2230 10690
rect 4290 10940 4430 10960
rect 4290 10690 4320 10940
rect 4400 10690 4430 10940
rect 4290 10660 4430 10690
rect 6490 10940 6630 10960
rect 6490 10690 6520 10940
rect 6600 10690 6630 10940
rect 6490 10660 6630 10690
rect 8690 10940 8830 10960
rect 8690 10690 8720 10940
rect 8800 10690 8830 10940
rect 8690 10660 8830 10690
rect 10890 10940 11030 10960
rect 10890 10690 10920 10940
rect 11000 10690 11030 10940
rect 10890 10660 11030 10690
rect 13090 10940 13230 10960
rect 13090 10690 13120 10940
rect 13200 10690 13230 10940
rect 13090 10660 13230 10690
rect 15290 10940 15430 10960
rect 15290 10690 15320 10940
rect 15400 10690 15430 10940
rect 15290 10660 15430 10690
rect 17490 10940 17630 10960
rect 17490 10690 17520 10940
rect 17600 10690 17630 10940
rect 17490 10660 17630 10690
rect 19690 10940 19830 10960
rect 19690 10690 19720 10940
rect 19800 10690 19830 10940
rect 19690 10660 19830 10690
rect 21890 10940 22030 10960
rect 21890 10690 21920 10940
rect 22000 10690 22030 10940
rect 30302 10932 30326 11060
rect 30682 10934 30824 11060
rect 31194 10934 31214 11060
rect 30682 10932 31214 10934
rect 30302 10912 31214 10932
rect 36880 11010 37060 11020
rect 36880 10850 36890 11010
rect 37050 10960 37060 11010
rect 37180 11010 37350 11020
rect 37180 10960 37190 11010
rect 37050 10900 37190 10960
rect 37050 10850 37060 10900
rect 37180 10860 37190 10900
rect 37340 10860 37350 11010
rect 37180 10850 37350 10860
rect 37980 10960 38130 10970
rect 36880 10840 37060 10850
rect 29270 10790 29520 10800
rect 33510 10790 33770 10800
rect 29200 10720 29280 10790
rect 29510 10720 33520 10790
rect 33760 10720 33770 10790
rect 37980 10780 37990 10960
rect 38120 10920 38130 10960
rect 38120 10820 39500 10920
rect 38120 10780 38130 10820
rect 37980 10770 38130 10780
rect 29270 10710 29520 10720
rect 33510 10710 33770 10720
rect 37080 10760 37260 10770
rect 21890 10660 22030 10690
rect 28950 10640 29200 10650
rect 2500 10610 4020 10620
rect 1620 10590 1820 10600
rect 1620 10580 1630 10590
rect 1600 10520 1630 10580
rect 1620 10510 1630 10520
rect 1810 10580 1820 10590
rect 2500 10580 2510 10610
rect 1810 10550 2510 10580
rect 4010 10580 4020 10610
rect 4700 10610 6220 10620
rect 4700 10580 4710 10610
rect 4010 10550 4710 10580
rect 6210 10580 6220 10610
rect 6900 10610 8420 10620
rect 6900 10580 6910 10610
rect 6210 10550 6910 10580
rect 8410 10580 8420 10610
rect 9100 10610 10620 10620
rect 9100 10580 9110 10610
rect 8410 10550 9110 10580
rect 10610 10580 10620 10610
rect 11300 10610 12820 10620
rect 11300 10580 11310 10610
rect 10610 10550 11310 10580
rect 12810 10580 12820 10610
rect 13500 10610 15020 10620
rect 13500 10580 13510 10610
rect 12810 10550 13510 10580
rect 15010 10580 15020 10610
rect 15700 10610 17220 10620
rect 15700 10580 15710 10610
rect 15010 10550 15710 10580
rect 17210 10580 17220 10610
rect 17900 10610 19420 10620
rect 17900 10580 17910 10610
rect 17210 10550 17910 10580
rect 19410 10580 19420 10610
rect 20100 10590 20300 10600
rect 20100 10580 20110 10590
rect 19410 10550 20110 10580
rect 1810 10520 20110 10550
rect 1810 10510 1820 10520
rect 1620 10500 1820 10510
rect 20100 10510 20110 10520
rect 20290 10580 20300 10590
rect 20290 10520 20320 10580
rect 28950 10570 28960 10640
rect 29190 10630 29200 10640
rect 32470 10630 32730 10640
rect 29190 10570 32480 10630
rect 28950 10560 32480 10570
rect 32720 10560 33768 10630
rect 37080 10600 37090 10760
rect 37250 10710 37260 10760
rect 37600 10750 37770 10760
rect 37600 10710 37610 10750
rect 37250 10650 37610 10710
rect 37250 10600 37260 10650
rect 37080 10590 37260 10600
rect 37600 10600 37610 10650
rect 37760 10600 37770 10750
rect 37600 10590 37770 10600
rect 32470 10550 32730 10560
rect 20290 10510 20300 10520
rect 20100 10500 20300 10510
rect 31670 10490 31930 10500
rect 28860 10480 31680 10490
rect 820 10450 1020 10460
rect 20500 10450 20700 10460
rect 820 10440 830 10450
rect -220 10380 830 10440
rect 820 10370 830 10380
rect 1010 10440 1020 10450
rect 2500 10440 2700 10450
rect 3160 10440 3360 10450
rect 3820 10440 4020 10450
rect 4700 10440 4900 10450
rect 5360 10440 5560 10450
rect 6020 10440 6220 10450
rect 6900 10440 7100 10450
rect 7560 10440 7760 10450
rect 8220 10440 8420 10450
rect 9100 10440 9300 10450
rect 9760 10440 9960 10450
rect 10420 10440 10620 10450
rect 11300 10440 11500 10450
rect 11960 10440 12160 10450
rect 12620 10440 12820 10450
rect 13500 10440 13700 10450
rect 14160 10440 14360 10450
rect 14820 10440 15020 10450
rect 15700 10440 15900 10450
rect 16360 10440 16560 10450
rect 17020 10440 17220 10450
rect 17900 10440 18100 10450
rect 18560 10440 18760 10450
rect 19220 10440 19420 10450
rect 20500 10440 20510 10450
rect 1010 10380 6910 10440
rect 7090 10380 7570 10440
rect 7750 10380 8230 10440
rect 8410 10380 9110 10440
rect 9290 10380 9770 10440
rect 9950 10380 10430 10440
rect 10610 10380 11310 10440
rect 11490 10380 11970 10440
rect 12150 10380 12630 10440
rect 12810 10380 13510 10440
rect 13690 10380 14170 10440
rect 14350 10380 14830 10440
rect 15010 10380 20510 10440
rect 1010 10370 1020 10380
rect 2500 10370 2700 10380
rect 3160 10370 3360 10380
rect 3820 10370 4020 10380
rect 4700 10370 4900 10380
rect 5360 10370 5560 10380
rect 6020 10370 6220 10380
rect 6900 10370 7100 10380
rect 7560 10370 7760 10380
rect 8220 10370 8420 10380
rect 9100 10370 9300 10380
rect 9760 10370 9960 10380
rect 10420 10370 10620 10380
rect 11300 10370 11500 10380
rect 11960 10370 12160 10380
rect 12620 10370 12820 10380
rect 13500 10370 13700 10380
rect 14160 10370 14360 10380
rect 14820 10370 15020 10380
rect 15700 10370 15900 10380
rect 16360 10370 16560 10380
rect 17020 10370 17220 10380
rect 17900 10370 18100 10380
rect 18560 10370 18760 10380
rect 19220 10370 19420 10380
rect 20500 10370 20510 10380
rect 20690 10440 20700 10450
rect 20690 10380 22180 10440
rect 20690 10370 20700 10380
rect 820 10360 1020 10370
rect 20500 10360 20700 10370
rect 1220 10310 1420 10320
rect 20900 10310 21100 10320
rect 1220 10300 1230 10310
rect -220 10240 1230 10300
rect 1220 10230 1230 10240
rect 1410 10300 1420 10310
rect 2500 10300 2700 10310
rect 3160 10300 3360 10310
rect 3820 10300 4020 10310
rect 4700 10300 4900 10310
rect 5360 10300 5560 10310
rect 6020 10300 6220 10310
rect 6900 10300 7100 10310
rect 7560 10300 7760 10310
rect 8220 10300 8420 10310
rect 9100 10300 9300 10310
rect 9760 10300 9960 10310
rect 10420 10300 10620 10310
rect 11300 10300 11500 10310
rect 11960 10300 12160 10310
rect 12620 10300 12820 10310
rect 13500 10300 13700 10310
rect 14160 10300 14360 10310
rect 14820 10300 15020 10310
rect 15700 10300 15900 10310
rect 16360 10300 16560 10310
rect 17020 10300 17220 10310
rect 17900 10300 18100 10310
rect 18560 10300 18760 10310
rect 19220 10300 19420 10310
rect 20900 10300 20910 10310
rect 1410 10240 2510 10300
rect 2690 10240 3170 10300
rect 3350 10240 3830 10300
rect 4010 10240 4710 10300
rect 4890 10240 5370 10300
rect 5550 10240 6030 10300
rect 6210 10240 15710 10300
rect 15890 10240 16370 10300
rect 16550 10240 17030 10300
rect 17210 10240 17910 10300
rect 18090 10240 18570 10300
rect 18750 10240 19230 10300
rect 19410 10240 20910 10300
rect 1410 10230 1420 10240
rect 2500 10230 2700 10240
rect 3160 10230 3360 10240
rect 3820 10230 4020 10240
rect 4700 10230 4900 10240
rect 5360 10230 5560 10240
rect 6020 10230 6220 10240
rect 6900 10230 7100 10240
rect 7560 10230 7760 10240
rect 8220 10230 8420 10240
rect 9100 10230 9300 10240
rect 9760 10230 9960 10240
rect 10420 10230 10620 10240
rect 11300 10230 11500 10240
rect 11960 10230 12160 10240
rect 12620 10230 12820 10240
rect 13500 10230 13700 10240
rect 14160 10230 14360 10240
rect 14820 10230 15020 10240
rect 15700 10230 15900 10240
rect 16360 10230 16560 10240
rect 17020 10230 17220 10240
rect 17900 10230 18100 10240
rect 18560 10230 18760 10240
rect 19220 10230 19420 10240
rect 20900 10230 20910 10240
rect 21090 10300 21100 10310
rect 28860 10310 28870 10480
rect 28930 10420 31680 10480
rect 31920 10420 33768 10490
rect 28930 10310 28940 10420
rect 31670 10410 31930 10420
rect 31320 10350 31580 10360
rect 28860 10300 28940 10310
rect 29010 10340 31330 10350
rect 21090 10240 22180 10300
rect 21090 10230 21100 10240
rect 1220 10220 1420 10230
rect 20900 10220 21100 10230
rect 29010 10170 29020 10340
rect 29080 10280 31330 10340
rect 31570 10280 33768 10350
rect 29080 10170 29090 10280
rect 31320 10270 31580 10280
rect 29010 10160 29090 10170
rect -110 10140 30 10160
rect -110 9890 -80 10140
rect 0 9890 30 10140
rect -110 9860 30 9890
rect 2090 10140 2230 10160
rect 2090 9890 2120 10140
rect 2200 9890 2230 10140
rect 2090 9860 2230 9890
rect 4290 10140 4430 10160
rect 4290 9890 4320 10140
rect 4400 9890 4430 10140
rect 4290 9860 4430 9890
rect 6490 10140 6630 10160
rect 6490 9890 6520 10140
rect 6600 9890 6630 10140
rect 6490 9860 6630 9890
rect 8690 10140 8830 10160
rect 8690 9890 8720 10140
rect 8800 9890 8830 10140
rect 8690 9860 8830 9890
rect 10890 10140 11030 10160
rect 10890 9890 10920 10140
rect 11000 9890 11030 10140
rect 10890 9860 11030 9890
rect 13090 10140 13230 10160
rect 13090 9890 13120 10140
rect 13200 9890 13230 10140
rect 13090 9860 13230 9890
rect 15290 10140 15430 10160
rect 15290 9890 15320 10140
rect 15400 9890 15430 10140
rect 15290 9860 15430 9890
rect 17490 10140 17630 10160
rect 17490 9890 17520 10140
rect 17600 9890 17630 10140
rect 17490 9860 17630 9890
rect 19690 10140 19830 10160
rect 19690 9890 19720 10140
rect 19800 9890 19830 10140
rect 19690 9860 19830 9890
rect 21890 10140 22030 10160
rect 21890 9890 21920 10140
rect 22000 9890 22030 10140
rect 21890 9860 22030 9890
rect 2500 9810 4020 9820
rect 1620 9790 1820 9800
rect 1620 9780 1630 9790
rect 1600 9720 1630 9780
rect 1620 9710 1630 9720
rect 1810 9780 1820 9790
rect 2500 9780 2510 9810
rect 1810 9750 2510 9780
rect 4010 9780 4020 9810
rect 4700 9810 6220 9820
rect 4700 9780 4710 9810
rect 4010 9750 4710 9780
rect 6210 9780 6220 9810
rect 6900 9810 8420 9820
rect 6900 9780 6910 9810
rect 6210 9750 6910 9780
rect 8410 9780 8420 9810
rect 9100 9810 10620 9820
rect 9100 9780 9110 9810
rect 8410 9750 9110 9780
rect 10610 9780 10620 9810
rect 11300 9810 12820 9820
rect 11300 9780 11310 9810
rect 10610 9750 11310 9780
rect 12810 9780 12820 9810
rect 13500 9810 15020 9820
rect 13500 9780 13510 9810
rect 12810 9750 13510 9780
rect 15010 9780 15020 9810
rect 15700 9810 17220 9820
rect 15700 9780 15710 9810
rect 15010 9750 15710 9780
rect 17210 9780 17220 9810
rect 17900 9810 19420 9820
rect 17900 9780 17910 9810
rect 17210 9750 17910 9780
rect 19410 9780 19420 9810
rect 20100 9790 20300 9800
rect 20100 9780 20110 9790
rect 19410 9750 20110 9780
rect 1810 9720 20110 9750
rect 1810 9710 1820 9720
rect 1620 9700 1820 9710
rect 20100 9710 20110 9720
rect 20290 9780 20300 9790
rect 20290 9720 20320 9780
rect 20290 9710 20300 9720
rect 20100 9700 20300 9710
rect 820 9650 1020 9660
rect 20500 9650 20700 9660
rect 820 9640 830 9650
rect -220 9580 830 9640
rect 820 9570 830 9580
rect 1010 9640 1020 9650
rect 2500 9640 2700 9650
rect 3160 9640 3360 9650
rect 3820 9640 4020 9650
rect 4700 9640 4900 9650
rect 5360 9640 5560 9650
rect 6020 9640 6220 9650
rect 6900 9640 7100 9650
rect 7560 9640 7760 9650
rect 8220 9640 8420 9650
rect 9100 9640 9300 9650
rect 9760 9640 9960 9650
rect 10420 9640 10620 9650
rect 11300 9640 11500 9650
rect 11960 9640 12160 9650
rect 12620 9640 12820 9650
rect 13500 9640 13700 9650
rect 14160 9640 14360 9650
rect 14820 9640 15020 9650
rect 15700 9640 15900 9650
rect 16360 9640 16560 9650
rect 17020 9640 17220 9650
rect 17900 9640 18100 9650
rect 18560 9640 18760 9650
rect 19220 9640 19420 9650
rect 20500 9640 20510 9650
rect 1010 9580 2510 9640
rect 2690 9580 3170 9640
rect 3350 9580 3830 9640
rect 4010 9580 4710 9640
rect 4890 9580 5370 9640
rect 5550 9580 6030 9640
rect 6210 9580 15710 9640
rect 15890 9580 16370 9640
rect 16550 9580 17030 9640
rect 17210 9580 17910 9640
rect 18090 9580 18570 9640
rect 18750 9580 19230 9640
rect 19410 9580 20510 9640
rect 1010 9570 1020 9580
rect 2500 9570 2700 9580
rect 3160 9570 3360 9580
rect 3820 9570 4020 9580
rect 4700 9570 4900 9580
rect 5360 9570 5560 9580
rect 6020 9570 6220 9580
rect 6900 9570 7100 9580
rect 7560 9570 7760 9580
rect 8220 9570 8420 9580
rect 9100 9570 9300 9580
rect 9760 9570 9960 9580
rect 10420 9570 10620 9580
rect 11300 9570 11500 9580
rect 11960 9570 12160 9580
rect 12620 9570 12820 9580
rect 13500 9570 13700 9580
rect 14160 9570 14360 9580
rect 14820 9570 15020 9580
rect 15700 9570 15900 9580
rect 16360 9570 16560 9580
rect 17020 9570 17220 9580
rect 17900 9570 18100 9580
rect 18560 9570 18760 9580
rect 19220 9570 19420 9580
rect 20500 9570 20510 9580
rect 20690 9640 20700 9650
rect 20690 9580 22180 9640
rect 20690 9570 20700 9580
rect 820 9560 1020 9570
rect 20500 9560 20700 9570
rect 1220 9510 1420 9520
rect 20900 9510 21100 9520
rect 1220 9500 1230 9510
rect -220 9440 1230 9500
rect 1220 9430 1230 9440
rect 1410 9500 1420 9510
rect 2500 9500 2700 9510
rect 3160 9500 3360 9510
rect 3820 9500 4020 9510
rect 4700 9500 4900 9510
rect 5360 9500 5560 9510
rect 6020 9500 6220 9510
rect 6900 9500 7100 9510
rect 7560 9500 7760 9510
rect 8220 9500 8420 9510
rect 9100 9500 9300 9510
rect 9760 9500 9960 9510
rect 10420 9500 10620 9510
rect 11300 9500 11500 9510
rect 11960 9500 12160 9510
rect 12620 9500 12820 9510
rect 13500 9500 13700 9510
rect 14160 9500 14360 9510
rect 14820 9500 15020 9510
rect 15700 9500 15900 9510
rect 16360 9500 16560 9510
rect 17020 9500 17220 9510
rect 17900 9500 18100 9510
rect 18560 9500 18760 9510
rect 19220 9500 19420 9510
rect 20900 9500 20910 9510
rect 1410 9440 6910 9500
rect 7090 9440 7570 9500
rect 7750 9440 8230 9500
rect 8410 9440 9110 9500
rect 9290 9440 9770 9500
rect 9950 9440 10430 9500
rect 10610 9440 11310 9500
rect 11490 9440 11970 9500
rect 12150 9440 12630 9500
rect 12810 9440 13510 9500
rect 13690 9440 14170 9500
rect 14350 9440 14830 9500
rect 15010 9440 20910 9500
rect 1410 9430 1420 9440
rect 2500 9430 2700 9440
rect 3160 9430 3360 9440
rect 3820 9430 4020 9440
rect 4700 9430 4900 9440
rect 5360 9430 5560 9440
rect 6020 9430 6220 9440
rect 6900 9430 7100 9440
rect 7560 9430 7760 9440
rect 8220 9430 8420 9440
rect 9100 9430 9300 9440
rect 9760 9430 9960 9440
rect 10420 9430 10620 9440
rect 11300 9430 11500 9440
rect 11960 9430 12160 9440
rect 12620 9430 12820 9440
rect 13500 9430 13700 9440
rect 14160 9430 14360 9440
rect 14820 9430 15020 9440
rect 15700 9430 15900 9440
rect 16360 9430 16560 9440
rect 17020 9430 17220 9440
rect 17900 9430 18100 9440
rect 18560 9430 18760 9440
rect 19220 9430 19420 9440
rect 20900 9430 20910 9440
rect 21090 9500 21100 9510
rect 21090 9440 22180 9500
rect 21090 9430 21100 9440
rect 1220 9420 1420 9430
rect 20900 9420 21100 9430
rect -110 9340 30 9360
rect -110 9090 -80 9340
rect 0 9090 30 9340
rect -110 9060 30 9090
rect 2090 9340 2230 9360
rect 2090 9090 2120 9340
rect 2200 9090 2230 9340
rect 2090 9060 2230 9090
rect 4290 9340 4430 9360
rect 4290 9090 4320 9340
rect 4400 9090 4430 9340
rect 4290 9060 4430 9090
rect 6490 9340 6630 9360
rect 6490 9090 6520 9340
rect 6600 9090 6630 9340
rect 6490 9060 6630 9090
rect 8690 9340 8830 9360
rect 8690 9090 8720 9340
rect 8800 9090 8830 9340
rect 8690 9060 8830 9090
rect 10890 9340 11030 9360
rect 10890 9090 10920 9340
rect 11000 9090 11030 9340
rect 10890 9060 11030 9090
rect 13090 9340 13230 9360
rect 13090 9090 13120 9340
rect 13200 9090 13230 9340
rect 13090 9060 13230 9090
rect 15290 9340 15430 9360
rect 15290 9090 15320 9340
rect 15400 9090 15430 9340
rect 15290 9060 15430 9090
rect 17490 9340 17630 9360
rect 17490 9090 17520 9340
rect 17600 9090 17630 9340
rect 17490 9060 17630 9090
rect 19690 9340 19830 9360
rect 19690 9090 19720 9340
rect 19800 9090 19830 9340
rect 19690 9060 19830 9090
rect 21890 9340 22030 9360
rect 21890 9090 21920 9340
rect 22000 9090 22030 9340
rect 21890 9060 22030 9090
rect 4700 9010 6220 9020
rect 420 8990 620 9000
rect 420 8910 430 8990
rect 610 8910 620 8990
rect 1620 8990 1820 9000
rect 1620 8980 1630 8990
rect 1600 8920 1630 8980
rect 420 8900 620 8910
rect 1620 8910 1630 8920
rect 1810 8980 1820 8990
rect 4700 8980 4710 9010
rect 1810 8950 4710 8980
rect 6210 8980 6220 9010
rect 6900 9010 8420 9020
rect 6900 8980 6910 9010
rect 6210 8950 6910 8980
rect 8410 8980 8420 9010
rect 9100 9010 10620 9020
rect 9100 8980 9110 9010
rect 8410 8950 9110 8980
rect 10610 8980 10620 9010
rect 11300 9010 12820 9020
rect 11300 8980 11310 9010
rect 10610 8950 11310 8980
rect 12810 8980 12820 9010
rect 13500 9010 15020 9020
rect 13500 8980 13510 9010
rect 12810 8950 13510 8980
rect 15010 8980 15020 9010
rect 15700 9010 17220 9020
rect 15700 8980 15710 9010
rect 15010 8950 15710 8980
rect 17210 8980 17220 9010
rect 20100 8990 20300 9000
rect 20100 8980 20110 8990
rect 17210 8950 20110 8980
rect 1810 8920 20110 8950
rect 1810 8910 1820 8920
rect 1620 8900 1820 8910
rect 20100 8910 20110 8920
rect 20290 8980 20300 8990
rect 21300 8990 21500 9000
rect 20290 8920 20320 8980
rect 20290 8910 20300 8920
rect 20100 8900 20300 8910
rect 21300 8910 21310 8990
rect 21490 8910 21500 8990
rect 21300 8900 21500 8910
rect 820 8850 1020 8860
rect 20500 8850 20700 8860
rect 820 8840 830 8850
rect -220 8780 830 8840
rect 820 8770 830 8780
rect 1010 8840 1020 8850
rect 2500 8840 2700 8850
rect 3160 8840 3360 8850
rect 3820 8840 4020 8850
rect 4700 8840 4900 8850
rect 5360 8840 5560 8850
rect 6020 8840 6220 8850
rect 6900 8840 7100 8850
rect 7560 8840 7760 8850
rect 8220 8840 8420 8850
rect 9100 8840 9300 8850
rect 9760 8840 9960 8850
rect 10420 8840 10620 8850
rect 11300 8840 11500 8850
rect 11960 8840 12160 8850
rect 12620 8840 12820 8850
rect 13500 8840 13700 8850
rect 14160 8840 14360 8850
rect 14820 8840 15020 8850
rect 15700 8840 15900 8850
rect 16360 8840 16560 8850
rect 17020 8840 17220 8850
rect 17900 8840 18100 8850
rect 18560 8840 18760 8850
rect 19220 8840 19420 8850
rect 20500 8840 20510 8850
rect 1010 8780 6910 8840
rect 7090 8780 7570 8840
rect 7750 8780 8230 8840
rect 8410 8780 9110 8840
rect 9290 8780 9770 8840
rect 9950 8780 10430 8840
rect 10610 8780 11310 8840
rect 11490 8780 11970 8840
rect 12150 8780 12630 8840
rect 12810 8780 13510 8840
rect 13690 8780 14170 8840
rect 14350 8780 14830 8840
rect 15010 8780 20510 8840
rect 1010 8770 1020 8780
rect 2500 8770 2700 8780
rect 3160 8770 3360 8780
rect 3820 8770 4020 8780
rect 4700 8770 4900 8780
rect 5360 8770 5560 8780
rect 6020 8770 6220 8780
rect 6900 8770 7100 8780
rect 7560 8770 7760 8780
rect 8220 8770 8420 8780
rect 9100 8770 9300 8780
rect 9760 8770 9960 8780
rect 10420 8770 10620 8780
rect 11300 8770 11500 8780
rect 11960 8770 12160 8780
rect 12620 8770 12820 8780
rect 13500 8770 13700 8780
rect 14160 8770 14360 8780
rect 14820 8770 15020 8780
rect 15700 8770 15900 8780
rect 16360 8770 16560 8780
rect 17020 8770 17220 8780
rect 17900 8770 18100 8780
rect 18560 8770 18760 8780
rect 19220 8770 19420 8780
rect 20500 8770 20510 8780
rect 20690 8840 20700 8850
rect 20690 8780 22180 8840
rect 20690 8770 20700 8780
rect 820 8760 1020 8770
rect 20500 8760 20700 8770
rect 1220 8710 1420 8720
rect 20900 8710 21100 8720
rect 1220 8700 1230 8710
rect -220 8640 1230 8700
rect 1220 8630 1230 8640
rect 1410 8700 1420 8710
rect 2500 8700 2700 8710
rect 3160 8700 3360 8710
rect 3820 8700 4020 8710
rect 4700 8700 4900 8710
rect 5360 8700 5560 8710
rect 6020 8700 6220 8710
rect 6900 8700 7100 8710
rect 7560 8700 7760 8710
rect 8220 8700 8420 8710
rect 9100 8700 9300 8710
rect 9760 8700 9960 8710
rect 10420 8700 10620 8710
rect 11300 8700 11500 8710
rect 11960 8700 12160 8710
rect 12620 8700 12820 8710
rect 13500 8700 13700 8710
rect 14160 8700 14360 8710
rect 14820 8700 15020 8710
rect 15700 8700 15900 8710
rect 16360 8700 16560 8710
rect 17020 8700 17220 8710
rect 17900 8700 18100 8710
rect 18560 8700 18760 8710
rect 19220 8700 19420 8710
rect 20900 8700 20910 8710
rect 1410 8640 2510 8700
rect 2690 8640 3170 8700
rect 3350 8640 3830 8700
rect 4010 8640 4710 8700
rect 4890 8640 5370 8700
rect 5550 8640 6030 8700
rect 6210 8640 15710 8700
rect 15890 8640 16370 8700
rect 16550 8640 17030 8700
rect 17210 8640 17910 8700
rect 18090 8640 18570 8700
rect 18750 8640 19230 8700
rect 19410 8640 20910 8700
rect 1410 8630 1420 8640
rect 2500 8630 2700 8640
rect 3160 8630 3360 8640
rect 3820 8630 4020 8640
rect 4700 8630 4900 8640
rect 5360 8630 5560 8640
rect 6020 8630 6220 8640
rect 6900 8630 7100 8640
rect 7560 8630 7760 8640
rect 8220 8630 8420 8640
rect 9100 8630 9300 8640
rect 9760 8630 9960 8640
rect 10420 8630 10620 8640
rect 11300 8630 11500 8640
rect 11960 8630 12160 8640
rect 12620 8630 12820 8640
rect 13500 8630 13700 8640
rect 14160 8630 14360 8640
rect 14820 8630 15020 8640
rect 15700 8630 15900 8640
rect 16360 8630 16560 8640
rect 17020 8630 17220 8640
rect 17900 8630 18100 8640
rect 18560 8630 18760 8640
rect 19220 8630 19420 8640
rect 20900 8630 20910 8640
rect 21090 8700 21100 8710
rect 21090 8640 22180 8700
rect 21090 8630 21100 8640
rect 1220 8620 1420 8630
rect 20900 8620 21100 8630
rect -110 8540 30 8560
rect -110 8290 -80 8540
rect 0 8290 30 8540
rect -110 8260 30 8290
rect 2090 8540 2230 8560
rect 2090 8290 2120 8540
rect 2200 8290 2230 8540
rect 2090 8260 2230 8290
rect 4290 8540 4430 8560
rect 4290 8290 4320 8540
rect 4400 8290 4430 8540
rect 4290 8260 4430 8290
rect 6490 8540 6630 8560
rect 6490 8290 6520 8540
rect 6600 8290 6630 8540
rect 6490 8260 6630 8290
rect 8690 8540 8830 8560
rect 8690 8290 8720 8540
rect 8800 8290 8830 8540
rect 8690 8260 8830 8290
rect 10890 8540 11030 8560
rect 10890 8290 10920 8540
rect 11000 8290 11030 8540
rect 10890 8260 11030 8290
rect 13090 8540 13230 8560
rect 13090 8290 13120 8540
rect 13200 8290 13230 8540
rect 13090 8260 13230 8290
rect 15290 8540 15430 8560
rect 15290 8290 15320 8540
rect 15400 8290 15430 8540
rect 15290 8260 15430 8290
rect 17490 8540 17630 8560
rect 17490 8290 17520 8540
rect 17600 8290 17630 8540
rect 17490 8260 17630 8290
rect 19690 8540 19830 8560
rect 19690 8290 19720 8540
rect 19800 8290 19830 8540
rect 19690 8260 19830 8290
rect 21890 8540 22030 8560
rect 21890 8290 21920 8540
rect 22000 8290 22030 8540
rect 21890 8260 22030 8290
rect 30510 8290 30650 8300
rect 4700 8210 6220 8220
rect 420 8190 620 8200
rect 420 8110 430 8190
rect 610 8110 620 8190
rect 1620 8190 1820 8200
rect 1620 8180 1630 8190
rect 1600 8120 1630 8180
rect 420 8100 620 8110
rect 1620 8110 1630 8120
rect 1810 8180 1820 8190
rect 4700 8180 4710 8210
rect 1810 8150 4710 8180
rect 6210 8180 6220 8210
rect 6900 8210 8420 8220
rect 6900 8180 6910 8210
rect 6210 8150 6910 8180
rect 8410 8180 8420 8210
rect 9100 8210 10620 8220
rect 9100 8180 9110 8210
rect 8410 8150 9110 8180
rect 10610 8180 10620 8210
rect 11300 8210 12820 8220
rect 11300 8180 11310 8210
rect 10610 8150 11310 8180
rect 12810 8180 12820 8210
rect 13500 8210 15020 8220
rect 13500 8180 13510 8210
rect 12810 8150 13510 8180
rect 15010 8180 15020 8210
rect 15700 8210 17220 8220
rect 15700 8180 15710 8210
rect 15010 8150 15710 8180
rect 17210 8180 17220 8210
rect 20100 8190 20300 8200
rect 20100 8180 20110 8190
rect 17210 8150 20110 8180
rect 1810 8120 20110 8150
rect 1810 8110 1820 8120
rect 1620 8100 1820 8110
rect 20100 8110 20110 8120
rect 20290 8180 20300 8190
rect 21300 8190 21500 8200
rect 20290 8120 20320 8180
rect 20290 8110 20300 8120
rect 20100 8100 20300 8110
rect 21300 8110 21310 8190
rect 21490 8110 21500 8190
rect 30510 8170 30520 8290
rect 30640 8270 30650 8290
rect 30640 8190 32602 8270
rect 30640 8170 30650 8190
rect 30510 8160 30650 8170
rect 21300 8100 21500 8110
rect 30900 8090 31040 8100
rect 820 8050 1020 8060
rect 20500 8050 20700 8060
rect 820 8040 830 8050
rect -220 7980 830 8040
rect 820 7970 830 7980
rect 1010 8040 1020 8050
rect 2500 8040 2700 8050
rect 3160 8040 3360 8050
rect 3820 8040 4020 8050
rect 4700 8040 4900 8050
rect 5360 8040 5560 8050
rect 6020 8040 6220 8050
rect 6900 8040 7100 8050
rect 7560 8040 7760 8050
rect 8220 8040 8420 8050
rect 9100 8040 9300 8050
rect 9760 8040 9960 8050
rect 10420 8040 10620 8050
rect 11300 8040 11500 8050
rect 11960 8040 12160 8050
rect 12620 8040 12820 8050
rect 13500 8040 13700 8050
rect 14160 8040 14360 8050
rect 14820 8040 15020 8050
rect 15700 8040 15900 8050
rect 16360 8040 16560 8050
rect 17020 8040 17220 8050
rect 17900 8040 18100 8050
rect 18560 8040 18760 8050
rect 19220 8040 19420 8050
rect 20500 8040 20510 8050
rect 1010 7980 6910 8040
rect 7090 7980 7570 8040
rect 7750 7980 8230 8040
rect 8410 7980 9110 8040
rect 9290 7980 9770 8040
rect 9950 7980 10430 8040
rect 10610 7980 11310 8040
rect 11490 7980 11970 8040
rect 12150 7980 12630 8040
rect 12810 7980 13510 8040
rect 13690 7980 14170 8040
rect 14350 7980 14830 8040
rect 15010 7980 20510 8040
rect 1010 7970 1020 7980
rect 2500 7970 2700 7980
rect 3160 7970 3360 7980
rect 3820 7970 4020 7980
rect 4700 7970 4900 7980
rect 5360 7970 5560 7980
rect 6020 7970 6220 7980
rect 6900 7970 7100 7980
rect 7560 7970 7760 7980
rect 8220 7970 8420 7980
rect 9100 7970 9300 7980
rect 9760 7970 9960 7980
rect 10420 7970 10620 7980
rect 11300 7970 11500 7980
rect 11960 7970 12160 7980
rect 12620 7970 12820 7980
rect 13500 7970 13700 7980
rect 14160 7970 14360 7980
rect 14820 7970 15020 7980
rect 15700 7970 15900 7980
rect 16360 7970 16560 7980
rect 17020 7970 17220 7980
rect 17900 7970 18100 7980
rect 18560 7970 18760 7980
rect 19220 7970 19420 7980
rect 20500 7970 20510 7980
rect 20690 8040 20700 8050
rect 20690 7980 22180 8040
rect 20690 7970 20700 7980
rect 820 7960 1020 7970
rect 20500 7960 20700 7970
rect 30900 7970 30910 8090
rect 31030 8070 31040 8090
rect 31030 7990 32366 8070
rect 31030 7970 31040 7990
rect 30900 7960 31040 7970
rect 1220 7910 1420 7920
rect 20900 7910 21100 7920
rect 1220 7900 1230 7910
rect -220 7840 1230 7900
rect 1220 7830 1230 7840
rect 1410 7900 1420 7910
rect 2500 7900 2700 7910
rect 3160 7900 3360 7910
rect 3820 7900 4020 7910
rect 4700 7900 4900 7910
rect 5360 7900 5560 7910
rect 6020 7900 6220 7910
rect 6900 7900 7100 7910
rect 7560 7900 7760 7910
rect 8220 7900 8420 7910
rect 9100 7900 9300 7910
rect 9760 7900 9960 7910
rect 10420 7900 10620 7910
rect 11300 7900 11500 7910
rect 11960 7900 12160 7910
rect 12620 7900 12820 7910
rect 13500 7900 13700 7910
rect 14160 7900 14360 7910
rect 14820 7900 15020 7910
rect 15700 7900 15900 7910
rect 16360 7900 16560 7910
rect 17020 7900 17220 7910
rect 17900 7900 18100 7910
rect 18560 7900 18760 7910
rect 19220 7900 19420 7910
rect 20900 7900 20910 7910
rect 1410 7840 2510 7900
rect 2690 7840 3170 7900
rect 3350 7840 3830 7900
rect 4010 7840 4710 7900
rect 4890 7840 5370 7900
rect 5550 7840 6030 7900
rect 6210 7840 15710 7900
rect 15890 7840 16370 7900
rect 16550 7840 17030 7900
rect 17210 7840 17910 7900
rect 18090 7840 18570 7900
rect 18750 7840 19230 7900
rect 19410 7840 20910 7900
rect 1410 7830 1420 7840
rect 2500 7830 2700 7840
rect 3160 7830 3360 7840
rect 3820 7830 4020 7840
rect 4700 7830 4900 7840
rect 5360 7830 5560 7840
rect 6020 7830 6220 7840
rect 6900 7830 7100 7840
rect 7560 7830 7760 7840
rect 8220 7830 8420 7840
rect 9100 7830 9300 7840
rect 9760 7830 9960 7840
rect 10420 7830 10620 7840
rect 11300 7830 11500 7840
rect 11960 7830 12160 7840
rect 12620 7830 12820 7840
rect 13500 7830 13700 7840
rect 14160 7830 14360 7840
rect 14820 7830 15020 7840
rect 15700 7830 15900 7840
rect 16360 7830 16560 7840
rect 17020 7830 17220 7840
rect 17900 7830 18100 7840
rect 18560 7830 18760 7840
rect 19220 7830 19420 7840
rect 20900 7830 20910 7840
rect 21090 7900 21100 7910
rect 21090 7840 22180 7900
rect 21090 7830 21100 7840
rect 1220 7820 1420 7830
rect 20900 7820 21100 7830
rect -110 7740 30 7760
rect -110 7490 -80 7740
rect 0 7490 30 7740
rect -110 7460 30 7490
rect 2090 7740 2230 7760
rect 2090 7490 2120 7740
rect 2200 7490 2230 7740
rect 2090 7460 2230 7490
rect 4290 7740 4430 7760
rect 4290 7490 4320 7740
rect 4400 7490 4430 7740
rect 4290 7460 4430 7490
rect 6490 7740 6630 7760
rect 6490 7490 6520 7740
rect 6600 7490 6630 7740
rect 6490 7460 6630 7490
rect 8690 7740 8830 7760
rect 8690 7490 8720 7740
rect 8800 7490 8830 7740
rect 8690 7460 8830 7490
rect 10890 7740 11030 7760
rect 10890 7490 10920 7740
rect 11000 7490 11030 7740
rect 10890 7460 11030 7490
rect 13090 7740 13230 7760
rect 13090 7490 13120 7740
rect 13200 7490 13230 7740
rect 13090 7460 13230 7490
rect 15290 7740 15430 7760
rect 15290 7490 15320 7740
rect 15400 7490 15430 7740
rect 15290 7460 15430 7490
rect 17490 7740 17630 7760
rect 17490 7490 17520 7740
rect 17600 7490 17630 7740
rect 17490 7460 17630 7490
rect 19690 7740 19830 7760
rect 19690 7490 19720 7740
rect 19800 7490 19830 7740
rect 19690 7460 19830 7490
rect 21890 7740 22030 7760
rect 21890 7490 21920 7740
rect 22000 7490 22030 7740
rect 21890 7460 22030 7490
rect 32286 7470 32366 7990
rect 32518 7670 32602 8190
rect 35340 7690 35480 7700
rect 35340 7670 35350 7690
rect 32518 7590 35350 7670
rect 35340 7570 35350 7590
rect 35470 7570 35480 7690
rect 35340 7560 35480 7570
rect 37500 7490 37640 7500
rect 37500 7470 37510 7490
rect 4700 7410 6220 7420
rect 420 7390 620 7400
rect 420 7310 430 7390
rect 610 7310 620 7390
rect 1620 7390 1820 7400
rect 1620 7380 1630 7390
rect 1600 7320 1630 7380
rect 420 7300 620 7310
rect 1620 7310 1630 7320
rect 1810 7380 1820 7390
rect 4700 7380 4710 7410
rect 1810 7350 4710 7380
rect 6210 7380 6220 7410
rect 6900 7410 8420 7420
rect 6900 7380 6910 7410
rect 6210 7350 6910 7380
rect 8410 7380 8420 7410
rect 9100 7410 10620 7420
rect 9100 7380 9110 7410
rect 8410 7350 9110 7380
rect 10610 7380 10620 7410
rect 11300 7410 12820 7420
rect 11300 7380 11310 7410
rect 10610 7350 11310 7380
rect 12810 7380 12820 7410
rect 13500 7410 15020 7420
rect 13500 7380 13510 7410
rect 12810 7350 13510 7380
rect 15010 7380 15020 7410
rect 15700 7410 17220 7420
rect 15700 7380 15710 7410
rect 15010 7350 15710 7380
rect 17210 7380 17220 7410
rect 20100 7390 20300 7400
rect 20100 7380 20110 7390
rect 17210 7350 20110 7380
rect 1810 7320 20110 7350
rect 1810 7310 1820 7320
rect 1620 7300 1820 7310
rect 20100 7310 20110 7320
rect 20290 7380 20300 7390
rect 21300 7390 21500 7400
rect 32286 7390 37510 7470
rect 20290 7320 20320 7380
rect 20290 7310 20300 7320
rect 20100 7300 20300 7310
rect 21300 7310 21310 7390
rect 21490 7310 21500 7390
rect 37500 7370 37510 7390
rect 37630 7370 37640 7490
rect 37500 7360 37640 7370
rect 21300 7300 21500 7310
rect 820 7250 1020 7260
rect 20500 7250 20700 7260
rect 820 7240 830 7250
rect -220 7180 830 7240
rect 820 7170 830 7180
rect 1010 7240 1020 7250
rect 2500 7240 2700 7250
rect 3160 7240 3360 7250
rect 3820 7240 4020 7250
rect 4700 7240 4900 7250
rect 5360 7240 5560 7250
rect 6020 7240 6220 7250
rect 6900 7240 7100 7250
rect 7560 7240 7760 7250
rect 8220 7240 8420 7250
rect 9100 7240 9300 7250
rect 9760 7240 9960 7250
rect 10420 7240 10620 7250
rect 11300 7240 11500 7250
rect 11960 7240 12160 7250
rect 12620 7240 12820 7250
rect 13500 7240 13700 7250
rect 14160 7240 14360 7250
rect 14820 7240 15020 7250
rect 15700 7240 15900 7250
rect 16360 7240 16560 7250
rect 17020 7240 17220 7250
rect 17900 7240 18100 7250
rect 18560 7240 18760 7250
rect 19220 7240 19420 7250
rect 20500 7240 20510 7250
rect 1010 7180 2510 7240
rect 2690 7180 3170 7240
rect 3350 7180 3830 7240
rect 4010 7180 4710 7240
rect 4890 7180 5370 7240
rect 5550 7180 6030 7240
rect 6210 7180 15710 7240
rect 15890 7180 16370 7240
rect 16550 7180 17030 7240
rect 17210 7180 17910 7240
rect 18090 7180 18570 7240
rect 18750 7180 19230 7240
rect 19410 7180 20510 7240
rect 1010 7170 1020 7180
rect 2500 7170 2700 7180
rect 3160 7170 3360 7180
rect 3820 7170 4020 7180
rect 4700 7170 4900 7180
rect 5360 7170 5560 7180
rect 6020 7170 6220 7180
rect 6900 7170 7100 7180
rect 7560 7170 7760 7180
rect 8220 7170 8420 7180
rect 9100 7170 9300 7180
rect 9760 7170 9960 7180
rect 10420 7170 10620 7180
rect 11300 7170 11500 7180
rect 11960 7170 12160 7180
rect 12620 7170 12820 7180
rect 13500 7170 13700 7180
rect 14160 7170 14360 7180
rect 14820 7170 15020 7180
rect 15700 7170 15900 7180
rect 16360 7170 16560 7180
rect 17020 7170 17220 7180
rect 17900 7170 18100 7180
rect 18560 7170 18760 7180
rect 19220 7170 19420 7180
rect 20500 7170 20510 7180
rect 20690 7240 20700 7250
rect 20690 7180 22180 7240
rect 33090 7186 37698 7198
rect 20690 7170 20700 7180
rect 820 7160 1020 7170
rect 20500 7160 20700 7170
rect 1220 7110 1420 7120
rect 20900 7110 21100 7120
rect 1220 7100 1230 7110
rect -220 7040 1230 7100
rect 1220 7030 1230 7040
rect 1410 7100 1420 7110
rect 2500 7100 2700 7110
rect 3160 7100 3360 7110
rect 3820 7100 4020 7110
rect 4700 7100 4900 7110
rect 5360 7100 5560 7110
rect 6020 7100 6220 7110
rect 6900 7100 7100 7110
rect 7560 7100 7760 7110
rect 8220 7100 8420 7110
rect 9100 7100 9300 7110
rect 9760 7100 9960 7110
rect 10420 7100 10620 7110
rect 11300 7100 11500 7110
rect 11960 7100 12160 7110
rect 12620 7100 12820 7110
rect 13500 7100 13700 7110
rect 14160 7100 14360 7110
rect 14820 7100 15020 7110
rect 15700 7100 15900 7110
rect 16360 7100 16560 7110
rect 17020 7100 17220 7110
rect 17900 7100 18100 7110
rect 18560 7100 18760 7110
rect 19220 7100 19420 7110
rect 20900 7100 20910 7110
rect 1410 7040 6910 7100
rect 7090 7040 7570 7100
rect 7750 7040 8230 7100
rect 8410 7040 9110 7100
rect 9290 7040 9770 7100
rect 9950 7040 10430 7100
rect 10610 7040 11310 7100
rect 11490 7040 11970 7100
rect 12150 7040 12630 7100
rect 12810 7040 13510 7100
rect 13690 7040 14170 7100
rect 14350 7040 14830 7100
rect 15010 7040 20910 7100
rect 1410 7030 1420 7040
rect 2500 7030 2700 7040
rect 3160 7030 3360 7040
rect 3820 7030 4020 7040
rect 4700 7030 4900 7040
rect 5360 7030 5560 7040
rect 6020 7030 6220 7040
rect 6900 7030 7100 7040
rect 7560 7030 7760 7040
rect 8220 7030 8420 7040
rect 9100 7030 9300 7040
rect 9760 7030 9960 7040
rect 10420 7030 10620 7040
rect 11300 7030 11500 7040
rect 11960 7030 12160 7040
rect 12620 7030 12820 7040
rect 13500 7030 13700 7040
rect 14160 7030 14360 7040
rect 14820 7030 15020 7040
rect 15700 7030 15900 7040
rect 16360 7030 16560 7040
rect 17020 7030 17220 7040
rect 17900 7030 18100 7040
rect 18560 7030 18760 7040
rect 19220 7030 19420 7040
rect 20900 7030 20910 7040
rect 21090 7100 21100 7110
rect 21090 7040 22180 7100
rect 21090 7030 21100 7040
rect 1220 7020 1420 7030
rect 20900 7020 21100 7030
rect 33090 6976 33108 7186
rect 33474 7176 37516 7186
rect 33474 6982 36128 7176
rect 36810 6982 37516 7176
rect 33474 6976 37516 6982
rect 33090 6974 37516 6976
rect 37684 6974 37698 7186
rect 33090 6960 37698 6974
rect -110 6940 30 6960
rect -110 6690 -80 6940
rect 0 6690 30 6940
rect -110 6660 30 6690
rect 2090 6940 2230 6960
rect 2090 6690 2120 6940
rect 2200 6690 2230 6940
rect 2090 6660 2230 6690
rect 4290 6940 4430 6960
rect 4290 6690 4320 6940
rect 4400 6690 4430 6940
rect 4290 6660 4430 6690
rect 6490 6940 6630 6960
rect 6490 6690 6520 6940
rect 6600 6690 6630 6940
rect 6490 6660 6630 6690
rect 8690 6940 8830 6960
rect 8690 6690 8720 6940
rect 8800 6690 8830 6940
rect 8690 6660 8830 6690
rect 10890 6940 11030 6960
rect 10890 6690 10920 6940
rect 11000 6690 11030 6940
rect 10890 6660 11030 6690
rect 13090 6940 13230 6960
rect 13090 6690 13120 6940
rect 13200 6690 13230 6940
rect 13090 6660 13230 6690
rect 15290 6940 15430 6960
rect 15290 6690 15320 6940
rect 15400 6690 15430 6940
rect 15290 6660 15430 6690
rect 17490 6940 17630 6960
rect 17490 6690 17520 6940
rect 17600 6690 17630 6940
rect 17490 6660 17630 6690
rect 19690 6940 19830 6960
rect 19690 6690 19720 6940
rect 19800 6690 19830 6940
rect 19690 6660 19830 6690
rect 21890 6940 22030 6960
rect 21890 6690 21920 6940
rect 22000 6690 22030 6940
rect 21890 6660 22030 6690
rect 4700 6610 6220 6620
rect 420 6590 620 6600
rect 420 6510 430 6590
rect 610 6510 620 6590
rect 1620 6590 1820 6600
rect 1620 6580 1630 6590
rect 1600 6520 1630 6580
rect 420 6500 620 6510
rect 1620 6510 1630 6520
rect 1810 6580 1820 6590
rect 4700 6580 4710 6610
rect 1810 6550 4710 6580
rect 6210 6580 6220 6610
rect 6900 6610 8420 6620
rect 6900 6580 6910 6610
rect 6210 6550 6910 6580
rect 8410 6580 8420 6610
rect 9100 6610 10620 6620
rect 9100 6580 9110 6610
rect 8410 6550 9110 6580
rect 10610 6580 10620 6610
rect 11300 6610 12820 6620
rect 11300 6580 11310 6610
rect 10610 6550 11310 6580
rect 12810 6580 12820 6610
rect 13500 6610 15020 6620
rect 13500 6580 13510 6610
rect 12810 6550 13510 6580
rect 15010 6580 15020 6610
rect 15700 6610 17220 6620
rect 15700 6580 15710 6610
rect 15010 6550 15710 6580
rect 17210 6580 17220 6610
rect 20100 6590 20300 6600
rect 20100 6580 20110 6590
rect 17210 6550 20110 6580
rect 1810 6520 20110 6550
rect 1810 6510 1820 6520
rect 1620 6500 1820 6510
rect 20100 6510 20110 6520
rect 20290 6580 20300 6590
rect 21300 6590 21500 6600
rect 20290 6520 20320 6580
rect 20290 6510 20300 6520
rect 20100 6500 20300 6510
rect 21300 6510 21310 6590
rect 21490 6510 21500 6590
rect 21300 6500 21500 6510
rect 820 6450 1020 6460
rect 20500 6450 20700 6460
rect 820 6440 830 6450
rect -220 6380 830 6440
rect 820 6370 830 6380
rect 1010 6440 1020 6450
rect 2500 6440 2700 6450
rect 3160 6440 3360 6450
rect 3820 6440 4020 6450
rect 4700 6440 4900 6450
rect 5360 6440 5560 6450
rect 6020 6440 6220 6450
rect 6900 6440 7100 6450
rect 7560 6440 7760 6450
rect 8220 6440 8420 6450
rect 9100 6440 9300 6450
rect 9760 6440 9960 6450
rect 10420 6440 10620 6450
rect 11300 6440 11500 6450
rect 11960 6440 12160 6450
rect 12620 6440 12820 6450
rect 13500 6440 13700 6450
rect 14160 6440 14360 6450
rect 14820 6440 15020 6450
rect 15700 6440 15900 6450
rect 16360 6440 16560 6450
rect 17020 6440 17220 6450
rect 17900 6440 18100 6450
rect 18560 6440 18760 6450
rect 19220 6440 19420 6450
rect 20500 6440 20510 6450
rect 1010 6380 6910 6440
rect 7090 6380 7570 6440
rect 7750 6380 8230 6440
rect 8410 6380 9110 6440
rect 9290 6380 9770 6440
rect 9950 6380 10430 6440
rect 10610 6380 11310 6440
rect 11490 6380 11970 6440
rect 12150 6380 12630 6440
rect 12810 6380 13510 6440
rect 13690 6380 14170 6440
rect 14350 6380 14830 6440
rect 15010 6380 20510 6440
rect 1010 6370 1020 6380
rect 2500 6370 2700 6380
rect 3160 6370 3360 6380
rect 3820 6370 4020 6380
rect 4700 6370 4900 6380
rect 5360 6370 5560 6380
rect 6020 6370 6220 6380
rect 6900 6370 7100 6380
rect 7560 6370 7760 6380
rect 8220 6370 8420 6380
rect 9100 6370 9300 6380
rect 9760 6370 9960 6380
rect 10420 6370 10620 6380
rect 11300 6370 11500 6380
rect 11960 6370 12160 6380
rect 12620 6370 12820 6380
rect 13500 6370 13700 6380
rect 14160 6370 14360 6380
rect 14820 6370 15020 6380
rect 15700 6370 15900 6380
rect 16360 6370 16560 6380
rect 17020 6370 17220 6380
rect 17900 6370 18100 6380
rect 18560 6370 18760 6380
rect 19220 6370 19420 6380
rect 20500 6370 20510 6380
rect 20690 6440 20700 6450
rect 20690 6380 22180 6440
rect 20690 6370 20700 6380
rect 820 6360 1020 6370
rect 20500 6360 20700 6370
rect 1220 6310 1420 6320
rect 20900 6310 21100 6320
rect 1220 6300 1230 6310
rect -220 6240 1230 6300
rect 1220 6230 1230 6240
rect 1410 6300 1420 6310
rect 2500 6300 2700 6310
rect 3160 6300 3360 6310
rect 3820 6300 4020 6310
rect 4700 6300 4900 6310
rect 5360 6300 5560 6310
rect 6020 6300 6220 6310
rect 6900 6300 7100 6310
rect 7560 6300 7760 6310
rect 8220 6300 8420 6310
rect 9100 6300 9300 6310
rect 9760 6300 9960 6310
rect 10420 6300 10620 6310
rect 11300 6300 11500 6310
rect 11960 6300 12160 6310
rect 12620 6300 12820 6310
rect 13500 6300 13700 6310
rect 14160 6300 14360 6310
rect 14820 6300 15020 6310
rect 15700 6300 15900 6310
rect 16360 6300 16560 6310
rect 17020 6300 17220 6310
rect 17900 6300 18100 6310
rect 18560 6300 18760 6310
rect 19220 6300 19420 6310
rect 20900 6300 20910 6310
rect 1410 6240 2510 6300
rect 2690 6240 3170 6300
rect 3350 6240 3830 6300
rect 4010 6240 4710 6300
rect 4890 6240 5370 6300
rect 5550 6240 6030 6300
rect 6210 6240 15710 6300
rect 15890 6240 16370 6300
rect 16550 6240 17030 6300
rect 17210 6240 17910 6300
rect 18090 6240 18570 6300
rect 18750 6240 19230 6300
rect 19410 6240 20910 6300
rect 1410 6230 1420 6240
rect 2500 6230 2700 6240
rect 3160 6230 3360 6240
rect 3820 6230 4020 6240
rect 4700 6230 4900 6240
rect 5360 6230 5560 6240
rect 6020 6230 6220 6240
rect 6900 6230 7100 6240
rect 7560 6230 7760 6240
rect 8220 6230 8420 6240
rect 9100 6230 9300 6240
rect 9760 6230 9960 6240
rect 10420 6230 10620 6240
rect 11300 6230 11500 6240
rect 11960 6230 12160 6240
rect 12620 6230 12820 6240
rect 13500 6230 13700 6240
rect 14160 6230 14360 6240
rect 14820 6230 15020 6240
rect 15700 6230 15900 6240
rect 16360 6230 16560 6240
rect 17020 6230 17220 6240
rect 17900 6230 18100 6240
rect 18560 6230 18760 6240
rect 19220 6230 19420 6240
rect 20900 6230 20910 6240
rect 21090 6300 21100 6310
rect 21090 6240 22180 6300
rect 36220 6260 36420 6270
rect 21090 6230 21100 6240
rect 1220 6220 1420 6230
rect 20900 6220 21100 6230
rect -110 6140 30 6160
rect -110 5890 -80 6140
rect 0 5890 30 6140
rect -110 5860 30 5890
rect 2090 6140 2230 6160
rect 2090 5890 2120 6140
rect 2200 5890 2230 6140
rect 2090 5860 2230 5890
rect 4290 6140 4430 6160
rect 4290 5890 4320 6140
rect 4400 5890 4430 6140
rect 4290 5860 4430 5890
rect 6490 6140 6630 6160
rect 6490 5890 6520 6140
rect 6600 5890 6630 6140
rect 6490 5860 6630 5890
rect 8690 6140 8830 6160
rect 8690 5890 8720 6140
rect 8800 5890 8830 6140
rect 8690 5860 8830 5890
rect 10890 6140 11030 6160
rect 10890 5890 10920 6140
rect 11000 5890 11030 6140
rect 10890 5860 11030 5890
rect 13090 6140 13230 6160
rect 13090 5890 13120 6140
rect 13200 5890 13230 6140
rect 13090 5860 13230 5890
rect 15290 6140 15430 6160
rect 15290 5890 15320 6140
rect 15400 5890 15430 6140
rect 15290 5860 15430 5890
rect 17490 6140 17630 6160
rect 17490 5890 17520 6140
rect 17600 5890 17630 6140
rect 17490 5860 17630 5890
rect 19690 6140 19830 6160
rect 19690 5890 19720 6140
rect 19800 5890 19830 6140
rect 19690 5860 19830 5890
rect 21890 6140 22030 6160
rect 21890 5890 21920 6140
rect 22000 5890 22030 6140
rect 36220 6080 36230 6260
rect 36410 6080 36420 6260
rect 36220 6070 36420 6080
rect 36520 6260 36720 6270
rect 36520 6080 36530 6260
rect 36710 6080 36720 6260
rect 36520 6070 36720 6080
rect 21890 5860 22030 5890
rect 2500 5810 4020 5820
rect 1620 5790 1820 5800
rect 1620 5780 1630 5790
rect 1600 5720 1630 5780
rect 1620 5710 1630 5720
rect 1810 5780 1820 5790
rect 2500 5780 2510 5810
rect 1810 5750 2510 5780
rect 4010 5780 4020 5810
rect 4700 5810 6220 5820
rect 4700 5780 4710 5810
rect 4010 5750 4710 5780
rect 6210 5780 6220 5810
rect 6900 5810 8420 5820
rect 6900 5780 6910 5810
rect 6210 5750 6910 5780
rect 8410 5780 8420 5810
rect 9100 5810 10620 5820
rect 9100 5780 9110 5810
rect 8410 5750 9110 5780
rect 10610 5780 10620 5810
rect 11300 5810 12820 5820
rect 11300 5780 11310 5810
rect 10610 5750 11310 5780
rect 12810 5780 12820 5810
rect 13500 5810 15020 5820
rect 13500 5780 13510 5810
rect 12810 5750 13510 5780
rect 15010 5780 15020 5810
rect 15700 5810 17220 5820
rect 15700 5780 15710 5810
rect 15010 5750 15710 5780
rect 17210 5780 17220 5810
rect 17900 5810 19420 5820
rect 17900 5780 17910 5810
rect 17210 5750 17910 5780
rect 19410 5780 19420 5810
rect 20100 5790 20300 5800
rect 20100 5780 20110 5790
rect 19410 5750 20110 5780
rect 1810 5720 20110 5750
rect 1810 5710 1820 5720
rect 1620 5700 1820 5710
rect 20100 5710 20110 5720
rect 20290 5780 20300 5790
rect 20290 5720 20320 5780
rect 20290 5710 20300 5720
rect 20100 5700 20300 5710
rect 820 5650 1020 5660
rect 20500 5650 20700 5660
rect 820 5640 830 5650
rect -220 5580 830 5640
rect 820 5570 830 5580
rect 1010 5640 1020 5650
rect 2500 5640 2700 5650
rect 3160 5640 3360 5650
rect 3820 5640 4020 5650
rect 4700 5640 4900 5650
rect 5360 5640 5560 5650
rect 6020 5640 6220 5650
rect 6900 5640 7100 5650
rect 7560 5640 7760 5650
rect 8220 5640 8420 5650
rect 9100 5640 9300 5650
rect 9760 5640 9960 5650
rect 10420 5640 10620 5650
rect 11300 5640 11500 5650
rect 11960 5640 12160 5650
rect 12620 5640 12820 5650
rect 13500 5640 13700 5650
rect 14160 5640 14360 5650
rect 14820 5640 15020 5650
rect 15700 5640 15900 5650
rect 16360 5640 16560 5650
rect 17020 5640 17220 5650
rect 17900 5640 18100 5650
rect 18560 5640 18760 5650
rect 19220 5640 19420 5650
rect 20500 5640 20510 5650
rect 1010 5580 2510 5640
rect 2690 5580 3170 5640
rect 3350 5580 3830 5640
rect 4010 5580 4710 5640
rect 4890 5580 5370 5640
rect 5550 5580 6030 5640
rect 6210 5580 15710 5640
rect 15890 5580 16370 5640
rect 16550 5580 17030 5640
rect 17210 5580 17910 5640
rect 18090 5580 18570 5640
rect 18750 5580 19230 5640
rect 19410 5580 20510 5640
rect 1010 5570 1020 5580
rect 2500 5570 2700 5580
rect 3160 5570 3360 5580
rect 3820 5570 4020 5580
rect 4700 5570 4900 5580
rect 5360 5570 5560 5580
rect 6020 5570 6220 5580
rect 6900 5570 7100 5580
rect 7560 5570 7760 5580
rect 8220 5570 8420 5580
rect 9100 5570 9300 5580
rect 9760 5570 9960 5580
rect 10420 5570 10620 5580
rect 11300 5570 11500 5580
rect 11960 5570 12160 5580
rect 12620 5570 12820 5580
rect 13500 5570 13700 5580
rect 14160 5570 14360 5580
rect 14820 5570 15020 5580
rect 15700 5570 15900 5580
rect 16360 5570 16560 5580
rect 17020 5570 17220 5580
rect 17900 5570 18100 5580
rect 18560 5570 18760 5580
rect 19220 5570 19420 5580
rect 20500 5570 20510 5580
rect 20690 5640 20700 5650
rect 20690 5580 22180 5640
rect 20690 5570 20700 5580
rect 820 5560 1020 5570
rect 20500 5560 20700 5570
rect 1220 5510 1420 5520
rect 20900 5510 21100 5520
rect 1220 5500 1230 5510
rect -220 5440 1230 5500
rect 1220 5430 1230 5440
rect 1410 5500 1420 5510
rect 2500 5500 2700 5510
rect 3160 5500 3360 5510
rect 3820 5500 4020 5510
rect 4700 5500 4900 5510
rect 5360 5500 5560 5510
rect 6020 5500 6220 5510
rect 6900 5500 7100 5510
rect 7560 5500 7760 5510
rect 8220 5500 8420 5510
rect 9100 5500 9300 5510
rect 9760 5500 9960 5510
rect 10420 5500 10620 5510
rect 11300 5500 11500 5510
rect 11960 5500 12160 5510
rect 12620 5500 12820 5510
rect 13500 5500 13700 5510
rect 14160 5500 14360 5510
rect 14820 5500 15020 5510
rect 15700 5500 15900 5510
rect 16360 5500 16560 5510
rect 17020 5500 17220 5510
rect 17900 5500 18100 5510
rect 18560 5500 18760 5510
rect 19220 5500 19420 5510
rect 20900 5500 20910 5510
rect 1410 5440 6910 5500
rect 7090 5440 7570 5500
rect 7750 5440 8230 5500
rect 8410 5440 9110 5500
rect 9290 5440 9770 5500
rect 9950 5440 10430 5500
rect 10610 5440 11310 5500
rect 11490 5440 11970 5500
rect 12150 5440 12630 5500
rect 12810 5440 13510 5500
rect 13690 5440 14170 5500
rect 14350 5440 14830 5500
rect 15010 5440 20910 5500
rect 1410 5430 1420 5440
rect 2500 5430 2700 5440
rect 3160 5430 3360 5440
rect 3820 5430 4020 5440
rect 4700 5430 4900 5440
rect 5360 5430 5560 5440
rect 6020 5430 6220 5440
rect 6900 5430 7100 5440
rect 7560 5430 7760 5440
rect 8220 5430 8420 5440
rect 9100 5430 9300 5440
rect 9760 5430 9960 5440
rect 10420 5430 10620 5440
rect 11300 5430 11500 5440
rect 11960 5430 12160 5440
rect 12620 5430 12820 5440
rect 13500 5430 13700 5440
rect 14160 5430 14360 5440
rect 14820 5430 15020 5440
rect 15700 5430 15900 5440
rect 16360 5430 16560 5440
rect 17020 5430 17220 5440
rect 17900 5430 18100 5440
rect 18560 5430 18760 5440
rect 19220 5430 19420 5440
rect 20900 5430 20910 5440
rect 21090 5500 21100 5510
rect 21090 5440 22180 5500
rect 21090 5430 21100 5440
rect 1220 5420 1420 5430
rect 20900 5420 21100 5430
rect 28490 5400 28670 5410
rect -110 5340 30 5360
rect -110 5090 -80 5340
rect 0 5090 30 5340
rect -110 5060 30 5090
rect 2090 5340 2230 5360
rect 2090 5090 2120 5340
rect 2200 5090 2230 5340
rect 2090 5060 2230 5090
rect 4290 5340 4430 5360
rect 4290 5090 4320 5340
rect 4400 5090 4430 5340
rect 4290 5060 4430 5090
rect 6490 5340 6630 5360
rect 6490 5090 6520 5340
rect 6600 5090 6630 5340
rect 6490 5060 6630 5090
rect 8690 5340 8830 5360
rect 8690 5090 8720 5340
rect 8800 5090 8830 5340
rect 8690 5060 8830 5090
rect 10890 5340 11030 5360
rect 10890 5090 10920 5340
rect 11000 5090 11030 5340
rect 10890 5060 11030 5090
rect 13090 5340 13230 5360
rect 13090 5090 13120 5340
rect 13200 5090 13230 5340
rect 13090 5060 13230 5090
rect 15290 5340 15430 5360
rect 15290 5090 15320 5340
rect 15400 5090 15430 5340
rect 15290 5060 15430 5090
rect 17490 5340 17630 5360
rect 17490 5090 17520 5340
rect 17600 5090 17630 5340
rect 17490 5060 17630 5090
rect 19690 5340 19830 5360
rect 19690 5090 19720 5340
rect 19800 5090 19830 5340
rect 19690 5060 19830 5090
rect 21890 5340 22030 5360
rect 21890 5090 21920 5340
rect 22000 5090 22030 5340
rect 28490 5240 28500 5400
rect 28660 5370 28670 5400
rect 36290 5370 36400 5380
rect 28660 5360 35120 5370
rect 28660 5280 34900 5360
rect 35110 5280 35120 5360
rect 28660 5270 35120 5280
rect 28660 5240 28670 5270
rect 28490 5230 28670 5240
rect 21890 5060 22030 5090
rect 36290 5040 36300 5370
rect 36390 5250 36400 5370
rect 37670 5370 37780 5380
rect 36860 5320 37020 5330
rect 36860 5250 36870 5320
rect 36390 5170 36870 5250
rect 36390 5040 36400 5170
rect 36860 5100 36870 5170
rect 37010 5100 37020 5320
rect 36860 5090 37020 5100
rect 37120 5320 37280 5330
rect 37120 5100 37130 5320
rect 37270 5250 37280 5320
rect 37670 5250 37680 5370
rect 37270 5170 37680 5250
rect 37270 5100 37280 5170
rect 37120 5090 37280 5100
rect 36290 5030 36400 5040
rect 37670 5040 37680 5170
rect 37770 5040 37780 5370
rect 37670 5030 37780 5040
rect 2500 5010 4020 5020
rect 1620 4990 1820 5000
rect 1620 4980 1630 4990
rect 1600 4920 1630 4980
rect 1620 4910 1630 4920
rect 1810 4980 1820 4990
rect 2500 4980 2510 5010
rect 1810 4950 2510 4980
rect 4010 4980 4020 5010
rect 4700 5010 6220 5020
rect 4700 4980 4710 5010
rect 4010 4950 4710 4980
rect 6210 4980 6220 5010
rect 6900 5010 8420 5020
rect 6900 4980 6910 5010
rect 6210 4950 6910 4980
rect 8410 4980 8420 5010
rect 9100 5010 10620 5020
rect 9100 4980 9110 5010
rect 8410 4950 9110 4980
rect 10610 4980 10620 5010
rect 11300 5010 12820 5020
rect 11300 4980 11310 5010
rect 10610 4950 11310 4980
rect 12810 4980 12820 5010
rect 13500 5010 15020 5020
rect 13500 4980 13510 5010
rect 12810 4950 13510 4980
rect 15010 4980 15020 5010
rect 15700 5010 17220 5020
rect 15700 4980 15710 5010
rect 15010 4950 15710 4980
rect 17210 4980 17220 5010
rect 17900 5010 19420 5020
rect 17900 4980 17910 5010
rect 17210 4950 17910 4980
rect 19410 4980 19420 5010
rect 20100 4990 20300 5000
rect 20100 4980 20110 4990
rect 19410 4950 20110 4980
rect 1810 4920 20110 4950
rect 1810 4910 1820 4920
rect 1620 4900 1820 4910
rect 20100 4910 20110 4920
rect 20290 4980 20300 4990
rect 20290 4920 20320 4980
rect 23040 4970 23590 4980
rect 20290 4910 20300 4920
rect 20100 4900 20300 4910
rect 23040 4710 23050 4970
rect 23580 4940 23590 4970
rect 23580 4930 27440 4940
rect 23580 4750 27250 4930
rect 27430 4750 27440 4930
rect 23580 4710 23590 4750
rect 27240 4740 27440 4750
rect 23040 4700 23590 4710
rect -300 4530 27560 4540
rect -300 4350 1290 4530
rect 1470 4350 20110 4530
rect 20290 4350 27370 4530
rect 27550 4350 27560 4530
rect -300 4340 27560 4350
rect 29130 4520 29210 4530
rect 29130 4290 29140 4520
rect 29200 4410 29210 4520
rect 32490 4480 32650 4490
rect 32490 4410 32500 4480
rect 29200 4340 32500 4410
rect 32640 4410 32650 4480
rect 34080 4480 34240 4490
rect 34080 4410 34090 4480
rect 32640 4340 34090 4410
rect 34230 4340 34240 4480
rect 29200 4290 29210 4340
rect 32490 4330 32650 4340
rect 34080 4330 34240 4340
rect 29130 4280 29210 4290
rect 35690 4290 35850 4300
rect 29270 4260 29520 4270
rect 35690 4260 35700 4290
rect 29270 4190 29280 4260
rect 29510 4190 35700 4260
rect 29270 4180 29520 4190
rect 35690 4150 35700 4190
rect 35840 4150 35850 4290
rect 35690 4140 35850 4150
rect -300 4130 27820 4140
rect -300 3950 1630 4130
rect 1810 3950 20450 4130
rect 20630 3950 27630 4130
rect 27810 3950 27820 4130
rect 33120 4110 33300 4120
rect -300 3940 27820 3950
rect 30070 4040 30270 4050
rect 30070 3860 30080 4040
rect 30260 3860 30270 4040
rect 30070 3850 30270 3860
rect 31670 4040 31870 4050
rect 31670 3860 31680 4040
rect 31860 3860 31870 4040
rect 33120 4010 33130 4110
rect 33290 4010 33300 4110
rect 33120 4000 33300 4010
rect 34860 4090 35200 4100
rect 34860 4010 34870 4090
rect 35190 4010 35200 4090
rect 34860 4000 35200 4010
rect 31670 3850 31870 3860
rect 32070 3740 32220 3750
rect -300 3730 31700 3740
rect -300 3550 430 3730
rect 610 3550 21310 3730
rect 21490 3550 31530 3730
rect 31690 3550 31700 3730
rect 32070 3610 32080 3740
rect 32210 3720 32220 3740
rect 32210 3710 38020 3720
rect 32210 3620 37880 3710
rect 32210 3610 32220 3620
rect 32070 3600 32220 3610
rect 37870 3580 37880 3620
rect 38010 3580 38020 3710
rect 37870 3570 38020 3580
rect -300 3540 31700 3550
rect 26200 3400 26380 3410
rect 26200 3370 26210 3400
rect 1160 3330 20300 3340
rect 1160 3150 1170 3330
rect 1330 3150 1630 3330
rect 1810 3150 2770 3330
rect 2930 3150 4370 3330
rect 4530 3150 5970 3330
rect 6130 3150 7570 3330
rect 7730 3150 9170 3330
rect 9330 3150 20110 3330
rect 20290 3150 20300 3330
rect 1160 3140 20300 3150
rect 20700 3270 26210 3370
rect 14180 3030 14360 3040
rect 10880 3010 11040 3020
rect 7800 2930 7940 2940
rect 7800 2810 7810 2930
rect 7930 2810 7940 2930
rect 10880 2870 10890 3010
rect 11030 3000 11040 3010
rect 14180 3000 14190 3030
rect 11030 2880 14190 3000
rect 11030 2870 11040 2880
rect 10880 2860 11040 2870
rect 14180 2870 14190 2880
rect 14350 2870 14360 3030
rect 14180 2860 14360 2870
rect 18050 3010 18210 3020
rect 18050 2870 18060 3010
rect 18200 2990 18210 3010
rect 20700 2990 20800 3270
rect 26200 3240 26210 3270
rect 26370 3370 26380 3400
rect 26370 3270 26410 3370
rect 26610 3360 26770 3370
rect 26370 3240 26380 3270
rect 26200 3230 26380 3240
rect 26610 3220 26620 3360
rect 26760 3340 26770 3360
rect 36580 3360 36740 3370
rect 36580 3340 36590 3360
rect 26760 3240 36590 3340
rect 26760 3220 26770 3240
rect 26610 3210 26770 3220
rect 36580 3220 36590 3240
rect 36730 3220 36740 3360
rect 36580 3210 36740 3220
rect 18200 2890 20800 2990
rect 23210 3090 32000 3100
rect 23210 2910 23220 3090
rect 23400 2910 31830 3090
rect 31990 2910 32000 3090
rect 23210 2900 32000 2910
rect 18200 2870 18210 2890
rect 18050 2860 18210 2870
rect 7800 2790 7940 2810
rect 16900 2780 17140 2790
rect 11690 2770 11850 2780
rect 11690 2620 11700 2770
rect 11840 2760 11850 2770
rect 16900 2760 16910 2780
rect 11840 2640 16910 2760
rect 17130 2760 17140 2780
rect 17370 2780 17500 2790
rect 17370 2760 17380 2780
rect 17130 2640 17380 2760
rect 17490 2760 17500 2780
rect 17730 2780 17970 2790
rect 17730 2760 17740 2780
rect 17490 2640 17740 2760
rect 17960 2760 17970 2780
rect 34770 2780 34940 2790
rect 34770 2760 34780 2780
rect 17960 2640 34780 2760
rect 11840 2630 34780 2640
rect 11840 2620 11850 2630
rect 11690 2610 11850 2620
rect 34770 2620 34780 2630
rect 34930 2620 34940 2780
rect 34770 2610 34940 2620
rect 33170 2550 33340 2560
rect 10990 2540 11150 2550
rect -1740 2400 11000 2540
rect 11140 2530 11150 2540
rect 12590 2540 12750 2550
rect 12590 2530 12600 2540
rect 11140 2400 12600 2530
rect 12740 2530 12750 2540
rect 13970 2540 14130 2550
rect 13970 2530 13980 2540
rect 12740 2400 13980 2530
rect 14120 2400 14130 2540
rect 33170 2530 33180 2550
rect 10990 2390 11150 2400
rect 12590 2390 12750 2400
rect 13970 2390 14130 2400
rect 14900 2400 33180 2530
rect 2090 2250 13440 2260
rect 470 2220 670 2240
rect 470 -4780 480 2220
rect 660 -4780 670 2220
rect 2090 2090 2110 2250
rect 2230 2090 3710 2250
rect 3830 2090 5310 2250
rect 5430 2090 6910 2250
rect 7030 2090 8510 2250
rect 8630 2090 10110 2250
rect 10230 2090 11710 2250
rect 11830 2090 13310 2250
rect 13430 2090 13440 2250
rect 2090 2080 13440 2090
rect 14900 1980 15040 2400
rect 33170 2390 33180 2400
rect 33330 2390 33340 2550
rect 33170 2380 33340 2390
rect 16500 2250 26240 2260
rect 16500 2090 16510 2250
rect 16630 2090 18110 2250
rect 18230 2090 19710 2250
rect 19830 2090 21310 2250
rect 21430 2090 22910 2250
rect 23030 2090 24510 2250
rect 24630 2090 26110 2250
rect 26230 2090 26240 2250
rect 16500 2080 26240 2090
rect 27700 2250 31040 2260
rect 27700 2070 27710 2250
rect 27830 2070 29310 2250
rect 29430 2070 30910 2250
rect 31030 2070 31040 2250
rect 27700 2060 31040 2070
rect 14900 1320 14910 1980
rect 15030 1320 15040 1980
rect 14900 1290 15040 1320
rect 32500 1150 32640 1160
rect 34100 1150 34240 1160
rect 34780 1150 34930 1160
rect 35700 1150 37440 1160
rect 32500 1030 32510 1150
rect 32630 1030 34110 1150
rect 34230 1030 34790 1150
rect 34920 1030 35710 1150
rect 35830 1030 37310 1150
rect 37430 1030 37440 1150
rect 32500 1020 32640 1030
rect 34100 1020 34240 1030
rect 34780 1020 34930 1030
rect 35700 1020 37440 1030
rect 2090 450 13440 460
rect 2090 290 2110 450
rect 2230 290 3710 450
rect 3830 290 5310 450
rect 5430 290 6910 450
rect 7030 290 8510 450
rect 8630 290 10110 450
rect 10230 290 11710 450
rect 11830 290 13310 450
rect 13430 290 13440 450
rect 2090 280 13440 290
rect 16500 450 26240 460
rect 16500 290 16510 450
rect 16630 290 18110 450
rect 18230 290 19710 450
rect 19830 290 21310 450
rect 21430 290 22910 450
rect 23030 290 24510 450
rect 24630 290 26110 450
rect 26230 290 26240 450
rect 16500 280 26240 290
rect 27700 450 31040 460
rect 27700 270 27710 450
rect 27830 270 29310 450
rect 29430 270 30910 450
rect 31030 270 31040 450
rect 27700 260 31040 270
rect 32500 440 35840 450
rect 32500 280 33180 440
rect 33330 280 35840 440
rect 32500 270 35840 280
rect 32500 190 32640 270
rect 32500 -490 32510 190
rect 32630 -490 32640 190
rect 32500 -500 32640 -490
rect 34100 190 34240 270
rect 34100 -490 34110 190
rect 34230 -490 34240 190
rect 34100 -500 34240 -490
rect 35700 190 35840 270
rect 35700 -490 35710 190
rect 35830 -490 35840 190
rect 35700 -500 35840 -490
rect 12870 -1110 13250 -1100
rect 12870 -1260 12880 -1110
rect 13240 -1260 13250 -1110
rect 12870 -1270 13250 -1260
rect 2090 -1350 15040 -1340
rect 2090 -1510 2110 -1350
rect 2230 -1510 3710 -1350
rect 3830 -1510 5310 -1350
rect 5430 -1510 6910 -1350
rect 7030 -1510 8510 -1350
rect 8630 -1510 10110 -1350
rect 10230 -1510 11710 -1350
rect 11830 -1510 13310 -1350
rect 13430 -1510 14910 -1350
rect 15030 -1510 15040 -1350
rect 2090 -1520 15040 -1510
rect 15240 -1350 26270 -1340
rect 15240 -1510 15250 -1350
rect 15370 -1510 16510 -1350
rect 16630 -1510 18110 -1350
rect 18230 -1510 19710 -1350
rect 19830 -1510 21310 -1350
rect 21430 -1510 22910 -1350
rect 23030 -1510 24510 -1350
rect 24630 -1510 26110 -1350
rect 26230 -1510 26270 -1350
rect 15240 -1520 26270 -1510
rect 27700 -1350 31040 -1340
rect 27700 -1530 27710 -1350
rect 27830 -1530 29310 -1350
rect 29430 -1530 30910 -1350
rect 31030 -1530 31040 -1350
rect 27700 -1540 31040 -1530
rect 32500 -2450 32640 -2440
rect 34100 -2450 34240 -2440
rect 34780 -2450 34930 -2440
rect 35700 -2450 35840 -2440
rect 32500 -2570 32510 -2450
rect 32630 -2570 34110 -2450
rect 34230 -2570 34790 -2450
rect 34920 -2570 35710 -2450
rect 35830 -2570 35840 -2450
rect 32500 -2580 32640 -2570
rect 34100 -2580 34240 -2570
rect 34780 -2580 34930 -2570
rect 35700 -2580 35840 -2570
rect 2090 -3150 15040 -3140
rect 2090 -3310 2110 -3150
rect 2230 -3310 3710 -3150
rect 3830 -3310 5310 -3150
rect 5430 -3310 6910 -3150
rect 7030 -3310 8510 -3150
rect 8630 -3310 10110 -3150
rect 10230 -3310 11710 -3150
rect 11830 -3310 13310 -3150
rect 13430 -3310 14910 -3150
rect 15030 -3310 15040 -3150
rect 2090 -3320 15040 -3310
rect 16500 -3150 26240 -3140
rect 16500 -3310 16510 -3150
rect 16630 -3310 18110 -3150
rect 18230 -3310 19710 -3150
rect 19830 -3310 21310 -3150
rect 21430 -3310 22910 -3150
rect 23030 -3310 24510 -3150
rect 24630 -3310 26110 -3150
rect 26230 -3310 26240 -3150
rect 16500 -3320 26240 -3310
rect 27700 -3150 31040 -3140
rect 27700 -3330 27710 -3150
rect 27830 -3330 29310 -3150
rect 29430 -3330 30910 -3150
rect 31030 -3330 31040 -3150
rect 27700 -3340 31040 -3330
rect 470 -4800 670 -4780
rect 680 -5170 37760 -5160
rect 680 -5350 2810 -5170
rect 2990 -5350 15570 -5170
rect 15730 -5350 18770 -5170
rect 18930 -5350 21280 -5170
rect 21460 -5350 21970 -5170
rect 22130 -5350 25170 -5170
rect 25330 -5350 28370 -5170
rect 28530 -5350 36030 -5170
rect 36210 -5350 37760 -5170
rect 680 -5360 37760 -5350
rect 680 -5570 37760 -5560
rect 80 -5750 280 -5740
rect 80 -5940 90 -5750
rect -1580 -6140 90 -5940
rect 80 -6330 90 -6140
rect 270 -6330 280 -5750
rect 680 -5750 1270 -5570
rect 1450 -5750 15570 -5570
rect 15730 -5750 18770 -5570
rect 18930 -5750 20510 -5570
rect 20690 -5750 21970 -5570
rect 22130 -5750 25170 -5570
rect 25330 -5750 28370 -5570
rect 28530 -5750 36230 -5570
rect 36410 -5750 37760 -5570
rect 680 -5760 37760 -5750
rect 15780 -5970 31990 -5960
rect 15780 -6150 15790 -5970
rect 15950 -6150 18990 -5970
rect 19150 -6150 22190 -5970
rect 22350 -6150 25390 -5970
rect 25550 -6150 27690 -5970
rect 27850 -6150 28590 -5970
rect 28750 -6150 29290 -5970
rect 29450 -6150 30890 -5970
rect 31050 -6150 31680 -5970
rect 31860 -6150 31990 -5970
rect 15780 -6160 31990 -6150
rect 80 -6340 280 -6330
rect 14900 -6490 15040 -6480
rect -360 -6590 -160 -6580
rect -360 -6780 -350 -6590
rect -1580 -6980 -350 -6780
rect -360 -7170 -350 -6980
rect -170 -6780 -160 -6590
rect 14900 -6610 14910 -6490
rect 15030 -6610 15040 -6490
rect 14900 -6620 15040 -6610
rect 17380 -6770 31990 -6760
rect -170 -6980 280 -6780
rect 12940 -6830 13120 -6820
rect -170 -7170 -160 -6980
rect 12940 -6990 12950 -6830
rect 13110 -6990 13120 -6830
rect 17380 -6950 17390 -6770
rect 17550 -6950 20590 -6770
rect 20750 -6950 23790 -6770
rect 23950 -6950 26990 -6770
rect 27150 -6950 30080 -6770
rect 30350 -6950 31990 -6770
rect 17380 -6960 31990 -6950
rect 12940 -7000 13120 -6990
rect -360 -7180 -160 -7170
rect 680 -7170 37760 -7160
rect 680 -7350 1260 -7170
rect 1440 -7350 17170 -7170
rect 17330 -7350 20370 -7170
rect 20690 -7350 23570 -7170
rect 23730 -7350 26770 -7170
rect 26930 -7350 29970 -7170
rect 30130 -7350 36530 -7170
rect 36710 -7350 37760 -7170
rect 680 -7360 37760 -7350
rect 680 -7570 37760 -7560
rect 680 -7750 2080 -7570
rect 2260 -7750 17170 -7570
rect 17330 -7750 20370 -7570
rect 20530 -7750 22070 -7570
rect 22250 -7750 23570 -7570
rect 23730 -7750 26770 -7570
rect 26930 -7750 29970 -7570
rect 30130 -7750 36230 -7570
rect 36410 -7750 37760 -7570
rect 680 -7760 37760 -7750
rect 7800 -7870 7940 -7860
rect 7800 -7990 7810 -7870
rect 7930 -7990 7940 -7870
rect 7800 -8000 7940 -7990
rect 480 -8090 680 -8080
rect 480 -22380 490 -8090
rect 670 -22380 680 -8090
rect 10800 -8260 16650 -8250
rect 10800 -8380 10810 -8260
rect 10930 -8380 13310 -8260
rect 13440 -8380 16510 -8260
rect 16640 -8380 16650 -8260
rect 10800 -8390 16650 -8380
rect 16500 -9570 26250 -9560
rect 2120 -9590 10240 -9580
rect 2120 -9750 2130 -9590
rect 2230 -9750 3730 -9590
rect 3830 -9750 5330 -9590
rect 5430 -9750 6930 -9590
rect 7030 -9750 8530 -9590
rect 8630 -9750 10130 -9590
rect 10230 -9750 10240 -9590
rect 16500 -9730 16510 -9570
rect 16640 -9730 18110 -9570
rect 18240 -9730 19710 -9570
rect 19840 -9730 21310 -9570
rect 21440 -9730 22910 -9570
rect 23040 -9730 24510 -9570
rect 24640 -9730 26110 -9570
rect 26240 -9730 26250 -9570
rect 16500 -9740 26250 -9730
rect 27700 -9570 35850 -9560
rect 27700 -9730 27710 -9570
rect 27840 -9730 29310 -9570
rect 29440 -9730 30910 -9570
rect 31040 -9730 32510 -9570
rect 32640 -9730 34110 -9570
rect 34240 -9730 35710 -9570
rect 35840 -9730 35850 -9570
rect 27700 -9740 35850 -9730
rect 2120 -9760 10240 -9750
rect 16500 -11370 26250 -11360
rect 2120 -11390 10240 -11380
rect 2120 -11550 2130 -11390
rect 2230 -11550 3730 -11390
rect 3830 -11550 5330 -11390
rect 5430 -11550 6930 -11390
rect 7030 -11550 8530 -11390
rect 8630 -11550 10130 -11390
rect 10230 -11550 10240 -11390
rect 16500 -11530 16510 -11370
rect 16640 -11530 18110 -11370
rect 18240 -11530 19710 -11370
rect 19840 -11530 21310 -11370
rect 21440 -11530 22910 -11370
rect 23040 -11530 24510 -11370
rect 24640 -11530 26110 -11370
rect 26240 -11530 26250 -11370
rect 16500 -11540 26250 -11530
rect 27700 -11370 35850 -11360
rect 27700 -11530 27710 -11370
rect 27840 -11530 29310 -11370
rect 29440 -11530 30910 -11370
rect 31040 -11530 32510 -11370
rect 32640 -11530 34110 -11370
rect 34240 -11530 35710 -11370
rect 35840 -11530 35850 -11370
rect 27700 -11540 35850 -11530
rect 2120 -11560 10240 -11550
rect 13280 -13170 26250 -13160
rect 2120 -13190 10240 -13180
rect 2120 -13350 2130 -13190
rect 2230 -13350 3730 -13190
rect 3830 -13350 5330 -13190
rect 5430 -13350 6930 -13190
rect 7030 -13350 8530 -13190
rect 8630 -13350 10130 -13190
rect 10230 -13350 10240 -13190
rect 2120 -13360 10240 -13350
rect 13280 -13330 13290 -13170
rect 13460 -13330 14890 -13170
rect 15060 -13330 16510 -13170
rect 16640 -13330 18110 -13170
rect 18240 -13330 19710 -13170
rect 19840 -13330 21310 -13170
rect 21440 -13330 22910 -13170
rect 23040 -13330 24510 -13170
rect 24640 -13330 26110 -13170
rect 26240 -13330 26250 -13170
rect 13280 -13340 26250 -13330
rect 27700 -13170 35850 -13160
rect 27700 -13330 27710 -13170
rect 27840 -13330 29310 -13170
rect 29440 -13330 30910 -13170
rect 31040 -13330 32510 -13170
rect 32640 -13330 34110 -13170
rect 34240 -13330 35710 -13170
rect 35840 -13330 35850 -13170
rect 27700 -13340 35850 -13330
rect 13280 -13360 15070 -13340
rect 13280 -14970 26250 -14960
rect 2120 -14990 10240 -14980
rect 2120 -15150 2130 -14990
rect 2230 -15150 3730 -14990
rect 3830 -15150 5330 -14990
rect 5430 -15150 6930 -14990
rect 7030 -15150 8530 -14990
rect 8630 -15150 10130 -14990
rect 10230 -15150 10240 -14990
rect 2120 -15160 10240 -15150
rect 13280 -15130 13290 -14970
rect 13460 -15130 14890 -14970
rect 15060 -15130 16510 -14970
rect 16640 -15130 18110 -14970
rect 18240 -15130 19710 -14970
rect 19840 -15130 21310 -14970
rect 21440 -15130 22910 -14970
rect 23040 -15130 24510 -14970
rect 24640 -15130 26110 -14970
rect 26240 -15130 26250 -14970
rect 13280 -15140 26250 -15130
rect 27700 -14970 31050 -14960
rect 27700 -15130 27710 -14970
rect 27840 -15130 29310 -14970
rect 29440 -15130 30910 -14970
rect 31040 -15130 31050 -14970
rect 27700 -15140 31050 -15130
rect 13280 -15160 15070 -15140
rect 16500 -16770 26250 -16760
rect 2120 -16790 15090 -16780
rect 2120 -16950 2130 -16790
rect 2230 -16950 3730 -16790
rect 3830 -16950 5330 -16790
rect 5430 -16950 6930 -16790
rect 7030 -16950 8530 -16790
rect 8630 -16950 10130 -16790
rect 10230 -16950 13300 -16790
rect 13450 -16950 14900 -16790
rect 15050 -16950 15090 -16790
rect 16500 -16930 16510 -16770
rect 16640 -16930 18110 -16770
rect 18240 -16930 19710 -16770
rect 19840 -16930 21310 -16770
rect 21440 -16930 22910 -16770
rect 23040 -16930 24510 -16770
rect 24640 -16930 26110 -16770
rect 26240 -16930 26250 -16770
rect 16500 -16940 26250 -16930
rect 27700 -16770 31050 -16760
rect 27700 -16930 27710 -16770
rect 27840 -16930 29310 -16770
rect 29440 -16930 30910 -16770
rect 31040 -16930 31050 -16770
rect 32510 -16770 35840 -16760
rect 32510 -16920 32520 -16770
rect 32630 -16920 34120 -16770
rect 34230 -16920 34910 -16770
rect 35050 -16920 35720 -16770
rect 35830 -16920 35840 -16770
rect 32510 -16930 35840 -16920
rect 27700 -16940 31050 -16930
rect 2120 -16960 15090 -16950
rect 16500 -18570 26250 -18560
rect 2120 -18590 15060 -18580
rect 2120 -18750 2130 -18590
rect 2230 -18750 3730 -18590
rect 3830 -18750 5330 -18590
rect 5430 -18750 6930 -18590
rect 7030 -18750 8530 -18590
rect 8630 -18750 10130 -18590
rect 10230 -18750 13300 -18590
rect 13450 -18750 14900 -18590
rect 15050 -18750 15060 -18590
rect 16500 -18730 16510 -18570
rect 16640 -18730 18110 -18570
rect 18240 -18730 19710 -18570
rect 19840 -18730 21310 -18570
rect 21440 -18730 22910 -18570
rect 23040 -18730 24510 -18570
rect 24640 -18730 26110 -18570
rect 26240 -18730 26250 -18570
rect 16500 -18740 26250 -18730
rect 27700 -18570 31050 -18560
rect 27700 -18730 27710 -18570
rect 27840 -18730 29310 -18570
rect 29440 -18730 30910 -18570
rect 31040 -18730 31050 -18570
rect 27700 -18740 31050 -18730
rect 2120 -18760 15060 -18750
rect 16500 -20370 26250 -20360
rect 2120 -20390 10240 -20380
rect 2120 -20550 2130 -20390
rect 2230 -20550 3730 -20390
rect 3830 -20550 5330 -20390
rect 5430 -20550 6930 -20390
rect 7030 -20550 8530 -20390
rect 8630 -20550 10130 -20390
rect 10230 -20550 10240 -20390
rect 16500 -20530 16510 -20370
rect 16640 -20530 18110 -20370
rect 18240 -20530 19710 -20370
rect 19840 -20530 21310 -20370
rect 21440 -20530 22910 -20370
rect 23040 -20530 24510 -20370
rect 24640 -20530 26110 -20370
rect 26240 -20530 26250 -20370
rect 16500 -20540 26250 -20530
rect 27700 -20370 35860 -20360
rect 27700 -20530 27710 -20370
rect 27840 -20530 29310 -20370
rect 29440 -20530 30910 -20370
rect 31040 -20530 32510 -20370
rect 32640 -20530 34110 -20370
rect 34240 -20530 35710 -20370
rect 35840 -20530 35860 -20370
rect 27700 -20540 35860 -20530
rect 2120 -20560 10240 -20550
rect 16500 -22170 26250 -22160
rect 2120 -22190 10240 -22180
rect 2120 -22350 2130 -22190
rect 2230 -22350 3730 -22190
rect 3830 -22350 5330 -22190
rect 5430 -22350 6930 -22190
rect 7030 -22350 8530 -22190
rect 8630 -22350 10130 -22190
rect 10230 -22350 10240 -22190
rect 16500 -22330 16510 -22170
rect 16640 -22330 18110 -22170
rect 18240 -22330 19710 -22170
rect 19840 -22330 21310 -22170
rect 21440 -22330 22910 -22170
rect 23040 -22330 24510 -22170
rect 24640 -22330 26110 -22170
rect 26240 -22330 26250 -22170
rect 16500 -22340 26250 -22330
rect 27700 -22170 31050 -22160
rect 27700 -22330 27710 -22170
rect 27840 -22330 29310 -22170
rect 29440 -22330 30910 -22170
rect 31040 -22330 31050 -22170
rect 27700 -22340 31050 -22330
rect 2120 -22360 10240 -22350
rect 480 -22400 680 -22380
rect 10120 -22440 10240 -22360
rect 10100 -22450 10260 -22440
rect 10100 -22590 10110 -22450
rect 10250 -22460 10260 -22450
rect 10250 -22470 35120 -22460
rect 10250 -22590 34910 -22470
rect 10100 -22600 10260 -22590
rect 34900 -22610 34910 -22590
rect 35050 -22590 35120 -22470
rect 35050 -22610 35060 -22590
rect 34900 -22620 35060 -22610
rect 28140 -22730 28380 -22720
rect 28990 -22730 29230 -22720
rect 11040 -22740 28150 -22730
rect 11040 -22850 11050 -22740
rect 11150 -22850 11720 -22740
rect 11820 -22850 27720 -22740
rect 27830 -22850 28150 -22740
rect 11040 -22860 28150 -22850
rect 28140 -22870 28150 -22860
rect 28370 -22740 29000 -22730
rect 28370 -22860 28630 -22740
rect 28370 -22870 28380 -22860
rect 28140 -22880 28380 -22870
rect 28620 -22870 28630 -22860
rect 28740 -22860 29000 -22740
rect 28740 -22870 28750 -22860
rect 28620 -22880 28750 -22870
rect 28990 -22870 29000 -22860
rect 29220 -22740 31040 -22730
rect 29220 -22850 29320 -22740
rect 29430 -22850 30920 -22740
rect 31030 -22850 31040 -22740
rect 29220 -22860 31040 -22850
rect 29220 -22870 29230 -22860
rect 28990 -22880 29230 -22870
rect 12410 -22980 26720 -22970
rect 12410 -23090 12420 -22980
rect 12520 -23090 26530 -22980
rect 12410 -23100 26530 -23090
rect 26520 -23160 26530 -23100
rect 26710 -23160 26720 -22980
rect 26520 -23170 26720 -23160
rect -300 -23270 20300 -23260
rect -300 -23450 1190 -23270
rect 1350 -23450 1630 -23270
rect 1810 -23450 2790 -23270
rect 2950 -23450 4390 -23270
rect 4550 -23450 5990 -23270
rect 6150 -23450 7590 -23270
rect 7750 -23450 9190 -23270
rect 9350 -23450 20110 -23270
rect 20290 -23450 20300 -23270
rect -300 -23460 20300 -23450
rect 23200 -23300 23400 -23290
rect 23200 -23480 23210 -23300
rect 23390 -23330 23400 -23300
rect 31550 -23300 31750 -23290
rect 31550 -23330 31560 -23300
rect 23390 -23460 31560 -23330
rect 23390 -23480 23400 -23460
rect 23200 -23490 23400 -23480
rect 31550 -23480 31560 -23460
rect 31740 -23480 31750 -23300
rect 31550 -23490 31750 -23480
rect -300 -23670 32010 -23660
rect -300 -23850 430 -23670
rect 610 -23850 21310 -23670
rect 21490 -23850 31820 -23670
rect 32000 -23850 32010 -23670
rect -300 -23860 32010 -23850
rect 28490 -24040 28670 -24030
rect -300 -24070 27820 -24060
rect -300 -24250 1630 -24070
rect 1810 -24250 20450 -24070
rect 20630 -24250 27630 -24070
rect 27810 -24250 27820 -24070
rect 28490 -24200 28500 -24040
rect 28660 -24200 28670 -24040
rect 28490 -24210 28670 -24200
rect 29970 -24140 30050 -24130
rect -300 -24260 27820 -24250
rect 29970 -24370 29980 -24140
rect 30040 -24210 30050 -24140
rect 30040 -24220 37030 -24210
rect 30040 -24280 34620 -24220
rect 34770 -24280 34990 -24220
rect 37020 -24280 37030 -24220
rect 30040 -24370 30050 -24280
rect 34610 -24290 37030 -24280
rect 29970 -24380 30050 -24370
rect -300 -24470 27590 -24460
rect -300 -24650 1290 -24470
rect 1470 -24650 20110 -24470
rect 20290 -24650 27400 -24470
rect 27580 -24650 27590 -24470
rect 32790 -24480 33040 -24470
rect -300 -24660 27590 -24650
rect 29370 -24490 32800 -24480
rect 29370 -24720 29380 -24490
rect 29440 -24550 32800 -24490
rect 33030 -24550 33040 -24480
rect 29440 -24720 29450 -24550
rect 32790 -24560 33040 -24550
rect 34110 -24630 34360 -24620
rect 29370 -24730 29450 -24720
rect 29520 -24640 34120 -24630
rect 23030 -24820 23570 -24810
rect 1620 -25030 1820 -25020
rect 1620 -25040 1630 -25030
rect 1600 -25100 1630 -25040
rect 1620 -25110 1630 -25100
rect 1810 -25040 1820 -25030
rect 20100 -25030 20300 -25020
rect 20100 -25040 20110 -25030
rect 1810 -25070 20110 -25040
rect 1810 -25100 2510 -25070
rect 1810 -25110 1820 -25100
rect 1620 -25120 1820 -25110
rect 2500 -25130 2510 -25100
rect 4010 -25100 4710 -25070
rect 4010 -25130 4020 -25100
rect 2500 -25140 4020 -25130
rect 4700 -25130 4710 -25100
rect 6210 -25100 6910 -25070
rect 6210 -25130 6220 -25100
rect 4700 -25140 6220 -25130
rect 6900 -25130 6910 -25100
rect 8410 -25100 9110 -25070
rect 8410 -25130 8420 -25100
rect 6900 -25140 8420 -25130
rect 9100 -25130 9110 -25100
rect 10610 -25100 11310 -25070
rect 10610 -25130 10620 -25100
rect 9100 -25140 10620 -25130
rect 11300 -25130 11310 -25100
rect 12810 -25100 13510 -25070
rect 12810 -25130 12820 -25100
rect 11300 -25140 12820 -25130
rect 13500 -25130 13510 -25100
rect 15010 -25100 15710 -25070
rect 15010 -25130 15020 -25100
rect 13500 -25140 15020 -25130
rect 15700 -25130 15710 -25100
rect 17210 -25100 17910 -25070
rect 17210 -25130 17220 -25100
rect 15700 -25140 17220 -25130
rect 17900 -25130 17910 -25100
rect 19410 -25100 20110 -25070
rect 19410 -25130 19420 -25100
rect 20100 -25110 20110 -25100
rect 20290 -25040 20300 -25030
rect 20290 -25100 20320 -25040
rect 23030 -25070 23040 -24820
rect 23560 -24880 23570 -24820
rect 29520 -24870 29530 -24640
rect 29590 -24700 34120 -24640
rect 34350 -24700 34360 -24630
rect 36860 -24640 37020 -24630
rect 36860 -24650 36870 -24640
rect 29590 -24870 29600 -24700
rect 34110 -24710 34360 -24700
rect 34800 -24660 36870 -24650
rect 30280 -24780 30520 -24770
rect 33550 -24780 33800 -24770
rect 30280 -24850 30290 -24780
rect 30510 -24850 33560 -24780
rect 33790 -24850 33800 -24780
rect 30280 -24860 30520 -24850
rect 33550 -24860 33800 -24850
rect 34800 -24860 34810 -24660
rect 34900 -24780 36870 -24660
rect 37010 -24780 37020 -24640
rect 34900 -24790 37020 -24780
rect 37120 -24640 37280 -24630
rect 37120 -24780 37130 -24640
rect 37270 -24780 37280 -24640
rect 37120 -24790 37280 -24780
rect 34900 -24860 34910 -24790
rect 34800 -24870 34910 -24860
rect 29520 -24880 29600 -24870
rect 23560 -24890 27440 -24880
rect 23560 -25070 27250 -24890
rect 27430 -25070 27440 -24890
rect 33020 -24930 33300 -24920
rect 23030 -25080 27440 -25070
rect 30120 -24940 33030 -24930
rect 20290 -25110 20300 -25100
rect 20100 -25120 20300 -25110
rect 17900 -25140 19420 -25130
rect 30120 -25170 30130 -24940
rect 30190 -25000 33030 -24940
rect 33290 -25000 33300 -24930
rect 30190 -25170 30200 -25000
rect 33020 -25010 33300 -25000
rect 33220 -25080 33500 -25070
rect 30120 -25180 30200 -25170
rect 30420 -25090 33230 -25080
rect 30420 -25320 30430 -25090
rect 30490 -25150 33230 -25090
rect 33490 -25150 33500 -25080
rect 30490 -25320 30500 -25150
rect 33220 -25160 33500 -25150
rect 30420 -25330 30500 -25320
rect 820 -25550 1020 -25540
rect 20500 -25550 20700 -25540
rect 820 -25560 830 -25550
rect -260 -25620 830 -25560
rect 820 -25630 830 -25620
rect 1010 -25560 1020 -25550
rect 2500 -25560 2700 -25550
rect 3160 -25560 3360 -25550
rect 3820 -25560 4020 -25550
rect 4700 -25560 4900 -25550
rect 5360 -25560 5560 -25550
rect 6020 -25560 6220 -25550
rect 6900 -25560 7100 -25550
rect 7560 -25560 7760 -25550
rect 8220 -25560 8420 -25550
rect 9100 -25560 9300 -25550
rect 9760 -25560 9960 -25550
rect 10420 -25560 10620 -25550
rect 11300 -25560 11500 -25550
rect 11960 -25560 12160 -25550
rect 12620 -25560 12820 -25550
rect 13500 -25560 13700 -25550
rect 14160 -25560 14360 -25550
rect 14820 -25560 15020 -25550
rect 15700 -25560 15900 -25550
rect 16360 -25560 16560 -25550
rect 17020 -25560 17220 -25550
rect 17900 -25560 18100 -25550
rect 18560 -25560 18760 -25550
rect 19220 -25560 19420 -25550
rect 20500 -25560 20510 -25550
rect 1010 -25620 6910 -25560
rect 7090 -25620 7570 -25560
rect 7750 -25620 8230 -25560
rect 8410 -25620 9110 -25560
rect 9290 -25620 9770 -25560
rect 9950 -25620 10430 -25560
rect 10610 -25620 11310 -25560
rect 11490 -25620 11970 -25560
rect 12150 -25620 12630 -25560
rect 12810 -25620 13510 -25560
rect 13690 -25620 14170 -25560
rect 14350 -25620 14830 -25560
rect 15010 -25620 20510 -25560
rect 1010 -25630 1020 -25620
rect 2500 -25630 2700 -25620
rect 3160 -25630 3360 -25620
rect 3820 -25630 4020 -25620
rect 4700 -25630 4900 -25620
rect 5360 -25630 5560 -25620
rect 6020 -25630 6220 -25620
rect 6900 -25630 7100 -25620
rect 7560 -25630 7760 -25620
rect 8220 -25630 8420 -25620
rect 9100 -25630 9300 -25620
rect 9760 -25630 9960 -25620
rect 10420 -25630 10620 -25620
rect 11300 -25630 11500 -25620
rect 11960 -25630 12160 -25620
rect 12620 -25630 12820 -25620
rect 13500 -25630 13700 -25620
rect 14160 -25630 14360 -25620
rect 14820 -25630 15020 -25620
rect 15700 -25630 15900 -25620
rect 16360 -25630 16560 -25620
rect 17020 -25630 17220 -25620
rect 17900 -25630 18100 -25620
rect 18560 -25630 18760 -25620
rect 19220 -25630 19420 -25620
rect 20500 -25630 20510 -25620
rect 20690 -25560 20700 -25550
rect 20690 -25620 22140 -25560
rect 20690 -25630 20700 -25620
rect 820 -25640 1020 -25630
rect 20500 -25640 20700 -25630
rect 1220 -25690 1420 -25680
rect 20900 -25690 21100 -25680
rect 1220 -25700 1230 -25690
rect -260 -25760 1230 -25700
rect 1220 -25770 1230 -25760
rect 1410 -25700 1420 -25690
rect 2500 -25700 2700 -25690
rect 3160 -25700 3360 -25690
rect 3820 -25700 4020 -25690
rect 4700 -25700 4900 -25690
rect 5360 -25700 5560 -25690
rect 6020 -25700 6220 -25690
rect 6900 -25700 7100 -25690
rect 7560 -25700 7760 -25690
rect 8220 -25700 8420 -25690
rect 9100 -25700 9300 -25690
rect 9760 -25700 9960 -25690
rect 10420 -25700 10620 -25690
rect 11300 -25700 11500 -25690
rect 11960 -25700 12160 -25690
rect 12620 -25700 12820 -25690
rect 13500 -25700 13700 -25690
rect 14160 -25700 14360 -25690
rect 14820 -25700 15020 -25690
rect 15700 -25700 15900 -25690
rect 16360 -25700 16560 -25690
rect 17020 -25700 17220 -25690
rect 17900 -25700 18100 -25690
rect 18560 -25700 18760 -25690
rect 19220 -25700 19420 -25690
rect 20900 -25700 20910 -25690
rect 1410 -25760 2510 -25700
rect 2690 -25760 3170 -25700
rect 3350 -25760 3830 -25700
rect 4010 -25760 4710 -25700
rect 4890 -25760 5370 -25700
rect 5550 -25760 6030 -25700
rect 6210 -25760 15710 -25700
rect 15890 -25760 16370 -25700
rect 16550 -25760 17030 -25700
rect 17210 -25760 17910 -25700
rect 18090 -25760 18570 -25700
rect 18750 -25760 19230 -25700
rect 19410 -25760 20910 -25700
rect 1410 -25770 1420 -25760
rect 2500 -25770 2700 -25760
rect 3160 -25770 3360 -25760
rect 3820 -25770 4020 -25760
rect 4700 -25770 4900 -25760
rect 5360 -25770 5560 -25760
rect 6020 -25770 6220 -25760
rect 6900 -25770 7100 -25760
rect 7560 -25770 7760 -25760
rect 8220 -25770 8420 -25760
rect 9100 -25770 9300 -25760
rect 9760 -25770 9960 -25760
rect 10420 -25770 10620 -25760
rect 11300 -25770 11500 -25760
rect 11960 -25770 12160 -25760
rect 12620 -25770 12820 -25760
rect 13500 -25770 13700 -25760
rect 14160 -25770 14360 -25760
rect 14820 -25770 15020 -25760
rect 15700 -25770 15900 -25760
rect 16360 -25770 16560 -25760
rect 17020 -25770 17220 -25760
rect 17900 -25770 18100 -25760
rect 18560 -25770 18760 -25760
rect 19220 -25770 19420 -25760
rect 20900 -25770 20910 -25760
rect 21090 -25700 21100 -25690
rect 21090 -25760 22140 -25700
rect 21090 -25770 21100 -25760
rect 1220 -25780 1420 -25770
rect 20900 -25780 21100 -25770
rect 1620 -25830 1820 -25820
rect 1620 -25840 1630 -25830
rect 1600 -25900 1630 -25840
rect 1620 -25910 1630 -25900
rect 1810 -25840 1820 -25830
rect 20100 -25830 20300 -25820
rect 20100 -25840 20110 -25830
rect 1810 -25870 20110 -25840
rect 1810 -25900 2510 -25870
rect 1810 -25910 1820 -25900
rect 1620 -25920 1820 -25910
rect 2500 -25930 2510 -25900
rect 4010 -25900 4710 -25870
rect 4010 -25930 4020 -25900
rect 2500 -25940 4020 -25930
rect 4700 -25930 4710 -25900
rect 6210 -25900 6910 -25870
rect 6210 -25930 6220 -25900
rect 4700 -25940 6220 -25930
rect 6900 -25930 6910 -25900
rect 8410 -25900 9110 -25870
rect 8410 -25930 8420 -25900
rect 6900 -25940 8420 -25930
rect 9100 -25930 9110 -25900
rect 10610 -25900 11310 -25870
rect 10610 -25930 10620 -25900
rect 9100 -25940 10620 -25930
rect 11300 -25930 11310 -25900
rect 12810 -25900 13510 -25870
rect 12810 -25930 12820 -25900
rect 11300 -25940 12820 -25930
rect 13500 -25930 13510 -25900
rect 15010 -25900 15710 -25870
rect 15010 -25930 15020 -25900
rect 13500 -25940 15020 -25930
rect 15700 -25930 15710 -25900
rect 17210 -25900 17910 -25870
rect 17210 -25930 17220 -25900
rect 15700 -25940 17220 -25930
rect 17900 -25930 17910 -25900
rect 19410 -25900 20110 -25870
rect 19410 -25930 19420 -25900
rect 20100 -25910 20110 -25900
rect 20290 -25840 20300 -25830
rect 20290 -25900 20320 -25840
rect 20290 -25910 20300 -25900
rect 20100 -25920 20300 -25910
rect 17900 -25940 19420 -25930
rect 820 -26350 1020 -26340
rect 20500 -26350 20700 -26340
rect 820 -26360 830 -26350
rect -260 -26420 830 -26360
rect 820 -26430 830 -26420
rect 1010 -26360 1020 -26350
rect 2500 -26360 2700 -26350
rect 3160 -26360 3360 -26350
rect 3820 -26360 4020 -26350
rect 4700 -26360 4900 -26350
rect 5360 -26360 5560 -26350
rect 6020 -26360 6220 -26350
rect 6900 -26360 7100 -26350
rect 7560 -26360 7760 -26350
rect 8220 -26360 8420 -26350
rect 9100 -26360 9300 -26350
rect 9760 -26360 9960 -26350
rect 10420 -26360 10620 -26350
rect 11300 -26360 11500 -26350
rect 11960 -26360 12160 -26350
rect 12620 -26360 12820 -26350
rect 13500 -26360 13700 -26350
rect 14160 -26360 14360 -26350
rect 14820 -26360 15020 -26350
rect 15700 -26360 15900 -26350
rect 16360 -26360 16560 -26350
rect 17020 -26360 17220 -26350
rect 17900 -26360 18100 -26350
rect 18560 -26360 18760 -26350
rect 19220 -26360 19420 -26350
rect 20500 -26360 20510 -26350
rect 1010 -26420 2510 -26360
rect 2690 -26420 3170 -26360
rect 3350 -26420 3830 -26360
rect 4010 -26420 4710 -26360
rect 4890 -26420 5370 -26360
rect 5550 -26420 6030 -26360
rect 6210 -26420 15710 -26360
rect 15890 -26420 16370 -26360
rect 16550 -26420 17030 -26360
rect 17210 -26420 17910 -26360
rect 18090 -26420 18570 -26360
rect 18750 -26420 19230 -26360
rect 19410 -26420 20510 -26360
rect 1010 -26430 1020 -26420
rect 2500 -26430 2700 -26420
rect 3160 -26430 3360 -26420
rect 3820 -26430 4020 -26420
rect 4700 -26430 4900 -26420
rect 5360 -26430 5560 -26420
rect 6020 -26430 6220 -26420
rect 6900 -26430 7100 -26420
rect 7560 -26430 7760 -26420
rect 8220 -26430 8420 -26420
rect 9100 -26430 9300 -26420
rect 9760 -26430 9960 -26420
rect 10420 -26430 10620 -26420
rect 11300 -26430 11500 -26420
rect 11960 -26430 12160 -26420
rect 12620 -26430 12820 -26420
rect 13500 -26430 13700 -26420
rect 14160 -26430 14360 -26420
rect 14820 -26430 15020 -26420
rect 15700 -26430 15900 -26420
rect 16360 -26430 16560 -26420
rect 17020 -26430 17220 -26420
rect 17900 -26430 18100 -26420
rect 18560 -26430 18760 -26420
rect 19220 -26430 19420 -26420
rect 20500 -26430 20510 -26420
rect 20690 -26360 20700 -26350
rect 20690 -26420 22140 -26360
rect 20690 -26430 20700 -26420
rect 820 -26440 1020 -26430
rect 20500 -26440 20700 -26430
rect 1220 -26490 1420 -26480
rect 20900 -26490 21100 -26480
rect 1220 -26500 1230 -26490
rect -260 -26560 1230 -26500
rect 1220 -26570 1230 -26560
rect 1410 -26500 1420 -26490
rect 2500 -26500 2700 -26490
rect 3160 -26500 3360 -26490
rect 3820 -26500 4020 -26490
rect 4700 -26500 4900 -26490
rect 5360 -26500 5560 -26490
rect 6020 -26500 6220 -26490
rect 6900 -26500 7100 -26490
rect 7560 -26500 7760 -26490
rect 8220 -26500 8420 -26490
rect 9100 -26500 9300 -26490
rect 9760 -26500 9960 -26490
rect 10420 -26500 10620 -26490
rect 11300 -26500 11500 -26490
rect 11960 -26500 12160 -26490
rect 12620 -26500 12820 -26490
rect 13500 -26500 13700 -26490
rect 14160 -26500 14360 -26490
rect 14820 -26500 15020 -26490
rect 15700 -26500 15900 -26490
rect 16360 -26500 16560 -26490
rect 17020 -26500 17220 -26490
rect 17900 -26500 18100 -26490
rect 18560 -26500 18760 -26490
rect 19220 -26500 19420 -26490
rect 20900 -26500 20910 -26490
rect 1410 -26560 6910 -26500
rect 7090 -26560 7570 -26500
rect 7750 -26560 8230 -26500
rect 8410 -26560 9110 -26500
rect 9290 -26560 9770 -26500
rect 9950 -26560 10430 -26500
rect 10610 -26560 11310 -26500
rect 11490 -26560 11970 -26500
rect 12150 -26560 12630 -26500
rect 12810 -26560 13510 -26500
rect 13690 -26560 14170 -26500
rect 14350 -26560 14830 -26500
rect 15010 -26560 20910 -26500
rect 1410 -26570 1420 -26560
rect 2500 -26570 2700 -26560
rect 3160 -26570 3360 -26560
rect 3820 -26570 4020 -26560
rect 4700 -26570 4900 -26560
rect 5360 -26570 5560 -26560
rect 6020 -26570 6220 -26560
rect 6900 -26570 7100 -26560
rect 7560 -26570 7760 -26560
rect 8220 -26570 8420 -26560
rect 9100 -26570 9300 -26560
rect 9760 -26570 9960 -26560
rect 10420 -26570 10620 -26560
rect 11300 -26570 11500 -26560
rect 11960 -26570 12160 -26560
rect 12620 -26570 12820 -26560
rect 13500 -26570 13700 -26560
rect 14160 -26570 14360 -26560
rect 14820 -26570 15020 -26560
rect 15700 -26570 15900 -26560
rect 16360 -26570 16560 -26560
rect 17020 -26570 17220 -26560
rect 17900 -26570 18100 -26560
rect 18560 -26570 18760 -26560
rect 19220 -26570 19420 -26560
rect 20900 -26570 20910 -26560
rect 21090 -26500 21100 -26490
rect 21090 -26560 22140 -26500
rect 21090 -26570 21100 -26560
rect 1220 -26580 1420 -26570
rect 20900 -26580 21100 -26570
rect 420 -26630 620 -26620
rect 420 -26710 430 -26630
rect 610 -26710 620 -26630
rect 1620 -26630 1820 -26620
rect 1620 -26640 1630 -26630
rect 1600 -26700 1630 -26640
rect 420 -26720 620 -26710
rect 1620 -26710 1630 -26700
rect 1810 -26640 1820 -26630
rect 20100 -26630 20300 -26620
rect 20100 -26640 20110 -26630
rect 1810 -26670 20110 -26640
rect 1810 -26700 4710 -26670
rect 1810 -26710 1820 -26700
rect 1620 -26720 1820 -26710
rect 4700 -26730 4710 -26700
rect 6210 -26700 6910 -26670
rect 6210 -26730 6220 -26700
rect 4700 -26740 6220 -26730
rect 6900 -26730 6910 -26700
rect 8410 -26700 9110 -26670
rect 8410 -26730 8420 -26700
rect 6900 -26740 8420 -26730
rect 9100 -26730 9110 -26700
rect 10610 -26700 11310 -26670
rect 10610 -26730 10620 -26700
rect 9100 -26740 10620 -26730
rect 11300 -26730 11310 -26700
rect 12810 -26700 13510 -26670
rect 12810 -26730 12820 -26700
rect 11300 -26740 12820 -26730
rect 13500 -26730 13510 -26700
rect 15010 -26700 15710 -26670
rect 15010 -26730 15020 -26700
rect 13500 -26740 15020 -26730
rect 15700 -26730 15710 -26700
rect 17210 -26700 20110 -26670
rect 17210 -26730 17220 -26700
rect 20100 -26710 20110 -26700
rect 20290 -26640 20300 -26630
rect 21300 -26630 21500 -26620
rect 20290 -26700 20320 -26640
rect 20290 -26710 20300 -26700
rect 20100 -26720 20300 -26710
rect 21300 -26710 21310 -26630
rect 21490 -26710 21500 -26630
rect 21300 -26720 21500 -26710
rect 15700 -26740 17220 -26730
rect 36020 -27010 36420 -27000
rect 36020 -27140 36030 -27010
rect 36410 -27140 36420 -27010
rect 820 -27150 1020 -27140
rect 20500 -27150 20700 -27140
rect 36020 -27150 36420 -27140
rect 36520 -27010 36920 -27000
rect 36520 -27140 36530 -27010
rect 36910 -27140 36920 -27010
rect 36520 -27150 36920 -27140
rect 820 -27160 830 -27150
rect -260 -27220 830 -27160
rect 820 -27230 830 -27220
rect 1010 -27160 1020 -27150
rect 2500 -27160 2700 -27150
rect 3160 -27160 3360 -27150
rect 3820 -27160 4020 -27150
rect 4700 -27160 4900 -27150
rect 5360 -27160 5560 -27150
rect 6020 -27160 6220 -27150
rect 6900 -27160 7100 -27150
rect 7560 -27160 7760 -27150
rect 8220 -27160 8420 -27150
rect 9100 -27160 9300 -27150
rect 9760 -27160 9960 -27150
rect 10420 -27160 10620 -27150
rect 11300 -27160 11500 -27150
rect 11960 -27160 12160 -27150
rect 12620 -27160 12820 -27150
rect 13500 -27160 13700 -27150
rect 14160 -27160 14360 -27150
rect 14820 -27160 15020 -27150
rect 15700 -27160 15900 -27150
rect 16360 -27160 16560 -27150
rect 17020 -27160 17220 -27150
rect 17900 -27160 18100 -27150
rect 18560 -27160 18760 -27150
rect 19220 -27160 19420 -27150
rect 20500 -27160 20510 -27150
rect 1010 -27220 6910 -27160
rect 7090 -27220 7570 -27160
rect 7750 -27220 8230 -27160
rect 8410 -27220 9110 -27160
rect 9290 -27220 9770 -27160
rect 9950 -27220 10430 -27160
rect 10610 -27220 11310 -27160
rect 11490 -27220 11970 -27160
rect 12150 -27220 12630 -27160
rect 12810 -27220 13510 -27160
rect 13690 -27220 14170 -27160
rect 14350 -27220 14830 -27160
rect 15010 -27220 20510 -27160
rect 1010 -27230 1020 -27220
rect 2500 -27230 2700 -27220
rect 3160 -27230 3360 -27220
rect 3820 -27230 4020 -27220
rect 4700 -27230 4900 -27220
rect 5360 -27230 5560 -27220
rect 6020 -27230 6220 -27220
rect 6900 -27230 7100 -27220
rect 7560 -27230 7760 -27220
rect 8220 -27230 8420 -27220
rect 9100 -27230 9300 -27220
rect 9760 -27230 9960 -27220
rect 10420 -27230 10620 -27220
rect 11300 -27230 11500 -27220
rect 11960 -27230 12160 -27220
rect 12620 -27230 12820 -27220
rect 13500 -27230 13700 -27220
rect 14160 -27230 14360 -27220
rect 14820 -27230 15020 -27220
rect 15700 -27230 15900 -27220
rect 16360 -27230 16560 -27220
rect 17020 -27230 17220 -27220
rect 17900 -27230 18100 -27220
rect 18560 -27230 18760 -27220
rect 19220 -27230 19420 -27220
rect 20500 -27230 20510 -27220
rect 20690 -27160 20700 -27150
rect 20690 -27220 22140 -27160
rect 20690 -27230 20700 -27220
rect 820 -27240 1020 -27230
rect 20500 -27240 20700 -27230
rect 1220 -27290 1420 -27280
rect 20900 -27290 21100 -27280
rect 1220 -27300 1230 -27290
rect -260 -27360 1230 -27300
rect 1220 -27370 1230 -27360
rect 1410 -27300 1420 -27290
rect 2500 -27300 2700 -27290
rect 3160 -27300 3360 -27290
rect 3820 -27300 4020 -27290
rect 4700 -27300 4900 -27290
rect 5360 -27300 5560 -27290
rect 6020 -27300 6220 -27290
rect 6900 -27300 7100 -27290
rect 7560 -27300 7760 -27290
rect 8220 -27300 8420 -27290
rect 9100 -27300 9300 -27290
rect 9760 -27300 9960 -27290
rect 10420 -27300 10620 -27290
rect 11300 -27300 11500 -27290
rect 11960 -27300 12160 -27290
rect 12620 -27300 12820 -27290
rect 13500 -27300 13700 -27290
rect 14160 -27300 14360 -27290
rect 14820 -27300 15020 -27290
rect 15700 -27300 15900 -27290
rect 16360 -27300 16560 -27290
rect 17020 -27300 17220 -27290
rect 17900 -27300 18100 -27290
rect 18560 -27300 18760 -27290
rect 19220 -27300 19420 -27290
rect 20900 -27300 20910 -27290
rect 1410 -27360 2510 -27300
rect 2690 -27360 3170 -27300
rect 3350 -27360 3830 -27300
rect 4010 -27360 4710 -27300
rect 4890 -27360 5370 -27300
rect 5550 -27360 6030 -27300
rect 6210 -27360 15710 -27300
rect 15890 -27360 16370 -27300
rect 16550 -27360 17030 -27300
rect 17210 -27360 17910 -27300
rect 18090 -27360 18570 -27300
rect 18750 -27360 19230 -27300
rect 19410 -27360 20910 -27300
rect 1410 -27370 1420 -27360
rect 2500 -27370 2700 -27360
rect 3160 -27370 3360 -27360
rect 3820 -27370 4020 -27360
rect 4700 -27370 4900 -27360
rect 5360 -27370 5560 -27360
rect 6020 -27370 6220 -27360
rect 6900 -27370 7100 -27360
rect 7560 -27370 7760 -27360
rect 8220 -27370 8420 -27360
rect 9100 -27370 9300 -27360
rect 9760 -27370 9960 -27360
rect 10420 -27370 10620 -27360
rect 11300 -27370 11500 -27360
rect 11960 -27370 12160 -27360
rect 12620 -27370 12820 -27360
rect 13500 -27370 13700 -27360
rect 14160 -27370 14360 -27360
rect 14820 -27370 15020 -27360
rect 15700 -27370 15900 -27360
rect 16360 -27370 16560 -27360
rect 17020 -27370 17220 -27360
rect 17900 -27370 18100 -27360
rect 18560 -27370 18760 -27360
rect 19220 -27370 19420 -27360
rect 20900 -27370 20910 -27360
rect 21090 -27300 21100 -27290
rect 21090 -27360 22140 -27300
rect 21090 -27370 21100 -27360
rect 1220 -27380 1420 -27370
rect 20900 -27380 21100 -27370
rect 420 -27430 620 -27420
rect 420 -27510 430 -27430
rect 610 -27510 620 -27430
rect 1620 -27430 1820 -27420
rect 1620 -27440 1630 -27430
rect 1600 -27500 1630 -27440
rect 420 -27520 620 -27510
rect 1620 -27510 1630 -27500
rect 1810 -27440 1820 -27430
rect 20100 -27430 20300 -27420
rect 20100 -27440 20110 -27430
rect 1810 -27470 20110 -27440
rect 1810 -27500 4710 -27470
rect 1810 -27510 1820 -27500
rect 1620 -27520 1820 -27510
rect 4700 -27530 4710 -27500
rect 6210 -27500 6910 -27470
rect 6210 -27530 6220 -27500
rect 4700 -27540 6220 -27530
rect 6900 -27530 6910 -27500
rect 8410 -27500 9110 -27470
rect 8410 -27530 8420 -27500
rect 6900 -27540 8420 -27530
rect 9100 -27530 9110 -27500
rect 10610 -27500 11310 -27470
rect 10610 -27530 10620 -27500
rect 9100 -27540 10620 -27530
rect 11300 -27530 11310 -27500
rect 12810 -27500 13510 -27470
rect 12810 -27530 12820 -27500
rect 11300 -27540 12820 -27530
rect 13500 -27530 13510 -27500
rect 15010 -27500 15710 -27470
rect 15010 -27530 15020 -27500
rect 13500 -27540 15020 -27530
rect 15700 -27530 15710 -27500
rect 17210 -27500 20110 -27470
rect 17210 -27530 17220 -27500
rect 20100 -27510 20110 -27500
rect 20290 -27440 20300 -27430
rect 21300 -27430 21500 -27420
rect 20290 -27500 20320 -27440
rect 20290 -27510 20300 -27500
rect 20100 -27520 20300 -27510
rect 21300 -27510 21310 -27430
rect 21490 -27510 21500 -27430
rect 21300 -27520 21500 -27510
rect 15700 -27540 17220 -27530
rect 36900 -27540 37700 -27520
rect 36900 -27900 36920 -27540
rect 37680 -27900 37700 -27540
rect 36900 -27920 37700 -27900
rect 820 -27950 1020 -27940
rect 20500 -27950 20700 -27940
rect 820 -27960 830 -27950
rect -260 -28020 830 -27960
rect 820 -28030 830 -28020
rect 1010 -27960 1020 -27950
rect 2500 -27960 2700 -27950
rect 3160 -27960 3360 -27950
rect 3820 -27960 4020 -27950
rect 4700 -27960 4900 -27950
rect 5360 -27960 5560 -27950
rect 6020 -27960 6220 -27950
rect 6900 -27960 7100 -27950
rect 7560 -27960 7760 -27950
rect 8220 -27960 8420 -27950
rect 9100 -27960 9300 -27950
rect 9760 -27960 9960 -27950
rect 10420 -27960 10620 -27950
rect 11300 -27960 11500 -27950
rect 11960 -27960 12160 -27950
rect 12620 -27960 12820 -27950
rect 13500 -27960 13700 -27950
rect 14160 -27960 14360 -27950
rect 14820 -27960 15020 -27950
rect 15700 -27960 15900 -27950
rect 16360 -27960 16560 -27950
rect 17020 -27960 17220 -27950
rect 17900 -27960 18100 -27950
rect 18560 -27960 18760 -27950
rect 19220 -27960 19420 -27950
rect 20500 -27960 20510 -27950
rect 1010 -28020 2510 -27960
rect 2690 -28020 3170 -27960
rect 3350 -28020 3830 -27960
rect 4010 -28020 4710 -27960
rect 4890 -28020 5370 -27960
rect 5550 -28020 6030 -27960
rect 6210 -28020 15710 -27960
rect 15890 -28020 16370 -27960
rect 16550 -28020 17030 -27960
rect 17210 -28020 17910 -27960
rect 18090 -28020 18570 -27960
rect 18750 -28020 19230 -27960
rect 19410 -28020 20510 -27960
rect 1010 -28030 1020 -28020
rect 2500 -28030 2700 -28020
rect 3160 -28030 3360 -28020
rect 3820 -28030 4020 -28020
rect 4700 -28030 4900 -28020
rect 5360 -28030 5560 -28020
rect 6020 -28030 6220 -28020
rect 6900 -28030 7100 -28020
rect 7560 -28030 7760 -28020
rect 8220 -28030 8420 -28020
rect 9100 -28030 9300 -28020
rect 9760 -28030 9960 -28020
rect 10420 -28030 10620 -28020
rect 11300 -28030 11500 -28020
rect 11960 -28030 12160 -28020
rect 12620 -28030 12820 -28020
rect 13500 -28030 13700 -28020
rect 14160 -28030 14360 -28020
rect 14820 -28030 15020 -28020
rect 15700 -28030 15900 -28020
rect 16360 -28030 16560 -28020
rect 17020 -28030 17220 -28020
rect 17900 -28030 18100 -28020
rect 18560 -28030 18760 -28020
rect 19220 -28030 19420 -28020
rect 20500 -28030 20510 -28020
rect 20690 -27960 20700 -27950
rect 20690 -28020 22140 -27960
rect 20690 -28030 20700 -28020
rect 820 -28040 1020 -28030
rect 20500 -28040 20700 -28030
rect 1220 -28090 1420 -28080
rect 20900 -28090 21100 -28080
rect 1220 -28100 1230 -28090
rect -260 -28160 1230 -28100
rect 1220 -28170 1230 -28160
rect 1410 -28100 1420 -28090
rect 2500 -28100 2700 -28090
rect 3160 -28100 3360 -28090
rect 3820 -28100 4020 -28090
rect 4700 -28100 4900 -28090
rect 5360 -28100 5560 -28090
rect 6020 -28100 6220 -28090
rect 6900 -28100 7100 -28090
rect 7560 -28100 7760 -28090
rect 8220 -28100 8420 -28090
rect 9100 -28100 9300 -28090
rect 9760 -28100 9960 -28090
rect 10420 -28100 10620 -28090
rect 11300 -28100 11500 -28090
rect 11960 -28100 12160 -28090
rect 12620 -28100 12820 -28090
rect 13500 -28100 13700 -28090
rect 14160 -28100 14360 -28090
rect 14820 -28100 15020 -28090
rect 15700 -28100 15900 -28090
rect 16360 -28100 16560 -28090
rect 17020 -28100 17220 -28090
rect 17900 -28100 18100 -28090
rect 18560 -28100 18760 -28090
rect 19220 -28100 19420 -28090
rect 20900 -28100 20910 -28090
rect 1410 -28160 6910 -28100
rect 7090 -28160 7570 -28100
rect 7750 -28160 8230 -28100
rect 8410 -28160 9110 -28100
rect 9290 -28160 9770 -28100
rect 9950 -28160 10430 -28100
rect 10610 -28160 11310 -28100
rect 11490 -28160 11970 -28100
rect 12150 -28160 12630 -28100
rect 12810 -28160 13510 -28100
rect 13690 -28160 14170 -28100
rect 14350 -28160 14830 -28100
rect 15010 -28160 20910 -28100
rect 1410 -28170 1420 -28160
rect 2500 -28170 2700 -28160
rect 3160 -28170 3360 -28160
rect 3820 -28170 4020 -28160
rect 4700 -28170 4900 -28160
rect 5360 -28170 5560 -28160
rect 6020 -28170 6220 -28160
rect 6900 -28170 7100 -28160
rect 7560 -28170 7760 -28160
rect 8220 -28170 8420 -28160
rect 9100 -28170 9300 -28160
rect 9760 -28170 9960 -28160
rect 10420 -28170 10620 -28160
rect 11300 -28170 11500 -28160
rect 11960 -28170 12160 -28160
rect 12620 -28170 12820 -28160
rect 13500 -28170 13700 -28160
rect 14160 -28170 14360 -28160
rect 14820 -28170 15020 -28160
rect 15700 -28170 15900 -28160
rect 16360 -28170 16560 -28160
rect 17020 -28170 17220 -28160
rect 17900 -28170 18100 -28160
rect 18560 -28170 18760 -28160
rect 19220 -28170 19420 -28160
rect 20900 -28170 20910 -28160
rect 21090 -28100 21100 -28090
rect 21090 -28160 22140 -28100
rect 36900 -28160 37700 -28140
rect 21090 -28170 21100 -28160
rect 1220 -28180 1420 -28170
rect 20900 -28180 21100 -28170
rect 420 -28230 620 -28220
rect 420 -28310 430 -28230
rect 610 -28310 620 -28230
rect 1620 -28230 1820 -28220
rect 1620 -28240 1630 -28230
rect 1600 -28300 1630 -28240
rect 420 -28320 620 -28310
rect 1620 -28310 1630 -28300
rect 1810 -28240 1820 -28230
rect 20100 -28230 20300 -28220
rect 20100 -28240 20110 -28230
rect 1810 -28270 20110 -28240
rect 1810 -28300 4710 -28270
rect 1810 -28310 1820 -28300
rect 1620 -28320 1820 -28310
rect 4700 -28330 4710 -28300
rect 6210 -28300 6910 -28270
rect 6210 -28330 6220 -28300
rect 4700 -28340 6220 -28330
rect 6900 -28330 6910 -28300
rect 8410 -28300 9110 -28270
rect 8410 -28330 8420 -28300
rect 6900 -28340 8420 -28330
rect 9100 -28330 9110 -28300
rect 10610 -28300 11310 -28270
rect 10610 -28330 10620 -28300
rect 9100 -28340 10620 -28330
rect 11300 -28330 11310 -28300
rect 12810 -28300 13510 -28270
rect 12810 -28330 12820 -28300
rect 11300 -28340 12820 -28330
rect 13500 -28330 13510 -28300
rect 15010 -28300 15710 -28270
rect 15010 -28330 15020 -28300
rect 13500 -28340 15020 -28330
rect 15700 -28330 15710 -28300
rect 17210 -28300 20110 -28270
rect 17210 -28330 17220 -28300
rect 20100 -28310 20110 -28300
rect 20290 -28240 20300 -28230
rect 21300 -28230 21500 -28220
rect 20290 -28300 20320 -28240
rect 20290 -28310 20300 -28300
rect 20100 -28320 20300 -28310
rect 21300 -28310 21310 -28230
rect 21490 -28310 21500 -28230
rect 21300 -28320 21500 -28310
rect 15700 -28340 17220 -28330
rect 36900 -28520 36920 -28160
rect 37680 -28520 37700 -28160
rect 36900 -28540 37700 -28520
rect 36020 -28710 36280 -28700
rect 29670 -28720 36030 -28710
rect 820 -28750 1020 -28740
rect 20500 -28750 20700 -28740
rect 820 -28760 830 -28750
rect -260 -28820 830 -28760
rect 820 -28830 830 -28820
rect 1010 -28760 1020 -28750
rect 2500 -28760 2700 -28750
rect 3160 -28760 3360 -28750
rect 3820 -28760 4020 -28750
rect 4700 -28760 4900 -28750
rect 5360 -28760 5560 -28750
rect 6020 -28760 6220 -28750
rect 6900 -28760 7100 -28750
rect 7560 -28760 7760 -28750
rect 8220 -28760 8420 -28750
rect 9100 -28760 9300 -28750
rect 9760 -28760 9960 -28750
rect 10420 -28760 10620 -28750
rect 11300 -28760 11500 -28750
rect 11960 -28760 12160 -28750
rect 12620 -28760 12820 -28750
rect 13500 -28760 13700 -28750
rect 14160 -28760 14360 -28750
rect 14820 -28760 15020 -28750
rect 15700 -28760 15900 -28750
rect 16360 -28760 16560 -28750
rect 17020 -28760 17220 -28750
rect 17900 -28760 18100 -28750
rect 18560 -28760 18760 -28750
rect 19220 -28760 19420 -28750
rect 20500 -28760 20510 -28750
rect 1010 -28820 2510 -28760
rect 2690 -28820 3170 -28760
rect 3350 -28820 3830 -28760
rect 4010 -28820 4710 -28760
rect 4890 -28820 5370 -28760
rect 5550 -28820 6030 -28760
rect 6210 -28820 15710 -28760
rect 15890 -28820 16370 -28760
rect 16550 -28820 17030 -28760
rect 17210 -28820 17910 -28760
rect 18090 -28820 18570 -28760
rect 18750 -28820 19230 -28760
rect 19410 -28820 20510 -28760
rect 1010 -28830 1020 -28820
rect 2500 -28830 2700 -28820
rect 3160 -28830 3360 -28820
rect 3820 -28830 4020 -28820
rect 4700 -28830 4900 -28820
rect 5360 -28830 5560 -28820
rect 6020 -28830 6220 -28820
rect 6900 -28830 7100 -28820
rect 7560 -28830 7760 -28820
rect 8220 -28830 8420 -28820
rect 9100 -28830 9300 -28820
rect 9760 -28830 9960 -28820
rect 10420 -28830 10620 -28820
rect 11300 -28830 11500 -28820
rect 11960 -28830 12160 -28820
rect 12620 -28830 12820 -28820
rect 13500 -28830 13700 -28820
rect 14160 -28830 14360 -28820
rect 14820 -28830 15020 -28820
rect 15700 -28830 15900 -28820
rect 16360 -28830 16560 -28820
rect 17020 -28830 17220 -28820
rect 17900 -28830 18100 -28820
rect 18560 -28830 18760 -28820
rect 19220 -28830 19420 -28820
rect 20500 -28830 20510 -28820
rect 20690 -28760 20700 -28750
rect 20690 -28820 22140 -28760
rect 20690 -28830 20700 -28820
rect 820 -28840 1020 -28830
rect 20500 -28840 20700 -28830
rect 1220 -28890 1420 -28880
rect 20900 -28890 21100 -28880
rect 1220 -28900 1230 -28890
rect -260 -28960 1230 -28900
rect 1220 -28970 1230 -28960
rect 1410 -28900 1420 -28890
rect 2500 -28900 2700 -28890
rect 3160 -28900 3360 -28890
rect 3820 -28900 4020 -28890
rect 4700 -28900 4900 -28890
rect 5360 -28900 5560 -28890
rect 6020 -28900 6220 -28890
rect 6900 -28900 7100 -28890
rect 7560 -28900 7760 -28890
rect 8220 -28900 8420 -28890
rect 9100 -28900 9300 -28890
rect 9760 -28900 9960 -28890
rect 10420 -28900 10620 -28890
rect 11300 -28900 11500 -28890
rect 11960 -28900 12160 -28890
rect 12620 -28900 12820 -28890
rect 13500 -28900 13700 -28890
rect 14160 -28900 14360 -28890
rect 14820 -28900 15020 -28890
rect 15700 -28900 15900 -28890
rect 16360 -28900 16560 -28890
rect 17020 -28900 17220 -28890
rect 17900 -28900 18100 -28890
rect 18560 -28900 18760 -28890
rect 19220 -28900 19420 -28890
rect 20900 -28900 20910 -28890
rect 1410 -28960 6910 -28900
rect 7090 -28960 7570 -28900
rect 7750 -28960 8230 -28900
rect 8410 -28960 9110 -28900
rect 9290 -28960 9770 -28900
rect 9950 -28960 10430 -28900
rect 10610 -28960 11310 -28900
rect 11490 -28960 11970 -28900
rect 12150 -28960 12630 -28900
rect 12810 -28960 13510 -28900
rect 13690 -28960 14170 -28900
rect 14350 -28960 14830 -28900
rect 15010 -28960 20910 -28900
rect 1410 -28970 1420 -28960
rect 2500 -28970 2700 -28960
rect 3160 -28970 3360 -28960
rect 3820 -28970 4020 -28960
rect 4700 -28970 4900 -28960
rect 5360 -28970 5560 -28960
rect 6020 -28970 6220 -28960
rect 6900 -28970 7100 -28960
rect 7560 -28970 7760 -28960
rect 8220 -28970 8420 -28960
rect 9100 -28970 9300 -28960
rect 9760 -28970 9960 -28960
rect 10420 -28970 10620 -28960
rect 11300 -28970 11500 -28960
rect 11960 -28970 12160 -28960
rect 12620 -28970 12820 -28960
rect 13500 -28970 13700 -28960
rect 14160 -28970 14360 -28960
rect 14820 -28970 15020 -28960
rect 15700 -28970 15900 -28960
rect 16360 -28970 16560 -28960
rect 17020 -28970 17220 -28960
rect 17900 -28970 18100 -28960
rect 18560 -28970 18760 -28960
rect 19220 -28970 19420 -28960
rect 20900 -28970 20910 -28960
rect 21090 -28900 21100 -28890
rect 21090 -28960 22140 -28900
rect 29670 -28940 29680 -28720
rect 29740 -28780 36030 -28720
rect 36270 -28780 38310 -28710
rect 29740 -28940 29750 -28780
rect 36020 -28790 36280 -28780
rect 35680 -28860 35940 -28850
rect 29670 -28950 29750 -28940
rect 29820 -28870 35690 -28860
rect 21090 -28970 21100 -28960
rect 1220 -28980 1420 -28970
rect 20900 -28980 21100 -28970
rect 420 -29030 620 -29020
rect 420 -29110 430 -29030
rect 610 -29110 620 -29030
rect 1620 -29030 1820 -29020
rect 1620 -29040 1630 -29030
rect 1600 -29100 1630 -29040
rect 420 -29120 620 -29110
rect 1620 -29110 1630 -29100
rect 1810 -29040 1820 -29030
rect 20100 -29030 20300 -29020
rect 20100 -29040 20110 -29030
rect 1810 -29070 20110 -29040
rect 1810 -29100 4710 -29070
rect 1810 -29110 1820 -29100
rect 1620 -29120 1820 -29110
rect 4700 -29130 4710 -29100
rect 6210 -29100 6910 -29070
rect 6210 -29130 6220 -29100
rect 4700 -29140 6220 -29130
rect 6900 -29130 6910 -29100
rect 8410 -29100 9110 -29070
rect 8410 -29130 8420 -29100
rect 6900 -29140 8420 -29130
rect 9100 -29130 9110 -29100
rect 10610 -29100 11310 -29070
rect 10610 -29130 10620 -29100
rect 9100 -29140 10620 -29130
rect 11300 -29130 11310 -29100
rect 12810 -29100 13510 -29070
rect 12810 -29130 12820 -29100
rect 11300 -29140 12820 -29130
rect 13500 -29130 13510 -29100
rect 15010 -29100 15710 -29070
rect 15010 -29130 15020 -29100
rect 13500 -29140 15020 -29130
rect 15700 -29130 15710 -29100
rect 17210 -29100 20110 -29070
rect 17210 -29130 17220 -29100
rect 20100 -29110 20110 -29100
rect 20290 -29040 20300 -29030
rect 21300 -29030 21500 -29020
rect 20290 -29100 20320 -29040
rect 20290 -29110 20300 -29100
rect 20100 -29120 20300 -29110
rect 21300 -29110 21310 -29030
rect 21490 -29110 21500 -29030
rect 29820 -29090 29830 -28870
rect 29890 -28930 35690 -28870
rect 35930 -28930 38310 -28860
rect 29890 -29090 29900 -28930
rect 35680 -28940 35940 -28930
rect 37020 -29010 37280 -29000
rect 29820 -29100 29900 -29090
rect 29970 -29020 37030 -29010
rect 21300 -29120 21500 -29110
rect 15700 -29140 17220 -29130
rect 29970 -29240 29980 -29020
rect 30040 -29080 37030 -29020
rect 37270 -29080 38310 -29010
rect 30040 -29240 30050 -29080
rect 37020 -29090 37280 -29080
rect 36690 -29160 36950 -29150
rect 29970 -29250 30050 -29240
rect 30120 -29170 36700 -29160
rect 30120 -29390 30130 -29170
rect 30190 -29230 36700 -29170
rect 36940 -29230 38310 -29160
rect 30190 -29390 30200 -29230
rect 36690 -29240 36950 -29230
rect 38020 -29310 38280 -29300
rect 30120 -29400 30200 -29390
rect 30270 -29320 38030 -29310
rect 30270 -29540 30280 -29320
rect 30340 -29380 38030 -29320
rect 38270 -29380 38310 -29310
rect 30340 -29540 30350 -29380
rect 38020 -29390 38280 -29380
rect 37690 -29460 37950 -29450
rect 820 -29550 1020 -29540
rect 20500 -29550 20700 -29540
rect 30270 -29550 30350 -29540
rect 30420 -29470 37700 -29460
rect 820 -29560 830 -29550
rect -260 -29620 830 -29560
rect 820 -29630 830 -29620
rect 1010 -29560 1020 -29550
rect 2500 -29560 2700 -29550
rect 3160 -29560 3360 -29550
rect 3820 -29560 4020 -29550
rect 4700 -29560 4900 -29550
rect 5360 -29560 5560 -29550
rect 6020 -29560 6220 -29550
rect 6900 -29560 7100 -29550
rect 7560 -29560 7760 -29550
rect 8220 -29560 8420 -29550
rect 9100 -29560 9300 -29550
rect 9760 -29560 9960 -29550
rect 10420 -29560 10620 -29550
rect 11300 -29560 11500 -29550
rect 11960 -29560 12160 -29550
rect 12620 -29560 12820 -29550
rect 13500 -29560 13700 -29550
rect 14160 -29560 14360 -29550
rect 14820 -29560 15020 -29550
rect 15700 -29560 15900 -29550
rect 16360 -29560 16560 -29550
rect 17020 -29560 17220 -29550
rect 17900 -29560 18100 -29550
rect 18560 -29560 18760 -29550
rect 19220 -29560 19420 -29550
rect 20500 -29560 20510 -29550
rect 1010 -29620 6910 -29560
rect 7090 -29620 7570 -29560
rect 7750 -29620 8230 -29560
rect 8410 -29620 9110 -29560
rect 9290 -29620 9770 -29560
rect 9950 -29620 10430 -29560
rect 10610 -29620 11310 -29560
rect 11490 -29620 11970 -29560
rect 12150 -29620 12630 -29560
rect 12810 -29620 13510 -29560
rect 13690 -29620 14170 -29560
rect 14350 -29620 14830 -29560
rect 15010 -29620 20510 -29560
rect 1010 -29630 1020 -29620
rect 2500 -29630 2700 -29620
rect 3160 -29630 3360 -29620
rect 3820 -29630 4020 -29620
rect 4700 -29630 4900 -29620
rect 5360 -29630 5560 -29620
rect 6020 -29630 6220 -29620
rect 6900 -29630 7100 -29620
rect 7560 -29630 7760 -29620
rect 8220 -29630 8420 -29620
rect 9100 -29630 9300 -29620
rect 9760 -29630 9960 -29620
rect 10420 -29630 10620 -29620
rect 11300 -29630 11500 -29620
rect 11960 -29630 12160 -29620
rect 12620 -29630 12820 -29620
rect 13500 -29630 13700 -29620
rect 14160 -29630 14360 -29620
rect 14820 -29630 15020 -29620
rect 15700 -29630 15900 -29620
rect 16360 -29630 16560 -29620
rect 17020 -29630 17220 -29620
rect 17900 -29630 18100 -29620
rect 18560 -29630 18760 -29620
rect 19220 -29630 19420 -29620
rect 20500 -29630 20510 -29620
rect 20690 -29560 20700 -29550
rect 20690 -29620 22140 -29560
rect 20690 -29630 20700 -29620
rect 820 -29640 1020 -29630
rect 20500 -29640 20700 -29630
rect 1220 -29690 1420 -29680
rect 20900 -29690 21100 -29680
rect 1220 -29700 1230 -29690
rect -260 -29760 1230 -29700
rect 1220 -29770 1230 -29760
rect 1410 -29700 1420 -29690
rect 2500 -29700 2700 -29690
rect 3160 -29700 3360 -29690
rect 3820 -29700 4020 -29690
rect 4700 -29700 4900 -29690
rect 5360 -29700 5560 -29690
rect 6020 -29700 6220 -29690
rect 6900 -29700 7100 -29690
rect 7560 -29700 7760 -29690
rect 8220 -29700 8420 -29690
rect 9100 -29700 9300 -29690
rect 9760 -29700 9960 -29690
rect 10420 -29700 10620 -29690
rect 11300 -29700 11500 -29690
rect 11960 -29700 12160 -29690
rect 12620 -29700 12820 -29690
rect 13500 -29700 13700 -29690
rect 14160 -29700 14360 -29690
rect 14820 -29700 15020 -29690
rect 15700 -29700 15900 -29690
rect 16360 -29700 16560 -29690
rect 17020 -29700 17220 -29690
rect 17900 -29700 18100 -29690
rect 18560 -29700 18760 -29690
rect 19220 -29700 19420 -29690
rect 20900 -29700 20910 -29690
rect 1410 -29760 2510 -29700
rect 2690 -29760 3170 -29700
rect 3350 -29760 3830 -29700
rect 4010 -29760 4710 -29700
rect 4890 -29760 5370 -29700
rect 5550 -29760 6030 -29700
rect 6210 -29760 15710 -29700
rect 15890 -29760 16370 -29700
rect 16550 -29760 17030 -29700
rect 17210 -29760 17910 -29700
rect 18090 -29760 18570 -29700
rect 18750 -29760 19230 -29700
rect 19410 -29760 20910 -29700
rect 1410 -29770 1420 -29760
rect 2500 -29770 2700 -29760
rect 3160 -29770 3360 -29760
rect 3820 -29770 4020 -29760
rect 4700 -29770 4900 -29760
rect 5360 -29770 5560 -29760
rect 6020 -29770 6220 -29760
rect 6900 -29770 7100 -29760
rect 7560 -29770 7760 -29760
rect 8220 -29770 8420 -29760
rect 9100 -29770 9300 -29760
rect 9760 -29770 9960 -29760
rect 10420 -29770 10620 -29760
rect 11300 -29770 11500 -29760
rect 11960 -29770 12160 -29760
rect 12620 -29770 12820 -29760
rect 13500 -29770 13700 -29760
rect 14160 -29770 14360 -29760
rect 14820 -29770 15020 -29760
rect 15700 -29770 15900 -29760
rect 16360 -29770 16560 -29760
rect 17020 -29770 17220 -29760
rect 17900 -29770 18100 -29760
rect 18560 -29770 18760 -29760
rect 19220 -29770 19420 -29760
rect 20900 -29770 20910 -29760
rect 21090 -29700 21100 -29690
rect 30420 -29690 30430 -29470
rect 30490 -29530 37700 -29470
rect 37940 -29530 38310 -29460
rect 30490 -29690 30500 -29530
rect 37690 -29540 37950 -29530
rect 30420 -29700 30500 -29690
rect 21090 -29760 22140 -29700
rect 21090 -29770 21100 -29760
rect 1220 -29780 1420 -29770
rect 20900 -29780 21100 -29770
rect 1620 -29830 1820 -29820
rect 1620 -29840 1630 -29830
rect 1600 -29900 1630 -29840
rect 1620 -29910 1630 -29900
rect 1810 -29840 1820 -29830
rect 20100 -29830 20300 -29820
rect 20100 -29840 20110 -29830
rect 1810 -29870 20110 -29840
rect 1810 -29900 2510 -29870
rect 1810 -29910 1820 -29900
rect 1620 -29920 1820 -29910
rect 2500 -29930 2510 -29900
rect 4010 -29900 4710 -29870
rect 4010 -29930 4020 -29900
rect 2500 -29940 4020 -29930
rect 4700 -29930 4710 -29900
rect 6210 -29900 6910 -29870
rect 6210 -29930 6220 -29900
rect 4700 -29940 6220 -29930
rect 6900 -29930 6910 -29900
rect 8410 -29900 9110 -29870
rect 8410 -29930 8420 -29900
rect 6900 -29940 8420 -29930
rect 9100 -29930 9110 -29900
rect 10610 -29900 11310 -29870
rect 10610 -29930 10620 -29900
rect 9100 -29940 10620 -29930
rect 11300 -29930 11310 -29900
rect 12810 -29900 13510 -29870
rect 12810 -29930 12820 -29900
rect 11300 -29940 12820 -29930
rect 13500 -29930 13510 -29900
rect 15010 -29900 15710 -29870
rect 15010 -29930 15020 -29900
rect 13500 -29940 15020 -29930
rect 15700 -29930 15710 -29900
rect 17210 -29900 17910 -29870
rect 17210 -29930 17220 -29900
rect 15700 -29940 17220 -29930
rect 17900 -29930 17910 -29900
rect 19410 -29900 20110 -29870
rect 19410 -29930 19420 -29900
rect 20100 -29910 20110 -29900
rect 20290 -29840 20300 -29830
rect 20290 -29900 20320 -29840
rect 20290 -29910 20300 -29900
rect 20100 -29920 20300 -29910
rect 17900 -29940 19420 -29930
rect 820 -30350 1020 -30340
rect 20500 -30350 20700 -30340
rect 820 -30360 830 -30350
rect -260 -30420 830 -30360
rect 820 -30430 830 -30420
rect 1010 -30360 1020 -30350
rect 2500 -30360 2700 -30350
rect 3160 -30360 3360 -30350
rect 3820 -30360 4020 -30350
rect 4700 -30360 4900 -30350
rect 5360 -30360 5560 -30350
rect 6020 -30360 6220 -30350
rect 6900 -30360 7100 -30350
rect 7560 -30360 7760 -30350
rect 8220 -30360 8420 -30350
rect 9100 -30360 9300 -30350
rect 9760 -30360 9960 -30350
rect 10420 -30360 10620 -30350
rect 11300 -30360 11500 -30350
rect 11960 -30360 12160 -30350
rect 12620 -30360 12820 -30350
rect 13500 -30360 13700 -30350
rect 14160 -30360 14360 -30350
rect 14820 -30360 15020 -30350
rect 15700 -30360 15900 -30350
rect 16360 -30360 16560 -30350
rect 17020 -30360 17220 -30350
rect 17900 -30360 18100 -30350
rect 18560 -30360 18760 -30350
rect 19220 -30360 19420 -30350
rect 20500 -30360 20510 -30350
rect 1010 -30420 2510 -30360
rect 2690 -30420 3170 -30360
rect 3350 -30420 3830 -30360
rect 4010 -30420 4710 -30360
rect 4890 -30420 5370 -30360
rect 5550 -30420 6030 -30360
rect 6210 -30420 15710 -30360
rect 15890 -30420 16370 -30360
rect 16550 -30420 17030 -30360
rect 17210 -30420 17910 -30360
rect 18090 -30420 18570 -30360
rect 18750 -30420 19230 -30360
rect 19410 -30420 20510 -30360
rect 1010 -30430 1020 -30420
rect 2500 -30430 2700 -30420
rect 3160 -30430 3360 -30420
rect 3820 -30430 4020 -30420
rect 4700 -30430 4900 -30420
rect 5360 -30430 5560 -30420
rect 6020 -30430 6220 -30420
rect 6900 -30430 7100 -30420
rect 7560 -30430 7760 -30420
rect 8220 -30430 8420 -30420
rect 9100 -30430 9300 -30420
rect 9760 -30430 9960 -30420
rect 10420 -30430 10620 -30420
rect 11300 -30430 11500 -30420
rect 11960 -30430 12160 -30420
rect 12620 -30430 12820 -30420
rect 13500 -30430 13700 -30420
rect 14160 -30430 14360 -30420
rect 14820 -30430 15020 -30420
rect 15700 -30430 15900 -30420
rect 16360 -30430 16560 -30420
rect 17020 -30430 17220 -30420
rect 17900 -30430 18100 -30420
rect 18560 -30430 18760 -30420
rect 19220 -30430 19420 -30420
rect 20500 -30430 20510 -30420
rect 20690 -30360 20700 -30350
rect 20690 -30420 22140 -30360
rect 28930 -30410 29170 -30400
rect 32600 -30410 32860 -30400
rect 20690 -30430 20700 -30420
rect 820 -30440 1020 -30430
rect 20500 -30440 20700 -30430
rect 28930 -30480 28940 -30410
rect 29160 -30480 32610 -30410
rect 32850 -30480 38300 -30410
rect 1220 -30490 1420 -30480
rect 20900 -30490 21100 -30480
rect 28930 -30490 29170 -30480
rect 32600 -30490 32860 -30480
rect 1220 -30500 1230 -30490
rect -260 -30560 1230 -30500
rect 1220 -30570 1230 -30560
rect 1410 -30500 1420 -30490
rect 2500 -30500 2700 -30490
rect 3160 -30500 3360 -30490
rect 3820 -30500 4020 -30490
rect 4700 -30500 4900 -30490
rect 5360 -30500 5560 -30490
rect 6020 -30500 6220 -30490
rect 6900 -30500 7100 -30490
rect 7560 -30500 7760 -30490
rect 8220 -30500 8420 -30490
rect 9100 -30500 9300 -30490
rect 9760 -30500 9960 -30490
rect 10420 -30500 10620 -30490
rect 11300 -30500 11500 -30490
rect 11960 -30500 12160 -30490
rect 12620 -30500 12820 -30490
rect 13500 -30500 13700 -30490
rect 14160 -30500 14360 -30490
rect 14820 -30500 15020 -30490
rect 15700 -30500 15900 -30490
rect 16360 -30500 16560 -30490
rect 17020 -30500 17220 -30490
rect 17900 -30500 18100 -30490
rect 18560 -30500 18760 -30490
rect 19220 -30500 19420 -30490
rect 20900 -30500 20910 -30490
rect 1410 -30560 6910 -30500
rect 7090 -30560 7570 -30500
rect 7750 -30560 8230 -30500
rect 8410 -30560 9110 -30500
rect 9290 -30560 9770 -30500
rect 9950 -30560 10430 -30500
rect 10610 -30560 11310 -30500
rect 11490 -30560 11970 -30500
rect 12150 -30560 12630 -30500
rect 12810 -30560 13510 -30500
rect 13690 -30560 14170 -30500
rect 14350 -30560 14830 -30500
rect 15010 -30560 20910 -30500
rect 1410 -30570 1420 -30560
rect 2500 -30570 2700 -30560
rect 3160 -30570 3360 -30560
rect 3820 -30570 4020 -30560
rect 4700 -30570 4900 -30560
rect 5360 -30570 5560 -30560
rect 6020 -30570 6220 -30560
rect 6900 -30570 7100 -30560
rect 7560 -30570 7760 -30560
rect 8220 -30570 8420 -30560
rect 9100 -30570 9300 -30560
rect 9760 -30570 9960 -30560
rect 10420 -30570 10620 -30560
rect 11300 -30570 11500 -30560
rect 11960 -30570 12160 -30560
rect 12620 -30570 12820 -30560
rect 13500 -30570 13700 -30560
rect 14160 -30570 14360 -30560
rect 14820 -30570 15020 -30560
rect 15700 -30570 15900 -30560
rect 16360 -30570 16560 -30560
rect 17020 -30570 17220 -30560
rect 17900 -30570 18100 -30560
rect 18560 -30570 18760 -30560
rect 19220 -30570 19420 -30560
rect 20900 -30570 20910 -30560
rect 21090 -30500 21100 -30490
rect 21090 -30560 22140 -30500
rect 29060 -30560 29300 -30550
rect 33310 -30560 33570 -30550
rect 21090 -30570 21100 -30560
rect 1220 -30580 1420 -30570
rect 20900 -30580 21100 -30570
rect 1620 -30630 1820 -30620
rect 1620 -30640 1630 -30630
rect 1600 -30700 1630 -30640
rect 1620 -30710 1630 -30700
rect 1810 -30640 1820 -30630
rect 20100 -30630 20300 -30620
rect 20100 -30640 20110 -30630
rect 1810 -30670 20110 -30640
rect 1810 -30700 2510 -30670
rect 1810 -30710 1820 -30700
rect 1620 -30720 1820 -30710
rect 2500 -30730 2510 -30700
rect 4010 -30700 4710 -30670
rect 4010 -30730 4020 -30700
rect 2500 -30740 4020 -30730
rect 4700 -30730 4710 -30700
rect 6210 -30700 6910 -30670
rect 6210 -30730 6220 -30700
rect 4700 -30740 6220 -30730
rect 6900 -30730 6910 -30700
rect 8410 -30700 9110 -30670
rect 8410 -30730 8420 -30700
rect 6900 -30740 8420 -30730
rect 9100 -30730 9110 -30700
rect 10610 -30700 11310 -30670
rect 10610 -30730 10620 -30700
rect 9100 -30740 10620 -30730
rect 11300 -30730 11310 -30700
rect 12810 -30700 13510 -30670
rect 12810 -30730 12820 -30700
rect 11300 -30740 12820 -30730
rect 13500 -30730 13510 -30700
rect 15010 -30700 15710 -30670
rect 15010 -30730 15020 -30700
rect 13500 -30740 15020 -30730
rect 15700 -30730 15710 -30700
rect 17210 -30700 17910 -30670
rect 17210 -30730 17220 -30700
rect 15700 -30740 17220 -30730
rect 17900 -30730 17910 -30700
rect 19410 -30700 20110 -30670
rect 19410 -30730 19420 -30700
rect 20100 -30710 20110 -30700
rect 20290 -30640 20300 -30630
rect 29060 -30630 29070 -30560
rect 29290 -30630 33320 -30560
rect 33560 -30630 38300 -30560
rect 29060 -30640 29300 -30630
rect 33310 -30640 33570 -30630
rect 20290 -30700 20320 -30640
rect 20290 -30710 20300 -30700
rect 20100 -30720 20300 -30710
rect 29210 -30710 29450 -30700
rect 34310 -30710 34570 -30700
rect 17900 -30740 19420 -30730
rect 29210 -30780 29220 -30710
rect 29440 -30712 38300 -30710
rect 29440 -30780 34320 -30712
rect 29210 -30790 29450 -30780
rect 34310 -30782 34320 -30780
rect 34560 -30780 38300 -30712
rect 34560 -30782 34570 -30780
rect 34310 -30790 34570 -30782
rect 29360 -30860 29600 -30850
rect 35310 -30860 35570 -30850
rect 29360 -30930 29370 -30860
rect 29590 -30930 35320 -30860
rect 35560 -30930 38300 -30860
rect 29360 -30940 29600 -30930
rect 35310 -30940 35570 -30930
rect 820 -31150 1020 -31140
rect 20500 -31150 20700 -31140
rect 820 -31160 830 -31150
rect -260 -31220 830 -31160
rect 820 -31230 830 -31220
rect 1010 -31160 1020 -31150
rect 2500 -31160 2700 -31150
rect 3160 -31160 3360 -31150
rect 3820 -31160 4020 -31150
rect 4700 -31160 4900 -31150
rect 5360 -31160 5560 -31150
rect 6020 -31160 6220 -31150
rect 6900 -31160 7100 -31150
rect 7560 -31160 7760 -31150
rect 8220 -31160 8420 -31150
rect 9100 -31160 9300 -31150
rect 9760 -31160 9960 -31150
rect 10420 -31160 10620 -31150
rect 11300 -31160 11500 -31150
rect 11960 -31160 12160 -31150
rect 12620 -31160 12820 -31150
rect 13500 -31160 13700 -31150
rect 14160 -31160 14360 -31150
rect 14820 -31160 15020 -31150
rect 15700 -31160 15900 -31150
rect 16360 -31160 16560 -31150
rect 17020 -31160 17220 -31150
rect 17900 -31160 18100 -31150
rect 18560 -31160 18760 -31150
rect 19220 -31160 19420 -31150
rect 20500 -31160 20510 -31150
rect 1010 -31220 6910 -31160
rect 7090 -31220 7570 -31160
rect 7750 -31220 8230 -31160
rect 8410 -31220 9110 -31160
rect 9290 -31220 9770 -31160
rect 9950 -31220 10430 -31160
rect 10610 -31220 11310 -31160
rect 11490 -31220 11970 -31160
rect 12150 -31220 12630 -31160
rect 12810 -31220 13510 -31160
rect 13690 -31220 14170 -31160
rect 14350 -31220 14830 -31160
rect 15010 -31220 20510 -31160
rect 1010 -31230 1020 -31220
rect 2500 -31230 2700 -31220
rect 3160 -31230 3360 -31220
rect 3820 -31230 4020 -31220
rect 4700 -31230 4900 -31220
rect 5360 -31230 5560 -31220
rect 6020 -31230 6220 -31220
rect 6900 -31230 7100 -31220
rect 7560 -31230 7760 -31220
rect 8220 -31230 8420 -31220
rect 9100 -31230 9300 -31220
rect 9760 -31230 9960 -31220
rect 10420 -31230 10620 -31220
rect 11300 -31230 11500 -31220
rect 11960 -31230 12160 -31220
rect 12620 -31230 12820 -31220
rect 13500 -31230 13700 -31220
rect 14160 -31230 14360 -31220
rect 14820 -31230 15020 -31220
rect 15700 -31230 15900 -31220
rect 16360 -31230 16560 -31220
rect 17020 -31230 17220 -31220
rect 17900 -31230 18100 -31220
rect 18560 -31230 18760 -31220
rect 19220 -31230 19420 -31220
rect 20500 -31230 20510 -31220
rect 20690 -31160 20700 -31150
rect 20690 -31220 22140 -31160
rect 20690 -31230 20700 -31220
rect 820 -31240 1020 -31230
rect 20500 -31240 20700 -31230
rect 1220 -31290 1420 -31280
rect 20900 -31290 21100 -31280
rect 1220 -31300 1230 -31290
rect -260 -31360 1230 -31300
rect 1220 -31370 1230 -31360
rect 1410 -31300 1420 -31290
rect 2500 -31300 2700 -31290
rect 3160 -31300 3360 -31290
rect 3820 -31300 4020 -31290
rect 4700 -31300 4900 -31290
rect 5360 -31300 5560 -31290
rect 6020 -31300 6220 -31290
rect 6900 -31300 7100 -31290
rect 7560 -31300 7760 -31290
rect 8220 -31300 8420 -31290
rect 9100 -31300 9300 -31290
rect 9760 -31300 9960 -31290
rect 10420 -31300 10620 -31290
rect 11300 -31300 11500 -31290
rect 11960 -31300 12160 -31290
rect 12620 -31300 12820 -31290
rect 13500 -31300 13700 -31290
rect 14160 -31300 14360 -31290
rect 14820 -31300 15020 -31290
rect 15700 -31300 15900 -31290
rect 16360 -31300 16560 -31290
rect 17020 -31300 17220 -31290
rect 17900 -31300 18100 -31290
rect 18560 -31300 18760 -31290
rect 19220 -31300 19420 -31290
rect 20900 -31300 20910 -31290
rect 1410 -31360 2510 -31300
rect 2690 -31360 3170 -31300
rect 3350 -31360 3830 -31300
rect 4010 -31360 4710 -31300
rect 4890 -31360 5370 -31300
rect 5550 -31360 6030 -31300
rect 6210 -31360 15710 -31300
rect 15890 -31360 16370 -31300
rect 16550 -31360 17030 -31300
rect 17210 -31360 17910 -31300
rect 18090 -31360 18570 -31300
rect 18750 -31360 19230 -31300
rect 19410 -31360 20910 -31300
rect 1410 -31370 1420 -31360
rect 2500 -31370 2700 -31360
rect 3160 -31370 3360 -31360
rect 3820 -31370 4020 -31360
rect 4700 -31370 4900 -31360
rect 5360 -31370 5560 -31360
rect 6020 -31370 6220 -31360
rect 6900 -31370 7100 -31360
rect 7560 -31370 7760 -31360
rect 8220 -31370 8420 -31360
rect 9100 -31370 9300 -31360
rect 9760 -31370 9960 -31360
rect 10420 -31370 10620 -31360
rect 11300 -31370 11500 -31360
rect 11960 -31370 12160 -31360
rect 12620 -31370 12820 -31360
rect 13500 -31370 13700 -31360
rect 14160 -31370 14360 -31360
rect 14820 -31370 15020 -31360
rect 15700 -31370 15900 -31360
rect 16360 -31370 16560 -31360
rect 17020 -31370 17220 -31360
rect 17900 -31370 18100 -31360
rect 18560 -31370 18760 -31360
rect 19220 -31370 19420 -31360
rect 20900 -31370 20910 -31360
rect 21090 -31300 21100 -31290
rect 21090 -31360 22140 -31300
rect 21090 -31370 21100 -31360
rect 1220 -31380 1420 -31370
rect 20900 -31380 21100 -31370
rect -360 -31450 570 -31440
rect -360 -31830 -350 -31450
rect -170 -31540 570 -31450
rect -170 -31830 -160 -31540
rect 460 -31720 570 -31540
rect 30820 -31680 31260 -31660
rect 1980 -31710 2120 -31700
rect 1980 -31720 1990 -31710
rect -360 -31840 -160 -31830
rect 80 -31730 280 -31720
rect 80 -32110 90 -31730
rect 270 -32020 280 -31730
rect 460 -31820 1990 -31720
rect 1980 -31830 1990 -31820
rect 2110 -31720 2120 -31710
rect 4180 -31710 4320 -31700
rect 4180 -31720 4190 -31710
rect 2110 -31820 4190 -31720
rect 2110 -31830 2120 -31820
rect 1980 -31840 2120 -31830
rect 4180 -31830 4190 -31820
rect 4310 -31720 4320 -31710
rect 6380 -31710 6520 -31700
rect 6380 -31720 6390 -31710
rect 4310 -31820 6390 -31720
rect 4310 -31830 4320 -31820
rect 4180 -31840 4320 -31830
rect 6380 -31830 6390 -31820
rect 6510 -31720 6520 -31710
rect 8580 -31710 8720 -31700
rect 8580 -31720 8590 -31710
rect 6510 -31820 8590 -31720
rect 6510 -31830 6520 -31820
rect 6380 -31840 6520 -31830
rect 8580 -31830 8590 -31820
rect 8710 -31720 8720 -31710
rect 10780 -31710 10920 -31700
rect 10780 -31720 10790 -31710
rect 8710 -31820 10790 -31720
rect 8710 -31830 8720 -31820
rect 8580 -31840 8720 -31830
rect 10780 -31830 10790 -31820
rect 10910 -31720 10920 -31710
rect 12980 -31710 13120 -31700
rect 12980 -31720 12990 -31710
rect 10910 -31820 12990 -31720
rect 10910 -31830 10920 -31820
rect 10780 -31840 10920 -31830
rect 12980 -31830 12990 -31820
rect 13110 -31720 13120 -31710
rect 15180 -31710 15320 -31700
rect 15180 -31720 15190 -31710
rect 13110 -31820 15190 -31720
rect 13110 -31830 13120 -31820
rect 12980 -31840 13120 -31830
rect 15180 -31830 15190 -31820
rect 15310 -31720 15320 -31710
rect 17380 -31710 17520 -31700
rect 17380 -31720 17390 -31710
rect 15310 -31820 17390 -31720
rect 15310 -31830 15320 -31820
rect 15180 -31840 15320 -31830
rect 17380 -31830 17390 -31820
rect 17510 -31720 17520 -31710
rect 19580 -31710 19720 -31700
rect 19580 -31720 19590 -31710
rect 17510 -31820 19590 -31720
rect 17510 -31830 17520 -31820
rect 17380 -31840 17520 -31830
rect 19580 -31830 19590 -31820
rect 19710 -31720 19720 -31710
rect 19710 -31820 22240 -31720
rect 19710 -31830 19720 -31820
rect 19580 -31840 19720 -31830
rect 2200 -32010 2340 -32000
rect 2200 -32020 2210 -32010
rect 270 -32110 2210 -32020
rect 80 -32120 2210 -32110
rect 2200 -32130 2210 -32120
rect 2330 -32020 2340 -32010
rect 4400 -32010 4540 -32000
rect 4400 -32020 4410 -32010
rect 2330 -32120 4410 -32020
rect 2330 -32130 2340 -32120
rect 2200 -32140 2340 -32130
rect 4400 -32130 4410 -32120
rect 4530 -32020 4540 -32010
rect 6600 -32010 6740 -32000
rect 6600 -32020 6610 -32010
rect 4530 -32120 6610 -32020
rect 4530 -32130 4540 -32120
rect 4400 -32140 4540 -32130
rect 6600 -32130 6610 -32120
rect 6730 -32020 6740 -32010
rect 8800 -32010 8940 -32000
rect 8800 -32020 8810 -32010
rect 6730 -32120 8810 -32020
rect 6730 -32130 6740 -32120
rect 6600 -32140 6740 -32130
rect 8800 -32130 8810 -32120
rect 8930 -32020 8940 -32010
rect 11000 -32010 11140 -32000
rect 11000 -32020 11010 -32010
rect 8930 -32120 11010 -32020
rect 8930 -32130 8940 -32120
rect 8800 -32140 8940 -32130
rect 11000 -32130 11010 -32120
rect 11130 -32020 11140 -32010
rect 13200 -32010 13340 -32000
rect 13200 -32020 13210 -32010
rect 11130 -32120 13210 -32020
rect 11130 -32130 11140 -32120
rect 11000 -32140 11140 -32130
rect 13200 -32130 13210 -32120
rect 13330 -32020 13340 -32010
rect 15400 -32010 15540 -32000
rect 15400 -32020 15410 -32010
rect 13330 -32120 15410 -32020
rect 13330 -32130 13340 -32120
rect 13200 -32140 13340 -32130
rect 15400 -32130 15410 -32120
rect 15530 -32020 15540 -32010
rect 17600 -32010 17740 -32000
rect 17600 -32020 17610 -32010
rect 15530 -32120 17610 -32020
rect 15530 -32130 15540 -32120
rect 15400 -32140 15540 -32130
rect 17600 -32130 17610 -32120
rect 17730 -32020 17740 -32010
rect 19800 -32010 19940 -32000
rect 19800 -32020 19810 -32010
rect 17730 -32120 19810 -32020
rect 17730 -32130 17740 -32120
rect 17600 -32140 17740 -32130
rect 19800 -32130 19810 -32120
rect 19930 -32020 19940 -32010
rect 19930 -32120 22240 -32020
rect 19930 -32130 19940 -32120
rect 19800 -32140 19940 -32130
rect 30820 -32440 30840 -31680
rect 31240 -32440 31260 -31680
rect 30820 -32460 31260 -32440
rect 38300 -32180 38540 -32160
rect 38300 -32690 38320 -32180
rect 38520 -32690 38540 -32180
rect 38300 -32910 38310 -32690
rect 38530 -32910 38540 -32690
rect 38300 -32920 38540 -32910
<< via3 >>
rect 36920 12280 38280 12540
rect 830 11170 1010 11250
rect 20510 11170 20690 11250
rect 1230 11030 1410 11110
rect 20910 11030 21090 11110
rect -80 10930 0 10940
rect -80 10870 -70 10930
rect -70 10870 -10 10930
rect -10 10870 0 10930
rect -80 10690 0 10870
rect 2120 10930 2200 10940
rect 2120 10870 2130 10930
rect 2130 10870 2190 10930
rect 2190 10870 2200 10930
rect 2120 10690 2200 10870
rect 4320 10930 4400 10940
rect 4320 10870 4330 10930
rect 4330 10870 4390 10930
rect 4390 10870 4400 10930
rect 4320 10690 4400 10870
rect 6520 10930 6600 10940
rect 6520 10870 6530 10930
rect 6530 10870 6590 10930
rect 6590 10870 6600 10930
rect 6520 10690 6600 10870
rect 8720 10930 8800 10940
rect 8720 10870 8730 10930
rect 8730 10870 8790 10930
rect 8790 10870 8800 10930
rect 8720 10690 8800 10870
rect 10920 10930 11000 10940
rect 10920 10870 10930 10930
rect 10930 10870 10990 10930
rect 10990 10870 11000 10930
rect 10920 10690 11000 10870
rect 13120 10930 13200 10940
rect 13120 10870 13130 10930
rect 13130 10870 13190 10930
rect 13190 10870 13200 10930
rect 13120 10690 13200 10870
rect 15320 10930 15400 10940
rect 15320 10870 15330 10930
rect 15330 10870 15390 10930
rect 15390 10870 15400 10930
rect 15320 10690 15400 10870
rect 17520 10930 17600 10940
rect 17520 10870 17530 10930
rect 17530 10870 17590 10930
rect 17590 10870 17600 10930
rect 17520 10690 17600 10870
rect 19720 10930 19800 10940
rect 19720 10870 19730 10930
rect 19730 10870 19790 10930
rect 19790 10870 19800 10930
rect 19720 10690 19800 10870
rect 21920 10930 22000 10940
rect 21920 10870 21930 10930
rect 21930 10870 21990 10930
rect 21990 10870 22000 10930
rect 21920 10690 22000 10870
rect 30326 10932 30682 11060
rect 36890 10850 37050 11010
rect 1630 10510 1810 10590
rect 20110 10510 20290 10590
rect 37090 10600 37250 10760
rect 830 10370 1010 10450
rect 20510 10370 20690 10450
rect 1230 10230 1410 10310
rect 20910 10230 21090 10310
rect -80 10130 0 10140
rect -80 10070 -70 10130
rect -70 10070 -10 10130
rect -10 10070 0 10130
rect -80 9890 0 10070
rect 2120 10130 2200 10140
rect 2120 10070 2130 10130
rect 2130 10070 2190 10130
rect 2190 10070 2200 10130
rect 2120 9890 2200 10070
rect 4320 10130 4400 10140
rect 4320 10070 4330 10130
rect 4330 10070 4390 10130
rect 4390 10070 4400 10130
rect 4320 9890 4400 10070
rect 6520 10130 6600 10140
rect 6520 10070 6530 10130
rect 6530 10070 6590 10130
rect 6590 10070 6600 10130
rect 6520 9890 6600 10070
rect 8720 10130 8800 10140
rect 8720 10070 8730 10130
rect 8730 10070 8790 10130
rect 8790 10070 8800 10130
rect 8720 9890 8800 10070
rect 10920 10130 11000 10140
rect 10920 10070 10930 10130
rect 10930 10070 10990 10130
rect 10990 10070 11000 10130
rect 10920 9890 11000 10070
rect 13120 10130 13200 10140
rect 13120 10070 13130 10130
rect 13130 10070 13190 10130
rect 13190 10070 13200 10130
rect 13120 9890 13200 10070
rect 15320 10130 15400 10140
rect 15320 10070 15330 10130
rect 15330 10070 15390 10130
rect 15390 10070 15400 10130
rect 15320 9890 15400 10070
rect 17520 10130 17600 10140
rect 17520 10070 17530 10130
rect 17530 10070 17590 10130
rect 17590 10070 17600 10130
rect 17520 9890 17600 10070
rect 19720 10130 19800 10140
rect 19720 10070 19730 10130
rect 19730 10070 19790 10130
rect 19790 10070 19800 10130
rect 19720 9890 19800 10070
rect 21920 10130 22000 10140
rect 21920 10070 21930 10130
rect 21930 10070 21990 10130
rect 21990 10070 22000 10130
rect 21920 9890 22000 10070
rect 1630 9710 1810 9790
rect 20110 9710 20290 9790
rect 830 9570 1010 9650
rect 20510 9570 20690 9650
rect 1230 9430 1410 9510
rect 20910 9430 21090 9510
rect -80 9330 0 9340
rect -80 9270 -70 9330
rect -70 9270 -10 9330
rect -10 9270 0 9330
rect -80 9090 0 9270
rect 2120 9330 2200 9340
rect 2120 9270 2130 9330
rect 2130 9270 2190 9330
rect 2190 9270 2200 9330
rect 2120 9090 2200 9270
rect 4320 9330 4400 9340
rect 4320 9270 4330 9330
rect 4330 9270 4390 9330
rect 4390 9270 4400 9330
rect 4320 9090 4400 9270
rect 6520 9330 6600 9340
rect 6520 9270 6530 9330
rect 6530 9270 6590 9330
rect 6590 9270 6600 9330
rect 6520 9090 6600 9270
rect 8720 9330 8800 9340
rect 8720 9270 8730 9330
rect 8730 9270 8790 9330
rect 8790 9270 8800 9330
rect 8720 9090 8800 9270
rect 10920 9330 11000 9340
rect 10920 9270 10930 9330
rect 10930 9270 10990 9330
rect 10990 9270 11000 9330
rect 10920 9090 11000 9270
rect 13120 9330 13200 9340
rect 13120 9270 13130 9330
rect 13130 9270 13190 9330
rect 13190 9270 13200 9330
rect 13120 9090 13200 9270
rect 15320 9330 15400 9340
rect 15320 9270 15330 9330
rect 15330 9270 15390 9330
rect 15390 9270 15400 9330
rect 15320 9090 15400 9270
rect 17520 9330 17600 9340
rect 17520 9270 17530 9330
rect 17530 9270 17590 9330
rect 17590 9270 17600 9330
rect 17520 9090 17600 9270
rect 19720 9330 19800 9340
rect 19720 9270 19730 9330
rect 19730 9270 19790 9330
rect 19790 9270 19800 9330
rect 19720 9090 19800 9270
rect 21920 9330 22000 9340
rect 21920 9270 21930 9330
rect 21930 9270 21990 9330
rect 21990 9270 22000 9330
rect 21920 9090 22000 9270
rect 430 8910 610 8990
rect 1630 8910 1810 8990
rect 20110 8910 20290 8990
rect 21310 8910 21490 8990
rect 830 8770 1010 8850
rect 20510 8770 20690 8850
rect 1230 8630 1410 8710
rect 20910 8630 21090 8710
rect -80 8530 0 8540
rect -80 8470 -70 8530
rect -70 8470 -10 8530
rect -10 8470 0 8530
rect -80 8290 0 8470
rect 2120 8530 2200 8540
rect 2120 8470 2130 8530
rect 2130 8470 2190 8530
rect 2190 8470 2200 8530
rect 2120 8290 2200 8470
rect 4320 8530 4400 8540
rect 4320 8470 4330 8530
rect 4330 8470 4390 8530
rect 4390 8470 4400 8530
rect 4320 8290 4400 8470
rect 6520 8530 6600 8540
rect 6520 8470 6530 8530
rect 6530 8470 6590 8530
rect 6590 8470 6600 8530
rect 6520 8290 6600 8470
rect 8720 8530 8800 8540
rect 8720 8470 8730 8530
rect 8730 8470 8790 8530
rect 8790 8470 8800 8530
rect 8720 8290 8800 8470
rect 10920 8530 11000 8540
rect 10920 8470 10930 8530
rect 10930 8470 10990 8530
rect 10990 8470 11000 8530
rect 10920 8290 11000 8470
rect 13120 8530 13200 8540
rect 13120 8470 13130 8530
rect 13130 8470 13190 8530
rect 13190 8470 13200 8530
rect 13120 8290 13200 8470
rect 15320 8530 15400 8540
rect 15320 8470 15330 8530
rect 15330 8470 15390 8530
rect 15390 8470 15400 8530
rect 15320 8290 15400 8470
rect 17520 8530 17600 8540
rect 17520 8470 17530 8530
rect 17530 8470 17590 8530
rect 17590 8470 17600 8530
rect 17520 8290 17600 8470
rect 19720 8530 19800 8540
rect 19720 8470 19730 8530
rect 19730 8470 19790 8530
rect 19790 8470 19800 8530
rect 19720 8290 19800 8470
rect 21920 8530 22000 8540
rect 21920 8470 21930 8530
rect 21930 8470 21990 8530
rect 21990 8470 22000 8530
rect 21920 8290 22000 8470
rect 430 8110 610 8190
rect 1630 8110 1810 8190
rect 20110 8110 20290 8190
rect 21310 8110 21490 8190
rect 830 7970 1010 8050
rect 20510 7970 20690 8050
rect 1230 7830 1410 7910
rect 20910 7830 21090 7910
rect -80 7730 0 7740
rect -80 7670 -70 7730
rect -70 7670 -10 7730
rect -10 7670 0 7730
rect -80 7490 0 7670
rect 2120 7730 2200 7740
rect 2120 7670 2130 7730
rect 2130 7670 2190 7730
rect 2190 7670 2200 7730
rect 2120 7490 2200 7670
rect 4320 7730 4400 7740
rect 4320 7670 4330 7730
rect 4330 7670 4390 7730
rect 4390 7670 4400 7730
rect 4320 7490 4400 7670
rect 6520 7730 6600 7740
rect 6520 7670 6530 7730
rect 6530 7670 6590 7730
rect 6590 7670 6600 7730
rect 6520 7490 6600 7670
rect 8720 7730 8800 7740
rect 8720 7670 8730 7730
rect 8730 7670 8790 7730
rect 8790 7670 8800 7730
rect 8720 7490 8800 7670
rect 10920 7730 11000 7740
rect 10920 7670 10930 7730
rect 10930 7670 10990 7730
rect 10990 7670 11000 7730
rect 10920 7490 11000 7670
rect 13120 7730 13200 7740
rect 13120 7670 13130 7730
rect 13130 7670 13190 7730
rect 13190 7670 13200 7730
rect 13120 7490 13200 7670
rect 15320 7730 15400 7740
rect 15320 7670 15330 7730
rect 15330 7670 15390 7730
rect 15390 7670 15400 7730
rect 15320 7490 15400 7670
rect 17520 7730 17600 7740
rect 17520 7670 17530 7730
rect 17530 7670 17590 7730
rect 17590 7670 17600 7730
rect 17520 7490 17600 7670
rect 19720 7730 19800 7740
rect 19720 7670 19730 7730
rect 19730 7670 19790 7730
rect 19790 7670 19800 7730
rect 19720 7490 19800 7670
rect 21920 7730 22000 7740
rect 21920 7670 21930 7730
rect 21930 7670 21990 7730
rect 21990 7670 22000 7730
rect 21920 7490 22000 7670
rect 430 7310 610 7390
rect 1630 7310 1810 7390
rect 20110 7310 20290 7390
rect 21310 7310 21490 7390
rect 830 7170 1010 7250
rect 20510 7170 20690 7250
rect 1230 7030 1410 7110
rect 20910 7030 21090 7110
rect 33108 6976 33474 7186
rect 37516 6974 37684 7186
rect -80 6930 0 6940
rect -80 6870 -70 6930
rect -70 6870 -10 6930
rect -10 6870 0 6930
rect -80 6690 0 6870
rect 2120 6930 2200 6940
rect 2120 6870 2130 6930
rect 2130 6870 2190 6930
rect 2190 6870 2200 6930
rect 2120 6690 2200 6870
rect 4320 6930 4400 6940
rect 4320 6870 4330 6930
rect 4330 6870 4390 6930
rect 4390 6870 4400 6930
rect 4320 6690 4400 6870
rect 6520 6930 6600 6940
rect 6520 6870 6530 6930
rect 6530 6870 6590 6930
rect 6590 6870 6600 6930
rect 6520 6690 6600 6870
rect 8720 6930 8800 6940
rect 8720 6870 8730 6930
rect 8730 6870 8790 6930
rect 8790 6870 8800 6930
rect 8720 6690 8800 6870
rect 10920 6930 11000 6940
rect 10920 6870 10930 6930
rect 10930 6870 10990 6930
rect 10990 6870 11000 6930
rect 10920 6690 11000 6870
rect 13120 6930 13200 6940
rect 13120 6870 13130 6930
rect 13130 6870 13190 6930
rect 13190 6870 13200 6930
rect 13120 6690 13200 6870
rect 15320 6930 15400 6940
rect 15320 6870 15330 6930
rect 15330 6870 15390 6930
rect 15390 6870 15400 6930
rect 15320 6690 15400 6870
rect 17520 6930 17600 6940
rect 17520 6870 17530 6930
rect 17530 6870 17590 6930
rect 17590 6870 17600 6930
rect 17520 6690 17600 6870
rect 19720 6930 19800 6940
rect 19720 6870 19730 6930
rect 19730 6870 19790 6930
rect 19790 6870 19800 6930
rect 19720 6690 19800 6870
rect 21920 6930 22000 6940
rect 21920 6870 21930 6930
rect 21930 6870 21990 6930
rect 21990 6870 22000 6930
rect 21920 6690 22000 6870
rect 430 6510 610 6590
rect 1630 6510 1810 6590
rect 20110 6510 20290 6590
rect 21310 6510 21490 6590
rect 830 6370 1010 6450
rect 20510 6370 20690 6450
rect 1230 6230 1410 6310
rect 20910 6230 21090 6310
rect -80 6130 0 6140
rect -80 6070 -70 6130
rect -70 6070 -10 6130
rect -10 6070 0 6130
rect -80 5890 0 6070
rect 2120 6130 2200 6140
rect 2120 6070 2130 6130
rect 2130 6070 2190 6130
rect 2190 6070 2200 6130
rect 2120 5890 2200 6070
rect 4320 6130 4400 6140
rect 4320 6070 4330 6130
rect 4330 6070 4390 6130
rect 4390 6070 4400 6130
rect 4320 5890 4400 6070
rect 6520 6130 6600 6140
rect 6520 6070 6530 6130
rect 6530 6070 6590 6130
rect 6590 6070 6600 6130
rect 6520 5890 6600 6070
rect 8720 6130 8800 6140
rect 8720 6070 8730 6130
rect 8730 6070 8790 6130
rect 8790 6070 8800 6130
rect 8720 5890 8800 6070
rect 10920 6130 11000 6140
rect 10920 6070 10930 6130
rect 10930 6070 10990 6130
rect 10990 6070 11000 6130
rect 10920 5890 11000 6070
rect 13120 6130 13200 6140
rect 13120 6070 13130 6130
rect 13130 6070 13190 6130
rect 13190 6070 13200 6130
rect 13120 5890 13200 6070
rect 15320 6130 15400 6140
rect 15320 6070 15330 6130
rect 15330 6070 15390 6130
rect 15390 6070 15400 6130
rect 15320 5890 15400 6070
rect 17520 6130 17600 6140
rect 17520 6070 17530 6130
rect 17530 6070 17590 6130
rect 17590 6070 17600 6130
rect 17520 5890 17600 6070
rect 19720 6130 19800 6140
rect 19720 6070 19730 6130
rect 19730 6070 19790 6130
rect 19790 6070 19800 6130
rect 19720 5890 19800 6070
rect 21920 6130 22000 6140
rect 21920 6070 21930 6130
rect 21930 6070 21990 6130
rect 21990 6070 22000 6130
rect 21920 5890 22000 6070
rect 36230 6080 36410 6260
rect 36530 6080 36710 6260
rect 1630 5710 1810 5790
rect 20110 5710 20290 5790
rect 830 5570 1010 5650
rect 20510 5570 20690 5650
rect 1230 5430 1410 5510
rect 20910 5430 21090 5510
rect -80 5330 0 5340
rect -80 5270 -70 5330
rect -70 5270 -10 5330
rect -10 5270 0 5330
rect -80 5090 0 5270
rect 2120 5330 2200 5340
rect 2120 5270 2130 5330
rect 2130 5270 2190 5330
rect 2190 5270 2200 5330
rect 2120 5090 2200 5270
rect 4320 5330 4400 5340
rect 4320 5270 4330 5330
rect 4330 5270 4390 5330
rect 4390 5270 4400 5330
rect 4320 5090 4400 5270
rect 6520 5330 6600 5340
rect 6520 5270 6530 5330
rect 6530 5270 6590 5330
rect 6590 5270 6600 5330
rect 6520 5090 6600 5270
rect 8720 5330 8800 5340
rect 8720 5270 8730 5330
rect 8730 5270 8790 5330
rect 8790 5270 8800 5330
rect 8720 5090 8800 5270
rect 10920 5330 11000 5340
rect 10920 5270 10930 5330
rect 10930 5270 10990 5330
rect 10990 5270 11000 5330
rect 10920 5090 11000 5270
rect 13120 5330 13200 5340
rect 13120 5270 13130 5330
rect 13130 5270 13190 5330
rect 13190 5270 13200 5330
rect 13120 5090 13200 5270
rect 15320 5330 15400 5340
rect 15320 5270 15330 5330
rect 15330 5270 15390 5330
rect 15390 5270 15400 5330
rect 15320 5090 15400 5270
rect 17520 5330 17600 5340
rect 17520 5270 17530 5330
rect 17530 5270 17590 5330
rect 17590 5270 17600 5330
rect 17520 5090 17600 5270
rect 19720 5330 19800 5340
rect 19720 5270 19730 5330
rect 19730 5270 19790 5330
rect 19790 5270 19800 5330
rect 19720 5090 19800 5270
rect 21920 5330 22000 5340
rect 21920 5270 21930 5330
rect 21930 5270 21990 5330
rect 21990 5270 22000 5330
rect 21920 5090 22000 5270
rect 28500 5240 28660 5400
rect 36870 5100 37010 5320
rect 37130 5100 37270 5320
rect 1630 4910 1810 4990
rect 20110 4910 20290 4990
rect 30080 3860 30260 4040
rect 31680 3860 31860 4040
rect 33130 4010 33290 4110
rect 34870 4010 35190 4090
rect 430 3550 610 3730
rect 21310 3550 21490 3730
rect 1630 3150 1810 3330
rect 20110 3150 20290 3330
rect 7810 2810 7930 2930
rect 26210 3240 26370 3400
rect 480 -4780 660 2220
rect 14910 1320 15030 1980
rect 12880 -1260 13240 -1110
rect 2810 -5350 2990 -5170
rect 21280 -5350 21460 -5170
rect 36030 -5350 36210 -5170
rect 1270 -5750 1450 -5570
rect 20510 -5750 20690 -5570
rect 36230 -5750 36410 -5570
rect 31680 -6150 31860 -5970
rect 14910 -6610 15030 -6490
rect 12950 -6990 13110 -6830
rect 30080 -6950 30190 -6770
rect 30190 -6950 30260 -6770
rect 1260 -7350 1440 -7170
rect 20510 -7350 20530 -7170
rect 20530 -7350 20690 -7170
rect 36530 -7350 36710 -7170
rect 2080 -7750 2260 -7570
rect 22070 -7750 22250 -7570
rect 36230 -7750 36410 -7570
rect 7810 -7990 7930 -7870
rect 490 -22380 670 -8090
rect 34910 -16920 35050 -16770
rect 34910 -22610 35050 -22470
rect 1630 -23450 1810 -23270
rect 20110 -23450 20290 -23270
rect 430 -23850 610 -23670
rect 21310 -23850 21490 -23670
rect 28500 -24200 28660 -24040
rect 1630 -25110 1810 -25030
rect 20110 -25110 20290 -25030
rect 36870 -24780 37010 -24640
rect 37130 -24780 37270 -24640
rect 33030 -25000 33290 -24930
rect 33230 -25150 33490 -25080
rect 830 -25630 1010 -25550
rect 20510 -25630 20690 -25550
rect 1230 -25770 1410 -25690
rect 20910 -25770 21090 -25690
rect 1630 -25910 1810 -25830
rect 20110 -25910 20290 -25830
rect 830 -26430 1010 -26350
rect 20510 -26430 20690 -26350
rect 1230 -26570 1410 -26490
rect 20910 -26570 21090 -26490
rect 430 -26710 610 -26630
rect 1630 -26710 1810 -26630
rect 20110 -26710 20290 -26630
rect 21310 -26710 21490 -26630
rect 36030 -27140 36410 -27010
rect 36530 -27140 36910 -27010
rect 830 -27230 1010 -27150
rect 20510 -27230 20690 -27150
rect 1230 -27370 1410 -27290
rect 20910 -27370 21090 -27290
rect 430 -27510 610 -27430
rect 1630 -27510 1810 -27430
rect 20110 -27510 20290 -27430
rect 21310 -27510 21490 -27430
rect 36920 -27900 37680 -27540
rect 830 -28030 1010 -27950
rect 20510 -28030 20690 -27950
rect 1230 -28170 1410 -28090
rect 20910 -28170 21090 -28090
rect 430 -28310 610 -28230
rect 1630 -28310 1810 -28230
rect 20110 -28310 20290 -28230
rect 21310 -28310 21490 -28230
rect 36920 -28520 37680 -28160
rect 830 -28830 1010 -28750
rect 20510 -28830 20690 -28750
rect 1230 -28970 1410 -28890
rect 20910 -28970 21090 -28890
rect 430 -29110 610 -29030
rect 1630 -29110 1810 -29030
rect 20110 -29110 20290 -29030
rect 21310 -29110 21490 -29030
rect 830 -29630 1010 -29550
rect 20510 -29630 20690 -29550
rect 1230 -29770 1410 -29690
rect 20910 -29770 21090 -29690
rect 1630 -29910 1810 -29830
rect 20110 -29910 20290 -29830
rect 830 -30430 1010 -30350
rect 20510 -30430 20690 -30350
rect 1230 -30570 1410 -30490
rect 20910 -30570 21090 -30490
rect 1630 -30710 1810 -30630
rect 20110 -30710 20290 -30630
rect 830 -31230 1010 -31150
rect 20510 -31230 20690 -31150
rect 1230 -31370 1410 -31290
rect 20910 -31370 21090 -31290
rect 30840 -32440 31240 -31680
rect 38320 -32314 38406 -32180
rect 38406 -32314 38520 -32180
rect 38320 -32690 38520 -32314
rect 38310 -32910 38530 -32690
<< metal4 >>
rect 28980 11900 29360 13520
rect 36900 12540 39520 12560
rect 36900 12280 36920 12540
rect 38280 12280 39520 12540
rect 36900 12260 39520 12280
rect -180 11500 30706 11900
rect -180 10940 100 11500
rect -180 10690 -80 10940
rect 0 10690 100 10940
rect -180 10140 100 10690
rect -180 9890 -80 10140
rect 0 9890 100 10140
rect -180 9340 100 9890
rect -180 9090 -80 9340
rect 0 9090 100 9340
rect -180 8540 100 9090
rect -180 8290 -80 8540
rect 0 8290 100 8540
rect -180 7740 100 8290
rect -180 7490 -80 7740
rect 0 7490 100 7740
rect -180 6940 100 7490
rect -180 6690 -80 6940
rect 0 6690 100 6940
rect -180 6140 100 6690
rect -180 5890 -80 6140
rect 0 5890 100 6140
rect -180 5340 100 5890
rect -180 5090 -80 5340
rect 0 5090 100 5340
rect -180 2240 100 5090
rect 420 8990 620 11300
rect 420 8910 430 8990
rect 610 8910 620 8990
rect 420 8190 620 8910
rect 420 8110 430 8190
rect 610 8110 620 8190
rect 420 7390 620 8110
rect 420 7310 430 7390
rect 610 7310 620 7390
rect 420 6590 620 7310
rect 420 6510 430 6590
rect 610 6510 620 6590
rect 420 3730 620 6510
rect 420 3550 430 3730
rect 610 3550 620 3730
rect 420 3540 620 3550
rect 820 11250 1020 11300
rect 820 11170 830 11250
rect 1010 11170 1020 11250
rect 820 10450 1020 11170
rect 820 10370 830 10450
rect 1010 10370 1020 10450
rect 820 9650 1020 10370
rect 820 9570 830 9650
rect 1010 9570 1020 9650
rect 820 8850 1020 9570
rect 820 8770 830 8850
rect 1010 8770 1020 8850
rect 820 8050 1020 8770
rect 820 7970 830 8050
rect 1010 7970 1020 8050
rect 820 7250 1020 7970
rect 820 7170 830 7250
rect 1010 7170 1020 7250
rect 820 6450 1020 7170
rect 820 6370 830 6450
rect 1010 6370 1020 6450
rect 820 5650 1020 6370
rect 820 5570 830 5650
rect 1010 5570 1020 5650
rect -180 2220 670 2240
rect -180 2000 480 2220
rect 470 -4780 480 2000
rect 660 -4780 670 2220
rect 820 2210 1020 5570
rect 1220 11110 1420 11300
rect 1220 11030 1230 11110
rect 1410 11030 1420 11110
rect 1220 10310 1420 11030
rect 1220 10230 1230 10310
rect 1410 10230 1420 10310
rect 1220 9510 1420 10230
rect 1220 9430 1230 9510
rect 1410 9430 1420 9510
rect 1220 8710 1420 9430
rect 1220 8630 1230 8710
rect 1410 8630 1420 8710
rect 1220 7910 1420 8630
rect 1220 7830 1230 7910
rect 1410 7830 1420 7910
rect 1220 7110 1420 7830
rect 1220 7030 1230 7110
rect 1410 7030 1420 7110
rect 1220 6310 1420 7030
rect 1220 6230 1230 6310
rect 1410 6230 1420 6310
rect 1220 5510 1420 6230
rect 1220 5430 1230 5510
rect 1410 5430 1420 5510
rect 1220 2600 1420 5430
rect 1620 10590 1820 11300
rect 1620 10510 1630 10590
rect 1810 10510 1820 10590
rect 1620 9790 1820 10510
rect 1620 9710 1630 9790
rect 1810 9710 1820 9790
rect 1620 8990 1820 9710
rect 1620 8910 1630 8990
rect 1810 8910 1820 8990
rect 1620 8190 1820 8910
rect 1620 8110 1630 8190
rect 1810 8110 1820 8190
rect 1620 7390 1820 8110
rect 1620 7310 1630 7390
rect 1810 7310 1820 7390
rect 1620 6590 1820 7310
rect 1620 6510 1630 6590
rect 1810 6510 1820 6590
rect 1620 5790 1820 6510
rect 1620 5710 1630 5790
rect 1810 5710 1820 5790
rect 1620 4990 1820 5710
rect 1620 4910 1630 4990
rect 1810 4910 1820 4990
rect 1620 3330 1820 4910
rect 2020 10940 2300 11500
rect 2020 10690 2120 10940
rect 2200 10690 2300 10940
rect 2020 10140 2300 10690
rect 2020 9890 2120 10140
rect 2200 9890 2300 10140
rect 2020 9340 2300 9890
rect 2020 9090 2120 9340
rect 2200 9090 2300 9340
rect 2020 8540 2300 9090
rect 2020 8290 2120 8540
rect 2200 8290 2300 8540
rect 2020 7740 2300 8290
rect 2020 7490 2120 7740
rect 2200 7490 2300 7740
rect 2020 6940 2300 7490
rect 2020 6690 2120 6940
rect 2200 6690 2300 6940
rect 2020 6140 2300 6690
rect 2020 5890 2120 6140
rect 2200 5890 2300 6140
rect 2020 5340 2300 5890
rect 2020 5090 2120 5340
rect 2200 5090 2300 5340
rect 2020 3660 2300 5090
rect 4220 10940 4500 11500
rect 4220 10690 4320 10940
rect 4400 10690 4500 10940
rect 4220 10140 4500 10690
rect 4220 9890 4320 10140
rect 4400 9890 4500 10140
rect 4220 9340 4500 9890
rect 4220 9090 4320 9340
rect 4400 9090 4500 9340
rect 4220 8540 4500 9090
rect 4220 8290 4320 8540
rect 4400 8290 4500 8540
rect 4220 7740 4500 8290
rect 4220 7490 4320 7740
rect 4400 7490 4500 7740
rect 4220 6940 4500 7490
rect 4220 6690 4320 6940
rect 4400 6690 4500 6940
rect 4220 6140 4500 6690
rect 4220 5890 4320 6140
rect 4400 5890 4500 6140
rect 4220 5340 4500 5890
rect 4220 5090 4320 5340
rect 4400 5090 4500 5340
rect 4220 3660 4500 5090
rect 6420 10940 6700 11500
rect 6420 10690 6520 10940
rect 6600 10690 6700 10940
rect 6420 10140 6700 10690
rect 6420 9890 6520 10140
rect 6600 9890 6700 10140
rect 6420 9340 6700 9890
rect 6420 9090 6520 9340
rect 6600 9090 6700 9340
rect 6420 8540 6700 9090
rect 6420 8290 6520 8540
rect 6600 8290 6700 8540
rect 6420 7740 6700 8290
rect 6420 7490 6520 7740
rect 6600 7490 6700 7740
rect 6420 6940 6700 7490
rect 6420 6690 6520 6940
rect 6600 6690 6700 6940
rect 6420 6140 6700 6690
rect 6420 5890 6520 6140
rect 6600 5890 6700 6140
rect 6420 5340 6700 5890
rect 6420 5090 6520 5340
rect 6600 5090 6700 5340
rect 6420 3660 6700 5090
rect 8620 10940 8900 11500
rect 8620 10690 8720 10940
rect 8800 10690 8900 10940
rect 8620 10140 8900 10690
rect 8620 9890 8720 10140
rect 8800 9890 8900 10140
rect 8620 9340 8900 9890
rect 8620 9090 8720 9340
rect 8800 9090 8900 9340
rect 8620 8540 8900 9090
rect 8620 8290 8720 8540
rect 8800 8290 8900 8540
rect 8620 7740 8900 8290
rect 8620 7490 8720 7740
rect 8800 7490 8900 7740
rect 8620 6940 8900 7490
rect 8620 6690 8720 6940
rect 8800 6690 8900 6940
rect 8620 6140 8900 6690
rect 8620 5890 8720 6140
rect 8800 5890 8900 6140
rect 8620 5340 8900 5890
rect 8620 5090 8720 5340
rect 8800 5090 8900 5340
rect 8620 3660 8900 5090
rect 10820 10940 11100 11500
rect 10820 10690 10920 10940
rect 11000 10690 11100 10940
rect 10820 10140 11100 10690
rect 10820 9890 10920 10140
rect 11000 9890 11100 10140
rect 10820 9340 11100 9890
rect 10820 9090 10920 9340
rect 11000 9090 11100 9340
rect 10820 8540 11100 9090
rect 10820 8290 10920 8540
rect 11000 8290 11100 8540
rect 10820 7740 11100 8290
rect 10820 7490 10920 7740
rect 11000 7490 11100 7740
rect 10820 6940 11100 7490
rect 10820 6690 10920 6940
rect 11000 6690 11100 6940
rect 10820 6140 11100 6690
rect 10820 5890 10920 6140
rect 11000 5890 11100 6140
rect 10820 5340 11100 5890
rect 10820 5090 10920 5340
rect 11000 5090 11100 5340
rect 10820 3660 11100 5090
rect 13020 10940 13300 11500
rect 13020 10690 13120 10940
rect 13200 10690 13300 10940
rect 13020 10140 13300 10690
rect 13020 9890 13120 10140
rect 13200 9890 13300 10140
rect 13020 9340 13300 9890
rect 13020 9090 13120 9340
rect 13200 9090 13300 9340
rect 13020 8540 13300 9090
rect 13020 8290 13120 8540
rect 13200 8290 13300 8540
rect 13020 7740 13300 8290
rect 13020 7490 13120 7740
rect 13200 7490 13300 7740
rect 13020 6940 13300 7490
rect 13020 6690 13120 6940
rect 13200 6690 13300 6940
rect 13020 6140 13300 6690
rect 13020 5890 13120 6140
rect 13200 5890 13300 6140
rect 13020 5340 13300 5890
rect 13020 5090 13120 5340
rect 13200 5090 13300 5340
rect 13020 3660 13300 5090
rect 15220 10940 15500 11500
rect 15220 10690 15320 10940
rect 15400 10690 15500 10940
rect 15220 10140 15500 10690
rect 15220 9890 15320 10140
rect 15400 9890 15500 10140
rect 15220 9340 15500 9890
rect 15220 9090 15320 9340
rect 15400 9090 15500 9340
rect 15220 8540 15500 9090
rect 15220 8290 15320 8540
rect 15400 8290 15500 8540
rect 15220 7740 15500 8290
rect 15220 7490 15320 7740
rect 15400 7490 15500 7740
rect 15220 6940 15500 7490
rect 15220 6690 15320 6940
rect 15400 6690 15500 6940
rect 15220 6140 15500 6690
rect 15220 5890 15320 6140
rect 15400 5890 15500 6140
rect 15220 5340 15500 5890
rect 15220 5090 15320 5340
rect 15400 5090 15500 5340
rect 15220 3660 15500 5090
rect 17420 10940 17700 11500
rect 17420 10690 17520 10940
rect 17600 10690 17700 10940
rect 17420 10140 17700 10690
rect 17420 9890 17520 10140
rect 17600 9890 17700 10140
rect 17420 9340 17700 9890
rect 17420 9090 17520 9340
rect 17600 9090 17700 9340
rect 17420 8540 17700 9090
rect 17420 8290 17520 8540
rect 17600 8290 17700 8540
rect 17420 7740 17700 8290
rect 17420 7490 17520 7740
rect 17600 7490 17700 7740
rect 17420 6940 17700 7490
rect 17420 6690 17520 6940
rect 17600 6690 17700 6940
rect 17420 6140 17700 6690
rect 17420 5890 17520 6140
rect 17600 5890 17700 6140
rect 17420 5340 17700 5890
rect 17420 5090 17520 5340
rect 17600 5090 17700 5340
rect 17420 3660 17700 5090
rect 19620 10940 19900 11500
rect 19620 10690 19720 10940
rect 19800 10690 19900 10940
rect 19620 10140 19900 10690
rect 19620 9890 19720 10140
rect 19800 9890 19900 10140
rect 19620 9340 19900 9890
rect 19620 9090 19720 9340
rect 19800 9090 19900 9340
rect 19620 8540 19900 9090
rect 19620 8290 19720 8540
rect 19800 8290 19900 8540
rect 19620 7740 19900 8290
rect 19620 7490 19720 7740
rect 19800 7490 19900 7740
rect 19620 6940 19900 7490
rect 19620 6690 19720 6940
rect 19800 6690 19900 6940
rect 19620 6140 19900 6690
rect 19620 5890 19720 6140
rect 19800 5890 19900 6140
rect 19620 5340 19900 5890
rect 19620 5090 19720 5340
rect 19800 5090 19900 5340
rect 19620 3660 19900 5090
rect 20100 10590 20300 11300
rect 20100 10510 20110 10590
rect 20290 10510 20300 10590
rect 20100 9790 20300 10510
rect 20100 9710 20110 9790
rect 20290 9710 20300 9790
rect 20100 8990 20300 9710
rect 20100 8910 20110 8990
rect 20290 8910 20300 8990
rect 20100 8190 20300 8910
rect 20100 8110 20110 8190
rect 20290 8110 20300 8190
rect 20100 7390 20300 8110
rect 20100 7310 20110 7390
rect 20290 7310 20300 7390
rect 20100 6590 20300 7310
rect 20100 6510 20110 6590
rect 20290 6510 20300 6590
rect 20100 5790 20300 6510
rect 20100 5710 20110 5790
rect 20290 5710 20300 5790
rect 20100 4990 20300 5710
rect 20100 4910 20110 4990
rect 20290 4910 20300 4990
rect 1620 3150 1630 3330
rect 1810 3150 1820 3330
rect 1620 3140 1820 3150
rect 20100 3330 20300 4910
rect 20100 3150 20110 3330
rect 20290 3150 20300 3330
rect 20100 3140 20300 3150
rect 20500 11250 20700 11300
rect 20500 11170 20510 11250
rect 20690 11170 20700 11250
rect 20500 10450 20700 11170
rect 20500 10370 20510 10450
rect 20690 10370 20700 10450
rect 20500 9650 20700 10370
rect 20500 9570 20510 9650
rect 20690 9570 20700 9650
rect 20500 8850 20700 9570
rect 20500 8770 20510 8850
rect 20690 8770 20700 8850
rect 20500 8050 20700 8770
rect 20500 7970 20510 8050
rect 20690 7970 20700 8050
rect 20500 7250 20700 7970
rect 20500 7170 20510 7250
rect 20690 7170 20700 7250
rect 20500 6450 20700 7170
rect 20500 6370 20510 6450
rect 20690 6370 20700 6450
rect 20500 5650 20700 6370
rect 20500 5570 20510 5650
rect 20690 5570 20700 5650
rect 7800 2930 7940 2940
rect 7800 2810 7810 2930
rect 7930 2810 7940 2930
rect 1220 2400 2270 2600
rect 820 2010 1460 2210
rect 470 -4800 670 -4780
rect 1260 -5570 1460 2010
rect 1260 -5750 1270 -5570
rect 1450 -5750 1460 -5570
rect 1260 -5760 1460 -5750
rect 1250 -7170 1450 -7160
rect 1250 -7350 1260 -7170
rect 1440 -7350 1450 -7170
rect 480 -8090 680 -8080
rect 480 -22200 490 -8090
rect -260 -22380 490 -22200
rect 670 -22380 680 -8090
rect -260 -22400 680 -22380
rect 1250 -22400 1450 -7350
rect 2070 -7570 2270 2400
rect 2070 -7750 2080 -7570
rect 2260 -7750 2270 -7570
rect 2070 -7760 2270 -7750
rect 2800 -5170 3000 -5160
rect 2800 -5350 2810 -5170
rect 2990 -5350 3000 -5170
rect -260 -31660 -60 -22400
rect 820 -22600 1460 -22400
rect 420 -23670 620 -23660
rect 420 -23850 430 -23670
rect 610 -23850 620 -23670
rect 420 -26630 620 -23850
rect 420 -26710 430 -26630
rect 610 -26710 620 -26630
rect 420 -27430 620 -26710
rect 420 -27510 430 -27430
rect 610 -27510 620 -27430
rect 420 -28230 620 -27510
rect 420 -28310 430 -28230
rect 610 -28310 620 -28230
rect 420 -29030 620 -28310
rect 420 -29110 430 -29030
rect 610 -29110 620 -29030
rect 420 -31420 620 -29110
rect 820 -25550 1020 -22600
rect 2800 -22800 3000 -5350
rect 7800 -7870 7940 2810
rect 14900 1980 15040 1990
rect 14900 1320 14910 1980
rect 15030 1320 15040 1980
rect 12870 -1110 13250 -1100
rect 12870 -1260 12880 -1110
rect 13240 -1260 13250 -1110
rect 12870 -1290 13250 -1260
rect 12980 -6820 13080 -1290
rect 14900 -6490 15040 1320
rect 20500 -5570 20700 5570
rect 20900 11110 21100 11300
rect 20900 11030 20910 11110
rect 21090 11030 21100 11110
rect 20900 10310 21100 11030
rect 20900 10230 20910 10310
rect 21090 10230 21100 10310
rect 20900 9510 21100 10230
rect 20900 9430 20910 9510
rect 21090 9430 21100 9510
rect 20900 8710 21100 9430
rect 20900 8630 20910 8710
rect 21090 8630 21100 8710
rect 20900 7910 21100 8630
rect 20900 7830 20910 7910
rect 21090 7830 21100 7910
rect 20900 7110 21100 7830
rect 20900 7030 20910 7110
rect 21090 7030 21100 7110
rect 20900 6310 21100 7030
rect 20900 6230 20910 6310
rect 21090 6230 21100 6310
rect 20900 5510 21100 6230
rect 20900 5430 20910 5510
rect 21090 5430 21100 5510
rect 20900 3340 21100 5430
rect 21300 8990 21500 11300
rect 21300 8910 21310 8990
rect 21490 8910 21500 8990
rect 21300 8190 21500 8910
rect 21300 8110 21310 8190
rect 21490 8110 21500 8190
rect 21300 7390 21500 8110
rect 21300 7310 21310 7390
rect 21490 7310 21500 7390
rect 21300 6590 21500 7310
rect 21300 6510 21310 6590
rect 21490 6510 21500 6590
rect 21300 3730 21500 6510
rect 21300 3550 21310 3730
rect 21490 3550 21500 3730
rect 21820 10940 22100 11500
rect 21820 10690 21920 10940
rect 22000 10690 22100 10940
rect 21820 10140 22100 10690
rect 21820 9890 21920 10140
rect 22000 9890 22100 10140
rect 21820 9340 22100 9890
rect 21820 9090 21920 9340
rect 22000 9090 22100 9340
rect 21820 8540 22100 9090
rect 21820 8290 21920 8540
rect 22000 8290 22100 8540
rect 30306 11060 30706 11500
rect 30306 10932 30326 11060
rect 30682 10932 30706 11060
rect 30306 8850 30706 10932
rect 36880 11010 37060 11020
rect 36880 10850 36890 11010
rect 37050 10850 37060 11010
rect 36880 10840 37060 10850
rect 30306 8450 33490 8850
rect 21820 7740 22100 8290
rect 21820 7490 21920 7740
rect 22000 7490 22100 7740
rect 21820 6940 22100 7490
rect 33090 7186 33490 8450
rect 33090 6976 33108 7186
rect 33474 6976 33490 7186
rect 33090 6960 33490 6976
rect 21820 6690 21920 6940
rect 22000 6690 22100 6940
rect 21820 6140 22100 6690
rect 21820 5890 21920 6140
rect 22000 5890 22100 6140
rect 36220 6260 36420 6270
rect 36220 6080 36230 6260
rect 36410 6080 36420 6260
rect 36220 6070 36420 6080
rect 21820 5340 22100 5890
rect 21820 5090 21920 5340
rect 22000 5090 22100 5340
rect 28490 5400 28670 5410
rect 28490 5240 28500 5400
rect 28660 5240 28670 5400
rect 28490 5230 28670 5240
rect 21820 3660 22100 5090
rect 21300 3540 21500 3550
rect 26200 3400 26380 3410
rect 20900 3140 22260 3340
rect 26200 3240 26210 3400
rect 26370 3370 26380 3400
rect 28530 3370 28630 5230
rect 33120 4110 33300 4120
rect 26370 3270 28630 3370
rect 26370 3240 26380 3270
rect 26200 3230 26380 3240
rect 20500 -5750 20510 -5570
rect 20690 -5750 20700 -5570
rect 20500 -5760 20700 -5750
rect 21270 -5170 21470 -5160
rect 21270 -5350 21280 -5170
rect 21460 -5350 21470 -5170
rect 14900 -6610 14910 -6490
rect 15030 -6610 15040 -6490
rect 14900 -6620 15040 -6610
rect 12940 -6830 13120 -6820
rect 12940 -6990 12950 -6830
rect 13110 -6990 13120 -6830
rect 12940 -7000 13120 -6990
rect 7800 -7990 7810 -7870
rect 7930 -7990 7940 -7870
rect 7800 -8000 7940 -7990
rect 20500 -7170 20700 -7160
rect 20500 -7350 20510 -7170
rect 20690 -7350 20700 -7170
rect 820 -25630 830 -25550
rect 1010 -25630 1020 -25550
rect 820 -26350 1020 -25630
rect 820 -26430 830 -26350
rect 1010 -26430 1020 -26350
rect 820 -27150 1020 -26430
rect 820 -27230 830 -27150
rect 1010 -27230 1020 -27150
rect 820 -27950 1020 -27230
rect 820 -28030 830 -27950
rect 1010 -28030 1020 -27950
rect 820 -28750 1020 -28030
rect 820 -28830 830 -28750
rect 1010 -28830 1020 -28750
rect 820 -29550 1020 -28830
rect 820 -29630 830 -29550
rect 1010 -29630 1020 -29550
rect 820 -30350 1020 -29630
rect 820 -30430 830 -30350
rect 1010 -30430 1020 -30350
rect 820 -31150 1020 -30430
rect 820 -31230 830 -31150
rect 1010 -31230 1020 -31150
rect 820 -31420 1020 -31230
rect 1220 -23000 3000 -22800
rect 1220 -25690 1420 -23000
rect 1220 -25770 1230 -25690
rect 1410 -25770 1420 -25690
rect 1220 -26490 1420 -25770
rect 1220 -26570 1230 -26490
rect 1410 -26570 1420 -26490
rect 1220 -27290 1420 -26570
rect 1220 -27370 1230 -27290
rect 1410 -27370 1420 -27290
rect 1220 -28090 1420 -27370
rect 1220 -28170 1230 -28090
rect 1410 -28170 1420 -28090
rect 1220 -28890 1420 -28170
rect 1220 -28970 1230 -28890
rect 1410 -28970 1420 -28890
rect 1220 -29690 1420 -28970
rect 1220 -29770 1230 -29690
rect 1410 -29770 1420 -29690
rect 1220 -30490 1420 -29770
rect 1220 -30570 1230 -30490
rect 1410 -30570 1420 -30490
rect 1220 -31290 1420 -30570
rect 1220 -31370 1230 -31290
rect 1410 -31370 1420 -31290
rect 1220 -31420 1420 -31370
rect 1620 -23270 1820 -23260
rect 1620 -23450 1630 -23270
rect 1810 -23450 1820 -23270
rect 1620 -25030 1820 -23450
rect 1620 -25110 1630 -25030
rect 1810 -25110 1820 -25030
rect 1620 -25830 1820 -25110
rect 1620 -25910 1630 -25830
rect 1810 -25910 1820 -25830
rect 1620 -26630 1820 -25910
rect 1620 -26710 1630 -26630
rect 1810 -26710 1820 -26630
rect 1620 -27430 1820 -26710
rect 1620 -27510 1630 -27430
rect 1810 -27510 1820 -27430
rect 1620 -28230 1820 -27510
rect 1620 -28310 1630 -28230
rect 1810 -28310 1820 -28230
rect 1620 -29030 1820 -28310
rect 1620 -29110 1630 -29030
rect 1810 -29110 1820 -29030
rect 1620 -29830 1820 -29110
rect 1620 -29910 1630 -29830
rect 1810 -29910 1820 -29830
rect 1620 -30630 1820 -29910
rect 1620 -30710 1630 -30630
rect 1810 -30710 1820 -30630
rect 1620 -31420 1820 -30710
rect 20100 -23270 20300 -23260
rect 20100 -23450 20110 -23270
rect 20290 -23450 20300 -23270
rect 20100 -25030 20300 -23450
rect 20100 -25110 20110 -25030
rect 20290 -25110 20300 -25030
rect 20100 -25830 20300 -25110
rect 20100 -25910 20110 -25830
rect 20290 -25910 20300 -25830
rect 20100 -26630 20300 -25910
rect 20100 -26710 20110 -26630
rect 20290 -26710 20300 -26630
rect 20100 -27430 20300 -26710
rect 20100 -27510 20110 -27430
rect 20290 -27510 20300 -27430
rect 20100 -28230 20300 -27510
rect 20100 -28310 20110 -28230
rect 20290 -28310 20300 -28230
rect 20100 -29030 20300 -28310
rect 20100 -29110 20110 -29030
rect 20290 -29110 20300 -29030
rect 20100 -29830 20300 -29110
rect 20100 -29910 20110 -29830
rect 20290 -29910 20300 -29830
rect 20100 -30630 20300 -29910
rect 20100 -30710 20110 -30630
rect 20290 -30710 20300 -30630
rect 20100 -31420 20300 -30710
rect 20500 -25550 20700 -7350
rect 21270 -22420 21470 -5350
rect 22060 -7570 22260 3140
rect 22060 -7750 22070 -7570
rect 22250 -7750 22260 -7570
rect 22060 -7760 22260 -7750
rect 20500 -25630 20510 -25550
rect 20690 -25630 20700 -25550
rect 20500 -26350 20700 -25630
rect 20500 -26430 20510 -26350
rect 20690 -26430 20700 -26350
rect 20500 -27150 20700 -26430
rect 20500 -27230 20510 -27150
rect 20690 -27230 20700 -27150
rect 20500 -27950 20700 -27230
rect 20500 -28030 20510 -27950
rect 20690 -28030 20700 -27950
rect 20500 -28750 20700 -28030
rect 20500 -28830 20510 -28750
rect 20690 -28830 20700 -28750
rect 20500 -29550 20700 -28830
rect 20500 -29630 20510 -29550
rect 20690 -29630 20700 -29550
rect 20500 -30350 20700 -29630
rect 20500 -30430 20510 -30350
rect 20690 -30430 20700 -30350
rect 20500 -31150 20700 -30430
rect 20500 -31230 20510 -31150
rect 20690 -31230 20700 -31150
rect 20500 -31420 20700 -31230
rect 20900 -22620 21470 -22420
rect 20900 -25690 21100 -22620
rect 20900 -25770 20910 -25690
rect 21090 -25770 21100 -25690
rect 20900 -26490 21100 -25770
rect 20900 -26570 20910 -26490
rect 21090 -26570 21100 -26490
rect 20900 -27290 21100 -26570
rect 20900 -27370 20910 -27290
rect 21090 -27370 21100 -27290
rect 20900 -28090 21100 -27370
rect 20900 -28170 20910 -28090
rect 21090 -28170 21100 -28090
rect 20900 -28890 21100 -28170
rect 20900 -28970 20910 -28890
rect 21090 -28970 21100 -28890
rect 20900 -29690 21100 -28970
rect 20900 -29770 20910 -29690
rect 21090 -29770 21100 -29690
rect 20900 -30490 21100 -29770
rect 20900 -30570 20910 -30490
rect 21090 -30570 21100 -30490
rect 20900 -31290 21100 -30570
rect 20900 -31370 20910 -31290
rect 21090 -31370 21100 -31290
rect 20900 -31420 21100 -31370
rect 21300 -23670 21500 -23660
rect 21300 -23850 21310 -23670
rect 21490 -23850 21500 -23670
rect 21300 -26630 21500 -23850
rect 28530 -24030 28630 3270
rect 30070 4040 30270 4050
rect 30070 3860 30080 4040
rect 30260 3860 30270 4040
rect 30070 -6770 30270 3860
rect 31670 4040 31870 4050
rect 31670 3860 31680 4040
rect 31860 3860 31870 4040
rect 33120 4010 33130 4110
rect 33290 4010 33300 4110
rect 33120 4000 33300 4010
rect 31670 -5970 31870 3860
rect 31670 -6150 31680 -5970
rect 31860 -6150 31870 -5970
rect 31670 -6160 31870 -6150
rect 30070 -6950 30080 -6770
rect 30260 -6950 30270 -6770
rect 30070 -6960 30270 -6950
rect 28490 -24040 28670 -24030
rect 28490 -24200 28500 -24040
rect 28660 -24200 28670 -24040
rect 28490 -24210 28670 -24200
rect 33200 -24920 33300 4000
rect 33020 -24930 33300 -24920
rect 33020 -25000 33030 -24930
rect 33290 -25000 33300 -24930
rect 33020 -25010 33300 -25000
rect 33400 4090 35200 4100
rect 33400 4010 34870 4090
rect 35190 4010 35200 4090
rect 33400 4000 35200 4010
rect 33400 -25070 33500 4000
rect 36020 -5170 36220 -5160
rect 36020 -5350 36030 -5170
rect 36210 -5350 36220 -5170
rect 36020 -5360 36220 -5350
rect 36020 -7870 36120 -5360
rect 36320 -5560 36420 6070
rect 36220 -5570 36420 -5560
rect 36220 -5750 36230 -5570
rect 36410 -5750 36420 -5570
rect 36220 -5760 36420 -5750
rect 36520 6260 36720 6270
rect 36520 6080 36530 6260
rect 36710 6080 36720 6260
rect 36520 6070 36720 6080
rect 36520 -6900 36620 6070
rect 36920 5330 37020 10840
rect 37080 10760 37260 10770
rect 37080 10600 37090 10760
rect 37250 10600 37260 10760
rect 37080 10590 37260 10600
rect 36860 5320 37020 5330
rect 36860 5100 36870 5320
rect 37010 5100 37020 5320
rect 36860 5090 37020 5100
rect 36320 -7000 36620 -6900
rect 36320 -7560 36420 -7000
rect 36220 -7570 36420 -7560
rect 36220 -7750 36230 -7570
rect 36410 -7750 36420 -7570
rect 36220 -7760 36420 -7750
rect 36520 -7170 36720 -7160
rect 36520 -7350 36530 -7170
rect 36710 -7350 36720 -7170
rect 36520 -7360 36720 -7350
rect 36020 -7970 36420 -7870
rect 34900 -16770 35060 -16740
rect 34900 -16920 34910 -16770
rect 35050 -16920 35060 -16770
rect 34900 -22470 35060 -16920
rect 34900 -22610 34910 -22470
rect 35050 -22610 35060 -22470
rect 34900 -22620 35060 -22610
rect 33220 -25080 33500 -25070
rect 33220 -25150 33230 -25080
rect 33490 -25150 33500 -25080
rect 33220 -25160 33500 -25150
rect 21300 -26710 21310 -26630
rect 21490 -26710 21500 -26630
rect 21300 -27430 21500 -26710
rect 36320 -27000 36420 -7970
rect 36020 -27010 36420 -27000
rect 36020 -27140 36030 -27010
rect 36410 -27140 36420 -27010
rect 36020 -27150 36420 -27140
rect 36520 -27000 36620 -7360
rect 36920 -24630 37020 5090
rect 36860 -24640 37020 -24630
rect 36860 -24780 36870 -24640
rect 37010 -24780 37020 -24640
rect 36860 -24790 37020 -24780
rect 37120 5330 37220 10590
rect 37500 7186 37700 7216
rect 37500 6974 37516 7186
rect 37684 6974 37700 7186
rect 37120 5320 37280 5330
rect 37120 5100 37130 5320
rect 37270 5100 37280 5320
rect 37120 5090 37280 5100
rect 37120 -24630 37220 5090
rect 37120 -24640 37280 -24630
rect 37120 -24780 37130 -24640
rect 37270 -24780 37280 -24640
rect 37120 -24790 37280 -24780
rect 36520 -27010 36920 -27000
rect 36520 -27140 36530 -27010
rect 36910 -27140 36920 -27010
rect 36520 -27150 36920 -27140
rect 21300 -27510 21310 -27430
rect 21490 -27510 21500 -27430
rect 21300 -28230 21500 -27510
rect 37500 -27520 37700 6974
rect 36900 -27540 37700 -27520
rect 36900 -27900 36920 -27540
rect 37680 -27900 37700 -27540
rect 36900 -27920 37700 -27900
rect 37900 -28140 38100 7212
rect 21300 -28310 21310 -28230
rect 21490 -28310 21500 -28230
rect 21300 -29030 21500 -28310
rect 21300 -29110 21310 -29030
rect 21490 -29110 21500 -29030
rect 21300 -31420 21500 -29110
rect 30820 -28160 38100 -28140
rect 30820 -28520 36920 -28160
rect 37680 -28520 38100 -28160
rect 30820 -28540 38100 -28520
rect 30820 -31660 31260 -28540
rect -260 -31680 31260 -31660
rect -260 -32060 30840 -31680
rect 30820 -32440 30840 -32060
rect 31240 -32440 31260 -31680
rect 30820 -33520 31260 -32440
rect 38300 -32160 38500 12260
rect 38300 -32180 38540 -32160
rect 38300 -32690 38320 -32180
rect 38520 -32690 38540 -32180
rect 38300 -32910 38310 -32690
rect 38530 -32910 38540 -32690
rect 38300 -32920 38540 -32910
use level_shifter_up  level_shifter_up_0
timestamp 1714698820
transform 1 0 32370 0 1 -31100
box 130 -1700 1108 1948
use level_shifter_up  level_shifter_up_1
timestamp 1714698820
transform 1 0 37370 0 1 -31100
box 130 -1700 1108 1948
use level_shifter_up  level_shifter_up_2
timestamp 1714698820
transform 1 0 36370 0 1 -31100
box 130 -1700 1108 1948
use level_shifter_up  level_shifter_up_3
timestamp 1714698820
transform 1 0 35370 0 1 -31100
box 130 -1700 1108 1948
use level_shifter_up  level_shifter_up_4
timestamp 1714698820
transform 1 0 34370 0 1 -31100
box 130 -1700 1108 1948
use level_shifter_up  level_shifter_up_5
timestamp 1714698820
transform 1 0 33370 0 1 -31100
box 130 -1700 1108 1948
use level_shifter_up  level_shifter_up_6
timestamp 1714698820
transform -1 0 33842 0 -1 11195
box 130 -1700 1108 1948
use level_shifter_up  level_shifter_up_7
timestamp 1714698820
transform -1 0 32242 0 -1 11195
box 130 -1700 1108 1948
use level_shifter_up  level_shifter_up_8
timestamp 1714698820
transform -1 0 33042 0 -1 11195
box 130 -1700 1108 1948
use sky130_fd_pr__nfet_01v8_HWT53N  sky130_fd_pr__nfet_01v8_HWT53N_0 paramcells
timestamp 1713548572
transform 1 0 37081 0 1 10410
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_HWT53N  sky130_fd_pr__nfet_01v8_HWT53N_1
timestamp 1713548572
transform 1 0 37921 0 1 10410
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_HWT53N  sky130_fd_pr__nfet_01v8_HWT53N_2
timestamp 1713548572
transform 1 0 37501 0 1 10410
box -211 -310 211 310
use sky130_fd_pr__nfet_g5v0d10v5_4RA4DJ  sky130_fd_pr__nfet_g5v0d10v5_4RA4DJ_0 paramcells
timestamp 1713585847
transform 1 0 33371 0 1 3758
box -831 -458 831 458
use sky130_fd_pr__nfet_g5v0d10v5_8TUSME  sky130_fd_pr__nfet_g5v0d10v5_8TUSME_0 paramcells
timestamp 1713589649
transform 1 0 36075 0 1 10378
box -515 -458 515 458
use sky130_fd_pr__nfet_g5v0d10v5_46Z5PG  sky130_fd_pr__nfet_g5v0d10v5_46Z5PG_0 paramcells
timestamp 1713585847
transform 1 0 32567 0 1 2828
box -357 -458 357 458
use sky130_fd_pr__nfet_g5v0d10v5_46Z5PG  sky130_fd_pr__nfet_g5v0d10v5_46Z5PG_1
timestamp 1713585847
transform 1 0 35767 0 1 2828
box -357 -458 357 458
use sky130_fd_pr__nfet_g5v0d10v5_46Z5PG  sky130_fd_pr__nfet_g5v0d10v5_46Z5PG_2
timestamp 1713585847
transform 1 0 34167 0 1 2828
box -357 -458 357 458
use sky130_fd_pr__nfet_g5v0d10v5_AUB4P8  sky130_fd_pr__nfet_g5v0d10v5_AUB4P8_0 paramcells
timestamp 1713548572
transform 0 1 9860 -1 0 4380
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_AUB4P8  sky130_fd_pr__nfet_g5v0d10v5_AUB4P8_1
timestamp 1713548572
transform 0 1 12060 -1 0 4380
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_CDNABP  sky130_fd_pr__nfet_g5v0d10v5_CDNABP_0 paramcells
array 0 3 -1800 0 23 1600
timestamp 1713548572
transform 0 1 568 -1 0 -4597
box -328 -767 328 767
use sky130_fd_pr__nfet_g5v0d10v5_EEFBWQ  sky130_fd_pr__nfet_g5v0d10v5_EEFBWQ_0 paramcells
timestamp 1713548572
transform 1 0 28368 0 1 -24912
box -628 -458 628 458
use sky130_fd_pr__nfet_g5v0d10v5_LHNF5N  sky130_fd_pr__nfet_g5v0d10v5_LHNF5N_0 paramcells
timestamp 1713548572
transform 0 1 28367 -1 0 -31075
box -515 -627 515 627
use sky130_fd_pr__nfet_g5v0d10v5_LHNF5N  sky130_fd_pr__nfet_g5v0d10v5_LHNF5N_1
timestamp 1713548572
transform 0 1 28367 -1 0 -28995
box -515 -627 515 627
use sky130_fd_pr__nfet_g5v0d10v5_LHNF5N  sky130_fd_pr__nfet_g5v0d10v5_LHNF5N_2
timestamp 1713548572
transform 0 1 28367 -1 0 -30035
box -515 -627 515 627
use sky130_fd_pr__nfet_g5v0d10v5_LHNF5N  sky130_fd_pr__nfet_g5v0d10v5_LHNF5N_3
timestamp 1713548572
transform 0 1 28367 -1 0 -26915
box -515 -627 515 627
use sky130_fd_pr__nfet_g5v0d10v5_LHNF5N  sky130_fd_pr__nfet_g5v0d10v5_LHNF5N_4
timestamp 1713548572
transform 0 1 28367 -1 0 -27955
box -515 -627 515 627
use sky130_fd_pr__nfet_g5v0d10v5_LHNF5N  sky130_fd_pr__nfet_g5v0d10v5_LHNF5N_5
timestamp 1713548572
transform 0 1 28367 -1 0 -25875
box -515 -627 515 627
use sky130_fd_pr__nfet_g5v0d10v5_LURNA9  sky130_fd_pr__nfet_g5v0d10v5_LURNA9_0 paramcells
timestamp 1713585847
transform 0 -1 36648 1 0 4951
box -1231 -458 1231 458
use sky130_fd_pr__nfet_g5v0d10v5_LURNA9  sky130_fd_pr__nfet_g5v0d10v5_LURNA9_1
timestamp 1713585847
transform 0 -1 37434 1 0 4951
box -1231 -458 1231 458
use sky130_fd_pr__nfet_g5v0d10v5_LUSSBJ  sky130_fd_pr__nfet_g5v0d10v5_LUSSBJ_0 paramcells
timestamp 1713585847
transform 1 0 35166 0 1 3758
box -436 -458 436 458
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_9 paramcells
timestamp 1713548572
transform 0 1 5458 -1 0 5178
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_10
timestamp 1713548572
transform 0 1 5458 -1 0 5978
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_11
timestamp 1713548572
transform 0 1 5458 -1 0 6778
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_12
timestamp 1713548572
transform 0 1 5458 -1 0 7578
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_13
timestamp 1713548572
transform 0 1 5458 -1 0 8378
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_14
timestamp 1713548572
transform 0 1 5458 -1 0 9178
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_15
timestamp 1713548572
transform 0 1 5458 -1 0 9978
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_17
timestamp 1713548572
transform 0 1 3258 -1 0 5178
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_18
timestamp 1713548572
transform 0 1 3258 -1 0 5978
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_19
timestamp 1713548572
transform 0 1 3258 -1 0 6778
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_20
timestamp 1713548572
transform 0 1 3258 -1 0 7578
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_21
timestamp 1713548572
transform 0 1 3258 -1 0 8378
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_22
timestamp 1713548572
transform 0 1 3258 -1 0 9178
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_23
timestamp 1713548572
transform 0 1 3258 -1 0 9978
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_25
timestamp 1713548572
transform 0 1 7658 -1 0 5178
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_26
timestamp 1713548572
transform 0 1 7658 -1 0 5978
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_27
timestamp 1713548572
transform 0 1 7658 -1 0 6778
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_28
timestamp 1713548572
transform 0 1 7658 -1 0 7578
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_29
timestamp 1713548572
transform 0 1 7658 -1 0 8378
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_30
timestamp 1713548572
transform 0 1 7658 -1 0 9178
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_31
timestamp 1713548572
transform 0 1 7658 -1 0 9978
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_32
timestamp 1713548572
transform 0 1 12058 -1 0 9978
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_33
timestamp 1713548572
transform 0 1 12058 -1 0 9178
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_34
timestamp 1713548572
transform 0 1 12058 -1 0 8378
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_35
timestamp 1713548572
transform 0 1 12058 -1 0 7578
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_36
timestamp 1713548572
transform 0 1 12058 -1 0 6778
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_37
timestamp 1713548572
transform 0 1 12058 -1 0 5978
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_38
timestamp 1713548572
transform 0 1 12058 -1 0 5178
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_40
timestamp 1713548572
transform 0 1 9858 -1 0 9978
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_41
timestamp 1713548572
transform 0 1 9858 -1 0 9178
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_42
timestamp 1713548572
transform 0 1 9858 -1 0 8378
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_43
timestamp 1713548572
transform 0 1 9858 -1 0 7578
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_44
timestamp 1713548572
transform 0 1 9858 -1 0 6778
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_45
timestamp 1713548572
transform 0 1 9858 -1 0 5978
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_46
timestamp 1713548572
transform 0 1 9858 -1 0 5178
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_49
timestamp 1713548572
transform 0 1 14258 -1 0 7578
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_50
timestamp 1713548572
transform 0 1 14258 -1 0 6778
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_51
timestamp 1713548572
transform 0 1 14258 -1 0 5978
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_52
timestamp 1713548572
transform 0 1 14258 -1 0 5178
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_53
timestamp 1713548572
transform 0 1 14258 -1 0 9978
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_54
timestamp 1713548572
transform 0 1 14258 -1 0 9178
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_55
timestamp 1713548572
transform 0 1 14258 -1 0 8378
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_57
timestamp 1713548572
transform 0 1 16458 -1 0 7578
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_58
timestamp 1713548572
transform 0 1 16458 -1 0 6778
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_59
timestamp 1713548572
transform 0 1 16458 -1 0 5978
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_60
timestamp 1713548572
transform 0 1 16458 -1 0 5178
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_61
timestamp 1713548572
transform 0 1 16458 -1 0 9978
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_62
timestamp 1713548572
transform 0 1 16458 -1 0 9178
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_63
timestamp 1713548572
transform 0 1 16458 -1 0 8378
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_73
timestamp 1713548572
transform 0 1 3258 -1 0 10778
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_74
timestamp 1713548572
transform 0 1 5458 -1 0 10778
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_75
timestamp 1713548572
transform 0 1 7658 -1 0 10778
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_76
timestamp 1713548572
transform 0 1 9858 -1 0 10778
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_77
timestamp 1713548572
transform 0 1 12058 -1 0 10778
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_78
timestamp 1713548572
transform 0 1 14258 -1 0 10778
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_79
timestamp 1713548572
transform 0 1 16458 -1 0 10778
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_81
timestamp 1713548572
transform 0 1 18658 -1 0 10778
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_82
timestamp 1713548572
transform 0 1 18658 -1 0 9978
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_83
timestamp 1713548572
transform 0 1 18658 -1 0 9178
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_84
timestamp 1713548572
transform 0 1 18658 -1 0 8378
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_85
timestamp 1713548572
transform 0 1 18658 -1 0 7578
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_86
timestamp 1713548572
transform 0 1 18658 -1 0 6778
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_87
timestamp 1713548572
transform 0 1 18658 -1 0 5978
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_M7X63G  sky130_fd_pr__nfet_g5v0d10v5_M7X63G_88
timestamp 1713548572
transform 0 1 18658 -1 0 5178
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_MMHSE7  sky130_fd_pr__nfet_g5v0d10v5_MMHSE7_0 paramcells
timestamp 1715629873
transform 0 1 35838 -1 0 8348
box -328 -658 328 658
use sky130_fd_pr__nfet_g5v0d10v5_MMHSE7  sky130_fd_pr__nfet_g5v0d10v5_MMHSE7_1
timestamp 1715629873
transform 0 1 35838 -1 0 9604
box -328 -658 328 658
use sky130_fd_pr__nfet_g5v0d10v5_MRHAE7  sky130_fd_pr__nfet_g5v0d10v5_MRHAE7_0 paramcells
timestamp 1715629873
transform 0 1 37138 -1 0 8348
box -328 -658 328 658
use sky130_fd_pr__nfet_g5v0d10v5_MRHAE7  sky130_fd_pr__nfet_g5v0d10v5_MRHAE7_1
timestamp 1715629873
transform 0 1 37138 -1 0 9604
box -328 -658 328 658
use sky130_fd_pr__nfet_g5v0d10v5_RM8L2M  sky130_fd_pr__nfet_g5v0d10v5_RM8L2M_0 paramcells
timestamp 1713587898
transform 1 0 36929 0 1 7709
box -428 -308 428 308
use sky130_fd_pr__nfet_g5v0d10v5_RRA4TL  sky130_fd_pr__nfet_g5v0d10v5_RRA4TL_0 paramcells
timestamp 1713587898
transform 1 0 36069 0 1 7709
box -428 -308 428 308
use sky130_fd_pr__nfet_g5v0d10v5_T8W2FW  sky130_fd_pr__nfet_g5v0d10v5_T8W2FW_0 paramcells
timestamp 1713548572
transform 0 1 1059 -1 0 9179
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_T8W2FW  sky130_fd_pr__nfet_g5v0d10v5_T8W2FW_1
timestamp 1713548572
transform 0 1 1059 -1 0 9979
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_T8W2FW  sky130_fd_pr__nfet_g5v0d10v5_T8W2FW_2
timestamp 1713548572
transform 0 1 1059 -1 0 10779
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_T8W2FW  sky130_fd_pr__nfet_g5v0d10v5_T8W2FW_3
timestamp 1713548572
transform 0 1 1059 -1 0 11579
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_T8W2FW  sky130_fd_pr__nfet_g5v0d10v5_T8W2FW_4
timestamp 1713548572
transform 0 1 1059 -1 0 8379
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_T8W2FW  sky130_fd_pr__nfet_g5v0d10v5_T8W2FW_5
timestamp 1713548572
transform 0 1 1059 -1 0 7579
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_T8W2FW  sky130_fd_pr__nfet_g5v0d10v5_T8W2FW_6
timestamp 1713548572
transform 0 1 1059 -1 0 4379
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_T8W2FW  sky130_fd_pr__nfet_g5v0d10v5_T8W2FW_7
timestamp 1713548572
transform 0 1 1059 -1 0 6779
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_T8W2FW  sky130_fd_pr__nfet_g5v0d10v5_T8W2FW_8
timestamp 1713548572
transform 0 1 1059 -1 0 5979
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_T8W2FW  sky130_fd_pr__nfet_g5v0d10v5_T8W2FW_9
timestamp 1713548572
transform 0 1 1059 -1 0 5179
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_T8W2FW  sky130_fd_pr__nfet_g5v0d10v5_T8W2FW_10
timestamp 1713548572
transform 0 1 3259 -1 0 4379
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_T8W2FW  sky130_fd_pr__nfet_g5v0d10v5_T8W2FW_11
timestamp 1713548572
transform 0 1 5459 -1 0 4379
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_T8W2FW  sky130_fd_pr__nfet_g5v0d10v5_T8W2FW_12
timestamp 1713548572
transform 0 1 7659 -1 0 4379
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_T8W2FW  sky130_fd_pr__nfet_g5v0d10v5_T8W2FW_15
timestamp 1713548572
transform 0 1 14259 -1 0 4379
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_T8W2FW  sky130_fd_pr__nfet_g5v0d10v5_T8W2FW_16
timestamp 1713548572
transform 0 1 16459 -1 0 4379
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_T8W2FW  sky130_fd_pr__nfet_g5v0d10v5_T8W2FW_17
timestamp 1713548572
transform 0 1 18659 -1 0 4379
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_T8W2FW  sky130_fd_pr__nfet_g5v0d10v5_T8W2FW_18
timestamp 1713548572
transform 0 1 3259 -1 0 11579
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_T8W2FW  sky130_fd_pr__nfet_g5v0d10v5_T8W2FW_19
timestamp 1713548572
transform 0 1 20859 -1 0 4379
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_T8W2FW  sky130_fd_pr__nfet_g5v0d10v5_T8W2FW_20
timestamp 1713548572
transform 0 1 20859 -1 0 5179
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_T8W2FW  sky130_fd_pr__nfet_g5v0d10v5_T8W2FW_21
timestamp 1713548572
transform 0 1 20859 -1 0 5979
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_T8W2FW  sky130_fd_pr__nfet_g5v0d10v5_T8W2FW_22
timestamp 1713548572
transform 0 1 20859 -1 0 6779
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_T8W2FW  sky130_fd_pr__nfet_g5v0d10v5_T8W2FW_23
timestamp 1713548572
transform 0 1 20859 -1 0 7579
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_T8W2FW  sky130_fd_pr__nfet_g5v0d10v5_T8W2FW_24
timestamp 1713548572
transform 0 1 20859 -1 0 8379
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_T8W2FW  sky130_fd_pr__nfet_g5v0d10v5_T8W2FW_25
timestamp 1713548572
transform 0 1 20859 -1 0 9179
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_T8W2FW  sky130_fd_pr__nfet_g5v0d10v5_T8W2FW_26
timestamp 1713548572
transform 0 1 20859 -1 0 9979
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_T8W2FW  sky130_fd_pr__nfet_g5v0d10v5_T8W2FW_27
timestamp 1713548572
transform 0 1 20859 -1 0 10779
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_T8W2FW  sky130_fd_pr__nfet_g5v0d10v5_T8W2FW_28
timestamp 1713548572
transform 0 1 20859 -1 0 11579
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_T8W2FW  sky130_fd_pr__nfet_g5v0d10v5_T8W2FW_29
timestamp 1713548572
transform 0 1 18659 -1 0 11579
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_T8W2FW  sky130_fd_pr__nfet_g5v0d10v5_T8W2FW_30
timestamp 1713548572
transform 0 1 16459 -1 0 11579
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_T8W2FW  sky130_fd_pr__nfet_g5v0d10v5_T8W2FW_31
timestamp 1713548572
transform 0 1 14259 -1 0 11579
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_T8W2FW  sky130_fd_pr__nfet_g5v0d10v5_T8W2FW_32
timestamp 1713548572
transform 0 1 12059 -1 0 11579
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_T8W2FW  sky130_fd_pr__nfet_g5v0d10v5_T8W2FW_33
timestamp 1713548572
transform 0 1 9859 -1 0 11579
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_T8W2FW  sky130_fd_pr__nfet_g5v0d10v5_T8W2FW_34
timestamp 1713548572
transform 0 1 7659 -1 0 11579
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_T8W2FW  sky130_fd_pr__nfet_g5v0d10v5_T8W2FW_35
timestamp 1713548572
transform 0 1 5459 -1 0 11579
box -378 -1058 378 1058
use sky130_fd_pr__nfet_g5v0d10v5_TAUUP3  sky130_fd_pr__nfet_g5v0d10v5_TAUUP3_0 paramcells
timestamp 1713548572
transform 1 0 17435 0 1 2947
box -515 -627 515 627
use sky130_fd_pr__nfet_g5v0d10v5_WGHV7X  sky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0 paramcells
array 0 3 -1800 0 23 1600
timestamp 1713585847
transform 0 1 568 -1 0 -3751
box -628 -767 628 767
use sky130_fd_pr__pfet_01v8_EPRAC4  sky130_fd_pr__pfet_01v8_EPRAC4_0 paramcells
timestamp 1713548572
transform 1 0 37921 0 1 11489
box -211 -419 211 419
use sky130_fd_pr__pfet_01v8_EPRAC4  sky130_fd_pr__pfet_01v8_EPRAC4_1
timestamp 1713548572
transform 1 0 37081 0 1 11489
box -211 -419 211 419
use sky130_fd_pr__pfet_01v8_EPRAC4  sky130_fd_pr__pfet_01v8_EPRAC4_2
timestamp 1713548572
transform 1 0 37501 0 1 11489
box -211 -419 211 419
use sky130_fd_pr__pfet_01v8_YTEHH6  sky130_fd_pr__pfet_01v8_YTEHH6_0 paramcells
timestamp 1713597193
transform 1 0 35595 0 1 11689
box -425 -619 425 619
use sky130_fd_pr__pfet_01v8_YTEHH6  sky130_fd_pr__pfet_01v8_YTEHH6_1
timestamp 1713597193
transform 1 0 36445 0 1 11689
box -425 -619 425 619
use sky130_fd_pr__pfet_g5v0d10v5_2CKAKF  sky130_fd_pr__pfet_g5v0d10v5_2CKAKF_0 paramcells
timestamp 1713548572
transform 1 0 35823 0 1 -23963
box -1493 -497 1493 497
use sky130_fd_pr__pfet_g5v0d10v5_6UJQA2  sky130_fd_pr__pfet_g5v0d10v5_6UJQA2_0 paramcells
timestamp 1713548572
transform -1 0 28685 0 -1 -23108
box -545 -662 545 662
use sky130_fd_pr__pfet_g5v0d10v5_8JQF8T  sky130_fd_pr__pfet_g5v0d10v5_8JQF8T_0 paramcells
timestamp 1713585847
transform 0 1 30775 -1 0 4998
box -358 -1215 358 1215
use sky130_fd_pr__pfet_g5v0d10v5_2432J2  sky130_fd_pr__pfet_g5v0d10v5_2432J2_1 paramcells
timestamp 1713548572
transform 1 0 32965 0 1 -22823
box -545 -497 545 497
use sky130_fd_pr__pfet_g5v0d10v5_9432CF  sky130_fd_pr__pfet_g5v0d10v5_9432CF_0 paramcells
timestamp 1713548572
transform 1 0 33661 0 1 -23965
box -703 -497 703 497
use sky130_fd_pr__pfet_g5v0d10v5_ASR39J  sky130_fd_pr__pfet_g5v0d10v5_ASR39J_0 paramcells
timestamp 1713548572
transform 1 0 38220 0 1 2040
box 0 0 1 1
use sky130_fd_pr__pfet_g5v0d10v5_CRL9SD  sky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0 paramcells
array 0 7 -800 0 7 2200
timestamp 1713548572
transform 0 1 3267 -1 0 -30902
box -408 -1097 408 1097
use sky130_fd_pr__pfet_g5v0d10v5_CS979Q  sky130_fd_pr__pfet_g5v0d10v5_CS979Q_0 paramcells
array 0 7 -1800 0 23 1600
timestamp 1713548572
transform 0 1 575 -1 0 -21742
box -658 -815 658 815
use sky130_fd_pr__pfet_g5v0d10v5_GHE6BF  sky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0 paramcells
array 0 7 -1800 0 23 1600
timestamp 1713548572
transform 0 1 575 -1 0 -20916
box -358 -815 358 815
use sky130_fd_pr__pfet_g5v0d10v5_N8ANR9  sky130_fd_pr__pfet_g5v0d10v5_N8ANR9_0 paramcells
timestamp 1713585847
transform 0 -1 28362 1 0 5925
box -545 -662 545 662
use sky130_fd_pr__pfet_g5v0d10v5_N8ANR9  sky130_fd_pr__pfet_g5v0d10v5_N8ANR9_1
timestamp 1713585847
transform 0 -1 28362 1 0 11125
box -545 -662 545 662
use sky130_fd_pr__pfet_g5v0d10v5_N8ANR9  sky130_fd_pr__pfet_g5v0d10v5_N8ANR9_2
timestamp 1713585847
transform 0 -1 28362 1 0 10085
box -545 -662 545 662
use sky130_fd_pr__pfet_g5v0d10v5_N8ANR9  sky130_fd_pr__pfet_g5v0d10v5_N8ANR9_3
timestamp 1713585847
transform 0 -1 28362 1 0 9045
box -545 -662 545 662
use sky130_fd_pr__pfet_g5v0d10v5_N8ANR9  sky130_fd_pr__pfet_g5v0d10v5_N8ANR9_4
timestamp 1713585847
transform 0 -1 28362 1 0 8005
box -545 -662 545 662
use sky130_fd_pr__pfet_g5v0d10v5_N8ANR9  sky130_fd_pr__pfet_g5v0d10v5_N8ANR9_5
timestamp 1713585847
transform 0 -1 28362 1 0 6965
box -545 -662 545 662
use sky130_fd_pr__pfet_g5v0d10v5_PNRDLC  sky130_fd_pr__pfet_g5v0d10v5_PNRDLC_0 paramcells
timestamp 1713548572
transform 0 1 20867 -1 0 -25302
box -408 -1097 408 1097
use sky130_fd_pr__pfet_g5v0d10v5_PNRDLC  sky130_fd_pr__pfet_g5v0d10v5_PNRDLC_1
timestamp 1713548572
transform 0 1 3267 -1 0 -31702
box -408 -1097 408 1097
use sky130_fd_pr__pfet_g5v0d10v5_PNRDLC  sky130_fd_pr__pfet_g5v0d10v5_PNRDLC_2
timestamp 1713548572
transform 0 1 5467 -1 0 -31702
box -408 -1097 408 1097
use sky130_fd_pr__pfet_g5v0d10v5_PNRDLC  sky130_fd_pr__pfet_g5v0d10v5_PNRDLC_3
timestamp 1713548572
transform 0 1 7667 -1 0 -31702
box -408 -1097 408 1097
use sky130_fd_pr__pfet_g5v0d10v5_PNRDLC  sky130_fd_pr__pfet_g5v0d10v5_PNRDLC_4
timestamp 1713548572
transform 0 1 9867 -1 0 -31702
box -408 -1097 408 1097
use sky130_fd_pr__pfet_g5v0d10v5_PNRDLC  sky130_fd_pr__pfet_g5v0d10v5_PNRDLC_5
timestamp 1713548572
transform 0 1 12067 -1 0 -31702
box -408 -1097 408 1097
use sky130_fd_pr__pfet_g5v0d10v5_PNRDLC  sky130_fd_pr__pfet_g5v0d10v5_PNRDLC_6
timestamp 1713548572
transform 0 1 14267 -1 0 -31702
box -408 -1097 408 1097
use sky130_fd_pr__pfet_g5v0d10v5_PNRDLC  sky130_fd_pr__pfet_g5v0d10v5_PNRDLC_7
timestamp 1713548572
transform 0 1 16467 -1 0 -31702
box -408 -1097 408 1097
use sky130_fd_pr__pfet_g5v0d10v5_PNRDLC  sky130_fd_pr__pfet_g5v0d10v5_PNRDLC_8
timestamp 1713548572
transform 0 1 18667 -1 0 -31702
box -408 -1097 408 1097
use sky130_fd_pr__pfet_g5v0d10v5_PNRDLC  sky130_fd_pr__pfet_g5v0d10v5_PNRDLC_9
timestamp 1713548572
transform 0 1 20867 -1 0 -31702
box -408 -1097 408 1097
use sky130_fd_pr__pfet_g5v0d10v5_PNRDLC  sky130_fd_pr__pfet_g5v0d10v5_PNRDLC_10
timestamp 1713548572
transform 0 1 20867 -1 0 -30902
box -408 -1097 408 1097
use sky130_fd_pr__pfet_g5v0d10v5_PNRDLC  sky130_fd_pr__pfet_g5v0d10v5_PNRDLC_11
timestamp 1713548572
transform 0 1 20867 -1 0 -30102
box -408 -1097 408 1097
use sky130_fd_pr__pfet_g5v0d10v5_PNRDLC  sky130_fd_pr__pfet_g5v0d10v5_PNRDLC_12
timestamp 1713548572
transform 0 1 20867 -1 0 -29302
box -408 -1097 408 1097
use sky130_fd_pr__pfet_g5v0d10v5_PNRDLC  sky130_fd_pr__pfet_g5v0d10v5_PNRDLC_13
timestamp 1713548572
transform 0 1 20867 -1 0 -28502
box -408 -1097 408 1097
use sky130_fd_pr__pfet_g5v0d10v5_PNRDLC  sky130_fd_pr__pfet_g5v0d10v5_PNRDLC_14
timestamp 1713548572
transform 0 1 20867 -1 0 -27702
box -408 -1097 408 1097
use sky130_fd_pr__pfet_g5v0d10v5_PNRDLC  sky130_fd_pr__pfet_g5v0d10v5_PNRDLC_15
timestamp 1713548572
transform 0 1 20867 -1 0 -26902
box -408 -1097 408 1097
use sky130_fd_pr__pfet_g5v0d10v5_PNRDLC  sky130_fd_pr__pfet_g5v0d10v5_PNRDLC_16
timestamp 1713548572
transform 0 1 20867 -1 0 -26102
box -408 -1097 408 1097
use sky130_fd_pr__pfet_g5v0d10v5_PNRDLC  sky130_fd_pr__pfet_g5v0d10v5_PNRDLC_17
timestamp 1713548572
transform 0 1 1067 -1 0 -31702
box -408 -1097 408 1097
use sky130_fd_pr__pfet_g5v0d10v5_PNRDLC  sky130_fd_pr__pfet_g5v0d10v5_PNRDLC_18
timestamp 1713548572
transform 0 1 20867 -1 0 -24502
box -408 -1097 408 1097
use sky130_fd_pr__pfet_g5v0d10v5_PNRDLC  sky130_fd_pr__pfet_g5v0d10v5_PNRDLC_19
timestamp 1713548572
transform 0 1 18667 -1 0 -24502
box -408 -1097 408 1097
use sky130_fd_pr__pfet_g5v0d10v5_PNRDLC  sky130_fd_pr__pfet_g5v0d10v5_PNRDLC_20
timestamp 1713548572
transform 0 1 16467 -1 0 -24502
box -408 -1097 408 1097
use sky130_fd_pr__pfet_g5v0d10v5_PNRDLC  sky130_fd_pr__pfet_g5v0d10v5_PNRDLC_21
timestamp 1713548572
transform 0 1 14267 -1 0 -24502
box -408 -1097 408 1097
use sky130_fd_pr__pfet_g5v0d10v5_PNRDLC  sky130_fd_pr__pfet_g5v0d10v5_PNRDLC_22
timestamp 1713548572
transform 0 1 12067 -1 0 -24502
box -408 -1097 408 1097
use sky130_fd_pr__pfet_g5v0d10v5_PNRDLC  sky130_fd_pr__pfet_g5v0d10v5_PNRDLC_23
timestamp 1713548572
transform 0 1 9867 -1 0 -24502
box -408 -1097 408 1097
use sky130_fd_pr__pfet_g5v0d10v5_PNRDLC  sky130_fd_pr__pfet_g5v0d10v5_PNRDLC_24
timestamp 1713548572
transform 0 1 7667 -1 0 -24502
box -408 -1097 408 1097
use sky130_fd_pr__pfet_g5v0d10v5_PNRDLC  sky130_fd_pr__pfet_g5v0d10v5_PNRDLC_25
timestamp 1713548572
transform 0 1 5467 -1 0 -24502
box -408 -1097 408 1097
use sky130_fd_pr__pfet_g5v0d10v5_PNRDLC  sky130_fd_pr__pfet_g5v0d10v5_PNRDLC_26
timestamp 1713548572
transform 0 1 3267 -1 0 -24502
box -408 -1097 408 1097
use sky130_fd_pr__pfet_g5v0d10v5_PNRDLC  sky130_fd_pr__pfet_g5v0d10v5_PNRDLC_27
timestamp 1713548572
transform 0 1 1067 -1 0 -24502
box -408 -1097 408 1097
use sky130_fd_pr__pfet_g5v0d10v5_PNRDLC  sky130_fd_pr__pfet_g5v0d10v5_PNRDLC_28
timestamp 1713548572
transform 0 1 1067 -1 0 -25302
box -408 -1097 408 1097
use sky130_fd_pr__pfet_g5v0d10v5_PNRDLC  sky130_fd_pr__pfet_g5v0d10v5_PNRDLC_29
timestamp 1713548572
transform 0 1 1067 -1 0 -26102
box -408 -1097 408 1097
use sky130_fd_pr__pfet_g5v0d10v5_PNRDLC  sky130_fd_pr__pfet_g5v0d10v5_PNRDLC_30
timestamp 1713548572
transform 0 1 1067 -1 0 -26902
box -408 -1097 408 1097
use sky130_fd_pr__pfet_g5v0d10v5_PNRDLC  sky130_fd_pr__pfet_g5v0d10v5_PNRDLC_31
timestamp 1713548572
transform 0 1 1067 -1 0 -27702
box -408 -1097 408 1097
use sky130_fd_pr__pfet_g5v0d10v5_PNRDLC  sky130_fd_pr__pfet_g5v0d10v5_PNRDLC_32
timestamp 1713548572
transform 0 1 1067 -1 0 -28502
box -408 -1097 408 1097
use sky130_fd_pr__pfet_g5v0d10v5_PNRDLC  sky130_fd_pr__pfet_g5v0d10v5_PNRDLC_33
timestamp 1713548572
transform 0 1 1067 -1 0 -29302
box -408 -1097 408 1097
use sky130_fd_pr__pfet_g5v0d10v5_PNRDLC  sky130_fd_pr__pfet_g5v0d10v5_PNRDLC_34
timestamp 1713548572
transform 0 1 1067 -1 0 -30102
box -408 -1097 408 1097
use sky130_fd_pr__pfet_g5v0d10v5_PNRDLC  sky130_fd_pr__pfet_g5v0d10v5_PNRDLC_35
timestamp 1713548572
transform 0 1 1067 -1 0 -30902
box -408 -1097 408 1097
use sky130_fd_pr__pfet_g5v0d10v5_Q8UPKT  sky130_fd_pr__pfet_g5v0d10v5_Q8UPKT_0 paramcells
timestamp 1713585847
transform 1 0 30767 0 1 6155
box -1087 -815 1087 815
use sky130_fd_pr__pfet_g5v0d10v5_REE66T  sky130_fd_pr__pfet_g5v0d10v5_REE66T_0 paramcells
timestamp 1713548572
transform 0 -1 35377 1 0 -25879
box -1261 -697 1261 697
use sky130_fd_pr__pfet_g5v0d10v5_REE66T  sky130_fd_pr__pfet_g5v0d10v5_REE66T_1
timestamp 1713548572
transform 0 -1 36717 1 0 -25879
box -1261 -697 1261 697
use sky130_fd_pr__pfet_g5v0d10v5_RJSTGP  sky130_fd_pr__pfet_g5v0d10v5_RJSTGP_0 paramcells
timestamp 1713585847
transform -1 0 30767 0 -1 7477
box -1087 -497 1087 497
use sky130_fd_pr__pfet_g5v0d10v5_RUG6CB  sky130_fd_pr__pfet_g5v0d10v5_RUG6CB_0 paramcells
timestamp 1713585847
transform 1 0 28358 0 1 4757
box -658 -697 658 697
use sky130_fd_pr__pfet_g5v0d10v5_X332GA  sky130_fd_pr__pfet_g5v0d10v5_X332GA_0 paramcells
timestamp 1713548572
transform 1 0 34177 0 1 -22843
box -387 -497 387 497
use sky130_fd_pr__res_high_po_2p85_EP2UD7  sky130_fd_pr__res_high_po_2p85_EP2UD7_0 paramcells
timestamp 1713601876
transform 1 0 24661 0 1 8202
box -2503 -3844 2503 3844
use sky130_fd_pr__res_high_po_2p85_EP2UD7  sky130_fd_pr__res_high_po_2p85_EP2UD7_1
timestamp 1713601876
transform 1 0 24621 0 1 -28298
box -2503 -3844 2503 3844
<< labels >>
flabel metal3 25908 -6132 26054 -5988 0 FreeSans 160 0 0 0 Vom
flabel metal3 25946 -6922 26060 -6808 0 FreeSans 160 0 0 0 Vop
flabel metal3 34058 -5336 34206 -5190 0 FreeSans 160 0 0 0 Vfold_bot_m
flabel metal3 5232 -23424 5384 -23282 0 FreeSans 160 0 0 0 Vxp
flabel metal3 5272 3160 5424 3302 0 FreeSans 160 0 0 0 Vxm
flabel metal2 11724 -850 11812 -754 0 FreeSans 160 0 0 0 bias_n
flabel metal1 12984 -776 13110 -652 0 FreeSans 160 0 0 0 casc_n
flabel metal1 16736 -8368 16836 -8274 0 FreeSans 160 0 0 0 casc_p
flabel metal1 11734 -10518 11822 -10426 0 FreeSans 160 0 0 0 bias_p
flabel metal2 15250 -1268 15372 -1144 0 FreeSans 160 0 0 0 bias_var_n
flabel metal3 31130 -28780 31200 -28710 0 FreeSans 160 0 0 0 enb_hv
flabel metal3 31130 -28930 31200 -28860 0 FreeSans 160 0 0 0 en_hv
flabel metal3 31130 -29080 31200 -29010 0 FreeSans 160 0 0 0 hyst1b_hv
flabel metal3 31130 -29230 31200 -29160 0 FreeSans 160 0 0 0 hyst1_hv
flabel metal3 31130 -29380 31200 -29310 0 FreeSans 160 0 0 0 hyst0b_hv
flabel metal3 31130 -29530 31200 -29460 0 FreeSans 160 0 0 0 hyst0_hv
flabel metal2 26540 -29250 26700 -29080 0 FreeSans 160 0 0 0 res_p_bot
flabel metal3 30640 -30480 30710 -30410 0 FreeSans 320 0 0 0 trim5_hv
flabel metal3 30640 -30630 30710 -30560 0 FreeSans 320 0 0 0 trim5b_hv
flabel metal3 30640 -30780 30710 -30710 0 FreeSans 320 0 0 0 trim4b_hv
flabel metal3 30640 -30930 30710 -30860 0 FreeSans 320 0 0 0 trim3b_hv
flabel metal3 -1580 -6980 -1380 -6780 0 FreeSans 320 0 0 0 Vinm
port 1 nsew
flabel metal3 -1580 -6140 -1380 -5940 0 FreeSans 320 0 0 0 Vinp
port 0 nsew
flabel metal2 33000 13310 33090 13400 0 FreeSans 320 0 0 0 trim[0]
port 12 nsew
flabel metal2 32200 13310 32290 13400 0 FreeSans 320 0 0 0 trim[1]
port 11 nsew
flabel metal2 31400 13310 31490 13400 0 FreeSans 320 0 0 0 trim[2]
port 10 nsew
flabel metal2 33120 -33520 33220 -33420 0 FreeSans 320 0 0 0 trim[5]
port 7 nsew
flabel metal2 34120 -33520 34220 -33420 0 FreeSans 320 0 0 0 trim[4]
port 8 nsew
flabel metal2 35120 -33520 35220 -33420 0 FreeSans 320 0 0 0 trim[3]
port 9 nsew
flabel metal2 36120 -33520 36220 -33420 0 FreeSans 320 0 0 0 en
port 4 nsew
flabel metal2 37120 -33520 37220 -33420 0 FreeSans 320 0 0 0 hyst[1]
port 5 nsew
flabel metal2 38120 -33520 38220 -33420 0 FreeSans 320 0 0 0 hyst[0]
port 6 nsew
flabel metal4 39260 12300 39480 12520 0 FreeSans 320 0 0 0 DVDD
port 14 nsew
flabel metal3 39400 10820 39500 10920 0 FreeSans 320 0 0 0 Vout
port 13 nsew
flabel metal4 29080 13320 29260 13500 0 FreeSans 320 0 0 0 AGND
port 3 nsew
flabel metal3 -1740 2400 -1600 2540 0 FreeSans 320 0 0 0 ibias
port 15 nsew
flabel metal4 30940 -33500 31140 -33340 0 FreeSans 320 0 0 0 AVDD
port 2 nsew
flabel metal1 38924 -31962 39430 -31470 0 FreeSans 480 0 0 0 DGND
port 16 nsew
<< properties >>
string MASKHINTS_HVI -200 -4926 38136 2278
<< end >>
