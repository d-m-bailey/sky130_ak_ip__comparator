magic
tech sky130A
magscale 1 2
timestamp 1713319068
<< pwell >>
rect -515 -627 515 627
<< mvnmos >>
rect -287 -369 -187 431
rect -129 -369 -29 431
rect 29 -369 129 431
rect 187 -369 287 431
<< mvndiff >>
rect -345 419 -287 431
rect -345 -357 -333 419
rect -299 -357 -287 419
rect -345 -369 -287 -357
rect -187 419 -129 431
rect -187 -357 -175 419
rect -141 -357 -129 419
rect -187 -369 -129 -357
rect -29 419 29 431
rect -29 -357 -17 419
rect 17 -357 29 419
rect -29 -369 29 -357
rect 129 419 187 431
rect 129 -357 141 419
rect 175 -357 187 419
rect 129 -369 187 -357
rect 287 419 345 431
rect 287 -357 299 419
rect 333 -357 345 419
rect 287 -369 345 -357
<< mvndiffc >>
rect -333 -357 -299 419
rect -175 -357 -141 419
rect -17 -357 17 419
rect 141 -357 175 419
rect 299 -357 333 419
<< mvpsubdiff >>
rect -479 579 479 591
rect -479 545 -371 579
rect 371 545 479 579
rect -479 533 479 545
rect -479 483 -421 533
rect -479 -483 -467 483
rect -433 -483 -421 483
rect 421 483 479 533
rect -479 -533 -421 -483
rect 421 -483 433 483
rect 467 -483 479 483
rect 421 -533 479 -483
rect -479 -545 479 -533
rect -479 -579 -371 -545
rect 371 -579 479 -545
rect -479 -591 479 -579
<< mvpsubdiffcont >>
rect -371 545 371 579
rect -467 -483 -433 483
rect 433 -483 467 483
rect -371 -579 371 -545
<< poly >>
rect -287 431 -187 457
rect -129 431 -29 457
rect 29 431 129 457
rect 187 431 287 457
rect -287 -407 -187 -369
rect -287 -441 -271 -407
rect -203 -441 -187 -407
rect -287 -457 -187 -441
rect -129 -407 -29 -369
rect -129 -441 -113 -407
rect -45 -441 -29 -407
rect -129 -457 -29 -441
rect 29 -407 129 -369
rect 29 -441 45 -407
rect 113 -441 129 -407
rect 29 -457 129 -441
rect 187 -407 287 -369
rect 187 -441 203 -407
rect 271 -441 287 -407
rect 187 -457 287 -441
<< polycont >>
rect -271 -441 -203 -407
rect -113 -441 -45 -407
rect 45 -441 113 -407
rect 203 -441 271 -407
<< locali >>
rect -467 545 -371 579
rect 371 545 467 579
rect -467 483 -433 545
rect 433 483 467 545
rect -333 419 -299 435
rect -333 -373 -299 -357
rect -175 419 -141 435
rect -175 -373 -141 -357
rect -17 419 17 435
rect -17 -373 17 -357
rect 141 419 175 435
rect 141 -373 175 -357
rect 299 419 333 435
rect 299 -373 333 -357
rect -287 -441 -271 -407
rect -203 -441 -187 -407
rect -129 -441 -113 -407
rect -45 -441 -29 -407
rect 29 -441 45 -407
rect 113 -441 129 -407
rect 187 -441 203 -407
rect 271 -441 287 -407
rect -467 -545 -433 -483
rect 433 -545 467 -483
rect -467 -579 -371 -545
rect 371 -579 467 -545
<< viali >>
rect -333 -357 -299 419
rect -175 -357 -141 419
rect -17 -357 17 419
rect 141 -357 175 419
rect 299 -357 333 419
rect -271 -441 -203 -407
rect -113 -441 -45 -407
rect 45 -441 113 -407
rect 203 -441 271 -407
<< metal1 >>
rect -339 419 -293 431
rect -339 -357 -333 419
rect -299 -357 -293 419
rect -339 -369 -293 -357
rect -181 419 -135 431
rect -181 -357 -175 419
rect -141 -357 -135 419
rect -181 -369 -135 -357
rect -23 419 23 431
rect -23 -357 -17 419
rect 17 -357 23 419
rect -23 -369 23 -357
rect 135 419 181 431
rect 135 -357 141 419
rect 175 -357 181 419
rect 135 -369 181 -357
rect 293 419 339 431
rect 293 -357 299 419
rect 333 -357 339 419
rect 293 -369 339 -357
rect -283 -407 -191 -401
rect -283 -441 -271 -407
rect -203 -441 -191 -407
rect -283 -447 -191 -441
rect -125 -407 -33 -401
rect -125 -441 -113 -407
rect -45 -441 -33 -407
rect -125 -447 -33 -441
rect 33 -407 125 -401
rect 33 -441 45 -407
rect 113 -441 125 -407
rect 33 -447 125 -441
rect 191 -407 283 -401
rect 191 -441 203 -407
rect 271 -441 283 -407
rect 191 -447 283 -441
<< properties >>
string FIXED_BBOX -450 -562 450 562
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 4 l 0.5 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
