magic
tech sky130A
magscale 1 2
timestamp 1713585847
<< error_p >>
rect -187 272 -129 278
rect -29 272 29 278
rect 129 272 187 278
rect -187 238 -175 272
rect -29 238 -17 272
rect 129 238 141 272
rect -187 232 -129 238
rect -29 232 29 238
rect 129 232 187 238
rect -187 -238 -129 -232
rect -29 -238 29 -232
rect 129 -238 187 -232
rect -187 -272 -175 -238
rect -29 -272 -17 -238
rect 129 -272 141 -238
rect -187 -278 -129 -272
rect -29 -278 29 -272
rect 129 -278 187 -272
<< pwell >>
rect -436 -458 436 458
<< mvnmos >>
rect -208 -200 -108 200
rect -50 -200 50 200
rect 108 -200 208 200
<< mvndiff >>
rect -266 188 -208 200
rect -266 -188 -254 188
rect -220 -188 -208 188
rect -266 -200 -208 -188
rect -108 188 -50 200
rect -108 -188 -96 188
rect -62 -188 -50 188
rect -108 -200 -50 -188
rect 50 188 108 200
rect 50 -188 62 188
rect 96 -188 108 188
rect 50 -200 108 -188
rect 208 188 266 200
rect 208 -188 220 188
rect 254 -188 266 188
rect 208 -200 266 -188
<< mvndiffc >>
rect -254 -188 -220 188
rect -96 -188 -62 188
rect 62 -188 96 188
rect 220 -188 254 188
<< mvpsubdiff >>
rect -400 410 400 422
rect -400 376 -292 410
rect 292 376 400 410
rect -400 364 400 376
rect -400 314 -342 364
rect -400 -314 -388 314
rect -354 -314 -342 314
rect 342 314 400 364
rect -400 -364 -342 -314
rect 342 -314 354 314
rect 388 -314 400 314
rect 342 -364 400 -314
rect -400 -376 400 -364
rect -400 -410 -292 -376
rect 292 -410 400 -376
rect -400 -422 400 -410
<< mvpsubdiffcont >>
rect -292 376 292 410
rect -388 -314 -354 314
rect 354 -314 388 314
rect -292 -410 292 -376
<< poly >>
rect -208 272 -108 288
rect -208 238 -192 272
rect -124 238 -108 272
rect -208 200 -108 238
rect -50 272 50 288
rect -50 238 -34 272
rect 34 238 50 272
rect -50 200 50 238
rect 108 272 208 288
rect 108 238 124 272
rect 192 238 208 272
rect 108 200 208 238
rect -208 -238 -108 -200
rect -208 -272 -192 -238
rect -124 -272 -108 -238
rect -208 -288 -108 -272
rect -50 -238 50 -200
rect -50 -272 -34 -238
rect 34 -272 50 -238
rect -50 -288 50 -272
rect 108 -238 208 -200
rect 108 -272 124 -238
rect 192 -272 208 -238
rect 108 -288 208 -272
<< polycont >>
rect -192 238 -124 272
rect -34 238 34 272
rect 124 238 192 272
rect -192 -272 -124 -238
rect -34 -272 34 -238
rect 124 -272 192 -238
<< locali >>
rect -388 376 -292 410
rect 292 376 388 410
rect -388 314 -354 376
rect 354 314 388 376
rect -208 238 -192 272
rect -124 238 -108 272
rect -50 238 -34 272
rect 34 238 50 272
rect 108 238 124 272
rect 192 238 208 272
rect -254 188 -220 204
rect -254 -204 -220 -188
rect -96 188 -62 204
rect -96 -204 -62 -188
rect 62 188 96 204
rect 62 -204 96 -188
rect 220 188 254 204
rect 220 -204 254 -188
rect -208 -272 -192 -238
rect -124 -272 -108 -238
rect -50 -272 -34 -238
rect 34 -272 50 -238
rect 108 -272 124 -238
rect 192 -272 208 -238
rect -388 -376 -354 -314
rect 354 -376 388 -314
rect -388 -410 -292 -376
rect 292 -410 388 -376
<< viali >>
rect -283 376 283 410
rect -388 -301 -354 301
rect -175 238 -141 272
rect -17 238 17 272
rect 141 238 175 272
rect -254 -188 -220 188
rect -96 -188 -62 188
rect 62 -188 96 188
rect 220 -188 254 188
rect -175 -272 -141 -238
rect -17 -272 17 -238
rect 141 -272 175 -238
rect 354 -301 388 301
<< metal1 >>
rect -295 410 295 416
rect -295 376 -283 410
rect 283 376 295 410
rect -295 370 295 376
rect -394 301 -348 313
rect -394 -301 -388 301
rect -354 -301 -348 301
rect 348 301 394 313
rect -187 272 -129 278
rect -187 238 -175 272
rect -141 238 -129 272
rect -187 232 -129 238
rect -29 272 29 278
rect -29 238 -17 272
rect 17 238 29 272
rect -29 232 29 238
rect 129 272 187 278
rect 129 238 141 272
rect 175 238 187 272
rect 129 232 187 238
rect -260 188 -214 200
rect -260 -188 -254 188
rect -220 -188 -214 188
rect -260 -200 -214 -188
rect -102 188 -56 200
rect -102 -188 -96 188
rect -62 -188 -56 188
rect -102 -200 -56 -188
rect 56 188 102 200
rect 56 -188 62 188
rect 96 -188 102 188
rect 56 -200 102 -188
rect 214 188 260 200
rect 214 -188 220 188
rect 254 -188 260 188
rect 214 -200 260 -188
rect -187 -238 -129 -232
rect -187 -272 -175 -238
rect -141 -272 -129 -238
rect -187 -278 -129 -272
rect -29 -238 29 -232
rect -29 -272 -17 -238
rect 17 -272 29 -238
rect -29 -278 29 -272
rect 129 -238 187 -232
rect 129 -272 141 -238
rect 175 -272 187 -238
rect 129 -278 187 -272
rect -394 -313 -348 -301
rect 348 -301 354 301
rect 388 -301 394 301
rect 348 -313 394 -301
<< properties >>
string FIXED_BBOX -371 -393 371 393
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 2 l 0.50 m 1 nf 3 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 80 viagl 80 viagt 80
<< end >>
