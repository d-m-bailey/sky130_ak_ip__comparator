magic
tech sky130A
magscale 1 2
timestamp 1713551257
<< error_p >>
rect -111 281 -47 287
rect 47 281 111 287
rect -111 247 -99 281
rect 47 247 59 281
rect -111 241 -47 247
rect 47 241 111 247
rect -111 -247 -47 -241
rect 47 -247 111 -241
rect -111 -281 -99 -247
rect 47 -281 59 -247
rect -111 -287 -47 -281
rect 47 -287 111 -281
<< nwell >>
rect -387 -497 387 497
<< mvpmos >>
rect -129 -200 -29 200
rect 29 -200 129 200
<< mvpdiff >>
rect -187 188 -129 200
rect -187 -188 -175 188
rect -141 -188 -129 188
rect -187 -200 -129 -188
rect -29 188 29 200
rect -29 -188 -17 188
rect 17 -188 29 188
rect -29 -200 29 -188
rect 129 188 187 200
rect 129 -188 141 188
rect 175 -188 187 188
rect 129 -200 187 -188
<< mvpdiffc >>
rect -175 -188 -141 188
rect -17 -188 17 188
rect 141 -188 175 188
<< mvnsubdiff >>
rect -321 419 321 431
rect -321 385 -213 419
rect 213 385 321 419
rect -321 373 321 385
rect -321 -373 -263 373
rect 263 -373 321 373
rect -321 -385 321 -373
rect -321 -419 -213 -385
rect 213 -419 321 -385
rect -321 -431 321 -419
<< mvnsubdiffcont >>
rect -213 385 213 419
rect -213 -419 213 -385
<< poly >>
rect -129 281 -29 297
rect -129 247 -113 281
rect -45 247 -29 281
rect -129 200 -29 247
rect 29 281 129 297
rect 29 247 45 281
rect 113 247 129 281
rect 29 200 129 247
rect -129 -247 -29 -200
rect -129 -281 -113 -247
rect -45 -281 -29 -247
rect -129 -297 -29 -281
rect 29 -247 129 -200
rect 29 -281 45 -247
rect 113 -281 129 -247
rect 29 -297 129 -281
<< polycont >>
rect -113 247 -45 281
rect 45 247 113 281
rect -113 -281 -45 -247
rect 45 -281 113 -247
<< locali >>
rect -309 385 -220 419
rect 220 385 309 419
rect -309 308 -275 385
rect 275 308 309 385
rect -129 247 -113 281
rect -45 247 -29 281
rect 29 247 45 281
rect 113 247 129 281
rect -175 188 -141 204
rect -175 -204 -141 -188
rect -17 188 17 204
rect -17 -204 17 -188
rect 141 188 175 204
rect 141 -204 175 -188
rect -129 -281 -113 -247
rect -45 -281 -29 -247
rect 29 -281 45 -247
rect 113 -281 129 -247
rect -309 -385 -275 -308
rect 275 -385 309 -308
rect -309 -419 -213 -385
rect 213 -419 309 -385
<< viali >>
rect -220 385 -213 419
rect -213 385 213 419
rect 213 385 220 419
rect -309 -308 -275 308
rect -99 247 -59 281
rect 59 247 99 281
rect -175 -188 -141 188
rect -17 -188 17 188
rect 141 -188 175 188
rect -99 -281 -59 -247
rect 59 -281 99 -247
rect 275 -308 309 308
<< metal1 >>
rect -232 419 232 425
rect -232 385 -220 419
rect 220 385 232 419
rect -232 379 232 385
rect -315 308 -269 320
rect -315 -308 -309 308
rect -275 -308 -269 308
rect 269 308 315 320
rect -111 281 -47 287
rect -111 247 -99 281
rect -59 247 -47 281
rect -111 241 -47 247
rect 47 281 111 287
rect 47 247 59 281
rect 99 247 111 281
rect 47 241 111 247
rect -181 188 -135 200
rect -181 -188 -175 188
rect -141 -188 -135 188
rect -181 -200 -135 -188
rect -23 188 23 200
rect -23 -188 -17 188
rect 17 -188 23 188
rect -23 -200 23 -188
rect 135 188 181 200
rect 135 -188 141 188
rect 175 -188 181 188
rect 135 -200 181 -188
rect -111 -247 -47 -241
rect -111 -281 -99 -247
rect -59 -281 -47 -247
rect -111 -287 -47 -281
rect 47 -247 111 -241
rect 47 -281 59 -247
rect 99 -281 111 -247
rect 47 -287 111 -281
rect -315 -320 -269 -308
rect 269 -308 275 308
rect 309 -308 315 308
rect 269 -320 315 -308
<< properties >>
string FIXED_BBOX -292 -402 292 402
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 2 l 0.50 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 0 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 60 viagb 0 viagr 80 viagl 80 viagt 80
<< end >>
