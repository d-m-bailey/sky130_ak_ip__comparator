magic
tech sky130A
magscale 1 2
timestamp 1713227719
<< nwell >>
rect -2374 -497 2374 497
<< mvpmos >>
rect -2116 -200 -1316 200
rect -1258 -200 -458 200
rect -400 -200 400 200
rect 458 -200 1258 200
rect 1316 -200 2116 200
<< mvpdiff >>
rect -2174 188 -2116 200
rect -2174 -188 -2162 188
rect -2128 -188 -2116 188
rect -2174 -200 -2116 -188
rect -1316 188 -1258 200
rect -1316 -188 -1304 188
rect -1270 -188 -1258 188
rect -1316 -200 -1258 -188
rect -458 188 -400 200
rect -458 -188 -446 188
rect -412 -188 -400 188
rect -458 -200 -400 -188
rect 400 188 458 200
rect 400 -188 412 188
rect 446 -188 458 188
rect 400 -200 458 -188
rect 1258 188 1316 200
rect 1258 -188 1270 188
rect 1304 -188 1316 188
rect 1258 -200 1316 -188
rect 2116 188 2174 200
rect 2116 -188 2128 188
rect 2162 -188 2174 188
rect 2116 -200 2174 -188
<< mvpdiffc >>
rect -2162 -188 -2128 188
rect -1304 -188 -1270 188
rect -446 -188 -412 188
rect 412 -188 446 188
rect 1270 -188 1304 188
rect 2128 -188 2162 188
<< mvnsubdiff >>
rect -2308 419 2308 431
rect -2308 385 -2200 419
rect 2200 385 2308 419
rect -2308 373 2308 385
rect -2308 323 -2250 373
rect -2308 -323 -2296 323
rect -2262 -323 -2250 323
rect 2250 323 2308 373
rect -2308 -373 -2250 -323
rect 2250 -323 2262 323
rect 2296 -323 2308 323
rect 2250 -373 2308 -323
rect -2308 -385 2308 -373
rect -2308 -419 -2200 -385
rect 2200 -419 2308 -385
rect -2308 -431 2308 -419
<< mvnsubdiffcont >>
rect -2200 385 2200 419
rect -2296 -323 -2262 323
rect 2262 -323 2296 323
rect -2200 -419 2200 -385
<< poly >>
rect -2116 281 -1316 297
rect -2116 247 -2100 281
rect -1332 247 -1316 281
rect -2116 200 -1316 247
rect -1258 281 -458 297
rect -1258 247 -1242 281
rect -474 247 -458 281
rect -1258 200 -458 247
rect -400 281 400 297
rect -400 247 -384 281
rect 384 247 400 281
rect -400 200 400 247
rect 458 281 1258 297
rect 458 247 474 281
rect 1242 247 1258 281
rect 458 200 1258 247
rect 1316 281 2116 297
rect 1316 247 1332 281
rect 2100 247 2116 281
rect 1316 200 2116 247
rect -2116 -247 -1316 -200
rect -2116 -281 -2100 -247
rect -1332 -281 -1316 -247
rect -2116 -297 -1316 -281
rect -1258 -247 -458 -200
rect -1258 -281 -1242 -247
rect -474 -281 -458 -247
rect -1258 -297 -458 -281
rect -400 -247 400 -200
rect -400 -281 -384 -247
rect 384 -281 400 -247
rect -400 -297 400 -281
rect 458 -247 1258 -200
rect 458 -281 474 -247
rect 1242 -281 1258 -247
rect 458 -297 1258 -281
rect 1316 -247 2116 -200
rect 1316 -281 1332 -247
rect 2100 -281 2116 -247
rect 1316 -297 2116 -281
<< polycont >>
rect -2100 247 -1332 281
rect -1242 247 -474 281
rect -384 247 384 281
rect 474 247 1242 281
rect 1332 247 2100 281
rect -2100 -281 -1332 -247
rect -1242 -281 -474 -247
rect -384 -281 384 -247
rect 474 -281 1242 -247
rect 1332 -281 2100 -247
<< locali >>
rect -2296 385 -2200 419
rect 2200 385 2296 419
rect -2296 323 -2262 385
rect 2262 323 2296 385
rect -2116 247 -2100 281
rect -1332 247 -1316 281
rect -1258 247 -1242 281
rect -474 247 -458 281
rect -400 247 -384 281
rect 384 247 400 281
rect 458 247 474 281
rect 1242 247 1258 281
rect 1316 247 1332 281
rect 2100 247 2116 281
rect -2162 188 -2128 204
rect -2162 -204 -2128 -188
rect -1304 188 -1270 204
rect -1304 -204 -1270 -188
rect -446 188 -412 204
rect -446 -204 -412 -188
rect 412 188 446 204
rect 412 -204 446 -188
rect 1270 188 1304 204
rect 1270 -204 1304 -188
rect 2128 188 2162 204
rect 2128 -204 2162 -188
rect -2116 -281 -2100 -247
rect -1332 -281 -1316 -247
rect -1258 -281 -1242 -247
rect -474 -281 -458 -247
rect -400 -281 -384 -247
rect 384 -281 400 -247
rect 458 -281 474 -247
rect 1242 -281 1258 -247
rect 1316 -281 1332 -247
rect 2100 -281 2116 -247
rect -2296 -385 -2262 -323
rect 2262 -385 2296 -323
rect -2296 -419 -2200 -385
rect 2200 -419 2296 -385
<< viali >>
rect -2100 247 -1332 281
rect -1242 247 -474 281
rect -384 247 384 281
rect 474 247 1242 281
rect 1332 247 2100 281
rect -2162 -188 -2128 188
rect -1304 -188 -1270 188
rect -446 -188 -412 188
rect 412 -188 446 188
rect 1270 -188 1304 188
rect 2128 -188 2162 188
rect -2100 -281 -1332 -247
rect -1242 -281 -474 -247
rect -384 -281 384 -247
rect 474 -281 1242 -247
rect 1332 -281 2100 -247
<< metal1 >>
rect -2112 281 -1320 287
rect -2112 247 -2100 281
rect -1332 247 -1320 281
rect -2112 241 -1320 247
rect -1254 281 -462 287
rect -1254 247 -1242 281
rect -474 247 -462 281
rect -1254 241 -462 247
rect -396 281 396 287
rect -396 247 -384 281
rect 384 247 396 281
rect -396 241 396 247
rect 462 281 1254 287
rect 462 247 474 281
rect 1242 247 1254 281
rect 462 241 1254 247
rect 1320 281 2112 287
rect 1320 247 1332 281
rect 2100 247 2112 281
rect 1320 241 2112 247
rect -2168 188 -2122 200
rect -2168 -188 -2162 188
rect -2128 -188 -2122 188
rect -2168 -200 -2122 -188
rect -1310 188 -1264 200
rect -1310 -188 -1304 188
rect -1270 -188 -1264 188
rect -1310 -200 -1264 -188
rect -452 188 -406 200
rect -452 -188 -446 188
rect -412 -188 -406 188
rect -452 -200 -406 -188
rect 406 188 452 200
rect 406 -188 412 188
rect 446 -188 452 188
rect 406 -200 452 -188
rect 1264 188 1310 200
rect 1264 -188 1270 188
rect 1304 -188 1310 188
rect 1264 -200 1310 -188
rect 2122 188 2168 200
rect 2122 -188 2128 188
rect 2162 -188 2168 188
rect 2122 -200 2168 -188
rect -2112 -247 -1320 -241
rect -2112 -281 -2100 -247
rect -1332 -281 -1320 -247
rect -2112 -287 -1320 -281
rect -1254 -247 -462 -241
rect -1254 -281 -1242 -247
rect -474 -281 -462 -247
rect -1254 -287 -462 -281
rect -396 -247 396 -241
rect -396 -281 -384 -247
rect 384 -281 396 -247
rect -396 -287 396 -281
rect 462 -247 1254 -241
rect 462 -281 474 -247
rect 1242 -281 1254 -247
rect 462 -287 1254 -281
rect 1320 -247 2112 -241
rect 1320 -281 1332 -247
rect 2100 -281 2112 -247
rect 1320 -287 2112 -281
<< properties >>
string FIXED_BBOX -2279 -402 2279 402
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 2 l 4 m 1 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
