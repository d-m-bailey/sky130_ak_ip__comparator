magic
tech sky130A
magscale 1 2
timestamp 1713585847
<< pwell >>
rect -1231 -458 1231 458
<< mvnmos >>
rect -1003 -200 -803 200
rect -745 -200 -545 200
rect -487 -200 -287 200
rect -229 -200 -29 200
rect 29 -200 229 200
rect 287 -200 487 200
rect 545 -200 745 200
rect 803 -200 1003 200
<< mvndiff >>
rect -1061 188 -1003 200
rect -1061 -188 -1049 188
rect -1015 -188 -1003 188
rect -1061 -200 -1003 -188
rect -803 188 -745 200
rect -803 -188 -791 188
rect -757 -188 -745 188
rect -803 -200 -745 -188
rect -545 188 -487 200
rect -545 -188 -533 188
rect -499 -188 -487 188
rect -545 -200 -487 -188
rect -287 188 -229 200
rect -287 -188 -275 188
rect -241 -188 -229 188
rect -287 -200 -229 -188
rect -29 188 29 200
rect -29 -188 -17 188
rect 17 -188 29 188
rect -29 -200 29 -188
rect 229 188 287 200
rect 229 -188 241 188
rect 275 -188 287 188
rect 229 -200 287 -188
rect 487 188 545 200
rect 487 -188 499 188
rect 533 -188 545 188
rect 487 -200 545 -188
rect 745 188 803 200
rect 745 -188 757 188
rect 791 -188 803 188
rect 745 -200 803 -188
rect 1003 188 1061 200
rect 1003 -188 1015 188
rect 1049 -188 1061 188
rect 1003 -200 1061 -188
<< mvndiffc >>
rect -1049 -188 -1015 188
rect -791 -188 -757 188
rect -533 -188 -499 188
rect -275 -188 -241 188
rect -17 -188 17 188
rect 241 -188 275 188
rect 499 -188 533 188
rect 757 -188 791 188
rect 1015 -188 1049 188
<< mvpsubdiff >>
rect -1195 410 1195 422
rect -1195 376 -1087 410
rect 1087 376 1195 410
rect -1195 364 1195 376
rect -1195 314 -1137 364
rect -1195 -314 -1183 314
rect -1149 -314 -1137 314
rect 1137 314 1195 364
rect -1195 -364 -1137 -314
rect 1137 -314 1149 314
rect 1183 -314 1195 314
rect 1137 -364 1195 -314
rect -1195 -376 1195 -364
rect -1195 -410 -1087 -376
rect 1087 -410 1195 -376
rect -1195 -422 1195 -410
<< mvpsubdiffcont >>
rect -1087 376 1087 410
rect -1183 -314 -1149 314
rect 1149 -314 1183 314
rect -1087 -410 1087 -376
<< poly >>
rect -1003 272 -803 288
rect -1003 238 -987 272
rect -819 238 -803 272
rect -1003 200 -803 238
rect -745 272 -545 288
rect -745 238 -729 272
rect -561 238 -545 272
rect -745 200 -545 238
rect -487 272 -287 288
rect -487 238 -471 272
rect -303 238 -287 272
rect -487 200 -287 238
rect -229 272 -29 288
rect -229 238 -213 272
rect -45 238 -29 272
rect -229 200 -29 238
rect 29 272 229 288
rect 29 238 45 272
rect 213 238 229 272
rect 29 200 229 238
rect 287 272 487 288
rect 287 238 303 272
rect 471 238 487 272
rect 287 200 487 238
rect 545 272 745 288
rect 545 238 561 272
rect 729 238 745 272
rect 545 200 745 238
rect 803 272 1003 288
rect 803 238 819 272
rect 987 238 1003 272
rect 803 200 1003 238
rect -1003 -238 -803 -200
rect -1003 -272 -987 -238
rect -819 -272 -803 -238
rect -1003 -288 -803 -272
rect -745 -238 -545 -200
rect -745 -272 -729 -238
rect -561 -272 -545 -238
rect -745 -288 -545 -272
rect -487 -238 -287 -200
rect -487 -272 -471 -238
rect -303 -272 -287 -238
rect -487 -288 -287 -272
rect -229 -238 -29 -200
rect -229 -272 -213 -238
rect -45 -272 -29 -238
rect -229 -288 -29 -272
rect 29 -238 229 -200
rect 29 -272 45 -238
rect 213 -272 229 -238
rect 29 -288 229 -272
rect 287 -238 487 -200
rect 287 -272 303 -238
rect 471 -272 487 -238
rect 287 -288 487 -272
rect 545 -238 745 -200
rect 545 -272 561 -238
rect 729 -272 745 -238
rect 545 -288 745 -272
rect 803 -238 1003 -200
rect 803 -272 819 -238
rect 987 -272 1003 -238
rect 803 -288 1003 -272
<< polycont >>
rect -987 238 -819 272
rect -729 238 -561 272
rect -471 238 -303 272
rect -213 238 -45 272
rect 45 238 213 272
rect 303 238 471 272
rect 561 238 729 272
rect 819 238 987 272
rect -987 -272 -819 -238
rect -729 -272 -561 -238
rect -471 -272 -303 -238
rect -213 -272 -45 -238
rect 45 -272 213 -238
rect 303 -272 471 -238
rect 561 -272 729 -238
rect 819 -272 987 -238
<< locali >>
rect -1183 376 -1087 410
rect 1087 376 1183 410
rect -1183 314 -1149 376
rect 1149 314 1183 376
rect -1003 238 -987 272
rect -819 238 -803 272
rect -745 238 -729 272
rect -561 238 -545 272
rect -487 238 -471 272
rect -303 238 -287 272
rect -229 238 -213 272
rect -45 238 -29 272
rect 29 238 45 272
rect 213 238 229 272
rect 287 238 303 272
rect 471 238 487 272
rect 545 238 561 272
rect 729 238 745 272
rect 803 238 819 272
rect 987 238 1003 272
rect -1049 188 -1015 204
rect -1049 -204 -1015 -188
rect -791 188 -757 204
rect -791 -204 -757 -188
rect -533 188 -499 204
rect -533 -204 -499 -188
rect -275 188 -241 204
rect -275 -204 -241 -188
rect -17 188 17 204
rect -17 -204 17 -188
rect 241 188 275 204
rect 241 -204 275 -188
rect 499 188 533 204
rect 499 -204 533 -188
rect 757 188 791 204
rect 757 -204 791 -188
rect 1015 188 1049 204
rect 1015 -204 1049 -188
rect -1003 -272 -987 -238
rect -819 -272 -803 -238
rect -745 -272 -729 -238
rect -561 -272 -545 -238
rect -487 -272 -471 -238
rect -303 -272 -287 -238
rect -229 -272 -213 -238
rect -45 -272 -29 -238
rect 29 -272 45 -238
rect 213 -272 229 -238
rect 287 -272 303 -238
rect 471 -272 487 -238
rect 545 -272 561 -238
rect 729 -272 745 -238
rect 803 -272 819 -238
rect 987 -272 1003 -238
rect -1183 -376 -1149 -314
rect 1149 -376 1183 -314
rect -1183 -410 -1087 -376
rect 1087 -410 1183 -376
<< viali >>
rect -970 238 -836 272
rect -712 238 -578 272
rect -454 238 -320 272
rect -196 238 -62 272
rect 62 238 196 272
rect 320 238 454 272
rect 578 238 712 272
rect 836 238 970 272
rect -1049 -188 -1015 188
rect -791 -188 -757 188
rect -533 -188 -499 188
rect -275 -188 -241 188
rect -17 -188 17 188
rect 241 -188 275 188
rect 499 -188 533 188
rect 757 -188 791 188
rect 1015 -188 1049 188
rect -970 -272 -836 -238
rect -712 -272 -578 -238
rect -454 -272 -320 -238
rect -196 -272 -62 -238
rect 62 -272 196 -238
rect 320 -272 454 -238
rect 578 -272 712 -238
rect 836 -272 970 -238
<< metal1 >>
rect -982 272 -824 278
rect -982 238 -970 272
rect -836 238 -824 272
rect -982 232 -824 238
rect -724 272 -566 278
rect -724 238 -712 272
rect -578 238 -566 272
rect -724 232 -566 238
rect -466 272 -308 278
rect -466 238 -454 272
rect -320 238 -308 272
rect -466 232 -308 238
rect -208 272 -50 278
rect -208 238 -196 272
rect -62 238 -50 272
rect -208 232 -50 238
rect 50 272 208 278
rect 50 238 62 272
rect 196 238 208 272
rect 50 232 208 238
rect 308 272 466 278
rect 308 238 320 272
rect 454 238 466 272
rect 308 232 466 238
rect 566 272 724 278
rect 566 238 578 272
rect 712 238 724 272
rect 566 232 724 238
rect 824 272 982 278
rect 824 238 836 272
rect 970 238 982 272
rect 824 232 982 238
rect -1055 188 -1009 200
rect -1055 -188 -1049 188
rect -1015 -188 -1009 188
rect -1055 -200 -1009 -188
rect -797 188 -751 200
rect -797 -188 -791 188
rect -757 -188 -751 188
rect -797 -200 -751 -188
rect -539 188 -493 200
rect -539 -188 -533 188
rect -499 -188 -493 188
rect -539 -200 -493 -188
rect -281 188 -235 200
rect -281 -188 -275 188
rect -241 -188 -235 188
rect -281 -200 -235 -188
rect -23 188 23 200
rect -23 -188 -17 188
rect 17 -188 23 188
rect -23 -200 23 -188
rect 235 188 281 200
rect 235 -188 241 188
rect 275 -188 281 188
rect 235 -200 281 -188
rect 493 188 539 200
rect 493 -188 499 188
rect 533 -188 539 188
rect 493 -200 539 -188
rect 751 188 797 200
rect 751 -188 757 188
rect 791 -188 797 188
rect 751 -200 797 -188
rect 1009 188 1055 200
rect 1009 -188 1015 188
rect 1049 -188 1055 188
rect 1009 -200 1055 -188
rect -982 -238 -824 -232
rect -982 -272 -970 -238
rect -836 -272 -824 -238
rect -982 -278 -824 -272
rect -724 -238 -566 -232
rect -724 -272 -712 -238
rect -578 -272 -566 -238
rect -724 -278 -566 -272
rect -466 -238 -308 -232
rect -466 -272 -454 -238
rect -320 -272 -308 -238
rect -466 -278 -308 -272
rect -208 -238 -50 -232
rect -208 -272 -196 -238
rect -62 -272 -50 -238
rect -208 -278 -50 -272
rect 50 -238 208 -232
rect 50 -272 62 -238
rect 196 -272 208 -238
rect 50 -278 208 -272
rect 308 -238 466 -232
rect 308 -272 320 -238
rect 454 -272 466 -238
rect 308 -278 466 -272
rect 566 -238 724 -232
rect 566 -272 578 -238
rect 712 -272 724 -238
rect 566 -278 724 -272
rect 824 -238 982 -232
rect 824 -272 836 -238
rect 970 -272 982 -238
rect 824 -278 982 -272
<< properties >>
string FIXED_BBOX -1166 -393 1166 393
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 2 l 1 m 1 nf 8 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 80 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
