magic
tech sky130A
magscale 1 2
timestamp 1713214796
<< nwell >>
rect -458 -347 458 347
<< mvpmos >>
rect -200 -50 200 50
<< mvpdiff >>
rect -258 38 -200 50
rect -258 -38 -246 38
rect -212 -38 -200 38
rect -258 -50 -200 -38
rect 200 38 258 50
rect 200 -38 212 38
rect 246 -38 258 38
rect 200 -50 258 -38
<< mvpdiffc >>
rect -246 -38 -212 38
rect 212 -38 246 38
<< mvnsubdiff >>
rect -392 269 392 281
rect -392 235 -284 269
rect 284 235 392 269
rect -392 223 392 235
rect -392 173 -334 223
rect -392 -173 -380 173
rect -346 -173 -334 173
rect 334 173 392 223
rect -392 -223 -334 -173
rect 334 -173 346 173
rect 380 -173 392 173
rect 334 -223 392 -173
rect -392 -235 392 -223
rect -392 -269 -284 -235
rect 284 -269 392 -235
rect -392 -281 392 -269
<< mvnsubdiffcont >>
rect -284 235 284 269
rect -380 -173 -346 173
rect 346 -173 380 173
rect -284 -269 284 -235
<< poly >>
rect -200 131 200 147
rect -200 97 -184 131
rect 184 97 200 131
rect -200 50 200 97
rect -200 -97 200 -50
rect -200 -131 -184 -97
rect 184 -131 200 -97
rect -200 -147 200 -131
<< polycont >>
rect -184 97 184 131
rect -184 -131 184 -97
<< locali >>
rect -380 173 -346 269
rect 346 173 380 269
rect -200 97 -184 131
rect 184 97 200 131
rect -246 38 -212 54
rect -246 -54 -212 -38
rect 212 38 246 54
rect 212 -54 246 -38
rect -200 -131 -184 -97
rect 184 -131 200 -97
rect -380 -235 -346 -173
rect 346 -235 380 -173
rect -380 -269 -284 -235
rect 284 -269 380 -235
<< viali >>
rect -346 235 -284 269
rect -284 235 284 269
rect 284 235 346 269
rect -110 97 110 131
rect -246 -38 -212 38
rect 212 -38 246 38
rect -110 -131 110 -97
<< metal1 >>
rect -358 269 358 275
rect -358 235 -346 269
rect 346 235 358 269
rect -358 229 358 235
rect -122 131 122 137
rect -122 97 -110 131
rect 110 97 122 131
rect -122 91 122 97
rect -252 38 -206 50
rect -252 -38 -246 38
rect -212 -38 -206 38
rect -252 -50 -206 -38
rect 206 38 252 50
rect 206 -38 212 38
rect 246 -38 252 38
rect 206 -50 252 -38
rect -122 -97 122 -91
rect -122 -131 -110 -97
rect 110 -131 122 -97
rect -122 -137 122 -131
<< properties >>
string FIXED_BBOX -363 -252 363 252
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 0.5 l 2 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 60 viagb 0 viagr 0 viagl 0 viagt 100
<< end >>
