magic
tech sky130A
magscale 1 2
timestamp 1713067540
<< pwell >>
rect -515 -3203 515 3203
<< mvnmos >>
rect -287 2145 -187 2945
rect -129 2145 -29 2945
rect 29 2145 129 2945
rect 187 2145 287 2945
rect -287 1127 -187 1927
rect -129 1127 -29 1927
rect 29 1127 129 1927
rect 187 1127 287 1927
rect -287 109 -187 909
rect -129 109 -29 909
rect 29 109 129 909
rect 187 109 287 909
rect -287 -909 -187 -109
rect -129 -909 -29 -109
rect 29 -909 129 -109
rect 187 -909 287 -109
rect -287 -1927 -187 -1127
rect -129 -1927 -29 -1127
rect 29 -1927 129 -1127
rect 187 -1927 287 -1127
rect -287 -2945 -187 -2145
rect -129 -2945 -29 -2145
rect 29 -2945 129 -2145
rect 187 -2945 287 -2145
<< mvndiff >>
rect -345 2933 -287 2945
rect -345 2157 -333 2933
rect -299 2157 -287 2933
rect -345 2145 -287 2157
rect -187 2933 -129 2945
rect -187 2157 -175 2933
rect -141 2157 -129 2933
rect -187 2145 -129 2157
rect -29 2933 29 2945
rect -29 2157 -17 2933
rect 17 2157 29 2933
rect -29 2145 29 2157
rect 129 2933 187 2945
rect 129 2157 141 2933
rect 175 2157 187 2933
rect 129 2145 187 2157
rect 287 2933 345 2945
rect 287 2157 299 2933
rect 333 2157 345 2933
rect 287 2145 345 2157
rect -345 1915 -287 1927
rect -345 1139 -333 1915
rect -299 1139 -287 1915
rect -345 1127 -287 1139
rect -187 1915 -129 1927
rect -187 1139 -175 1915
rect -141 1139 -129 1915
rect -187 1127 -129 1139
rect -29 1915 29 1927
rect -29 1139 -17 1915
rect 17 1139 29 1915
rect -29 1127 29 1139
rect 129 1915 187 1927
rect 129 1139 141 1915
rect 175 1139 187 1915
rect 129 1127 187 1139
rect 287 1915 345 1927
rect 287 1139 299 1915
rect 333 1139 345 1915
rect 287 1127 345 1139
rect -345 897 -287 909
rect -345 121 -333 897
rect -299 121 -287 897
rect -345 109 -287 121
rect -187 897 -129 909
rect -187 121 -175 897
rect -141 121 -129 897
rect -187 109 -129 121
rect -29 897 29 909
rect -29 121 -17 897
rect 17 121 29 897
rect -29 109 29 121
rect 129 897 187 909
rect 129 121 141 897
rect 175 121 187 897
rect 129 109 187 121
rect 287 897 345 909
rect 287 121 299 897
rect 333 121 345 897
rect 287 109 345 121
rect -345 -121 -287 -109
rect -345 -897 -333 -121
rect -299 -897 -287 -121
rect -345 -909 -287 -897
rect -187 -121 -129 -109
rect -187 -897 -175 -121
rect -141 -897 -129 -121
rect -187 -909 -129 -897
rect -29 -121 29 -109
rect -29 -897 -17 -121
rect 17 -897 29 -121
rect -29 -909 29 -897
rect 129 -121 187 -109
rect 129 -897 141 -121
rect 175 -897 187 -121
rect 129 -909 187 -897
rect 287 -121 345 -109
rect 287 -897 299 -121
rect 333 -897 345 -121
rect 287 -909 345 -897
rect -345 -1139 -287 -1127
rect -345 -1915 -333 -1139
rect -299 -1915 -287 -1139
rect -345 -1927 -287 -1915
rect -187 -1139 -129 -1127
rect -187 -1915 -175 -1139
rect -141 -1915 -129 -1139
rect -187 -1927 -129 -1915
rect -29 -1139 29 -1127
rect -29 -1915 -17 -1139
rect 17 -1915 29 -1139
rect -29 -1927 29 -1915
rect 129 -1139 187 -1127
rect 129 -1915 141 -1139
rect 175 -1915 187 -1139
rect 129 -1927 187 -1915
rect 287 -1139 345 -1127
rect 287 -1915 299 -1139
rect 333 -1915 345 -1139
rect 287 -1927 345 -1915
rect -345 -2157 -287 -2145
rect -345 -2933 -333 -2157
rect -299 -2933 -287 -2157
rect -345 -2945 -287 -2933
rect -187 -2157 -129 -2145
rect -187 -2933 -175 -2157
rect -141 -2933 -129 -2157
rect -187 -2945 -129 -2933
rect -29 -2157 29 -2145
rect -29 -2933 -17 -2157
rect 17 -2933 29 -2157
rect -29 -2945 29 -2933
rect 129 -2157 187 -2145
rect 129 -2933 141 -2157
rect 175 -2933 187 -2157
rect 129 -2945 187 -2933
rect 287 -2157 345 -2145
rect 287 -2933 299 -2157
rect 333 -2933 345 -2157
rect 287 -2945 345 -2933
<< mvndiffc >>
rect -333 2157 -299 2933
rect -175 2157 -141 2933
rect -17 2157 17 2933
rect 141 2157 175 2933
rect 299 2157 333 2933
rect -333 1139 -299 1915
rect -175 1139 -141 1915
rect -17 1139 17 1915
rect 141 1139 175 1915
rect 299 1139 333 1915
rect -333 121 -299 897
rect -175 121 -141 897
rect -17 121 17 897
rect 141 121 175 897
rect 299 121 333 897
rect -333 -897 -299 -121
rect -175 -897 -141 -121
rect -17 -897 17 -121
rect 141 -897 175 -121
rect 299 -897 333 -121
rect -333 -1915 -299 -1139
rect -175 -1915 -141 -1139
rect -17 -1915 17 -1139
rect 141 -1915 175 -1139
rect 299 -1915 333 -1139
rect -333 -2933 -299 -2157
rect -175 -2933 -141 -2157
rect -17 -2933 17 -2157
rect 141 -2933 175 -2157
rect 299 -2933 333 -2157
<< mvpsubdiff >>
rect -479 3155 479 3167
rect -479 3121 -371 3155
rect 371 3121 479 3155
rect -479 3109 479 3121
rect -479 3059 -421 3109
rect -479 -3059 -467 3059
rect -433 -3059 -421 3059
rect 421 3059 479 3109
rect -479 -3109 -421 -3059
rect 421 -3059 433 3059
rect 467 -3059 479 3059
rect 421 -3109 479 -3059
rect -479 -3121 479 -3109
rect -479 -3155 -371 -3121
rect 371 -3155 479 -3121
rect -479 -3167 479 -3155
<< mvpsubdiffcont >>
rect -371 3121 371 3155
rect -467 -3059 -433 3059
rect 433 -3059 467 3059
rect -371 -3155 371 -3121
<< poly >>
rect -287 3017 -187 3033
rect -287 2983 -271 3017
rect -203 2983 -187 3017
rect -287 2945 -187 2983
rect -129 3017 -29 3033
rect -129 2983 -113 3017
rect -45 2983 -29 3017
rect -129 2945 -29 2983
rect 29 3017 129 3033
rect 29 2983 45 3017
rect 113 2983 129 3017
rect 29 2945 129 2983
rect 187 3017 287 3033
rect 187 2983 203 3017
rect 271 2983 287 3017
rect 187 2945 287 2983
rect -287 2107 -187 2145
rect -287 2073 -271 2107
rect -203 2073 -187 2107
rect -287 2057 -187 2073
rect -129 2107 -29 2145
rect -129 2073 -113 2107
rect -45 2073 -29 2107
rect -129 2057 -29 2073
rect 29 2107 129 2145
rect 29 2073 45 2107
rect 113 2073 129 2107
rect 29 2057 129 2073
rect 187 2107 287 2145
rect 187 2073 203 2107
rect 271 2073 287 2107
rect 187 2057 287 2073
rect -287 1999 -187 2015
rect -287 1965 -271 1999
rect -203 1965 -187 1999
rect -287 1927 -187 1965
rect -129 1999 -29 2015
rect -129 1965 -113 1999
rect -45 1965 -29 1999
rect -129 1927 -29 1965
rect 29 1999 129 2015
rect 29 1965 45 1999
rect 113 1965 129 1999
rect 29 1927 129 1965
rect 187 1999 287 2015
rect 187 1965 203 1999
rect 271 1965 287 1999
rect 187 1927 287 1965
rect -287 1089 -187 1127
rect -287 1055 -271 1089
rect -203 1055 -187 1089
rect -287 1039 -187 1055
rect -129 1089 -29 1127
rect -129 1055 -113 1089
rect -45 1055 -29 1089
rect -129 1039 -29 1055
rect 29 1089 129 1127
rect 29 1055 45 1089
rect 113 1055 129 1089
rect 29 1039 129 1055
rect 187 1089 287 1127
rect 187 1055 203 1089
rect 271 1055 287 1089
rect 187 1039 287 1055
rect -287 981 -187 997
rect -287 947 -271 981
rect -203 947 -187 981
rect -287 909 -187 947
rect -129 981 -29 997
rect -129 947 -113 981
rect -45 947 -29 981
rect -129 909 -29 947
rect 29 981 129 997
rect 29 947 45 981
rect 113 947 129 981
rect 29 909 129 947
rect 187 981 287 997
rect 187 947 203 981
rect 271 947 287 981
rect 187 909 287 947
rect -287 71 -187 109
rect -287 37 -271 71
rect -203 37 -187 71
rect -287 21 -187 37
rect -129 71 -29 109
rect -129 37 -113 71
rect -45 37 -29 71
rect -129 21 -29 37
rect 29 71 129 109
rect 29 37 45 71
rect 113 37 129 71
rect 29 21 129 37
rect 187 71 287 109
rect 187 37 203 71
rect 271 37 287 71
rect 187 21 287 37
rect -287 -37 -187 -21
rect -287 -71 -271 -37
rect -203 -71 -187 -37
rect -287 -109 -187 -71
rect -129 -37 -29 -21
rect -129 -71 -113 -37
rect -45 -71 -29 -37
rect -129 -109 -29 -71
rect 29 -37 129 -21
rect 29 -71 45 -37
rect 113 -71 129 -37
rect 29 -109 129 -71
rect 187 -37 287 -21
rect 187 -71 203 -37
rect 271 -71 287 -37
rect 187 -109 287 -71
rect -287 -947 -187 -909
rect -287 -981 -271 -947
rect -203 -981 -187 -947
rect -287 -997 -187 -981
rect -129 -947 -29 -909
rect -129 -981 -113 -947
rect -45 -981 -29 -947
rect -129 -997 -29 -981
rect 29 -947 129 -909
rect 29 -981 45 -947
rect 113 -981 129 -947
rect 29 -997 129 -981
rect 187 -947 287 -909
rect 187 -981 203 -947
rect 271 -981 287 -947
rect 187 -997 287 -981
rect -287 -1055 -187 -1039
rect -287 -1089 -271 -1055
rect -203 -1089 -187 -1055
rect -287 -1127 -187 -1089
rect -129 -1055 -29 -1039
rect -129 -1089 -113 -1055
rect -45 -1089 -29 -1055
rect -129 -1127 -29 -1089
rect 29 -1055 129 -1039
rect 29 -1089 45 -1055
rect 113 -1089 129 -1055
rect 29 -1127 129 -1089
rect 187 -1055 287 -1039
rect 187 -1089 203 -1055
rect 271 -1089 287 -1055
rect 187 -1127 287 -1089
rect -287 -1965 -187 -1927
rect -287 -1999 -271 -1965
rect -203 -1999 -187 -1965
rect -287 -2015 -187 -1999
rect -129 -1965 -29 -1927
rect -129 -1999 -113 -1965
rect -45 -1999 -29 -1965
rect -129 -2015 -29 -1999
rect 29 -1965 129 -1927
rect 29 -1999 45 -1965
rect 113 -1999 129 -1965
rect 29 -2015 129 -1999
rect 187 -1965 287 -1927
rect 187 -1999 203 -1965
rect 271 -1999 287 -1965
rect 187 -2015 287 -1999
rect -287 -2073 -187 -2057
rect -287 -2107 -271 -2073
rect -203 -2107 -187 -2073
rect -287 -2145 -187 -2107
rect -129 -2073 -29 -2057
rect -129 -2107 -113 -2073
rect -45 -2107 -29 -2073
rect -129 -2145 -29 -2107
rect 29 -2073 129 -2057
rect 29 -2107 45 -2073
rect 113 -2107 129 -2073
rect 29 -2145 129 -2107
rect 187 -2073 287 -2057
rect 187 -2107 203 -2073
rect 271 -2107 287 -2073
rect 187 -2145 287 -2107
rect -287 -2983 -187 -2945
rect -287 -3017 -271 -2983
rect -203 -3017 -187 -2983
rect -287 -3033 -187 -3017
rect -129 -2983 -29 -2945
rect -129 -3017 -113 -2983
rect -45 -3017 -29 -2983
rect -129 -3033 -29 -3017
rect 29 -2983 129 -2945
rect 29 -3017 45 -2983
rect 113 -3017 129 -2983
rect 29 -3033 129 -3017
rect 187 -2983 287 -2945
rect 187 -3017 203 -2983
rect 271 -3017 287 -2983
rect 187 -3033 287 -3017
<< polycont >>
rect -271 2983 -203 3017
rect -113 2983 -45 3017
rect 45 2983 113 3017
rect 203 2983 271 3017
rect -271 2073 -203 2107
rect -113 2073 -45 2107
rect 45 2073 113 2107
rect 203 2073 271 2107
rect -271 1965 -203 1999
rect -113 1965 -45 1999
rect 45 1965 113 1999
rect 203 1965 271 1999
rect -271 1055 -203 1089
rect -113 1055 -45 1089
rect 45 1055 113 1089
rect 203 1055 271 1089
rect -271 947 -203 981
rect -113 947 -45 981
rect 45 947 113 981
rect 203 947 271 981
rect -271 37 -203 71
rect -113 37 -45 71
rect 45 37 113 71
rect 203 37 271 71
rect -271 -71 -203 -37
rect -113 -71 -45 -37
rect 45 -71 113 -37
rect 203 -71 271 -37
rect -271 -981 -203 -947
rect -113 -981 -45 -947
rect 45 -981 113 -947
rect 203 -981 271 -947
rect -271 -1089 -203 -1055
rect -113 -1089 -45 -1055
rect 45 -1089 113 -1055
rect 203 -1089 271 -1055
rect -271 -1999 -203 -1965
rect -113 -1999 -45 -1965
rect 45 -1999 113 -1965
rect 203 -1999 271 -1965
rect -271 -2107 -203 -2073
rect -113 -2107 -45 -2073
rect 45 -2107 113 -2073
rect 203 -2107 271 -2073
rect -271 -3017 -203 -2983
rect -113 -3017 -45 -2983
rect 45 -3017 113 -2983
rect 203 -3017 271 -2983
<< locali >>
rect -467 3121 -371 3155
rect 371 3121 467 3155
rect -467 3059 -433 3121
rect 433 3059 467 3121
rect -287 2983 -271 3017
rect -203 2983 -187 3017
rect -129 2983 -113 3017
rect -45 2983 -29 3017
rect 29 2983 45 3017
rect 113 2983 129 3017
rect 187 2983 203 3017
rect 271 2983 287 3017
rect -333 2933 -299 2949
rect -333 2141 -299 2157
rect -175 2933 -141 2949
rect -175 2141 -141 2157
rect -17 2933 17 2949
rect -17 2141 17 2157
rect 141 2933 175 2949
rect 141 2141 175 2157
rect 299 2933 333 2949
rect 299 2141 333 2157
rect -287 2073 -271 2107
rect -203 2073 -187 2107
rect -129 2073 -113 2107
rect -45 2073 -29 2107
rect 29 2073 45 2107
rect 113 2073 129 2107
rect 187 2073 203 2107
rect 271 2073 287 2107
rect -287 1965 -271 1999
rect -203 1965 -187 1999
rect -129 1965 -113 1999
rect -45 1965 -29 1999
rect 29 1965 45 1999
rect 113 1965 129 1999
rect 187 1965 203 1999
rect 271 1965 287 1999
rect -333 1915 -299 1931
rect -333 1123 -299 1139
rect -175 1915 -141 1931
rect -175 1123 -141 1139
rect -17 1915 17 1931
rect -17 1123 17 1139
rect 141 1915 175 1931
rect 141 1123 175 1139
rect 299 1915 333 1931
rect 299 1123 333 1139
rect -287 1055 -271 1089
rect -203 1055 -187 1089
rect -129 1055 -113 1089
rect -45 1055 -29 1089
rect 29 1055 45 1089
rect 113 1055 129 1089
rect 187 1055 203 1089
rect 271 1055 287 1089
rect -287 947 -271 981
rect -203 947 -187 981
rect -129 947 -113 981
rect -45 947 -29 981
rect 29 947 45 981
rect 113 947 129 981
rect 187 947 203 981
rect 271 947 287 981
rect -333 897 -299 913
rect -333 105 -299 121
rect -175 897 -141 913
rect -175 105 -141 121
rect -17 897 17 913
rect -17 105 17 121
rect 141 897 175 913
rect 141 105 175 121
rect 299 897 333 913
rect 299 105 333 121
rect -287 37 -271 71
rect -203 37 -187 71
rect -129 37 -113 71
rect -45 37 -29 71
rect 29 37 45 71
rect 113 37 129 71
rect 187 37 203 71
rect 271 37 287 71
rect -287 -71 -271 -37
rect -203 -71 -187 -37
rect -129 -71 -113 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 113 -71 129 -37
rect 187 -71 203 -37
rect 271 -71 287 -37
rect -333 -121 -299 -105
rect -333 -913 -299 -897
rect -175 -121 -141 -105
rect -175 -913 -141 -897
rect -17 -121 17 -105
rect -17 -913 17 -897
rect 141 -121 175 -105
rect 141 -913 175 -897
rect 299 -121 333 -105
rect 299 -913 333 -897
rect -287 -981 -271 -947
rect -203 -981 -187 -947
rect -129 -981 -113 -947
rect -45 -981 -29 -947
rect 29 -981 45 -947
rect 113 -981 129 -947
rect 187 -981 203 -947
rect 271 -981 287 -947
rect -287 -1089 -271 -1055
rect -203 -1089 -187 -1055
rect -129 -1089 -113 -1055
rect -45 -1089 -29 -1055
rect 29 -1089 45 -1055
rect 113 -1089 129 -1055
rect 187 -1089 203 -1055
rect 271 -1089 287 -1055
rect -333 -1139 -299 -1123
rect -333 -1931 -299 -1915
rect -175 -1139 -141 -1123
rect -175 -1931 -141 -1915
rect -17 -1139 17 -1123
rect -17 -1931 17 -1915
rect 141 -1139 175 -1123
rect 141 -1931 175 -1915
rect 299 -1139 333 -1123
rect 299 -1931 333 -1915
rect -287 -1999 -271 -1965
rect -203 -1999 -187 -1965
rect -129 -1999 -113 -1965
rect -45 -1999 -29 -1965
rect 29 -1999 45 -1965
rect 113 -1999 129 -1965
rect 187 -1999 203 -1965
rect 271 -1999 287 -1965
rect -287 -2107 -271 -2073
rect -203 -2107 -187 -2073
rect -129 -2107 -113 -2073
rect -45 -2107 -29 -2073
rect 29 -2107 45 -2073
rect 113 -2107 129 -2073
rect 187 -2107 203 -2073
rect 271 -2107 287 -2073
rect -333 -2157 -299 -2141
rect -333 -2949 -299 -2933
rect -175 -2157 -141 -2141
rect -175 -2949 -141 -2933
rect -17 -2157 17 -2141
rect -17 -2949 17 -2933
rect 141 -2157 175 -2141
rect 141 -2949 175 -2933
rect 299 -2157 333 -2141
rect 299 -2949 333 -2933
rect -287 -3017 -271 -2983
rect -203 -3017 -187 -2983
rect -129 -3017 -113 -2983
rect -45 -3017 -29 -2983
rect 29 -3017 45 -2983
rect 113 -3017 129 -2983
rect 187 -3017 203 -2983
rect 271 -3017 287 -2983
rect -467 -3121 -433 -3059
rect 433 -3121 467 -3059
rect -467 -3155 -371 -3121
rect 371 -3155 467 -3121
<< viali >>
rect -271 2983 -203 3017
rect -113 2983 -45 3017
rect 45 2983 113 3017
rect 203 2983 271 3017
rect -333 2157 -299 2933
rect -175 2157 -141 2933
rect -17 2157 17 2933
rect 141 2157 175 2933
rect 299 2157 333 2933
rect -271 2073 -203 2107
rect -113 2073 -45 2107
rect 45 2073 113 2107
rect 203 2073 271 2107
rect -271 1965 -203 1999
rect -113 1965 -45 1999
rect 45 1965 113 1999
rect 203 1965 271 1999
rect -333 1139 -299 1915
rect -175 1139 -141 1915
rect -17 1139 17 1915
rect 141 1139 175 1915
rect 299 1139 333 1915
rect -271 1055 -203 1089
rect -113 1055 -45 1089
rect 45 1055 113 1089
rect 203 1055 271 1089
rect -271 947 -203 981
rect -113 947 -45 981
rect 45 947 113 981
rect 203 947 271 981
rect -333 121 -299 897
rect -175 121 -141 897
rect -17 121 17 897
rect 141 121 175 897
rect 299 121 333 897
rect -271 37 -203 71
rect -113 37 -45 71
rect 45 37 113 71
rect 203 37 271 71
rect -271 -71 -203 -37
rect -113 -71 -45 -37
rect 45 -71 113 -37
rect 203 -71 271 -37
rect -333 -897 -299 -121
rect -175 -897 -141 -121
rect -17 -897 17 -121
rect 141 -897 175 -121
rect 299 -897 333 -121
rect -271 -981 -203 -947
rect -113 -981 -45 -947
rect 45 -981 113 -947
rect 203 -981 271 -947
rect -271 -1089 -203 -1055
rect -113 -1089 -45 -1055
rect 45 -1089 113 -1055
rect 203 -1089 271 -1055
rect -333 -1915 -299 -1139
rect -175 -1915 -141 -1139
rect -17 -1915 17 -1139
rect 141 -1915 175 -1139
rect 299 -1915 333 -1139
rect -271 -1999 -203 -1965
rect -113 -1999 -45 -1965
rect 45 -1999 113 -1965
rect 203 -1999 271 -1965
rect -271 -2107 -203 -2073
rect -113 -2107 -45 -2073
rect 45 -2107 113 -2073
rect 203 -2107 271 -2073
rect -333 -2933 -299 -2157
rect -175 -2933 -141 -2157
rect -17 -2933 17 -2157
rect 141 -2933 175 -2157
rect 299 -2933 333 -2157
rect -271 -3017 -203 -2983
rect -113 -3017 -45 -2983
rect 45 -3017 113 -2983
rect 203 -3017 271 -2983
<< metal1 >>
rect -283 3017 -191 3023
rect -283 2983 -271 3017
rect -203 2983 -191 3017
rect -283 2977 -191 2983
rect -125 3017 -33 3023
rect -125 2983 -113 3017
rect -45 2983 -33 3017
rect -125 2977 -33 2983
rect 33 3017 125 3023
rect 33 2983 45 3017
rect 113 2983 125 3017
rect 33 2977 125 2983
rect 191 3017 283 3023
rect 191 2983 203 3017
rect 271 2983 283 3017
rect 191 2977 283 2983
rect -339 2933 -293 2945
rect -339 2157 -333 2933
rect -299 2157 -293 2933
rect -339 2145 -293 2157
rect -181 2933 -135 2945
rect -181 2157 -175 2933
rect -141 2157 -135 2933
rect -181 2145 -135 2157
rect -23 2933 23 2945
rect -23 2157 -17 2933
rect 17 2157 23 2933
rect -23 2145 23 2157
rect 135 2933 181 2945
rect 135 2157 141 2933
rect 175 2157 181 2933
rect 135 2145 181 2157
rect 293 2933 339 2945
rect 293 2157 299 2933
rect 333 2157 339 2933
rect 293 2145 339 2157
rect -283 2107 -191 2113
rect -283 2073 -271 2107
rect -203 2073 -191 2107
rect -283 2067 -191 2073
rect -125 2107 -33 2113
rect -125 2073 -113 2107
rect -45 2073 -33 2107
rect -125 2067 -33 2073
rect 33 2107 125 2113
rect 33 2073 45 2107
rect 113 2073 125 2107
rect 33 2067 125 2073
rect 191 2107 283 2113
rect 191 2073 203 2107
rect 271 2073 283 2107
rect 191 2067 283 2073
rect -283 1999 -191 2005
rect -283 1965 -271 1999
rect -203 1965 -191 1999
rect -283 1959 -191 1965
rect -125 1999 -33 2005
rect -125 1965 -113 1999
rect -45 1965 -33 1999
rect -125 1959 -33 1965
rect 33 1999 125 2005
rect 33 1965 45 1999
rect 113 1965 125 1999
rect 33 1959 125 1965
rect 191 1999 283 2005
rect 191 1965 203 1999
rect 271 1965 283 1999
rect 191 1959 283 1965
rect -339 1915 -293 1927
rect -339 1139 -333 1915
rect -299 1139 -293 1915
rect -339 1127 -293 1139
rect -181 1915 -135 1927
rect -181 1139 -175 1915
rect -141 1139 -135 1915
rect -181 1127 -135 1139
rect -23 1915 23 1927
rect -23 1139 -17 1915
rect 17 1139 23 1915
rect -23 1127 23 1139
rect 135 1915 181 1927
rect 135 1139 141 1915
rect 175 1139 181 1915
rect 135 1127 181 1139
rect 293 1915 339 1927
rect 293 1139 299 1915
rect 333 1139 339 1915
rect 293 1127 339 1139
rect -283 1089 -191 1095
rect -283 1055 -271 1089
rect -203 1055 -191 1089
rect -283 1049 -191 1055
rect -125 1089 -33 1095
rect -125 1055 -113 1089
rect -45 1055 -33 1089
rect -125 1049 -33 1055
rect 33 1089 125 1095
rect 33 1055 45 1089
rect 113 1055 125 1089
rect 33 1049 125 1055
rect 191 1089 283 1095
rect 191 1055 203 1089
rect 271 1055 283 1089
rect 191 1049 283 1055
rect -283 981 -191 987
rect -283 947 -271 981
rect -203 947 -191 981
rect -283 941 -191 947
rect -125 981 -33 987
rect -125 947 -113 981
rect -45 947 -33 981
rect -125 941 -33 947
rect 33 981 125 987
rect 33 947 45 981
rect 113 947 125 981
rect 33 941 125 947
rect 191 981 283 987
rect 191 947 203 981
rect 271 947 283 981
rect 191 941 283 947
rect -339 897 -293 909
rect -339 121 -333 897
rect -299 121 -293 897
rect -339 109 -293 121
rect -181 897 -135 909
rect -181 121 -175 897
rect -141 121 -135 897
rect -181 109 -135 121
rect -23 897 23 909
rect -23 121 -17 897
rect 17 121 23 897
rect -23 109 23 121
rect 135 897 181 909
rect 135 121 141 897
rect 175 121 181 897
rect 135 109 181 121
rect 293 897 339 909
rect 293 121 299 897
rect 333 121 339 897
rect 293 109 339 121
rect -283 71 -191 77
rect -283 37 -271 71
rect -203 37 -191 71
rect -283 31 -191 37
rect -125 71 -33 77
rect -125 37 -113 71
rect -45 37 -33 71
rect -125 31 -33 37
rect 33 71 125 77
rect 33 37 45 71
rect 113 37 125 71
rect 33 31 125 37
rect 191 71 283 77
rect 191 37 203 71
rect 271 37 283 71
rect 191 31 283 37
rect -283 -37 -191 -31
rect -283 -71 -271 -37
rect -203 -71 -191 -37
rect -283 -77 -191 -71
rect -125 -37 -33 -31
rect -125 -71 -113 -37
rect -45 -71 -33 -37
rect -125 -77 -33 -71
rect 33 -37 125 -31
rect 33 -71 45 -37
rect 113 -71 125 -37
rect 33 -77 125 -71
rect 191 -37 283 -31
rect 191 -71 203 -37
rect 271 -71 283 -37
rect 191 -77 283 -71
rect -339 -121 -293 -109
rect -339 -897 -333 -121
rect -299 -897 -293 -121
rect -339 -909 -293 -897
rect -181 -121 -135 -109
rect -181 -897 -175 -121
rect -141 -897 -135 -121
rect -181 -909 -135 -897
rect -23 -121 23 -109
rect -23 -897 -17 -121
rect 17 -897 23 -121
rect -23 -909 23 -897
rect 135 -121 181 -109
rect 135 -897 141 -121
rect 175 -897 181 -121
rect 135 -909 181 -897
rect 293 -121 339 -109
rect 293 -897 299 -121
rect 333 -897 339 -121
rect 293 -909 339 -897
rect -283 -947 -191 -941
rect -283 -981 -271 -947
rect -203 -981 -191 -947
rect -283 -987 -191 -981
rect -125 -947 -33 -941
rect -125 -981 -113 -947
rect -45 -981 -33 -947
rect -125 -987 -33 -981
rect 33 -947 125 -941
rect 33 -981 45 -947
rect 113 -981 125 -947
rect 33 -987 125 -981
rect 191 -947 283 -941
rect 191 -981 203 -947
rect 271 -981 283 -947
rect 191 -987 283 -981
rect -283 -1055 -191 -1049
rect -283 -1089 -271 -1055
rect -203 -1089 -191 -1055
rect -283 -1095 -191 -1089
rect -125 -1055 -33 -1049
rect -125 -1089 -113 -1055
rect -45 -1089 -33 -1055
rect -125 -1095 -33 -1089
rect 33 -1055 125 -1049
rect 33 -1089 45 -1055
rect 113 -1089 125 -1055
rect 33 -1095 125 -1089
rect 191 -1055 283 -1049
rect 191 -1089 203 -1055
rect 271 -1089 283 -1055
rect 191 -1095 283 -1089
rect -339 -1139 -293 -1127
rect -339 -1915 -333 -1139
rect -299 -1915 -293 -1139
rect -339 -1927 -293 -1915
rect -181 -1139 -135 -1127
rect -181 -1915 -175 -1139
rect -141 -1915 -135 -1139
rect -181 -1927 -135 -1915
rect -23 -1139 23 -1127
rect -23 -1915 -17 -1139
rect 17 -1915 23 -1139
rect -23 -1927 23 -1915
rect 135 -1139 181 -1127
rect 135 -1915 141 -1139
rect 175 -1915 181 -1139
rect 135 -1927 181 -1915
rect 293 -1139 339 -1127
rect 293 -1915 299 -1139
rect 333 -1915 339 -1139
rect 293 -1927 339 -1915
rect -283 -1965 -191 -1959
rect -283 -1999 -271 -1965
rect -203 -1999 -191 -1965
rect -283 -2005 -191 -1999
rect -125 -1965 -33 -1959
rect -125 -1999 -113 -1965
rect -45 -1999 -33 -1965
rect -125 -2005 -33 -1999
rect 33 -1965 125 -1959
rect 33 -1999 45 -1965
rect 113 -1999 125 -1965
rect 33 -2005 125 -1999
rect 191 -1965 283 -1959
rect 191 -1999 203 -1965
rect 271 -1999 283 -1965
rect 191 -2005 283 -1999
rect -283 -2073 -191 -2067
rect -283 -2107 -271 -2073
rect -203 -2107 -191 -2073
rect -283 -2113 -191 -2107
rect -125 -2073 -33 -2067
rect -125 -2107 -113 -2073
rect -45 -2107 -33 -2073
rect -125 -2113 -33 -2107
rect 33 -2073 125 -2067
rect 33 -2107 45 -2073
rect 113 -2107 125 -2073
rect 33 -2113 125 -2107
rect 191 -2073 283 -2067
rect 191 -2107 203 -2073
rect 271 -2107 283 -2073
rect 191 -2113 283 -2107
rect -339 -2157 -293 -2145
rect -339 -2933 -333 -2157
rect -299 -2933 -293 -2157
rect -339 -2945 -293 -2933
rect -181 -2157 -135 -2145
rect -181 -2933 -175 -2157
rect -141 -2933 -135 -2157
rect -181 -2945 -135 -2933
rect -23 -2157 23 -2145
rect -23 -2933 -17 -2157
rect 17 -2933 23 -2157
rect -23 -2945 23 -2933
rect 135 -2157 181 -2145
rect 135 -2933 141 -2157
rect 175 -2933 181 -2157
rect 135 -2945 181 -2933
rect 293 -2157 339 -2145
rect 293 -2933 299 -2157
rect 333 -2933 339 -2157
rect 293 -2945 339 -2933
rect -283 -2983 -191 -2977
rect -283 -3017 -271 -2983
rect -203 -3017 -191 -2983
rect -283 -3023 -191 -3017
rect -125 -2983 -33 -2977
rect -125 -3017 -113 -2983
rect -45 -3017 -33 -2983
rect -125 -3023 -33 -3017
rect 33 -2983 125 -2977
rect 33 -3017 45 -2983
rect 113 -3017 125 -2983
rect 33 -3023 125 -3017
rect 191 -2983 283 -2977
rect 191 -3017 203 -2983
rect 271 -3017 283 -2983
rect 191 -3023 283 -3017
<< properties >>
string FIXED_BBOX -450 -3138 450 3138
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 4 l 0.5 m 6 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
