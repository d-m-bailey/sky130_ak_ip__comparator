magic
tech sky130A
magscale 1 2
timestamp 1715629873
<< pwell >>
rect -328 -658 328 658
<< mvnmos >>
rect -100 -400 100 400
<< mvndiff >>
rect -158 388 -100 400
rect -158 -388 -146 388
rect -112 -388 -100 388
rect -158 -400 -100 -388
rect 100 388 158 400
rect 100 -388 112 388
rect 146 -388 158 388
rect 100 -400 158 -388
<< mvndiffc >>
rect -146 -388 -112 388
rect 112 -388 146 388
<< mvpsubdiff >>
rect -292 610 292 622
rect -292 576 -184 610
rect 184 576 292 610
rect -292 564 292 576
rect -292 514 -234 564
rect -292 -514 -280 514
rect -246 -514 -234 514
rect 234 514 292 564
rect -292 -564 -234 -514
rect 234 -514 246 514
rect 280 -514 292 514
rect 234 -564 292 -514
rect -292 -576 292 -564
rect -292 -610 -184 -576
rect 184 -610 292 -576
rect -292 -622 292 -610
<< mvpsubdiffcont >>
rect -184 576 184 610
rect -280 -514 -246 514
rect 246 -514 280 514
rect -184 -610 184 -576
<< poly >>
rect -100 472 100 488
rect -100 438 -84 472
rect 84 438 100 472
rect -100 400 100 438
rect -100 -438 100 -400
rect -100 -472 -84 -438
rect 84 -472 100 -438
rect -100 -488 100 -472
<< polycont >>
rect -84 438 84 472
rect -84 -472 84 -438
<< locali >>
rect -280 576 -184 610
rect 184 576 280 610
rect -280 514 -246 576
rect 246 514 280 576
rect -100 438 -84 472
rect 84 438 100 472
rect -146 388 -112 404
rect -146 -404 -112 -388
rect 112 388 146 404
rect 112 -404 146 -388
rect -100 -472 -84 -438
rect 84 -472 100 -438
rect -280 -576 -246 -514
rect 246 -576 280 -514
rect -280 -610 -197 -576
rect 197 -610 280 -576
<< viali >>
rect -67 438 67 472
rect -146 -388 -112 388
rect 112 -388 146 388
rect -67 -472 67 -438
rect -197 -610 -184 -576
rect -184 -610 184 -576
rect 184 -610 197 -576
<< metal1 >>
rect -79 472 79 478
rect -79 438 -67 472
rect 67 438 79 472
rect -79 432 79 438
rect -152 388 -106 400
rect -152 -388 -146 388
rect -112 -388 -106 388
rect -152 -400 -106 -388
rect 106 388 152 400
rect 106 -388 112 388
rect 146 -388 152 388
rect 106 -400 152 -388
rect -79 -438 79 -432
rect -79 -472 -67 -438
rect 67 -472 79 -438
rect -79 -478 79 -472
rect -209 -576 209 -570
rect -209 -610 -197 -576
rect 197 -610 209 -576
rect -209 -616 209 -610
<< properties >>
string FIXED_BBOX -263 -593 263 593
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 4 l 1 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 80 viagb 80 viagr 0 viagl 0 viagt 0
<< end >>
