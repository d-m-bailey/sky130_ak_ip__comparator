magic
tech sky130A
magscale 1 2
timestamp 1713548572
<< error_p >>
rect -424 281 -366 287
rect -266 281 -208 287
rect -108 281 -50 287
rect 50 281 108 287
rect 208 281 266 287
rect 366 281 424 287
rect -424 247 -412 281
rect -266 247 -254 281
rect -108 247 -96 281
rect 50 247 62 281
rect 208 247 220 281
rect 366 247 378 281
rect -424 241 -366 247
rect -266 241 -208 247
rect -108 241 -50 247
rect 50 241 108 247
rect 208 241 266 247
rect 366 241 424 247
rect -424 -247 -366 -241
rect -266 -247 -208 -241
rect -108 -247 -50 -241
rect 50 -247 108 -241
rect 208 -247 266 -241
rect 366 -247 424 -241
rect -424 -281 -412 -247
rect -266 -281 -254 -247
rect -108 -281 -96 -247
rect 50 -281 62 -247
rect 208 -281 220 -247
rect 366 -281 378 -247
rect -424 -287 -366 -281
rect -266 -287 -208 -281
rect -108 -287 -50 -281
rect 50 -287 108 -281
rect 208 -287 266 -281
rect 366 -287 424 -281
<< nwell >>
rect -703 -497 703 497
<< mvpmos >>
rect -445 -200 -345 200
rect -287 -200 -187 200
rect -129 -200 -29 200
rect 29 -200 129 200
rect 187 -200 287 200
rect 345 -200 445 200
<< mvpdiff >>
rect -503 188 -445 200
rect -503 -188 -491 188
rect -457 -188 -445 188
rect -503 -200 -445 -188
rect -345 188 -287 200
rect -345 -188 -333 188
rect -299 -188 -287 188
rect -345 -200 -287 -188
rect -187 188 -129 200
rect -187 -188 -175 188
rect -141 -188 -129 188
rect -187 -200 -129 -188
rect -29 188 29 200
rect -29 -188 -17 188
rect 17 -188 29 188
rect -29 -200 29 -188
rect 129 188 187 200
rect 129 -188 141 188
rect 175 -188 187 188
rect 129 -200 187 -188
rect 287 188 345 200
rect 287 -188 299 188
rect 333 -188 345 188
rect 287 -200 345 -188
rect 445 188 503 200
rect 445 -188 457 188
rect 491 -188 503 188
rect 445 -200 503 -188
<< mvpdiffc >>
rect -491 -188 -457 188
rect -333 -188 -299 188
rect -175 -188 -141 188
rect -17 -188 17 188
rect 141 -188 175 188
rect 299 -188 333 188
rect 457 -188 491 188
<< mvnsubdiff >>
rect -637 419 637 431
rect -637 385 -529 419
rect 529 385 637 419
rect -637 373 637 385
rect -637 323 -579 373
rect -637 -323 -625 323
rect -591 -323 -579 323
rect 579 323 637 373
rect -637 -373 -579 -323
rect 579 -323 591 323
rect 625 -323 637 323
rect 579 -373 637 -323
rect -637 -385 637 -373
rect -637 -419 -529 -385
rect 529 -419 637 -385
rect -637 -431 637 -419
<< mvnsubdiffcont >>
rect -529 385 529 419
rect -625 -323 -591 323
rect 591 -323 625 323
rect -529 -419 529 -385
<< poly >>
rect -445 281 -345 297
rect -445 247 -429 281
rect -361 247 -345 281
rect -445 200 -345 247
rect -287 281 -187 297
rect -287 247 -271 281
rect -203 247 -187 281
rect -287 200 -187 247
rect -129 281 -29 297
rect -129 247 -113 281
rect -45 247 -29 281
rect -129 200 -29 247
rect 29 281 129 297
rect 29 247 45 281
rect 113 247 129 281
rect 29 200 129 247
rect 187 281 287 297
rect 187 247 203 281
rect 271 247 287 281
rect 187 200 287 247
rect 345 281 445 297
rect 345 247 361 281
rect 429 247 445 281
rect 345 200 445 247
rect -445 -247 -345 -200
rect -445 -281 -429 -247
rect -361 -281 -345 -247
rect -445 -297 -345 -281
rect -287 -247 -187 -200
rect -287 -281 -271 -247
rect -203 -281 -187 -247
rect -287 -297 -187 -281
rect -129 -247 -29 -200
rect -129 -281 -113 -247
rect -45 -281 -29 -247
rect -129 -297 -29 -281
rect 29 -247 129 -200
rect 29 -281 45 -247
rect 113 -281 129 -247
rect 29 -297 129 -281
rect 187 -247 287 -200
rect 187 -281 203 -247
rect 271 -281 287 -247
rect 187 -297 287 -281
rect 345 -247 445 -200
rect 345 -281 361 -247
rect 429 -281 445 -247
rect 345 -297 445 -281
<< polycont >>
rect -429 247 -361 281
rect -271 247 -203 281
rect -113 247 -45 281
rect 45 247 113 281
rect 203 247 271 281
rect 361 247 429 281
rect -429 -281 -361 -247
rect -271 -281 -203 -247
rect -113 -281 -45 -247
rect 45 -281 113 -247
rect 203 -281 271 -247
rect 361 -281 429 -247
<< locali >>
rect -625 385 -529 419
rect 529 385 625 419
rect -625 323 -591 385
rect 591 323 625 385
rect -445 247 -429 281
rect -361 247 -345 281
rect -287 247 -271 281
rect -203 247 -187 281
rect -129 247 -113 281
rect -45 247 -29 281
rect 29 247 45 281
rect 113 247 129 281
rect 187 247 203 281
rect 271 247 287 281
rect 345 247 361 281
rect 429 247 445 281
rect -491 188 -457 204
rect -491 -204 -457 -188
rect -333 188 -299 204
rect -333 -204 -299 -188
rect -175 188 -141 204
rect -175 -204 -141 -188
rect -17 188 17 204
rect -17 -204 17 -188
rect 141 188 175 204
rect 141 -204 175 -188
rect 299 188 333 204
rect 299 -204 333 -188
rect 457 188 491 204
rect 457 -204 491 -188
rect -445 -281 -429 -247
rect -361 -281 -345 -247
rect -287 -281 -271 -247
rect -203 -281 -187 -247
rect -129 -281 -113 -247
rect -45 -281 -29 -247
rect 29 -281 45 -247
rect 113 -281 129 -247
rect 187 -281 203 -247
rect 271 -281 287 -247
rect 345 -281 361 -247
rect 429 -281 445 -247
rect -625 -385 -591 -323
rect 591 -385 625 -323
rect -625 -419 -529 -385
rect 529 -419 625 -385
<< viali >>
rect -625 -308 -591 308
rect -412 247 -378 281
rect -254 247 -220 281
rect -96 247 -62 281
rect 62 247 96 281
rect 220 247 254 281
rect 378 247 412 281
rect -491 -188 -457 188
rect -333 -188 -299 188
rect -175 -188 -141 188
rect -17 -188 17 188
rect 141 -188 175 188
rect 299 -188 333 188
rect 457 -188 491 188
rect -412 -281 -378 -247
rect -254 -281 -220 -247
rect -96 -281 -62 -247
rect 62 -281 96 -247
rect 220 -281 254 -247
rect 378 -281 412 -247
rect 591 -308 625 308
rect -473 -419 473 -385
<< metal1 >>
rect -631 308 -585 320
rect -631 -308 -625 308
rect -591 -308 -585 308
rect 585 308 631 320
rect -424 281 -366 287
rect -424 247 -412 281
rect -378 247 -366 281
rect -424 241 -366 247
rect -266 281 -208 287
rect -266 247 -254 281
rect -220 247 -208 281
rect -266 241 -208 247
rect -108 281 -50 287
rect -108 247 -96 281
rect -62 247 -50 281
rect -108 241 -50 247
rect 50 281 108 287
rect 50 247 62 281
rect 96 247 108 281
rect 50 241 108 247
rect 208 281 266 287
rect 208 247 220 281
rect 254 247 266 281
rect 208 241 266 247
rect 366 281 424 287
rect 366 247 378 281
rect 412 247 424 281
rect 366 241 424 247
rect -497 188 -451 200
rect -497 -188 -491 188
rect -457 -188 -451 188
rect -497 -200 -451 -188
rect -339 188 -293 200
rect -339 -188 -333 188
rect -299 -188 -293 188
rect -339 -200 -293 -188
rect -181 188 -135 200
rect -181 -188 -175 188
rect -141 -188 -135 188
rect -181 -200 -135 -188
rect -23 188 23 200
rect -23 -188 -17 188
rect 17 -188 23 188
rect -23 -200 23 -188
rect 135 188 181 200
rect 135 -188 141 188
rect 175 -188 181 188
rect 135 -200 181 -188
rect 293 188 339 200
rect 293 -188 299 188
rect 333 -188 339 188
rect 293 -200 339 -188
rect 451 188 497 200
rect 451 -188 457 188
rect 491 -188 497 188
rect 451 -200 497 -188
rect -424 -247 -366 -241
rect -424 -281 -412 -247
rect -378 -281 -366 -247
rect -424 -287 -366 -281
rect -266 -247 -208 -241
rect -266 -281 -254 -247
rect -220 -281 -208 -247
rect -266 -287 -208 -281
rect -108 -247 -50 -241
rect -108 -281 -96 -247
rect -62 -281 -50 -247
rect -108 -287 -50 -281
rect 50 -247 108 -241
rect 50 -281 62 -247
rect 96 -281 108 -247
rect 50 -287 108 -281
rect 208 -247 266 -241
rect 208 -281 220 -247
rect 254 -281 266 -247
rect 208 -287 266 -281
rect 366 -247 424 -241
rect 366 -281 378 -247
rect 412 -281 424 -247
rect 366 -287 424 -281
rect -631 -320 -585 -308
rect 585 -308 591 308
rect 625 -308 631 308
rect 585 -320 631 -308
rect -485 -385 485 -379
rect -485 -419 -473 -385
rect 473 -419 485 -385
rect -485 -425 485 -419
<< properties >>
string FIXED_BBOX -608 -402 608 402
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 2 l 0.5 m 1 nf 6 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 80 viagr 80 viagl 80 viagt 0
<< end >>
