magic
tech sky130A
magscale 1 2
timestamp 1713076297
<< nwell >>
rect -545 -662 545 662
<< mvpmos >>
rect -287 -436 -187 364
rect -129 -436 -29 364
rect 29 -436 129 364
rect 187 -436 287 364
<< mvpdiff >>
rect -345 352 -287 364
rect -345 -424 -333 352
rect -299 -424 -287 352
rect -345 -436 -287 -424
rect -187 352 -129 364
rect -187 -424 -175 352
rect -141 -424 -129 352
rect -187 -436 -129 -424
rect -29 352 29 364
rect -29 -424 -17 352
rect 17 -424 29 352
rect -29 -436 29 -424
rect 129 352 187 364
rect 129 -424 141 352
rect 175 -424 187 352
rect 129 -436 187 -424
rect 287 352 345 364
rect 287 -424 299 352
rect 333 -424 345 352
rect 287 -436 345 -424
<< mvpdiffc >>
rect -333 -424 -299 352
rect -175 -424 -141 352
rect -17 -424 17 352
rect 141 -424 175 352
rect 299 -424 333 352
<< mvnsubdiff >>
rect -479 584 479 596
rect -479 550 -371 584
rect 371 550 479 584
rect -479 538 479 550
rect -479 488 -421 538
rect -479 -488 -467 488
rect -433 -488 -421 488
rect 421 488 479 538
rect -479 -538 -421 -488
rect 421 -488 433 488
rect 467 -488 479 488
rect 421 -538 479 -488
rect -479 -550 479 -538
rect -479 -584 -371 -550
rect 371 -584 479 -550
rect -479 -596 479 -584
<< mvnsubdiffcont >>
rect -371 550 371 584
rect -467 -488 -433 488
rect 433 -488 467 488
rect -371 -584 371 -550
<< poly >>
rect -287 445 -187 461
rect -287 411 -271 445
rect -203 411 -187 445
rect -287 364 -187 411
rect -129 445 -29 461
rect -129 411 -113 445
rect -45 411 -29 445
rect -129 364 -29 411
rect 29 445 129 461
rect 29 411 45 445
rect 113 411 129 445
rect 29 364 129 411
rect 187 445 287 461
rect 187 411 203 445
rect 271 411 287 445
rect 187 364 287 411
rect -287 -462 -187 -436
rect -129 -462 -29 -436
rect 29 -462 129 -436
rect 187 -462 287 -436
<< polycont >>
rect -271 411 -203 445
rect -113 411 -45 445
rect 45 411 113 445
rect 203 411 271 445
<< locali >>
rect -467 550 -371 584
rect 371 550 467 584
rect -467 488 -433 550
rect 433 488 467 550
rect -287 411 -271 445
rect -203 411 -187 445
rect -129 411 -113 445
rect -45 411 -29 445
rect 29 411 45 445
rect 113 411 129 445
rect 187 411 203 445
rect 271 411 287 445
rect -333 352 -299 368
rect -333 -440 -299 -424
rect -175 352 -141 368
rect -175 -440 -141 -424
rect -17 352 17 368
rect -17 -440 17 -424
rect 141 352 175 368
rect 141 -440 175 -424
rect 299 352 333 368
rect 299 -440 333 -424
rect -467 -550 -433 -488
rect 433 -550 467 -488
rect -467 -584 -371 -550
rect 371 -584 467 -550
<< viali >>
rect -264 411 -210 445
rect -106 411 -52 445
rect 52 411 106 445
rect 210 411 264 445
rect -333 -424 -299 352
rect -175 -424 -141 352
rect -17 -424 17 352
rect 141 -424 175 352
rect 299 -424 333 352
<< metal1 >>
rect -276 445 -198 451
rect -276 411 -264 445
rect -210 411 -198 445
rect -276 405 -198 411
rect -118 445 -40 451
rect -118 411 -106 445
rect -52 411 -40 445
rect -118 405 -40 411
rect 40 445 118 451
rect 40 411 52 445
rect 106 411 118 445
rect 40 405 118 411
rect 198 445 276 451
rect 198 411 210 445
rect 264 411 276 445
rect 198 405 276 411
rect -339 352 -293 364
rect -339 -424 -333 352
rect -299 -424 -293 352
rect -339 -436 -293 -424
rect -181 352 -135 364
rect -181 -424 -175 352
rect -141 -424 -135 352
rect -181 -436 -135 -424
rect -23 352 23 364
rect -23 -424 -17 352
rect 17 -424 23 352
rect -23 -436 23 -424
rect 135 352 181 364
rect 135 -424 141 352
rect 175 -424 181 352
rect 135 -436 181 -424
rect 293 352 339 364
rect 293 -424 299 352
rect 333 -424 339 352
rect 293 -436 339 -424
<< properties >>
string FIXED_BBOX -450 -567 450 567
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 4 l 0.5 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 80 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
