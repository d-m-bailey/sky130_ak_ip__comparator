magic
tech sky130A
magscale 1 2
timestamp 1713589649
<< error_p >>
rect -269 272 -205 278
rect -111 272 -47 278
rect 47 272 111 278
rect 205 272 269 278
rect -269 238 -257 272
rect -111 238 -99 272
rect 47 238 59 272
rect 205 238 217 272
rect -269 232 -205 238
rect -111 232 -47 238
rect 47 232 111 238
rect 205 232 269 238
rect -269 -238 -205 -232
rect -111 -238 -47 -232
rect 47 -238 111 -232
rect 205 -238 269 -232
rect -269 -272 -257 -238
rect -111 -272 -99 -238
rect 47 -272 59 -238
rect 205 -272 217 -238
rect -269 -278 -205 -272
rect -111 -278 -47 -272
rect 47 -278 111 -272
rect 205 -278 269 -272
<< pwell >>
rect -515 -458 515 458
<< mvnmos >>
rect -287 -200 -187 200
rect -129 -200 -29 200
rect 29 -200 129 200
rect 187 -200 287 200
<< mvndiff >>
rect -345 188 -287 200
rect -345 -188 -333 188
rect -299 -188 -287 188
rect -345 -200 -287 -188
rect -187 188 -129 200
rect -187 -188 -175 188
rect -141 -188 -129 188
rect -187 -200 -129 -188
rect -29 188 29 200
rect -29 -188 -17 188
rect 17 -188 29 188
rect -29 -200 29 -188
rect 129 188 187 200
rect 129 -188 141 188
rect 175 -188 187 188
rect 129 -200 187 -188
rect 287 188 345 200
rect 287 -188 299 188
rect 333 -188 345 188
rect 287 -200 345 -188
<< mvndiffc >>
rect -333 -188 -299 188
rect -175 -188 -141 188
rect -17 -188 17 188
rect 141 -188 175 188
rect 299 -188 333 188
<< mvpsubdiff >>
rect -479 410 479 422
rect -479 376 -371 410
rect 371 376 479 410
rect -479 364 479 376
rect -479 314 -421 364
rect -479 -314 -467 314
rect -433 -314 -421 314
rect 421 314 479 364
rect -479 -364 -421 -314
rect 421 -314 433 314
rect 467 -314 479 314
rect 421 -364 479 -314
rect -479 -376 479 -364
rect -479 -410 -371 -376
rect 371 -410 479 -376
rect -479 -422 479 -410
<< mvpsubdiffcont >>
rect -371 376 371 410
rect -467 -314 -433 314
rect 433 -314 467 314
rect -371 -410 371 -376
<< poly >>
rect -287 272 -187 288
rect -287 238 -271 272
rect -203 238 -187 272
rect -287 200 -187 238
rect -129 272 -29 288
rect -129 238 -113 272
rect -45 238 -29 272
rect -129 200 -29 238
rect 29 272 129 288
rect 29 238 45 272
rect 113 238 129 272
rect 29 200 129 238
rect 187 272 287 288
rect 187 238 203 272
rect 271 238 287 272
rect 187 200 287 238
rect -287 -238 -187 -200
rect -287 -272 -271 -238
rect -203 -272 -187 -238
rect -287 -288 -187 -272
rect -129 -238 -29 -200
rect -129 -272 -113 -238
rect -45 -272 -29 -238
rect -129 -288 -29 -272
rect 29 -238 129 -200
rect 29 -272 45 -238
rect 113 -272 129 -238
rect 29 -288 129 -272
rect 187 -238 287 -200
rect 187 -272 203 -238
rect 271 -272 287 -238
rect 187 -288 287 -272
<< polycont >>
rect -271 238 -203 272
rect -113 238 -45 272
rect 45 238 113 272
rect 203 238 271 272
rect -271 -272 -203 -238
rect -113 -272 -45 -238
rect 45 -272 113 -238
rect 203 -272 271 -238
<< locali >>
rect -467 376 -371 410
rect 371 376 467 410
rect -467 314 -433 376
rect 433 314 467 376
rect -287 238 -271 272
rect -203 238 -187 272
rect -129 238 -113 272
rect -45 238 -29 272
rect 29 238 45 272
rect 113 238 129 272
rect 187 238 203 272
rect 271 238 287 272
rect -333 188 -299 204
rect -333 -204 -299 -188
rect -175 188 -141 204
rect -175 -204 -141 -188
rect -17 188 17 204
rect -17 -204 17 -188
rect 141 188 175 204
rect 141 -204 175 -188
rect 299 188 333 204
rect 299 -204 333 -188
rect -287 -272 -271 -238
rect -203 -272 -187 -238
rect -129 -272 -113 -238
rect -45 -272 -29 -238
rect 29 -272 45 -238
rect 113 -272 129 -238
rect 187 -272 203 -238
rect 271 -272 287 -238
rect -467 -376 -433 -314
rect 433 -376 467 -314
rect -467 -410 -371 -376
rect 371 -410 467 -376
<< viali >>
rect -467 -301 -433 301
rect -257 238 -217 272
rect -99 238 -59 272
rect 59 238 99 272
rect 217 238 257 272
rect -333 -188 -299 188
rect -175 -188 -141 188
rect -17 -188 17 188
rect 141 -188 175 188
rect 299 -188 333 188
rect -257 -272 -217 -238
rect -99 -272 -59 -238
rect 59 -272 99 -238
rect 217 -272 257 -238
rect 433 -301 467 301
rect -346 -410 346 -376
<< metal1 >>
rect -473 301 -427 313
rect -473 -301 -467 301
rect -433 -301 -427 301
rect 427 301 473 313
rect -269 272 -205 278
rect -269 238 -257 272
rect -217 238 -205 272
rect -269 232 -205 238
rect -111 272 -47 278
rect -111 238 -99 272
rect -59 238 -47 272
rect -111 232 -47 238
rect 47 272 111 278
rect 47 238 59 272
rect 99 238 111 272
rect 47 232 111 238
rect 205 272 269 278
rect 205 238 217 272
rect 257 238 269 272
rect 205 232 269 238
rect -339 188 -293 200
rect -339 -188 -333 188
rect -299 -188 -293 188
rect -339 -200 -293 -188
rect -181 188 -135 200
rect -181 -188 -175 188
rect -141 -188 -135 188
rect -181 -200 -135 -188
rect -23 188 23 200
rect -23 -188 -17 188
rect 17 -188 23 188
rect -23 -200 23 -188
rect 135 188 181 200
rect 135 -188 141 188
rect 175 -188 181 188
rect 135 -200 181 -188
rect 293 188 339 200
rect 293 -188 299 188
rect 333 -188 339 188
rect 293 -200 339 -188
rect -269 -238 -205 -232
rect -269 -272 -257 -238
rect -217 -272 -205 -238
rect -269 -278 -205 -272
rect -111 -238 -47 -232
rect -111 -272 -99 -238
rect -59 -272 -47 -238
rect -111 -278 -47 -272
rect 47 -238 111 -232
rect 47 -272 59 -238
rect 99 -272 111 -238
rect 47 -278 111 -272
rect 205 -238 269 -232
rect 205 -272 217 -238
rect 257 -272 269 -238
rect 205 -278 269 -272
rect -473 -313 -427 -301
rect 427 -301 433 301
rect 467 -301 473 301
rect 427 -313 473 -301
rect -358 -376 358 -370
rect -358 -410 -346 -376
rect 346 -410 358 -376
rect -358 -416 358 -410
<< properties >>
string FIXED_BBOX -450 -393 450 393
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 2 l 0.50 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 60 viagb 80 viagr 80 viagl 80 viagt 0
<< end >>
