magic
tech sky130A
timestamp 1713550110
<< pwell >>
rect -139 -388 139 388
<< mvnmos >>
rect -25 159 25 259
rect -25 -50 25 50
rect -25 -259 25 -159
<< mvndiff >>
rect -54 253 -25 259
rect -54 165 -48 253
rect -31 165 -25 253
rect -54 159 -25 165
rect 25 253 54 259
rect 25 165 31 253
rect 48 165 54 253
rect 25 159 54 165
rect -54 44 -25 50
rect -54 -44 -48 44
rect -31 -44 -25 44
rect -54 -50 -25 -44
rect 25 44 54 50
rect 25 -44 31 44
rect 48 -44 54 44
rect 25 -50 54 -44
rect -54 -165 -25 -159
rect -54 -253 -48 -165
rect -31 -253 -25 -165
rect -54 -259 -25 -253
rect 25 -165 54 -159
rect 25 -253 31 -165
rect 48 -253 54 -165
rect 25 -259 54 -253
<< mvndiffc >>
rect -48 165 -31 253
rect 31 165 48 253
rect -48 -44 -31 44
rect 31 -44 48 44
rect -48 -253 -31 -165
rect 31 -253 48 -165
<< mvpsubdiff >>
rect -121 364 121 370
rect -121 347 -67 364
rect 67 347 121 364
rect -121 341 121 347
rect -121 316 -92 341
rect -121 -316 -115 316
rect -98 -316 -92 316
rect 92 316 121 341
rect -121 -341 -92 -316
rect 92 -316 98 316
rect 115 -316 121 316
rect 92 -341 121 -316
rect -121 -347 121 -341
rect -121 -364 -67 -347
rect 67 -364 121 -347
rect -121 -370 121 -364
<< mvpsubdiffcont >>
rect -67 347 67 364
rect -115 -316 -98 316
rect 98 -316 115 316
rect -67 -364 67 -347
<< poly >>
rect -25 295 25 303
rect -25 278 -17 295
rect 17 278 25 295
rect -25 259 25 278
rect -25 140 25 159
rect -25 123 -17 140
rect 17 123 25 140
rect -25 115 25 123
rect -25 86 25 94
rect -25 69 -17 86
rect 17 69 25 86
rect -25 50 25 69
rect -25 -69 25 -50
rect -25 -86 -17 -69
rect 17 -86 25 -69
rect -25 -94 25 -86
rect -25 -123 25 -115
rect -25 -140 -17 -123
rect 17 -140 25 -123
rect -25 -159 25 -140
rect -25 -278 25 -259
rect -25 -295 -17 -278
rect 17 -295 25 -278
rect -25 -303 25 -295
<< polycont >>
rect -17 278 17 295
rect -17 123 17 140
rect -17 69 17 86
rect -17 -86 17 -69
rect -17 -140 17 -123
rect -17 -295 17 -278
<< locali >>
rect -115 347 -67 364
rect 67 347 115 364
rect -115 316 -98 347
rect 98 316 115 347
rect -25 278 -17 295
rect 17 278 25 295
rect -48 253 -31 261
rect -48 157 -31 165
rect 31 253 48 261
rect 31 157 48 165
rect -25 123 -17 140
rect 17 123 25 140
rect -25 69 -17 86
rect 17 69 25 86
rect -48 44 -31 52
rect -48 -52 -31 -44
rect 31 44 48 52
rect 31 -52 48 -44
rect -25 -86 -17 -69
rect 17 -86 25 -69
rect -25 -140 -17 -123
rect 17 -140 25 -123
rect -48 -165 -31 -157
rect -48 -261 -31 -253
rect 31 -165 48 -157
rect 31 -261 48 -253
rect -25 -295 -17 -278
rect 17 -295 25 -278
rect -115 -347 -98 -316
rect 98 -347 115 -316
rect -115 -364 -67 -347
rect 67 -364 115 -347
<< viali >>
rect -17 278 17 295
rect -48 165 -31 253
rect 31 165 48 253
rect -17 123 17 140
rect -17 69 17 86
rect -48 -44 -31 44
rect 31 -44 48 44
rect -17 -86 17 -69
rect -17 -140 17 -123
rect -48 -253 -31 -165
rect 31 -253 48 -165
rect -17 -295 17 -278
<< metal1 >>
rect -23 295 23 298
rect -23 278 -17 295
rect 17 278 23 295
rect -23 275 23 278
rect -51 253 -28 259
rect -51 165 -48 253
rect -31 165 -28 253
rect -51 159 -28 165
rect 28 253 51 259
rect 28 165 31 253
rect 48 165 51 253
rect 28 159 51 165
rect -23 140 23 143
rect -23 123 -17 140
rect 17 123 23 140
rect -23 120 23 123
rect -23 86 23 89
rect -23 69 -17 86
rect 17 69 23 86
rect -23 66 23 69
rect -51 44 -28 50
rect -51 -44 -48 44
rect -31 -44 -28 44
rect -51 -50 -28 -44
rect 28 44 51 50
rect 28 -44 31 44
rect 48 -44 51 44
rect 28 -50 51 -44
rect -23 -69 23 -66
rect -23 -86 -17 -69
rect 17 -86 23 -69
rect -23 -89 23 -86
rect -23 -123 23 -120
rect -23 -140 -17 -123
rect 17 -140 23 -123
rect -23 -143 23 -140
rect -51 -165 -28 -159
rect -51 -253 -48 -165
rect -31 -253 -28 -165
rect -51 -259 -28 -253
rect 28 -165 51 -159
rect 28 -253 31 -165
rect 48 -253 51 -165
rect 28 -259 51 -253
rect -23 -278 23 -275
rect -23 -295 -17 -278
rect 17 -295 23 -278
rect -23 -298 23 -295
<< properties >>
string FIXED_BBOX -106 -355 106 355
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 1 l 0.50 m 3 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
