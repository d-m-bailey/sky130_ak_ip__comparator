magic
tech sky130A
magscale 1 2
timestamp 1713072694
<< pwell >>
rect -3115 -2878 3115 2878
<< psubdiff >>
rect -3079 2808 -2983 2842
rect 2983 2808 3079 2842
rect -3079 2746 -3045 2808
rect 3045 2746 3079 2808
rect -3079 -2808 -3045 -2746
rect 3045 -2808 3079 -2746
rect -3079 -2842 -2983 -2808
rect 2983 -2842 3079 -2808
<< psubdiffcont >>
rect -2983 2808 2983 2842
rect -3079 -2746 -3045 2746
rect 3045 -2746 3079 2746
rect -2983 -2842 2983 -2808
<< xpolycontact >>
rect -2949 2280 -2379 2712
rect -2949 -2712 -2379 -2280
rect -2283 2280 -1713 2712
rect -2283 -2712 -1713 -2280
rect -1617 2280 -1047 2712
rect -1617 -2712 -1047 -2280
rect -951 2280 -381 2712
rect -951 -2712 -381 -2280
rect -285 2280 285 2712
rect -285 -2712 285 -2280
rect 381 2280 951 2712
rect 381 -2712 951 -2280
rect 1047 2280 1617 2712
rect 1047 -2712 1617 -2280
rect 1713 2280 2283 2712
rect 1713 -2712 2283 -2280
rect 2379 2280 2949 2712
rect 2379 -2712 2949 -2280
<< ppolyres >>
rect -2949 -2280 -2379 2280
rect -2283 -2280 -1713 2280
rect -1617 -2280 -1047 2280
rect -951 -2280 -381 2280
rect -285 -2280 285 2280
rect 381 -2280 951 2280
rect 1047 -2280 1617 2280
rect 1713 -2280 2283 2280
rect 2379 -2280 2949 2280
<< locali >>
rect -3079 2808 -2983 2842
rect 2983 2808 3079 2842
rect -3079 2746 -3045 2808
rect 3045 2746 3079 2808
rect -3079 -2808 -3045 -2746
rect 3045 -2808 3079 -2746
rect -3079 -2842 -2983 -2808
rect 2983 -2842 3079 -2808
<< viali >>
rect -2741 2808 2741 2842
rect -3079 -2527 -3045 2527
rect -2933 2297 -2395 2694
rect -2267 2297 -1729 2694
rect -1601 2297 -1063 2694
rect -935 2297 -397 2694
rect -269 2297 269 2694
rect 397 2297 935 2694
rect 1063 2297 1601 2694
rect 1729 2297 2267 2694
rect 2395 2297 2933 2694
rect -2933 -2694 -2395 -2297
rect -2267 -2694 -1729 -2297
rect -1601 -2694 -1063 -2297
rect -935 -2694 -397 -2297
rect -269 -2694 269 -2297
rect 397 -2694 935 -2297
rect 1063 -2694 1601 -2297
rect 1729 -2694 2267 -2297
rect 2395 -2694 2933 -2297
rect 3045 -2527 3079 2527
rect -2741 -2842 2741 -2808
<< metal1 >>
rect -2753 2842 2753 2848
rect -2753 2808 -2741 2842
rect 2741 2808 2753 2842
rect -2753 2802 2753 2808
rect -2945 2694 -2383 2700
rect -3085 2527 -3039 2539
rect -3085 -2527 -3079 2527
rect -3045 -2527 -3039 2527
rect -2945 2297 -2933 2694
rect -2395 2297 -2383 2694
rect -2945 2291 -2383 2297
rect -2279 2694 -1717 2700
rect -2279 2297 -2267 2694
rect -1729 2297 -1717 2694
rect -2279 2291 -1717 2297
rect -1613 2694 -1051 2700
rect -1613 2297 -1601 2694
rect -1063 2297 -1051 2694
rect -1613 2291 -1051 2297
rect -947 2694 -385 2700
rect -947 2297 -935 2694
rect -397 2297 -385 2694
rect -947 2291 -385 2297
rect -281 2694 281 2700
rect -281 2297 -269 2694
rect 269 2297 281 2694
rect -281 2291 281 2297
rect 385 2694 947 2700
rect 385 2297 397 2694
rect 935 2297 947 2694
rect 385 2291 947 2297
rect 1051 2694 1613 2700
rect 1051 2297 1063 2694
rect 1601 2297 1613 2694
rect 1051 2291 1613 2297
rect 1717 2694 2279 2700
rect 1717 2297 1729 2694
rect 2267 2297 2279 2694
rect 1717 2291 2279 2297
rect 2383 2694 2945 2700
rect 2383 2297 2395 2694
rect 2933 2297 2945 2694
rect 2383 2291 2945 2297
rect 3039 2527 3085 2539
rect -3085 -2539 -3039 -2527
rect -2945 -2297 -2383 -2291
rect -2945 -2694 -2933 -2297
rect -2395 -2694 -2383 -2297
rect -2945 -2700 -2383 -2694
rect -2279 -2297 -1717 -2291
rect -2279 -2694 -2267 -2297
rect -1729 -2694 -1717 -2297
rect -2279 -2700 -1717 -2694
rect -1613 -2297 -1051 -2291
rect -1613 -2694 -1601 -2297
rect -1063 -2694 -1051 -2297
rect -1613 -2700 -1051 -2694
rect -947 -2297 -385 -2291
rect -947 -2694 -935 -2297
rect -397 -2694 -385 -2297
rect -947 -2700 -385 -2694
rect -281 -2297 281 -2291
rect -281 -2694 -269 -2297
rect 269 -2694 281 -2297
rect -281 -2700 281 -2694
rect 385 -2297 947 -2291
rect 385 -2694 397 -2297
rect 935 -2694 947 -2297
rect 385 -2700 947 -2694
rect 1051 -2297 1613 -2291
rect 1051 -2694 1063 -2297
rect 1601 -2694 1613 -2297
rect 1051 -2700 1613 -2694
rect 1717 -2297 2279 -2291
rect 1717 -2694 1729 -2297
rect 2267 -2694 2279 -2297
rect 1717 -2700 2279 -2694
rect 2383 -2297 2945 -2291
rect 2383 -2694 2395 -2297
rect 2933 -2694 2945 -2297
rect 3039 -2527 3045 2527
rect 3079 -2527 3085 2527
rect 3039 -2539 3085 -2527
rect 2383 -2700 2945 -2694
rect -2753 -2808 2753 -2802
rect -2753 -2842 -2741 -2808
rect 2741 -2842 2753 -2808
rect -2753 -2848 2753 -2842
<< res2p85 >>
rect -2951 -2282 -2377 2282
rect -2285 -2282 -1711 2282
rect -1619 -2282 -1045 2282
rect -953 -2282 -379 2282
rect -287 -2282 287 2282
rect 379 -2282 953 2282
rect 1045 -2282 1619 2282
rect 1711 -2282 2285 2282
rect 2377 -2282 2951 2282
<< properties >>
string FIXED_BBOX -3062 -2825 3062 2825
string gencell sky130_fd_pr__res_high_po_2p85
string library sky130
string parameters w 2.85 l 22.8 m 1 nx 9 wmin 2.850 lmin 0.50 rho 319.8 val 2.695k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 2.850 n_guard 0 hv_guard 0 vias 1 viagb 90 viagt 90 viagl 90 viagr 90
<< end >>
