* NGSPICE file created from comparator_rcx.ext - technology: sky130A

.subckt comparator_rcx Vinp Vinm AGND en hyst[1] hyst[0] trim[5] trim[4] trim[3] trim[2]
+ trim[1] trim[0] Vout ibias DVDD AVDD DGND
X0 a_1659_n4497.t93 casc_n.t37 Vxm.t67 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1 AVDD.t706 AVDD.t704 AVDD.t705 AVDD.t401 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2 a_1657_n21342.t154 a_1560_n22142.t10 AVDD.t327 AVDD.t203 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X3 Vom.t79 casc_p.t70 a_2458_5328.t113 AVDD.t68 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X4 a_1659_n4497.t92 casc_n.t38 Vxm.t68 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5 a_2458_5328.t67 a_12760_n20342.t5 AVDD.t251 AVDD.t68 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X6 casc_p.t63 casc_p.t61 casc_p.t62 AVDD.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7 a_2467_n29152.t5 a_2370_n29452.t8 Vfold_bot_m.t18 AVDD.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X8 a_1659_n4497.t91 casc_n.t39 Vxm.t69 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9 Vom.t78 casc_p.t71 a_2458_5328.t112 AVDD.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10 Vop.t79 casc_p.t72 a_2458_6128.t159 AVDD.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X11 Vxp.t136 casc_p.t73 a_1657_n21342.t155 AVDD.t155 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12 level_shifter_up_8.x_hv a_34648_11527# DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=3.103e+14p ps=2.34242e+09u w=1e+06u l=500000u
X13 a_23013_n25097.t15 casc_p.t74 a_33657_n21342.t2 AVDD.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14 a_2458_6128.t86 bias_p.t11 AVDD.t277 AVDD.t148 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X15 a_2458_6128.t87 bias_p.t12 AVDD.t278 AVDD.t5 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X16 Vop.t78 casc_p.t75 a_2458_6128.t158 AVDD.t74 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X17 Vxp.t135 casc_p.t76 a_1657_n21342.t156 AVDD.t172 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X18 a_2467_n30310.t108 casc_n.t40 Vop.t109 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X19 Vfold_bot_m.t104 casc_n.t41 Vom.t119 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X20 a_32057_n15000.t33 level_shifter_up_0.xb_hv.t2 AVDD.t288 AVDD.t287 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X21 a_32059_n897.t11 casc_n.t42 a_2458_6570.t11 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X22 casc_n.t36 casc_n.t34 casc_n.t35 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X23 a_1657_n21342.t153 a_1560_n22142.t11 AVDD.t328 AVDD.t163 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X24 AVDD.t703 AVDD.t701 AVDD.t702 AVDD.t366 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X25 a_2458_5328.t193 bias_p.t13 AVDD.t805 AVDD.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X26 Vop.t77 casc_p.t77 a_2458_6128.t136 AVDD.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X27 AVDD.t700 AVDD.t698 AVDD.t699 AVDD.t374 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X28 a_2458_5328.t0 Vinp.t0 Vxm.t0 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X29 AVDD.t697 AVDD.t695 AVDD.t696 AVDD.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X30 a_2458_6128.t61 a_12760_n20342.t6 AVDD.t252 AVDD.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X31 AVDD.t694 AVDD.t692 AVDD.t693 AVDD.t374 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X32 AVDD.t691 AVDD.t689 AVDD.t690 AVDD.t370 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X33 Vom.t77 casc_p.t78 a_2458_5328.t111 AVDD.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X34 DGND bias_var_n bias_var_n DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.16e+12p ps=9.16e+06u w=2e+06u l=4e+06u
X35 a_32057_n13616.t16 casc_p.t79 a_32057_n8742.t10 AVDD.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X36 a_11160_n9542.t3 a_11160_n9542.t2 a_11257_n8742.t5 AVDD.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X37 AVDD.t688 AVDD.t686 AVDD.t687 AVDD.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X38 Vop.t76 casc_p.t80 a_2458_6128.t135 AVDD.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X39 bias_p bias_p.t1 AVDD.t45 AVDD.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=5.8e+12p pd=4.406e+07u as=0p ps=0u w=2e+06u l=4e+06u
X40 a_23032_4566.t7 level_shifter_up_8.xb_hv.t1 a_2370_6628.t1 AVDD.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X41 Vop.t75 casc_p.t81 a_2458_6128.t134 AVDD.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X42 AVDD.t60 level_shifter_up_5.xb_hv.t2 a_32057_n9600.t11 AVDD.t59 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X43 a_31928_n30483# trim[5].t0 DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=500000u
X44 DGND bias_n.t8 casc_n.t1 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X45 a_36328_n30483# trim[3].t0 DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=500000u
X46 a_32057_n14142.t17 bias_p.t14 a_32057_n15000.t5 AVDD.t147 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X47 a_23013_n25097.t21 level_shifter_up_3.x_hv.t2 a_2370_n28652.t3 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X48 casc_n.t33 casc_n.t31 casc_n.t32 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X49 Vxp.t3 Vinm.t0 a_2467_n30310.t0 AVDD.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X50 a_1657_n21342.t152 a_1560_n22142.t12 AVDD.t329 AVDD.t159 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X51 Vom.t76 casc_p.t82 a_2458_5328.t151 AVDD.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X52 Vom.t75 casc_p.t83 a_2458_5328.t150 AVDD.t15 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X53 bias_n.t7 level_shifter_up_4.xb_hv.t2 DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X54 a_2458_6128.t189 a_35086_7130.t2 a_32059_n4755.t24 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X55 res_p_bot.t6 a_25011_n25097# DGND sky130_fd_pr__res_high_po_2p85 l=3.192e+07u
X56 level_shifter_up_2.x_hv a_34128_n30483# DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X57 a_2458_6128.t60 a_12760_n20342.t7 AVDD.t253 AVDD.t113 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X58 a_1659_n4497.t90 casc_n.t43 Vxm.t70 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X59 a_2458_5328.t197 a_2370_6628.t8 a_2458_6570.t13 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X60 a_1659_n4497.t89 casc_n.t44 Vxm.t71 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X61 DGND bias_var_n.t7 Vfold_bot_m.t55 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X62 Vxp.t4 Vinm.t1 a_2467_n30310.t1 AVDD.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X63 DGND a_36699_n29829# a_36259_n29829# DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X64 a_2370_6628.t0 level_shifter_up_8.xb_hv.t2 a_23032_4566.t6 AVDD.t37 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X65 a_2458_6128.t5 Vinm.t2 Vxm.t4 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X66 Vop.t74 casc_p.t84 a_2458_6128.t133 AVDD.t148 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X67 AVDD.t685 AVDD.t683 AVDD.t684 AVDD.t394 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X68 Vop.t73 casc_p.t85 a_2458_6128.t132 AVDD.t125 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X69 Vop.t72 casc_p.t86 a_2458_6128.t106 AVDD.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X70 a_2458_6128.t59 a_12760_n20342.t8 AVDD.t254 AVDD.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X71 DGND.t146 Vop_stg2.t3 a_31098_4670.t2 DGND.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X72 a_2467_n30310.t15 a_35086_7130.t3 a_32057_n13616.t1 AVDD.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X73 a_2458_5328.t45 bias_p.t15 AVDD.t183 AVDD.t5 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X74 a_29757_7018.t0 Vop.t120 Vom_stg2 AVDD.t185 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1.16e+12p ps=8.58e+06u w=4e+06u l=1e+06u
X75 DGND bias_var_n.t8 Vfold_bot_m.t56 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X76 DGND bias_n.t9 a_1659_n4497.t17 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X77 AVDD.t682 AVDD.t680 AVDD.t681 AVDD.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X78 Vop.t71 casc_p.t87 a_2458_6128.t105 AVDD.t74 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X79 a_2467_n30310.t16 a_35086_7130.t4 a_32057_n13616.t2 AVDD.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X80 a_32059_n4497.t7 casc_n.t45 a_32059_n4755.t15 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X81 a_11259_n4497# casc_n.t46 casc_p.t69 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=2.32e+12p pd=1.832e+07u as=0p ps=0u w=2e+06u l=1e+06u
X82 a_2458_6128.t58 a_12760_n20342.t9 AVDD.t255 AVDD.t74 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X83 a_1657_n21342.t151 a_1560_n22142.t13 AVDD.t330 AVDD.t163 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X84 DGND bias_var_n.t9 a_2467_n30310.t22 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X85 AVDD.t815 level_shifter_up_0.xb_hv.t3 a_32057_n15000.t32 AVDD.t814 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X86 a_2458_5328.t46 bias_p.t16 AVDD.t184 AVDD.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X87 a_27936_n27260.t3 level_shifter_up_1.xb_hv.t1 a_23013_n25097.t2 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X88 a_12857_n14142.t3 a_12760_n20342.t10 AVDD.t256 AVDD.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X89 a_32057_n14142.t16 bias_p.t17 a_32057_n15000.t4 AVDD.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X90 a_2458_6128.t69 Vinm.t3 Vxm.t18 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X91 a_1659_n4497.t88 casc_n.t47 Vxm.t72 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X92 Vxp.t0 Vinp.t1 Vfold_bot_m.t0 AVDD.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X93 DGND bias_var_n.t10 Vfold_bot_m.t15 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X94 a_2458_5328.t1 Vinp.t2 Vxm.t1 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X95 a_1657_n21342.t150 a_1560_n22142.t14 AVDD.t331 AVDD.t168 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X96 a_1657_n21342.t149 a_1560_n22142.t15 AVDD.t332 AVDD.t159 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X97 a_2370_6628.t4 level_shifter_up_8.x_hv.t1 a_25696_11382.t15 AVDD.t3 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X98 Vop.t70 casc_p.t88 a_2458_6128.t104 AVDD.t85 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X99 a_11257_n14142.t3 bias_p.t18 AVDD.t268 AVDD.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X100 a_1657_n21342.t148 a_1560_n22142.t16 AVDD.t333 AVDD.t168 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X101 Vop.t69 casc_p.t89 a_2458_6128.t103 AVDD.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X102 Vop.t68 casc_p.t90 a_2458_6128.t102 AVDD.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X103 a_9060_4530.t3 a_12760_n20342.t11 AVDD.t257 AVDD.t93 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X104 a_1659_n4497.t87 casc_n.t48 Vxm.t73 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X105 a_2458_5328.t185 Vinp.t3 Vxm.t94 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X106 a_2458_6128.t57 a_12760_n20342.t12 AVDD.t258 AVDD.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X107 casc_n.t30 casc_n.t28 casc_n.t29 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X108 AVDD.t679 AVDD.t677 AVDD.t678 AVDD.t381 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X109 a_32057_n14142.t15 bias_p.t19 a_32057_n15000.t3 AVDD.t147 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X110 a_34883_n30483# a_34128_n30483# AVDD.t730 AVDD.t729 sky130_fd_pr__pfet_g5v0d10v5 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=500000u
X111 a_9060_4530.t4 Vinm.t4 a_9060_4172.t0 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X112 Vom.t74 casc_p.t91 a_2458_5328.t149 AVDD.t113 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X113 a_1657_n21342.t147 a_1560_n22142.t17 AVDD.t334 AVDD.t159 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X114 a_32059_n4497.t6 casc_n.t49 a_32059_n4755.t14 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X115 a_1657_n21342.t146 a_1560_n22142.t18 AVDD.t335 AVDD.t155 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X116 AVDD.t676 AVDD.t674 AVDD.t675 AVDD.t401 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X117 a_2467_n30310.t107 casc_n.t50 Vop.t108 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X118 AVDD.t673 AVDD.t671 AVDD.t672 AVDD.t46 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X119 a_1659_n4497.t86 casc_n.t51 Vxm.t66 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X120 a_32057_n8742.t2 bias_p.t20 a_32057_n9600.t5 AVDD.t48 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X121 a_32057_n14142.t14 bias_p.t21 a_32057_n15000.t11 AVDD.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X122 a_2458_6128.t56 a_12760_n20342.t13 AVDD.t259 AVDD.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X123 a_32057_n8742.t1 bias_p.t22 a_32057_n9600.t4 AVDD.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X124 casc_p.t3 casc_p.t2 a_11257_n8742.t11 AVDD.t93 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X125 a_2458_5328.t68 a_12760_n20342.t14 AVDD.t260 AVDD.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X126 DGND level_shifter_up_5.x_hv.t2 a_33659_n1551.t5 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X127 a_11257_n8742.t7 a_11160_n9542.t13 AVDD.t139 AVDD.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X128 a_2467_n30310.t106 casc_n.t52 Vop.t107 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X129 a_2458_5328.t97 a_34666_7130.t2 a_32059_n4755.t4 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X130 a_1657_n21342.t145 a_1560_n22142.t19 AVDD.t336 AVDD.t157 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X131 Vfold_bot_m.t103 casc_n.t53 Vom.t91 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X132 DGND bias_n.t10 a_1659_n4497.t18 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X133 Vop.t67 casc_p.t92 a_2458_6128.t118 AVDD.t148 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X134 a_2458_5328.t69 a_12760_n20342.t15 AVDD.t261 AVDD.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X135 Vop.t66 casc_p.t93 a_2458_6128.t117 AVDD.t5 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X136 a_1659_n4497.t85 casc_n.t54 Vxm.t87 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X137 DGND bias_n.t11 a_1659_n4497.t19 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X138 Vxp.t19 Vinm.t5 a_2467_n30310.t21 AVDD.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X139 a_1657_n21342.t144 a_1560_n22142.t20 AVDD.t337 AVDD.t203 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X140 a_23698_4566.t0 a_24364_11382.t0 DGND sky130_fd_pr__res_high_po_2p85 l=3.192e+07u
X141 a_2458_6128.t81 bias_p.t23 AVDD.t269 AVDD.t148 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X142 Vxp.t134 casc_p.t94 a_1657_n21342.t176 AVDD.t163 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X143 DGND bias_n.t12 a_1659_n4497.t28 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X144 DGND bias_n.t13 a_1659_n4497.t29 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X145 DGND DGND DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X146 Vom.t73 casc_p.t95 a_2458_5328.t148 AVDD.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X147 Vom.t72 casc_p.t96 a_2458_5328.t147 AVDD.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X148 a_9060_4530.t7 bias_p.t24 a_11257_n14142.t1 AVDD.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X149 DGND DGND DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X150 DGND DGND DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X151 a_29758_4670.t3 a_29758_4670.t2 DVDD.t7 DVDD.t6 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X152 a_30248_11527# trim[0].t0 AVDD.t740 AVDD.t739 sky130_fd_pr__pfet_g5v0d10v5 ad=1.45e+11p pd=1.58e+06u as=0p ps=0u w=500000u l=2e+06u
X153 a_32057_n14142.t13 bias_p.t25 a_32057_n15000.t10 AVDD.t48 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X154 a_2458_5328.t58 a_12760_n20342.t16 AVDD.t232 AVDD.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X155 Vxp.t139 Vinm.t6 a_2467_n30310.t66 AVDD.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X156 DGND DGND DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X157 AVDD.t670 AVDD.t668 AVDD.t669 AVDD.t366 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X158 a_32057_n14142.t12 bias_p.t26 a_32057_n15000.t9 AVDD.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X159 DGND DGND DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X160 DGND trim[2].t0 a_34648_11527# DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=500000u
X161 a_32057_n13616.t7 a_34666_7130.t3 Vfold_bot_m.t60 AVDD.t344 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X162 a_1657_n21342.t143 a_1560_n22142.t21 AVDD.t338 AVDD.t168 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X163 a_32059_n3351.t15 bias_n.t14 a_32059_n4497.t12 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X164 DGND bias_var_n.t11 a_2467_n30310.t23 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X165 DGND en.t0 a_32299_n29829# DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=500000u
X166 DGND bias_n.t15 a_12859_n4209# DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.16e+12p ps=9.16e+06u w=2e+06u l=4e+06u
X167 DGND bias_n.t16 a_12859_n2697# DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=2.32e+12p ps=1.832e+07u w=2e+06u l=4e+06u
X168 a_12857_n15942.t3 a_1560_n22142.t22 AVDD.t840 AVDD.t93 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X169 Vop.t65 casc_p.t97 a_2458_6128.t116 AVDD.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X170 AVDD.t667 AVDD.t665 AVDD.t666 AVDD.t374 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X171 a_2458_6128.t66 bias_p.t27 AVDD.t50 AVDD.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X172 a_1659_n4497.t84 casc_n.t55 Vxm.t88 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X173 DGND level_shifter_up_0.x_hv.t2 a_32059_n3351.t0 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X174 a_1659_n4497.t83 casc_n.t56 Vxm.t89 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X175 a_23032_4566.t5 level_shifter_up_8.xb_hv.t3 a_2370_6628.t3 AVDD.t38 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X176 a_1657_n21342.t142 a_1560_n22142.t23 AVDD.t841 AVDD.t166 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X177 Vop.t64 casc_p.t98 a_2458_6128.t115 AVDD.t113 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X178 AVDD.t664 AVDD.t662 AVDD.t663 AVDD.t111 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X179 DGND bias_var_n.t12 a_2467_n30310.t24 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X180 a_2458_6128.t188 Vinm.t7 Vxm.t45 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X181 casc_n.t27 casc_n.t25 casc_n.t26 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X182 AVDD.t1 level_shifter_up_3.x_hv.t3 level_shifter_up_3.xb_hv.t0 AVDD.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X183 Vxp.t140 Vinm.t8 a_2467_n30310.t67 AVDD.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X184 a_1657_n21342.t141 a_1560_n22142.t24 AVDD.t842 AVDD.t155 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X185 a_2458_6128.t55 a_12760_n20342.t17 AVDD.t233 AVDD.t113 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X186 DGND level_shifter_up_4.xb_hv.t3 bias_n.t1 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X187 Vout.t0 a_35086_7130.t5 DVDD.t13 DVDD.t12 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X188 a_2458_6128.t82 Vinm.t9 Vxm.t32 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X189 a_32057_n15000.t31 level_shifter_up_0.xb_hv.t4 AVDD.t817 AVDD.t816 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X190 Vxp.t133 casc_p.t99 a_1657_n21342.t177 AVDD.t196 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X191 a_32057_n17742.t11 a_1560_n22142.t25 AVDD.t843 AVDD.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X192 DGND bias_var_n.t13 Vfold_bot_m.t58 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X193 AVDD.t819 level_shifter_up_0.xb_hv.t5 level_shifter_up_0.x_hv.t1 AVDD.t818 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X194 DGND DGND DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X195 DGND DGND DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X196 Vxp.t132 casc_p.t100 a_1657_n21342.t178 AVDD.t203 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X197 DGND a_31003_11527# level_shifter_up_6.xb_hv DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X198 a_2467_n30310.t105 casc_n.t57 Vop.t106 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X199 a_1657_n21342.t140 a_1560_n22142.t26 AVDD.t844 AVDD.t157 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X200 Vfold_bot_m.t102 casc_n.t58 Vom.t90 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X201 Vfold_bot_m.t101 casc_n.t59 Vom.t89 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X202 a_2458_6128.t83 Vinm.t10 Vxm.t33 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X203 a_1657_n21342.t139 a_1560_n22142.t27 AVDD.t845 AVDD.t194 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X204 Vop.t63 casc_p.t101 a_2458_6128.t114 AVDD.t125 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X205 a_2467_n30310.t104 casc_n.t60 Vop.t100 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X206 a_2458_5328.t59 a_12760_n20342.t18 AVDD.t234 AVDD.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X207 a_33659_n1551.t1 bias_n.t17 a_33659_n2697.t5 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X208 Vom.t71 casc_p.t102 a_2458_5328.t146 AVDD.t15 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X209 Vop.t62 casc_p.t103 a_2458_6128.t131 AVDD.t5 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X210 a_2458_6128.t54 a_12760_n20342.t19 AVDD.t235 AVDD.t103 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X211 a_32057_n14142.t11 bias_p.t28 a_32057_n15000.t17 AVDD.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X212 DGND bias_var_n.t14 Vfold_bot_m.t59 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X213 a_2467_n29152.t4 a_2370_n29452.t9 Vfold_bot_m.t16 AVDD.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X214 DGND a_12857_n19016.t8 a_32059_n897.t0 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X215 a_1659_n4497.t82 casc_n.t61 Vxm.t90 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X216 a_2458_5328.t12 bias_p.t29 AVDD.t51 AVDD.t15 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X217 a_1657_n21342.t138 a_1560_n22142.t28 AVDD.t846 AVDD.t196 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X218 Vxp.t131 casc_p.t104 a_1657_n21342.t179 AVDD.t163 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X219 a_29757_7018.t2 bias_stg2.t5 AVDD.t762 AVDD.t709 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X220 DGND Vom.t120 Vfold_bot_m.t52 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X221 Vom.t70 casc_p.t105 a_2458_5328.t145 AVDD.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X222 a_1657_n21342.t137 a_1560_n22142.t29 AVDD.t847 AVDD.t194 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X223 a_11160_n9542.t1 a_11160_n9542.t0 a_11257_n8742.t4 AVDD.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X224 Vfold_bot_m.t100 casc_n.t62 Vom.t88 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X225 AVDD.t661 AVDD.t659 AVDD.t660 AVDD.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X226 Vop.t61 casc_p.t106 a_2458_6128.t130 AVDD.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X227 a_32057_n14142.t10 bias_p.t30 a_32057_n15000.t16 AVDD.t48 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X228 AVDD.t658 AVDD.t656 AVDD.t657 AVDD.t370 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X229 a_23013_n25097.t3 level_shifter_up_1.xb_hv.t2 a_27936_n27260.t2 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X230 casc_p.t60 casc_p.t58 casc_p.t59 AVDD.t93 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X231 Vop.t60 casc_p.t107 a_2458_6128.t129 AVDD.t74 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X232 Vxp.t141 Vinp.t4 Vfold_bot_m.t105 AVDD.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X233 a_23013_n31913# a_23679_n25097# DGND sky130_fd_pr__res_high_po_2p85 l=3.192e+07u
X234 Vxp.t142 Vinp.t5 Vfold_bot_m.t106 AVDD.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X235 a_1657_n21342.t136 a_1560_n22142.t30 AVDD.t848 AVDD.t161 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X236 DGND DGND DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X237 DGND level_shifter_up_0.x_hv.t3 a_32059_n3351.t5 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X238 Vfold_bot_m.t99 casc_n.t63 Vom.t87 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X239 a_2458_6128.t192 a_2370_7428.t8 a_2458_6570.t12 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X240 a_14459_n2697# casc_n.t64 a_1560_n22142.t8 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=2.32e+12p pd=1.832e+07u as=0p ps=0u w=2e+06u l=1e+06u
X241 DGND bias_n.t18 a_1659_n4497.t5 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X242 Vfold_bot_m.t98 casc_n.t65 Vom.t86 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X243 a_2458_5328.t3 bias_p.t31 AVDD.t16 AVDD.t15 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X244 a_2458_6128.t53 a_12760_n20342.t20 AVDD.t236 AVDD.t103 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X245 a_2458_5328.t4 bias_p.t32 AVDD.t17 AVDD.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X246 a_12857_n17742.t3 a_1560_n22142.t31 AVDD.t849 AVDD.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X247 a_2458_6128.t3 bias_p.t33 AVDD.t18 AVDD.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X248 a_2458_5328.t60 a_12760_n20342.t21 AVDD.t237 AVDD.t66 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X249 DGND bias_n.t19 a_1659_n4497.t6 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X250 a_34648_11527# trim[2].t1 DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X251 Vxp.t130 casc_p.t108 a_1657_n21342.t180 AVDD.t155 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X252 a_1659_n4497.t81 casc_n.t66 Vxm.t63 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X253 a_1657_n21342.t135 a_1560_n22142.t32 AVDD.t850 AVDD.t166 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X254 Vxp.t143 Vinp.t6 Vfold_bot_m.t107 AVDD.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X255 a_32057_n13616.t28 casc_p.t109 a_32057_n14142.t35 AVDD.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X256 AVDD.t655 AVDD.t653 AVDD.t654 AVDD.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X257 a_12857_n14142.t2 a_12760_n20342.t22 AVDD.t238 AVDD.t111 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X258 Vop.t59 casc_p.t110 a_2458_6128.t128 AVDD.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X259 a_2458_5328.t61 a_12760_n20342.t23 AVDD.t239 AVDD.t66 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X260 Vxp.t20 Vinp.t7 Vfold_bot_m.t20 AVDD.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X261 Vxp.t129 casc_p.t111 a_1657_n21342.t181 AVDD.t157 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X262 DGND bias_n.t20 a_1659_n4497.t42 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X263 a_2458_6128.t4 bias_p.t34 AVDD.t19 AVDD.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X264 a_32059_2049.t3 level_shifter_up_7.x_hv.t1 DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X265 a_32057_n17742.t10 a_1560_n22142.t33 AVDD.t851 AVDD.t147 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X266 DGND DGND DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X267 Vxp.t128 casc_p.t112 a_1657_n21342.t8 AVDD.t203 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X268 a_9060_4530.t2 a_12760_n20342.t24 AVDD.t240 AVDD.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X269 DGND a_12857_n19016.t6 a_12857_n19016.t7 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X270 a_1657_n21342.t134 a_1560_n22142.t34 AVDD.t852 AVDD.t159 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X271 a_30248_11527# trim[0].t1 DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=500000u
X272 a_1657_n21342.t133 a_1560_n22142.t35 AVDD.t853 AVDD.t194 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X273 a_1657_n21342.t132 a_1560_n22142.t36 AVDD.t854 AVDD.t203 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X274 a_2467_n30310.t103 casc_n.t67 Vop.t99 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X275 AVDD.t276 hyst[1].t0 a_34499_n29829# AVDD.t275 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1.45e+11p ps=1.58e+06u w=500000u l=2e+06u
X276 a_32057_n14142.t9 bias_p.t35 a_32057_n15000.t15 AVDD.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X277 a_2458_6128.t52 a_12760_n20342.t25 AVDD.t241 AVDD.t103 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X278 a_32057_n14142.t8 bias_p.t36 a_32057_n15000.t14 AVDD.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X279 a_12859_2049# ibias.t0 ibias.t1 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=1.16e+12p pd=9.16e+06u as=0p ps=0u w=2e+06u l=4e+06u
X280 a_35086_7130.t1 a_34666_7130.t4 DGND.t518 DGND.t517 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X281 casc_p.t57 casc_p.t55 casc_p.t56 AVDD.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X282 a_2458_6128.t84 Vinm.t11 Vxm.t34 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X283 a_1657_n21342.t131 a_1560_n22142.t37 AVDD.t855 AVDD.t196 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X284 a_2370_7428.t3 level_shifter_up_8.xb_hv.t4 a_25696_11382.t4 AVDD.t716 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X285 a_1657_n21342.t130 a_1560_n22142.t38 AVDD.t856 AVDD.t172 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X286 a_24345_n31913# a_25011_n25097# DGND sky130_fd_pr__res_high_po_2p85 l=3.192e+07u
X287 DGND Vom.t121 Vfold_bot_m.t51 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X288 DGND Vom.t122 Vfold_bot_m.t50 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X289 a_2458_5328.t40 Vinp.t8 Vxm.t25 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X290 a_34883_n30483# a_34128_n30483# DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X291 DGND bias_var_n.t15 a_2467_n30310.t62 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X292 DGND bias_var_n.t16 a_2467_n30310.t63 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X293 Vop.t58 casc_p.t113 a_2458_6128.t127 AVDD.t148 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X294 AVDD.t652 AVDD.t650 AVDD.t651 AVDD.t366 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X295 a_2458_5328.t62 a_12760_n20342.t26 AVDD.t242 AVDD.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X296 a_32059_n4755.t23 a_35086_7130.t6 a_2458_6128.t64 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X297 DGND bias_n.t21 a_1659_n4497.t43 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X298 DGND bias_var_n.t17 Vfold_bot_m.t3 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X299 DGND a_36699_n29829# level_shifter_up_5.x_hv.t1 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X300 a_1659_n4497.t80 casc_n.t68 Vxm.t64 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X301 AVDD.t649 AVDD.t647 AVDD.t648 AVDD.t370 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X302 DGND bias_n.t22 a_1659_n4497.t44 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X303 a_32059_n4755.t3 a_34666_7130.t5 a_2458_5328.t96 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X304 a_2467_n30310.t102 casc_n.t69 Vop.t98 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X305 DGND bias_var_n.t18 a_2467_n30310.t4 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X306 a_1560_n22142.t0 casc_p.t114 a_12857_n14142.t7 AVDD.t93 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X307 Vxp.t25 Vinm.t12 a_2467_n30310.t25 AVDD.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X308 a_12760_n20342.t0 casc_p.t115 a_9060_4530.t11 AVDD.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X309 Vop.t57 casc_p.t116 a_2458_6128.t126 AVDD.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X310 a_1657_n21342.t129 a_1560_n22142.t39 AVDD.t857 AVDD.t161 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X311 AVDD.t646 AVDD.t644 AVDD.t645 AVDD.t374 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X312 Vop.t56 casc_p.t117 a_2458_6128.t101 AVDD.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X313 Vxp.t127 casc_p.t118 a_1657_n21342.t9 AVDD.t166 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X314 Vxp.t126 casc_p.t119 a_1657_n21342.t10 AVDD.t208 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X315 a_2467_n30310.t101 casc_n.t70 Vop.t97 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X316 a_2467_n30310.t100 casc_n.t71 Vop.t96 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X317 a_32057_n13616.t0 a_35086_7130.t7 a_2467_n30310.t3 AVDD.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X318 DGND hyst[1].t1 a_34499_n29829# DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=500000u
X319 casc_p.t54 casc_p.t52 casc_p.t53 AVDD.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X320 a_32057_n17742.t9 a_1560_n22142.t40 AVDD.t787 AVDD.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X321 AVDD.t839 a_32299_n29829# a_31859_n29829# AVDD.t838 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X322 a_1657_n21342.t128 a_1560_n22142.t41 AVDD.t788 AVDD.t208 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X323 Vxp.t125 casc_p.t120 a_1657_n21342.t11 AVDD.t155 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X324 DGND DGND DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X325 a_2467_n30310.t99 casc_n.t72 Vop.t85 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X326 a_1657_n21342.t127 a_1560_n22142.t42 AVDD.t789 AVDD.t168 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X327 a_2458_5328.t63 a_12760_n20342.t27 AVDD.t243 AVDD.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X328 a_32057_n13616.t27 casc_p.t121 a_32057_n14142.t34 AVDD.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X329 casc_n.t24 casc_n.t22 casc_n.t23 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X330 a_32057_n13616.t26 casc_p.t122 a_32057_n14142.t33 AVDD.t147 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X331 DGND bias_var_n.t19 Vfold_bot_m.t4 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X332 a_2458_5328.t64 a_12760_n20342.t28 AVDD.t244 AVDD.t66 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X333 Vxp.t26 Vinm.t13 a_2467_n30310.t26 AVDD.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X334 Vxp.t124 casc_p.t123 a_1657_n21342.t12 AVDD.t157 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X335 DGND bias_var_n.t20 a_2467_n30310.t5 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X336 a_2458_6128.t181 a_2370_7428.t9 a_2458_6570.t3 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X337 Vxp.t123 casc_p.t124 a_1657_n21342.t13 AVDD.t159 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X338 AVDD.t643 AVDD.t641 AVDD.t642 AVDD.t381 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X339 AVDD.t761 bias_stg2.t3 bias_stg2.t4 AVDD.t760 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X340 Vom.t69 casc_p.t125 a_2458_5328.t144 AVDD.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X341 a_32059_903.t3 casc_n.t73 a_23032_4566.t14 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X342 DGND bias_n.t23 a_1659_n4497.t45 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X343 Vop.t55 casc_p.t126 a_2458_6128.t100 AVDD.t103 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X344 Vom.t68 casc_p.t127 a_2458_5328.t143 AVDD.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X345 a_2458_5328.t41 Vinp.t9 Vxm.t26 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X346 a_12857_n15942.t2 a_1560_n22142.t43 AVDD.t790 AVDD.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X347 Vop.t54 casc_p.t128 a_2458_6128.t99 AVDD.t85 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X348 Vop.t53 casc_p.t129 a_2458_6128.t98 AVDD.t113 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X349 a_32057_n22200.t3 level_shifter_up_2.xb_hv.t2 AVDD.t88 AVDD.t87 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X350 AVDD.t821 level_shifter_up_0.xb_hv.t6 a_32057_n15000.t30 AVDD.t820 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X351 AVDD.t640 AVDD.t638 AVDD.t639 AVDD.t394 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X352 a_27936_n27260.t1 level_shifter_up_1.xb_hv.t3 a_23013_n25097.t23 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X353 DGND Vom.t123 a_2467_n30310.t57 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X354 a_32057_n17742.t8 a_1560_n22142.t44 AVDD.t791 AVDD.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X355 a_23013_n25097.t4 level_shifter_up_3.xb_hv.t2 a_2370_n29452.t0 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X356 Vxp.t27 Vinm.t14 a_2467_n30310.t27 AVDD.t46 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X357 casc_p.t51 casc_p.t49 casc_p.t50 AVDD.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X358 Vxp.t21 Vinp.t10 Vfold_bot_m.t21 AVDD.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X359 DGND bias_var_n.t21 a_2467_n30310.t19 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X360 a_1657_n21342.t126 a_1560_n22142.t45 AVDD.t792 AVDD.t172 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X361 a_34128_n30483# trim[4].t0 AVDD.t263 AVDD.t262 sky130_fd_pr__pfet_g5v0d10v5 ad=1.45e+11p pd=1.58e+06u as=0p ps=0u w=500000u l=2e+06u
X362 AVDD.t637 AVDD.t635 AVDD.t636 AVDD.t370 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X363 Vop.t52 casc_p.t130 a_2458_6128.t97 AVDD.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X364 DGND DGND DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X365 a_2458_5328.t65 a_12760_n20342.t29 AVDD.t245 AVDD.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X366 a_2458_5328.t66 a_12760_n20342.t30 AVDD.t246 AVDD.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X367 a_32059_n3351.t14 bias_n.t24 a_32059_n4497.t11 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X368 Vom.t67 casc_p.t131 a_2458_5328.t142 AVDD.t5 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X369 DGND bias_var_n.t22 Vfold_bot_m.t13 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X370 DGND bias_n.t25 a_11259_n4497# DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X371 DGND a_32683_n30483# level_shifter_up_3.xb_hv.t1 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X372 Vxp.t122 casc_p.t132 a_1657_n21342.t14 AVDD.t161 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X373 Vfold_bot_m.t97 casc_n.t74 Vom.t85 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X374 a_1659_n4497.t79 casc_n.t75 Vxm.t65 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X375 a_2458_5328.t5 bias_p.t37 AVDD.t22 AVDD.t5 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X376 Vxp.t121 casc_p.t133 a_1657_n21342.t15 AVDD.t163 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X377 Vop.t51 casc_p.t134 a_2458_6128.t96 AVDD.t74 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X378 DGND bias_n.t26 a_1659_n4497.t35 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X379 Vom.t66 casc_p.t135 a_2458_5328.t141 AVDD.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X380 Vop.t50 casc_p.t136 a_2458_6128.t95 AVDD.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X381 a_2458_6128.t51 a_12760_n20342.t31 AVDD.t217 AVDD.t85 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X382 a_1560_n22142.t1 casc_p.t137 a_12857_n15942.t7 AVDD.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X383 a_1657_n21342.t125 a_1560_n22142.t46 AVDD.t793 AVDD.t163 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X384 a_32057_n13616.t31 casc_p.t138 a_32057_n14142.t32 AVDD.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X385 a_2458_6128.t78 Vinm.t15 Vxm.t28 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X386 a_23013_n25097.t24 level_shifter_up_1.xb_hv.t4 a_27936_n27260.t0 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X387 a_2458_5328.t70 bias_p.t38 AVDD.t272 AVDD.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X388 a_12857_n19542.t3 a_12760_n20342.t32 AVDD.t218 AVDD.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X389 DGND bias_n.t27 casc_n.t3 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X390 AVDD.t634 AVDD.t632 AVDD.t633 AVDD.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X391 Vxp.t120 casc_p.t139 a_1657_n21342.t16 AVDD.t166 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X392 a_32057_n17742.t7 a_1560_n22142.t47 AVDD.t794 AVDD.t48 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X393 Vxp.t119 casc_p.t140 a_1657_n21342.t17 AVDD.t168 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X394 level_shifter_up_7.x_hv a_32448_11527# DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X395 casc_p.t48 casc_p.t46 casc_p.t47 AVDD.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X396 DGND bias_n.t6 bias_n.t5 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X397 Vom.t65 casc_p.t141 a_2458_5328.t140 AVDD.t66 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X398 a_1657_n21342.t124 a_1560_n22142.t48 AVDD.t795 AVDD.t208 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X399 AVDD.t631 AVDD.t629 AVDD.t630 AVDD.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X400 DGND DGND DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X401 Vfold_bot_m.t96 casc_n.t76 Vom.t84 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X402 a_2458_5328.t52 a_12760_n20342.t33 AVDD.t219 AVDD.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X403 a_14459_n4497# casc_n.t77 a_14459_n4755.t0 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=1.16e+12p pd=9.16e+06u as=0p ps=0u w=2e+06u l=1e+06u
X404 AVDD.t628 AVDD.t626 AVDD.t627 AVDD.t401 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X405 a_2467_n29152.t17 casc_p.t142 a_32057_n17742.t23 AVDD.t147 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X406 a_2458_5328.t53 a_12760_n20342.t34 AVDD.t220 AVDD.t68 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X407 Vxp.t145 Vinp.t11 Vfold_bot_m.t111 AVDD.t46 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X408 Vxp.t28 Vinm.t16 a_2467_n30310.t29 AVDD.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X409 casc_p.t45 casc_p.t43 casc_p.t44 AVDD.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X410 a_2467_n29152.t18 a_2370_n28652.t8 a_2467_n30310.t68 AVDD.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X411 a_32059_n3351.t13 bias_n.t28 a_32059_n4497.t10 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X412 DGND bias_n.t29 a_11259_n2697# DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=2.32e+12p ps=1.832e+07u w=2e+06u l=4e+06u
X413 a_32059_903.t2 casc_n.t78 a_23032_4566.t13 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X414 a_32057_n21342.t7 bias_p.t39 a_32057_n22200.t5 AVDD.t147 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X415 a_2458_6128.t79 Vinm.t17 Vxm.t29 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X416 Vxp.t118 casc_p.t143 a_1657_n21342.t49 AVDD.t159 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X417 AVDD.t625 AVDD.t623 AVDD.t624 AVDD.t381 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X418 Vop.t49 casc_p.t144 a_2458_6128.t173 AVDD.t103 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X419 a_1657_n21342.t123 a_1560_n22142.t49 AVDD.t796 AVDD.t159 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X420 a_32057_n13616.t30 casc_p.t145 a_32057_n14142.t31 AVDD.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X421 a_12857_n17742.t2 a_1560_n22142.t50 AVDD.t797 AVDD.t111 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X422 Vxp.t117 casc_p.t146 a_1657_n21342.t50 AVDD.t172 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X423 a_35259_903# casc_n.t79 a_23032_4566.t10 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=2.32e+12p pd=1.832e+07u as=0p ps=0u w=2e+06u l=1e+06u
X424 DGND a_34499_n29829# a_34059_n29829# DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X425 a_32057_n15000.t29 level_shifter_up_0.xb_hv.t7 AVDD.t280 AVDD.t279 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X426 Vom.t64 casc_p.t147 a_2458_5328.t139 AVDD.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X427 Vxp.t116 casc_p.t148 a_1657_n21342.t51 AVDD.t203 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X428 Vop.t48 casc_p.t149 a_2458_6128.t172 AVDD.t148 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X429 a_32057_n9600.t10 level_shifter_up_5.xb_hv.t3 AVDD.t352 AVDD.t351 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X430 a_1657_n21342.t122 a_1560_n22142.t51 AVDD.t798 AVDD.t194 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X431 AVDD.t622 AVDD.t620 AVDD.t621 AVDD.t370 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X432 a_33659_n2697.t2 casc_n.t80 a_32059_n4755.t13 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X433 a_2467_n30310.t98 casc_n.t81 Vop.t84 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X434 a_29757_7018.t1 Vom.t124 Vop_stg2 AVDD.t192 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1.16e+12p ps=8.58e+06u w=4e+06u l=1e+06u
X435 a_32057_n17742.t6 a_1560_n22142.t52 AVDD.t799 AVDD.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X436 DGND bias_var_n.t23 a_2467_n30310.t20 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X437 a_2458_6128.t67 Vinm.t18 Vxm.t11 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X438 DGND DGND DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X439 a_32057_n15000.t28 level_shifter_up_0.xb_hv.t8 AVDD.t282 AVDD.t281 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X440 Vxp.t115 casc_p.t150 a_1657_n21342.t52 AVDD.t161 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X441 DGND DGND DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X442 a_1657_n21342.t121 a_1560_n22142.t53 AVDD.t800 AVDD.t196 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X443 DGND bias_var_n.t24 Vfold_bot_m.t14 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X444 a_32057_n13616.t29 casc_p.t151 a_32057_n14142.t30 AVDD.t48 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X445 a_31098_4670.t6 level_shifter_up_4.xb_hv.t4 DGND.t474 DGND.t473 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X446 Vfold_bot_m.t95 casc_n.t82 Vom.t83 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X447 AVDD.t835 bias_stg2.t6 a_29757_7018.t3 AVDD.t760 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X448 a_2458_6128.t50 a_12760_n20342.t35 AVDD.t221 AVDD.t85 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X449 a_32057_n13616.t15 casc_p.t152 a_32057_n8742.t9 AVDD.t147 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X450 a_2467_n29152.t16 casc_p.t153 a_32057_n17742.t22 AVDD.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X451 Vom.t63 casc_p.t154 a_2458_5328.t177 AVDD.t68 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X452 a_32057_n13616.t14 casc_p.t155 a_32057_n8742.t8 AVDD.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X453 level_shifter_up_0.xb_hv.t1 a_34059_n29829# DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X454 a_32057_n21342.t6 bias_p.t40 a_32057_n22200.t4 AVDD.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X455 Vxp.t114 casc_p.t156 a_1657_n21342.t53 AVDD.t168 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X456 Vom.t62 casc_p.t157 a_2458_5328.t176 AVDD.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X457 AVDD.t216 level_shifter_up_7.x_hv.t2 level_shifter_up_7.xb_hv AVDD.t215 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X458 a_34499_n29829# hyst[1].t2 DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X459 DGND bias_n.t30 a_1659_n4497.t27 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X460 a_32059_2049.t7 bias_n.t31 a_32059_903.t7 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X461 bias_var_n.t5 casc_p.t158 a_12857_n17742.t7 AVDD.t93 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X462 Vom.t61 casc_p.t159 a_2458_5328.t175 AVDD.t66 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X463 DGND DGND DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X464 a_1657_n21342.t120 a_1560_n22142.t54 AVDD.t801 AVDD.t168 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X465 DGND level_shifter_up_0.x_hv.t4 a_32059_n3351.t6 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X466 AVDD.t619 AVDD.t617 AVDD.t618 AVDD.t93 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X467 DGND Vom.t125 Vfold_bot_m.t49 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X468 AVDD.t616 AVDD.t614 AVDD.t615 AVDD.t401 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X469 a_2370_n29452.t3 level_shifter_up_3.xb_hv.t3 a_23013_n25097.t5 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X470 a_2458_5328.t54 a_12760_n20342.t36 AVDD.t222 AVDD.t68 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X471 a_23013_n31913# a_23013_n25097.t22 DGND sky130_fd_pr__res_high_po_2p85 l=3.192e+07u
X472 a_1560_n22142.t6 casc_p.t160 a_12857_n14142.t6 AVDD.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X473 a_12760_n20342.t3 casc_p.t161 a_9060_4530.t10 AVDD.t111 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X474 a_31003_11527# a_30248_11527# AVDD.t807 AVDD.t806 sky130_fd_pr__pfet_g5v0d10v5 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=500000u
X475 DGND DGND DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X476 Vxp.t113 casc_p.t162 a_1657_n21342.t54 AVDD.t155 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X477 Vop.t47 casc_p.t163 a_2458_6128.t171 AVDD.t113 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X478 AVDD.t613 AVDD.t611 AVDD.t612 AVDD.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X479 a_2458_6128.t68 Vinm.t19 Vxm.t12 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X480 a_2467_n29152.t15 casc_p.t164 a_32057_n17742.t21 AVDD.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X481 a_32057_n13616.t10 casc_p.t165 a_32057_n14142.t29 AVDD.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X482 a_2458_6128.t49 a_12760_n20342.t37 AVDD.t223 AVDD.t125 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X483 a_32059_903.t1 casc_n.t83 a_23032_4566.t12 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X484 a_1657_n21342.t119 a_1560_n22142.t55 AVDD.t802 AVDD.t155 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X485 AVDD.t610 AVDD.t608 AVDD.t609 AVDD.t366 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X486 DGND Vom.t126 a_2467_n30310.t56 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X487 AVDD.t98 level_shifter_up_2.xb_hv.t3 a_32057_n22200.t2 AVDD.t97 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X488 DGND bias_var_n.t25 Vfold_bot_m.t33 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X489 a_32057_n13616.t3 a_34666_7130.t6 Vfold_bot_m.t53 AVDD.t344 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X490 a_32057_n21342.t5 bias_p.t41 a_32057_n22200.t11 AVDD.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X491 res_p_bot.t5 level_shifter_up_3.xb_hv.t4 a_2370_n28652.t4 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X492 Vxp.t112 casc_p.t166 a_1657_n21342.t55 AVDD.t157 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X493 DGND bias_n.t32 a_1659_n4497.t12 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X494 Vxp.t111 casc_p.t167 a_1657_n21342.t56 AVDD.t172 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X495 Vxp.t110 casc_p.t168 a_1657_n21342.t57 AVDD.t194 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X496 a_2458_5328.t190 Vinp.t12 Vxm.t98 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X497 level_shifter_up_1.x_hv level_shifter_up_1.xb_hv.t5 AVDD.t768 AVDD.t767 sky130_fd_pr__pfet_g5v0d10v5 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=500000u
X498 DGND bias_n.t33 a_1659_n4497.t13 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X499 a_31098_4670.t0 a_29758_4670.t5 DVDD.t5 DVDD.t4 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X500 Vom.t60 casc_p.t169 a_2458_5328.t174 AVDD.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X501 a_1657_n21342.t118 a_1560_n22142.t56 AVDD.t803 AVDD.t157 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X502 a_32057_n13616.t9 casc_p.t170 a_32057_n14142.t28 AVDD.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X503 AVDD.t607 AVDD.t605 AVDD.t606 AVDD.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X504 DGND bias_n.t34 a_1659_n4497.t14 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X505 Vxp.t16 Vinm.t20 a_2467_n30310.t12 AVDD.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X506 a_2458_5328.t55 a_12760_n20342.t38 AVDD.t224 AVDD.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X507 a_23013_n25097.t6 level_shifter_up_3.xb_hv.t5 a_2370_n29452.t4 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X508 Vxp.t109 casc_p.t171 a_1657_n21342.t58 AVDD.t196 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X509 Vop.t46 casc_p.t172 a_2458_6128.t170 AVDD.t85 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X510 casc_p.t42 casc_p.t40 casc_p.t41 AVDD.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X511 a_2467_n29152.t3 a_2370_n29452.t10 Vfold_bot_m.t17 AVDD.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X512 a_2467_n29152.t14 casc_p.t173 a_32057_n17742.t20 AVDD.t48 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X513 Vfold_bot_m.t94 casc_n.t84 Vom.t82 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X514 a_2458_5328.t8 a_2370_6628.t9 a_2458_6570.t0 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X515 a_2458_6128.t48 a_12760_n20342.t39 AVDD.t225 AVDD.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X516 a_11257_n21342# bias_p.t42 AVDD.t273 AVDD.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=2.32e+12p pd=1.832e+07u as=0p ps=0u w=2e+06u l=4e+06u
X517 DGND Vom.t127 a_2467_n30310.t55 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X518 a_2458_5328.t56 a_12760_n20342.t40 AVDD.t226 AVDD.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X519 DGND bias_var_n.t26 Vfold_bot_m.t34 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X520 a_32057_n21342.t4 bias_p.t43 a_32057_n22200.t10 AVDD.t48 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X521 a_1657_n21342.t117 a_1560_n22142.t57 AVDD.t804 AVDD.t163 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X522 a_32057_n13616.t4 a_34666_7130.t7 Vfold_bot_m.t54 AVDD.t344 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X523 AVDD.t284 level_shifter_up_0.xb_hv.t9 a_32057_n15000.t27 AVDD.t283 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X524 a_2458_6128.t65 a_35086_7130.t8 a_32059_n4755.t22 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X525 a_2458_6128.t73 Vinm.t21 Vxm.t22 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X526 a_2458_6128.t74 Vinm.t22 Vxm.t23 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X527 a_1659_n4497.t78 casc_n.t85 Vxm.t86 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X528 Vom.t59 casc_p.t174 a_2458_5328.t173 AVDD.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X529 AVDD.t604 AVDD.t602 AVDD.t603 AVDD.t401 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X530 a_23032_4566.t3 a_23032_11382.t0 DGND sky130_fd_pr__res_high_po_2p85 l=3.192e+07u
X531 a_2458_5328.t191 Vinp.t13 Vxm.t99 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X532 a_12857_n19016.t1 casc_p.t175 a_12857_n19542.t7 AVDD.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X533 Vom.t58 casc_p.t176 a_2458_5328.t172 AVDD.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X534 a_2458_5328.t192 Vinp.t14 Vxm.t100 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X535 a_2458_5328.t91 a_34666_7130.t8 a_32059_n4755.t2 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X536 a_2458_5328.t71 bias_p.t44 AVDD.t274 AVDD.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X537 DGND DGND DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X538 Vxp.t108 casc_p.t177 a_1657_n21342.t28 AVDD.t166 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X539 AVDD.t601 AVDD.t599 AVDD.t600 AVDD.t394 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X540 DGND bias_n.t35 a_1659_n4497.t15 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X541 casc_p.t39 casc_p.t37 casc_p.t38 AVDD.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X542 a_1560_n22142.t4 casc_p.t178 a_12857_n15942.t6 AVDD.t111 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X543 DGND bias_var_n.t27 Vfold_bot_m.t35 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X544 a_1657_n21342.t116 a_1560_n22142.t58 AVDD.t769 AVDD.t166 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X545 a_2370_7428.t2 level_shifter_up_8.xb_hv.t5 a_25696_11382.t6 AVDD.t717 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X546 a_32057_n8742.t0 bias_p.t45 a_32057_n9600.t3 AVDD.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X547 AVDD.t598 AVDD.t596 AVDD.t597 AVDD.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X548 a_2458_6128.t47 a_12760_n20342.t41 AVDD.t227 AVDD.t125 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X549 a_1657_n21342.t115 a_1560_n22142.t59 AVDD.t770 AVDD.t208 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X550 a_1657_n21342.t114 a_1560_n22142.t60 AVDD.t771 AVDD.t203 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X551 DGND bias_n.t36 a_1659_n4497.t2 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X552 DGND trim[1].t0 a_32448_11527# DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=500000u
X553 a_12857_n19542.t2 a_12760_n20342.t42 AVDD.t228 AVDD.t111 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X554 a_2458_6128.t193 bias_p.t46 AVDD.t822 AVDD.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X555 Vfold_bot_m.t93 casc_n.t86 Vom.t81 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X556 a_1659_n4497.t77 casc_n.t87 Vxm.t79 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X557 a_32059_n897.t10 casc_n.t88 a_2458_6570.t10 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X558 DGND bias_var_n.t28 a_2467_n30310.t34 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X559 a_2458_6128.t46 a_12760_n20342.t43 AVDD.t229 AVDD.t125 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X560 a_2467_n30310.t97 casc_n.t89 Vop.t83 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X561 a_23013_n25097.t16 casc_p.t179 a_32057_n21342.t15 AVDD.t147 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X562 casc_n.t2 ibias.t2 AVDD.t343 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X563 a_27926_9740.t3 level_shifter_up_6.x_hv.t1 a_25696_11382.t0 AVDD.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X564 Vxp.t107 casc_p.t180 a_1657_n21342.t29 AVDD.t159 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X565 Vxp.t106 casc_p.t181 a_1657_n21342.t30 AVDD.t194 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X566 AVDD.t595 AVDD.t593 AVDD.t594 AVDD.t381 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X567 Vxp.t105 casc_p.t182 a_1657_n21342.t31 AVDD.t203 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X568 a_2467_n29152.t13 casc_p.t183 a_32057_n17742.t19 AVDD.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X569 a_2458_5328.t57 a_12760_n20342.t44 AVDD.t230 AVDD.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X570 Vop.t45 casc_p.t184 a_2458_6128.t169 AVDD.t103 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X571 a_1657_n21342.t113 a_1560_n22142.t61 AVDD.t772 AVDD.t194 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X572 DGND bias_n.t37 a_1659_n4497.t3 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X573 DGND bias_n.t38 a_1659_n4497.t4 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X574 DGND Vom.t128 Vfold_bot_m.t48 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X575 bias_n.t2 level_shifter_up_4.xb_hv.t5 DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X576 a_35403_11527# a_34648_11527# DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X577 a_32057_n21342.t3 bias_p.t47 a_32057_n22200.t9 AVDD.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X578 a_2458_6128.t45 a_12760_n20342.t45 AVDD.t231 AVDD.t103 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X579 Vxp.t104 casc_p.t185 a_1657_n21342.t32 AVDD.t196 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X580 AVDD.t342 a_36699_n29829# a_36259_n29829# AVDD.t341 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X581 a_25696_11382.t3 level_shifter_up_8.xb_hv.t6 a_2370_7428.t1 AVDD.t718 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X582 Vop.t44 casc_p.t186 a_2458_6128.t168 AVDD.t85 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X583 a_1657_n21342.t112 a_1560_n22142.t62 AVDD.t773 AVDD.t196 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X584 Vom.t57 casc_p.t187 a_2458_5328.t171 AVDD.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X585 Vom_stg2.t1 Vom_stg2.t0 DGND.t615 DGND.t529 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X586 DGND DGND DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X587 a_2458_6128.t44 a_12760_n20342.t46 AVDD.t63 AVDD.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X588 AVDD.t592 AVDD.t590 AVDD.t591 AVDD.t394 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X589 AVDD.t589 AVDD.t587 AVDD.t588 AVDD.t370 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X590 AVDD.t586 AVDD.t584 AVDD.t585 AVDD.t374 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X591 a_2458_5328.t21 a_12760_n20342.t47 AVDD.t65 AVDD.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X592 AVDD.t286 level_shifter_up_0.xb_hv.t10 a_32057_n15000.t26 AVDD.t285 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X593 Vxp.t31 Vinp.t15 Vfold_bot_m.t30 AVDD.t46 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X594 a_32059_n3351.t12 bias_n.t39 a_32059_n4497.t9 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X595 AVDD.t583 AVDD.t581 AVDD.t582 AVDD.t370 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X596 DGND bias_var_n.t29 a_2467_n30310.t112 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X597 Vxp.t103 casc_p.t188 a_1657_n21342.t33 AVDD.t161 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X598 DGND bias_var_n.t30 a_2467_n30310.t113 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X599 DGND bias_n.t40 a_1659_n4497.t39 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X600 DGND Vom.t129 a_2467_n30310.t54 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X601 a_1659_n4497.t76 casc_n.t90 Vxm.t80 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X602 a_1659_n4497.t75 casc_n.t91 Vxm.t81 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X603 AVDD.t580 AVDD.t578 AVDD.t579 AVDD.t401 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X604 a_1657_n21342.t111 a_1560_n22142.t63 AVDD.t774 AVDD.t161 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X605 a_23013_n25097.t11 casc_p.t189 a_32057_n21342.t14 AVDD.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X606 DGND bias_var_n.t31 a_2467_n30310.t114 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X607 Vxp.t102 casc_p.t190 a_1657_n21342.t34 AVDD.t208 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X608 DGND DGND DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X609 Vxp.t32 Vinp.t16 Vfold_bot_m.t31 AVDD.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X610 Vxp.t101 casc_p.t191 a_1657_n21342.t35 AVDD.t168 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X611 Vop.t43 casc_p.t192 a_2458_6128.t167 AVDD.t125 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X612 Vxp.t100 casc_p.t193 a_1657_n21342.t36 AVDD.t157 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X613 DGND DGND DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X614 a_32059_n3351.t7 level_shifter_up_0.x_hv.t5 DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X615 Vom.t56 casc_p.t194 a_2458_5328.t170 AVDD.t66 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X616 Vxp.t99 casc_p.t195 a_1657_n21342.t37 AVDD.t166 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X617 DGND a_12857_n19016.t9 a_32059_n897.t3 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X618 a_2458_5328.t196 bias_p.t48 AVDD.t823 AVDD.t15 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X619 a_2458_5328.t22 a_12760_n20342.t48 AVDD.t67 AVDD.t66 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X620 AVDD.t577 AVDD.t575 AVDD.t576 AVDD.t381 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X621 a_32059_n4497.t5 casc_n.t92 a_32059_n4755.t8 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X622 a_2467_n30310.t96 casc_n.t93 Vop.t82 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X623 a_2458_5328.t23 a_12760_n20342.t49 AVDD.t69 AVDD.t68 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X624 a_12859_n4497# casc_n.t94 a_11160_n9542.t12 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=1.16e+12p pd=9.16e+06u as=0p ps=0u w=2e+06u l=1e+06u
X625 a_12859_n2697# casc_n.t95 a_9060_4172.t3 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X626 a_2458_6128.t75 Vinm.t23 Vxm.t24 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X627 bias_var_n.t4 casc_p.t196 a_12857_n17742.t6 AVDD.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X628 DGND a_12857_n19016.t10 a_32059_n897.t4 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X629 DGND Vom.t130 a_2467_n30310.t53 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X630 a_12859_2049# ibias.t3 a_11877_1191# DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.16e+12p ps=9.16e+06u w=2e+06u l=4e+06u
X631 a_1659_n4497.t74 casc_n.t96 Vxm.t82 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X632 AVDD.t574 AVDD.t572 AVDD.t573 AVDD.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X633 a_32448_11527# trim[1].t1 DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X634 a_32057_n13616.t5 a_35086_7130.t9 a_2467_n30310.t59 AVDD.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X635 AVDD.t571 AVDD.t569 AVDD.t570 AVDD.t374 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X636 a_2458_5328.t24 a_12760_n20342.t50 AVDD.t71 AVDD.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X637 a_11259_2049# ibias.t4 a_11877_1191# DGND sky130_fd_pr__nfet_g5v0d10v5 ad=1.16e+12p pd=9.16e+06u as=0p ps=0u w=2e+06u l=4e+06u
X638 bias_p.t5 level_shifter_up_4.x_hv.t2 AVDD.t141 AVDD.t140 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X639 a_2467_n29152.t12 casc_p.t197 a_32057_n17742.t18 AVDD.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X640 a_2458_6128.t43 a_12760_n20342.t51 AVDD.t73 AVDD.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X641 a_1657_n21342.t110 a_1560_n22142.t64 AVDD.t775 AVDD.t155 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X642 level_shifter_up_8.x_hv.t0 level_shifter_up_8.xb_hv.t7 AVDD.t720 AVDD.t719 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X643 a_11160_n9542.t7 a_11160_n9542.t6 a_11257_n8742.t3 AVDD.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X644 a_33657_n21342.t7 bias_p.t49 a_33657_n22200.t5 AVDD.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X645 AVDD.t568 AVDD.t566 AVDD.t567 AVDD.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X646 a_2370_n29452.t5 level_shifter_up_3.xb_hv.t6 a_23013_n25097.t7 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X647 Vop.t42 casc_p.t198 a_2458_6128.t143 AVDD.t74 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X648 Vxp.t98 casc_p.t199 a_1657_n21342.t38 AVDD.t172 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X649 a_1659_n4497.t73 casc_n.t97 Vxm.t83 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X650 a_34128_n30483# trim[4].t1 DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=500000u
X651 Vom.t55 casc_p.t200 a_2458_5328.t169 AVDD.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X652 a_2458_6128.t42 a_12760_n20342.t52 AVDD.t75 AVDD.t74 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X653 Vom.t54 casc_p.t201 a_2458_5328.t168 AVDD.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X654 a_1657_n21342.t109 a_1560_n22142.t65 AVDD.t776 AVDD.t172 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X655 DGND bias_var_n.t32 a_2467_n30310.t115 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X656 a_2458_5328.t25 a_12760_n20342.t53 AVDD.t77 AVDD.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X657 a_2458_5328.t51 Vinp.t17 Vxm.t31 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X658 AVDD.t565 AVDD.t563 AVDD.t564 AVDD.t374 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X659 DGND DGND DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X660 a_2458_6128.t41 a_12760_n20342.t54 AVDD.t78 AVDD.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X661 a_33659_n2697.t1 casc_n.t98 a_32059_n4755.t12 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X662 Vfold_bot_m.t92 casc_n.t99 Vom.t80 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X663 a_32057_n15000.t25 level_shifter_up_0.xb_hv.t11 AVDD.t358 AVDD.t357 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X664 AVDD.t562 AVDD.t560 AVDD.t561 AVDD.t370 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X665 a_2458_5328.t26 a_12760_n20342.t55 AVDD.t79 AVDD.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X666 casc_p.t1 casc_p.t0 a_11257_n8742.t10 AVDD.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X667 a_32057_n8742.t3 bias_p.t50 a_32057_n9600.t2 AVDD.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X668 casc_p.t36 casc_p.t34 casc_p.t35 AVDD.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X669 a_32057_n13616.t6 a_35086_7130.t10 a_2467_n30310.t60 AVDD.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X670 a_2458_6128.t40 a_12760_n20342.t56 AVDD.t80 AVDD.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X671 level_shifter_up_1.x_hv a_36328_n30483# DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X672 a_23013_n25097.t10 casc_p.t202 a_32057_n21342.t13 AVDD.t48 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X673 a_2458_6128.t194 bias_p.t51 AVDD.t824 AVDD.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X674 Vfold_bot_m.t91 casc_n.t100 Vom.t106 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X675 a_2467_n30310.t95 casc_n.t101 Vop.t81 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X676 a_34666_7130.t0 a_31098_4670.t7 DGND.t219 DGND.t218 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X677 a_35259_2049# level_shifter_up_6.x_hv.t2 DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=1.74e+12p pd=1.374e+07u as=0p ps=0u w=2e+06u l=500000u
X678 Vxp.t13 Vinm.t24 a_2467_n30310.t9 AVDD.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X679 Vxp.t97 casc_p.t203 a_1657_n21342.t168 AVDD.t208 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X680 casc_n.t21 casc_n.t19 casc_n.t20 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X681 res_p_bot.t15 casc_p.t204 a_11257_n21342# AVDD.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X682 Vom.t53 casc_p.t205 a_2458_5328.t167 AVDD.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X683 Vop.t41 casc_p.t206 a_2458_6128.t142 AVDD.t125 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X684 DGND bias_var_n.t33 a_2467_n30310.t35 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X685 a_1657_n21342.t108 a_1560_n22142.t66 AVDD.t777 AVDD.t208 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X686 Vom.t52 casc_p.t207 a_2458_5328.t166 AVDD.t68 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X687 DGND bias_n.t41 a_1659_n4497.t40 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X688 DGND bias_n.t42 a_1659_n4497.t41 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X689 a_2458_5328.t27 a_12760_n20342.t57 AVDD.t82 AVDD.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X690 DGND DGND DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X691 a_23013_n25097.t14 casc_p.t208 a_33657_n21342.t4 AVDD.t147 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X692 DGND bias_var_n.t34 Vfold_bot_m.t36 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X693 a_2458_5328.t182 bias_p.t52 AVDD.t751 AVDD.t15 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X694 AVDD.t559 AVDD.t557 AVDD.t558 AVDD.t381 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X695 a_2467_n30310.t94 casc_n.t102 Vop.t90 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X696 a_1659_n4497.t72 casc_n.t103 Vxm.t84 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X697 Vxp.t96 casc_p.t209 a_1657_n21342.t169 AVDD.t159 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X698 AVDD.t556 AVDD.t554 AVDD.t555 AVDD.t381 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X699 a_12857_n19016.t0 casc_p.t210 a_12857_n19542.t6 AVDD.t111 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X700 a_25696_11382.t9 level_shifter_up_6.x_hv.t3 a_27926_9740.t2 AVDD.t747 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X701 DGND DGND DGND sky130_fd_pr__res_high_po_2p85 l=3.192e+07u
X702 a_2467_n29152.t0 a_2370_n28652.t9 a_2467_n30310.t17 AVDD.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X703 a_2458_6128.t184 bias_p.t53 AVDD.t752 AVDD.t148 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X704 DGND bias_var_n.t35 a_2467_n30310.t36 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X705 DGND DGND DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X706 a_2458_6128.t39 a_12760_n20342.t58 AVDD.t83 AVDD.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X707 Vxp.t14 Vinm.t25 a_2467_n30310.t10 AVDD.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X708 DGND DGND DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X709 a_1659_n4497.t71 casc_n.t104 Vxm.t85 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X710 DGND DGND DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X711 DGND bias_var_n.t36 Vfold_bot_m.t37 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X712 DGND bias_var_n.t37 Vfold_bot_m.t38 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X713 DGND bias_var_n.t38 a_2467_n30310.t37 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X714 DGND DGND DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X715 DGND bias_n.t43 a_14459_n4209# DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.16e+12p ps=9.16e+06u w=2e+06u l=4e+06u
X716 DGND bias_n.t44 a_14459_n2697# DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X717 a_2467_n30310.t93 casc_n.t105 Vop.t89 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X718 DGND level_shifter_up_7.x_hv.t3 a_32059_2049.t2 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X719 DGND DGND DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X720 a_31928_n30483# trim[5].t1 AVDD.t732 AVDD.t731 sky130_fd_pr__pfet_g5v0d10v5 ad=1.45e+11p pd=1.58e+06u as=0p ps=0u w=500000u l=2e+06u
X721 a_1659_n4497.t70 casc_n.t106 Vxm.t78 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X722 Vxp.t95 casc_p.t211 a_1657_n21342.t170 AVDD.t194 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X723 Vom.t51 casc_p.t212 a_2458_5328.t165 AVDD.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X724 AVDD.t553 AVDD.t551 AVDD.t552 AVDD.t374 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X725 DGND DGND DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X726 a_2458_6128.t38 a_12760_n20342.t59 AVDD.t84 AVDD.t74 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X727 a_1659_n4497.t69 casc_n.t107 Vxm.t60 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X728 a_23013_n25097.t9 casc_p.t213 a_32057_n21342.t12 AVDD.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X729 AVDD.t550 AVDD.t548 AVDD.t549 AVDD.t366 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X730 a_37083_n30483# a_36328_n30483# AVDD.t834 AVDD.t833 sky130_fd_pr__pfet_g5v0d10v5 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=500000u
X731 Vxp.t15 Vinm.t26 a_2467_n30310.t11 AVDD.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X732 Vxp.t94 casc_p.t214 a_1657_n21342.t171 AVDD.t196 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X733 Vxp.t93 casc_p.t215 a_1657_n21342.t172 AVDD.t161 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X734 AVDD.t547 AVDD.t545 AVDD.t546 AVDD.t394 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X735 Vop.t40 casc_p.t216 a_2458_6128.t141 AVDD.t85 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X736 Vxp.t92 casc_p.t217 a_1657_n21342.t173 AVDD.t172 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X737 a_2458_6128.t37 a_12760_n20342.t60 AVDD.t86 AVDD.t85 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X738 AVDD.t100 level_shifter_up_2.xb_hv.t4 a_32057_n22200.t1 AVDD.t99 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X739 a_23013_n25097.t19 casc_p.t218 a_32057_n21342.t11 AVDD.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X740 a_2458_6128.t36 a_12760_n20342.t61 AVDD.t120 AVDD.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X741 a_2458_6128.t185 bias_p.t54 AVDD.t753 AVDD.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X742 Vfold_bot_m.t90 casc_n.t108 Vom.t105 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X743 Vfold_bot_m.t89 casc_n.t109 Vom.t104 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X744 a_1659_n4497.t68 casc_n.t110 Vxm.t61 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X745 a_2467_n30310.t92 casc_n.t111 Vop.t88 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X746 a_2467_n30310.t91 casc_n.t112 Vop.t87 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X747 res_p_bot.t10 level_shifter_up_3.xb_hv.t7 a_2370_n28652.t5 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X748 a_32059_n897.t9 casc_n.t113 a_2458_6570.t9 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X749 Vfold_bot_m.t88 casc_n.t114 Vom.t103 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X750 Vxp.t91 casc_p.t219 a_1657_n21342.t174 AVDD.t168 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X751 casc_n.t18 casc_n.t16 casc_n.t17 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X752 Vfold_bot_m.t108 a_34666_7130.t9 a_32057_n13616.t34 AVDD.t344 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X753 Vxp.t33 Vinp.t18 Vfold_bot_m.t32 AVDD.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X754 AVDD.t544 AVDD.t542 AVDD.t543 AVDD.t401 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X755 a_2458_5328.t35 a_12760_n20342.t62 AVDD.t121 AVDD.t113 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X756 Vom.t50 casc_p.t220 a_2458_5328.t138 AVDD.t68 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X757 a_2458_5328.t178 Vinp.t19 Vxm.t43 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X758 a_2458_5328.t179 Vinp.t20 Vxm.t44 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X759 Vop.t39 casc_p.t221 a_2458_6128.t140 AVDD.t148 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X760 Vfold_bot_m.t87 casc_n.t115 Vom.t102 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X761 AVDD.t541 AVDD.t539 AVDD.t540 AVDD.t401 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X762 AVDD.t538 AVDD.t536 AVDD.t537 AVDD.t401 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X763 Vom.t49 casc_p.t222 a_2458_5328.t137 AVDD.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X764 a_2458_5328.t36 a_12760_n20342.t63 AVDD.t122 AVDD.t68 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X765 Vom.t48 casc_p.t223 a_2458_5328.t136 AVDD.t113 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X766 a_11160_n9542.t5 a_11160_n9542.t4 a_11257_n8742.t2 AVDD.t111 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X767 DGND res_p_bot.t7 res_p_bot.t8 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X768 DGND a_32299_n29829# level_shifter_up_4.x_hv.t1 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X769 bias_stg2.t2 bias_stg2.t1 AVDD.t710 AVDD.t709 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X770 DGND Vom.t131 Vfold_bot_m.t47 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X771 a_2458_6128.t174 Vinm.t27 Vxm.t40 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X772 Vop.t38 casc_p.t224 a_2458_6128.t139 AVDD.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X773 AVDD.t360 level_shifter_up_0.xb_hv.t12 a_32057_n15000.t24 AVDD.t359 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X774 level_shifter_up_6.x_hv a_30248_11527# DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X775 a_32059_n4755.t16 a_34666_7130.t10 a_2458_5328.t186 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X776 Vxp.t137 Vinp.t21 Vfold_bot_m.t61 AVDD.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X777 Vxp.t138 Vinp.t22 Vfold_bot_m.t62 AVDD.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X778 a_2458_5328.t187 Vinp.t23 Vxm.t95 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X779 Vfold_bot_m.t86 casc_n.t116 Vom.t101 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X780 DGND DGND DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X781 a_2458_6128.t186 bias_p.t55 AVDD.t754 AVDD.t148 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X782 AVDD.t248 level_shifter_up_4.x_hv.t3 bias_p.t6 AVDD.t247 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X783 a_2370_n28652.t6 level_shifter_up_3.xb_hv.t8 res_p_bot.t11 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X784 a_2458_6128.t187 bias_p.t56 AVDD.t755 AVDD.t5 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X785 Vop.t37 casc_p.t225 a_2458_6128.t138 AVDD.t74 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X786 a_1657_n21342.t107 a_1560_n22142.t67 AVDD.t778 AVDD.t163 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X787 Vom.t47 casc_p.t226 a_2458_5328.t135 AVDD.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X788 DGND Vom.t132 a_2467_n30310.t52 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X789 DGND hyst[1].t3 a_34499_n29829# DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X790 a_2458_5328.t183 bias_p.t57 AVDD.t756 AVDD.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X791 a_2458_6128.t175 Vinm.t28 Vxm.t41 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X792 Vom.t46 casc_p.t227 a_2458_5328.t134 AVDD.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X793 AVDD.t535 AVDD.t533 AVDD.t534 AVDD.t374 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X794 a_1659_n4497.t67 casc_n.t117 Vxm.t62 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X795 a_2458_5328.t37 a_12760_n20342.t64 AVDD.t123 AVDD.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X796 res_p_bot.t0 level_shifter_up_2.xb_hv.t5 a_27936_n27260.t4 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X797 Vop.t36 casc_p.t228 a_2458_6128.t137 AVDD.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X798 a_2458_6128.t176 Vinm.t29 Vxm.t42 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X799 AVDD.t145 level_shifter_up_2.x_hv level_shifter_up_2.xb_hv.t0 AVDD.t144 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X800 Vom.t45 casc_p.t229 a_2458_5328.t133 AVDD.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X801 Vxp.t29 Vinm.t30 a_2467_n30310.t32 AVDD.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X802 a_23013_n25097.t13 casc_p.t230 a_33657_n21342.t3 AVDD.t48 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X803 a_2458_5328.t188 Vinp.t24 Vxm.t96 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X804 Vfold_bot_m.t109 a_34666_7130.t11 a_32057_n13616.t35 AVDD.t344 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X805 level_shifter_up_4.xb_hv.t0 a_31859_n29829# DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X806 Vfold_bot_m.t85 casc_n.t118 Vom.t100 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X807 AVDD.t354 level_shifter_up_5.xb_hv.t4 level_shifter_up_5.x_hv.t0 AVDD.t353 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X808 DGND DGND DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X809 a_32057_n22200.t0 level_shifter_up_2.xb_hv.t6 AVDD.t715 AVDD.t714 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X810 DGND Vom.t133 Vfold_bot_m.t46 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X811 a_32059_n4497.t4 casc_n.t119 a_32059_n4755.t7 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X812 a_27926_9740.t1 level_shifter_up_6.x_hv.t4 a_25696_11382.t10 AVDD.t748 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X813 Vfold_bot_m.t84 casc_n.t120 Vom.t99 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X814 a_11259_n4497# casc_n.t121 casc_p.t68 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X815 DGND.t524 level_shifter_up_4.xb_hv.t6 a_31098_4670.t5 DGND.t523 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X816 AVDD.t726 level_shifter_up_1.xb_hv.t6 a_33657_n22200.t1 AVDD.t725 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X817 a_2458_6128.t35 a_12760_n20342.t65 AVDD.t124 AVDD.t113 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X818 a_1659_n4497.t66 casc_n.t122 Vxm.t74 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X819 a_27936_n27260.t6 level_shifter_up_2.xb_hv.t7 res_p_bot.t12 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X820 DGND bias_var_n.t39 Vfold_bot_m.t39 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X821 a_1657_n21342.t106 a_1560_n22142.t68 AVDD.t779 AVDD.t196 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X822 Vxp.t90 casc_p.t231 a_1657_n21342.t175 AVDD.t208 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X823 Vop.t35 casc_p.t232 a_2458_6128.t166 AVDD.t148 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X824 a_25696_11382.t5 level_shifter_up_8.xb_hv.t8 a_2370_7428.t0 AVDD.t721 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X825 casc_p.t33 casc_p.t31 casc_p.t32 AVDD.t111 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X826 a_1659_n4497.t65 casc_n.t123 Vxm.t75 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X827 a_2467_n30310.t90 casc_n.t124 Vop.t86 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X828 DGND DGND DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X829 Vop.t34 casc_p.t233 a_2458_6128.t165 AVDD.t125 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X830 Vop.t33 casc_p.t234 a_2458_6128.t164 AVDD.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X831 a_1657_n21342.t105 a_1560_n22142.t69 AVDD.t780 AVDD.t203 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X832 AVDD.t750 level_shifter_up_6.x_hv.t5 level_shifter_up_6.xb_hv AVDD.t749 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X833 a_2458_6128.t80 Vinm.t31 Vxm.t30 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X834 a_2458_6128.t34 a_12760_n20342.t66 AVDD.t126 AVDD.t125 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X835 a_2458_5328.t189 Vinp.t25 Vxm.t97 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X836 a_2458_5328.t184 bias_p.t58 AVDD.t757 AVDD.t15 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X837 a_25696_11382.t2 level_shifter_up_6.x_hv.t6 a_27926_9740.t0 AVDD.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X838 AVDD.t532 AVDD.t530 AVDD.t531 AVDD.t381 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X839 a_2458_6128.t0 bias_p.t59 AVDD.t6 AVDD.t5 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X840 Vxp.t144 Vinp.t26 Vfold_bot_m.t110 AVDD.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X841 Vop.t32 casc_p.t235 a_2458_6128.t163 AVDD.t74 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X842 DGND bias_var_n.t40 Vfold_bot_m.t40 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X843 Vom.t44 casc_p.t236 a_2458_5328.t132 AVDD.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X844 Vxp.t89 casc_p.t237 a_1657_n21342.t3 AVDD.t194 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X845 a_32059_n4497.t3 casc_n.t125 a_32059_n4755.t6 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X846 a_11259_n2697# casc_n.t126 bias_p.t10 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X847 a_1657_n21342.t104 a_1560_n22142.t70 AVDD.t781 AVDD.t163 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X848 a_23013_n25097.t12 casc_p.t238 a_33657_n21342.t5 AVDD.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X849 a_2467_n30310.t89 casc_n.t127 Vop.t119 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X850 a_2458_5328.t2 bias_p.t60 AVDD.t8 AVDD.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X851 casc_p.t67 casc_p.t66 a_11257_n8742.t9 AVDD.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X852 AVDD.t529 AVDD.t527 AVDD.t528 AVDD.t394 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X853 Vxp.t88 casc_p.t239 a_1657_n21342.t4 AVDD.t196 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X854 a_2467_n30310.t88 casc_n.t128 Vop.t118 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X855 Vxp.t30 Vinm.t32 a_2467_n30310.t33 AVDD.t46 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X856 Vfold_bot_m.t83 casc_n.t129 Vom.t98 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X857 a_35259_2049# bias_n.t45 a_35259_903# DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X858 Vxp.t6 Vinp.t27 Vfold_bot_m.t5 AVDD.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X859 Vop.t31 casc_p.t240 a_2458_6128.t162 AVDD.t5 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X860 a_33659_n1551.t4 level_shifter_up_5.x_hv.t3 DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X861 Vop.t30 casc_p.t241 a_2458_6128.t161 AVDD.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X862 bias_p bias_p AVDD.t94 AVDD.t93 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X863 a_2467_n30310.t87 casc_n.t130 Vop.t117 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X864 a_29757_7018.t4 bias_stg2.t7 AVDD.t836 AVDD.t709 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X865 Vxp.t7 Vinp.t28 Vfold_bot_m.t6 AVDD.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X866 a_32059_2049.t6 bias_n.t46 a_32059_903.t6 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X867 a_2458_6128.t91 a_35086_7130.t11 a_32059_n4755.t21 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X868 a_2458_6128.t33 a_12760_n20342.t67 AVDD.t127 AVDD.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X869 Vom.t43 casc_p.t242 a_2458_5328.t131 AVDD.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X870 Vom.t42 casc_p.t243 a_2458_5328.t130 AVDD.t113 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X871 a_23698_4566.t1 a_23032_11382.t1 DGND sky130_fd_pr__res_high_po_2p85 l=3.192e+07u
X872 a_1657_n21342.t103 a_1560_n22142.t71 AVDD.t782 AVDD.t155 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X873 AVDD.t53 hyst[0].t0 a_36699_n29829# AVDD.t52 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1.45e+11p ps=1.58e+06u w=500000u l=2e+06u
X874 Vfold_bot_m.t82 casc_n.t131 Vom.t97 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X875 a_32057_n14142.t7 bias_p.t62 a_32057_n15000.t13 AVDD.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X876 a_2458_6128.t1 bias_p.t63 AVDD.t11 AVDD.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X877 DGND bias_var_n.t41 a_2467_n30310.t40 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X878 a_1657_n21342.t102 a_1560_n22142.t72 AVDD.t783 AVDD.t157 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X879 a_2467_n30310.t116 a_35086_7130.t12 a_32057_n13616.t38 AVDD.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X880 a_2458_5328.t11 Vinp.t29 Vxm.t7 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X881 a_37083_n30483# a_36328_n30483# DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X882 a_32059_n3351.t11 bias_n.t47 a_32059_n4497.t8 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X883 AVDD.t713 a_25696_11382.t7 a_25696_11382.t8 AVDD.t712 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=4e+06u
X884 Vop.t29 casc_p.t244 a_2458_6128.t160 AVDD.t148 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X885 DGND bias_var_n.t42 a_2467_n30310.t41 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X886 Vom.t41 casc_p.t245 a_2458_5328.t129 AVDD.t15 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X887 a_1659_n4497.t64 casc_n.t132 Vxm.t76 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X888 a_1657_n21342.t101 a_1560_n22142.t73 AVDD.t784 AVDD.t203 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X889 Vom.t40 casc_p.t246 a_2458_5328.t128 AVDD.t68 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X890 DGND bias_n.t48 a_1659_n4497.t94 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X891 a_2370_n28652.t2 level_shifter_up_3.x_hv.t4 a_23013_n25097.t0 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X892 Vxp.t36 Vinm.t33 a_2467_n30310.t44 AVDD.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X893 Vom.t39 casc_p.t247 a_2458_5328.t127 AVDD.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X894 bias_p.t2 bias_p.t1 AVDD.t44 AVDD.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X895 DGND DGND DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X896 a_2458_5328.t38 a_12760_n20342.t68 AVDD.t128 AVDD.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X897 AVDD.t89 AVDD.t90 DGND sky130_fd_pr__res_high_po_2p85 l=3.192e+07u
X898 DGND hyst[0].t1 a_36699_n29829# DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=500000u
X899 a_33659_n1551.t3 level_shifter_up_5.x_hv.t4 DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X900 AVDD.t96 a_34499_n29829# a_34059_n29829# AVDD.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X901 DGND trim[0].t2 a_30248_11527# DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X902 Vop_stg2.t1 Vop_stg2.t0 DGND.t23 DGND.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X903 DGND a_35403_11527# level_shifter_up_8.xb_hv DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X904 a_2467_n30310.t86 casc_n.t133 Vop.t116 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X905 Vfold_bot_m.t81 casc_n.t134 Vom.t96 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X906 a_32057_n9600.t9 level_shifter_up_5.xb_hv.t5 AVDD.t356 AVDD.t355 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X907 DGND DGND DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X908 DGND.t528 Vom_stg2.t3 Vop_stg2.t2 DGND.t527 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X909 Vom.t38 casc_p.t248 a_2458_5328.t126 AVDD.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X910 DGND bias_var_n.t43 a_2467_n30310.t42 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X911 DGND bias_n.t49 a_12859_n2697# DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X912 res_p_bot.t13 level_shifter_up_2.xb_hv.t8 a_27936_n27260.t7 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X913 a_12857_n14142.t1 a_12760_n20342.t69 AVDD.t129 AVDD.t93 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X914 Vop.t28 casc_p.t249 a_2458_6128.t157 AVDD.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X915 AVDD.t526 AVDD.t524 AVDD.t525 AVDD.t374 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X916 a_2458_6128.t2 bias_p.t64 AVDD.t13 AVDD.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X917 a_1659_n4497.t63 casc_n.t135 Vxm.t77 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X918 a_9060_4530.t1 a_12760_n20342.t70 AVDD.t131 AVDD.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X919 AVDD.t523 AVDD.t521 AVDD.t522 AVDD.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X920 Vxp.t8 Vinp.t30 Vfold_bot_m.t7 AVDD.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X921 a_1659_n4497.t62 casc_n.t136 Vxm.t59 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X922 a_2458_5328.t9 a_2370_6628.t10 a_2458_6570.t1 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X923 AVDD.t520 AVDD.t518 AVDD.t519 AVDD.t374 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X924 a_2458_6128.t32 a_12760_n20342.t71 AVDD.t132 AVDD.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X925 a_1657_n21342.t100 a_1560_n22142.t74 AVDD.t785 AVDD.t166 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X926 a_1657_n21342.t99 a_1560_n22142.t75 AVDD.t786 AVDD.t208 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X927 DGND bias_var_n.t44 a_2467_n30310.t43 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X928 Vfold_bot_m.t80 casc_n.t137 Vom.t95 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X929 a_33203_11527# a_32448_11527# DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X930 DGND DGND DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X931 AVDD.t517 AVDD.t515 AVDD.t516 AVDD.t366 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X932 a_2467_n30310.t117 a_35086_7130.t13 a_32057_n13616.t39 AVDD.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X933 Vom.t37 casc_p.t250 a_2458_5328.t110 AVDD.t113 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X934 a_9060_4530.t6 bias_p.t65 a_11257_n14142.t0 AVDD.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X935 DGND DGND DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X936 Vop.t27 casc_p.t251 a_2458_6128.t156 AVDD.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X937 level_shifter_up_3.x_hv.t1 level_shifter_up_3.xb_hv.t9 AVDD.t764 AVDD.t763 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X938 DGND bias_var_n.t45 a_2467_n30310.t30 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X939 a_1657_n21342.t98 a_1560_n22142.t76 AVDD.t156 AVDD.t155 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X940 Vxp.t1 Vinp.t31 Vfold_bot_m.t1 AVDD.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X941 a_32057_n14142.t6 bias_p.t66 a_32057_n15000.t12 AVDD.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X942 level_shifter_up_0.xb_hv.t0 level_shifter_up_0.x_hv.t6 AVDD.t265 AVDD.t264 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X943 a_32057_n14142.t5 bias_p.t67 a_32057_n15000.t2 AVDD.t147 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X944 Vxp.t87 casc_p.t252 a_1657_n21342.t5 AVDD.t203 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X945 Vxp.t86 casc_p.t253 a_1657_n21342.t6 AVDD.t208 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X946 Vxp.t37 Vinm.t34 a_2467_n30310.t45 AVDD.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X947 a_2467_n30310.t85 casc_n.t138 Vop.t115 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X948 a_1657_n21342.t97 a_1560_n22142.t77 AVDD.t158 AVDD.t157 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X949 Vfold_bot_m.t79 casc_n.t139 Vom.t118 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X950 a_32059_903.t0 casc_n.t140 a_23032_4566.t11 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X951 a_36328_n30483# trim[3].t1 AVDD.t143 AVDD.t142 sky130_fd_pr__pfet_g5v0d10v5 ad=1.45e+11p pd=1.58e+06u as=0p ps=0u w=500000u l=2e+06u
X952 a_1657_n21342.t96 a_1560_n22142.t78 AVDD.t160 AVDD.t159 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X953 a_27926_9740.t7 level_shifter_up_7.x_hv.t4 a_23032_4566.t8 AVDD.t711 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X954 a_32059_n897.t8 casc_n.t141 a_2458_6570.t8 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X955 a_2467_n30310.t84 casc_n.t142 Vop.t114 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X956 DGND a_12857_n19016.t11 a_32059_n897.t5 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X957 a_2458_5328.t39 a_12760_n20342.t72 AVDD.t133 AVDD.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X958 a_1659_n4497.t61 casc_n.t143 Vxm.t52 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X959 DGND trim[4].t2 a_34128_n30483# DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X960 Vom.t36 casc_p.t254 a_2458_5328.t109 AVDD.t15 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X961 a_2458_6128.t31 a_12760_n20342.t73 AVDD.t134 AVDD.t103 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X962 a_2458_5328.t92 bias_p.t68 AVDD.t345 AVDD.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X963 DGND level_shifter_up_0.x_hv.t7 a_32059_n3351.t3 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X964 a_2458_6128.t30 a_12760_n20342.t74 AVDD.t135 AVDD.t85 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X965 DGND a_34883_n30483# level_shifter_up_2.xb_hv.t1 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X966 DGND a_12857_n19016.t12 a_32059_n897.t1 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X967 a_2458_5328.t93 bias_p.t69 AVDD.t346 AVDD.t15 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X968 AVDD.t514 AVDD.t512 AVDD.t513 AVDD.t381 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X969 a_11257_n14142.t2 bias_p.t70 AVDD.t347 AVDD.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X970 AVDD.t362 level_shifter_up_0.xb_hv.t13 a_32057_n15000.t23 AVDD.t361 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X971 Vop.t26 casc_p.t255 a_2458_6128.t155 AVDD.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X972 AVDD.t511 AVDD.t509 AVDD.t510 AVDD.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X973 a_2458_5328.t6 Vinp.t32 Vxm.t2 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X974 AVDD.t508 AVDD.t506 AVDD.t507 AVDD.t370 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X975 a_2458_6128.t29 a_12760_n20342.t75 AVDD.t136 AVDD.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X976 AVDD.t505 AVDD.t503 AVDD.t504 AVDD.t366 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X977 a_2458_5328.t43 a_34666_7130.t12 a_32059_n4755.t0 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X978 a_2458_5328.t94 bias_p.t71 AVDD.t348 AVDD.t5 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X979 Vop.t25 casc_p.t256 a_2458_6128.t154 AVDD.t74 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X980 a_1657_n21342.t95 a_1560_n22142.t79 AVDD.t162 AVDD.t161 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X981 Vout.t1 a_35086_7130.t14 DGND.t676 DGND.t675 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X982 a_2458_6128.t28 a_12760_n20342.t76 AVDD.t101 AVDD.t74 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X983 a_1657_n21342.t94 a_1560_n22142.t80 AVDD.t164 AVDD.t163 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X984 DGND Vom.t134 Vfold_bot_m.t45 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X985 Vxp.t2 Vinp.t33 Vfold_bot_m.t2 AVDD.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X986 a_2458_5328.t95 bias_p.t72 AVDD.t349 AVDD.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X987 a_12857_n15942.t1 a_1560_n22142.t81 AVDD.t165 AVDD.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X988 a_2458_6128.t92 bias_p.t73 AVDD.t350 AVDD.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X989 a_32057_n14142.t4 bias_p.t74 a_32057_n15000.t1 AVDD.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X990 a_30248_11527# trim[0].t3 DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X991 a_1659_n4497.t60 casc_n.t144 Vxm.t53 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X992 a_1659_n4497.t59 casc_n.t145 Vxm.t54 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X993 a_23032_4566.t18 level_shifter_up_8.x_hv.t2 a_2370_7428.t7 AVDD.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X994 a_1657_n21342.t93 a_1560_n22142.t82 AVDD.t167 AVDD.t166 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X995 DGND bias_var_n.t46 Vfold_bot_m.t28 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X996 a_1657_n21342.t92 a_1560_n22142.t83 AVDD.t169 AVDD.t168 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X997 level_shifter_up_7.x_hv.t0 level_shifter_up_7.xb_hv AVDD.t271 AVDD.t270 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X998 AVDD.t502 AVDD.t500 AVDD.t501 AVDD.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X999 Vop.t24 casc_p.t257 a_2458_6128.t153 AVDD.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1000 Vop.t23 casc_p.t258 a_2458_6128.t152 AVDD.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1001 a_2458_5328.t28 a_12760_n20342.t77 AVDD.t102 AVDD.t66 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1002 a_2458_6128.t190 bias_p.t75 AVDD.t758 AVDD.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1003 DGND DGND DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1004 a_2370_n28652.t7 level_shifter_up_3.xb_hv.t10 res_p_bot.t16 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X1005 a_32057_n17742.t5 a_1560_n22142.t84 AVDD.t170 AVDD.t147 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1006 DGND DGND DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1007 Vfold_bot_m.t78 casc_n.t146 Vom.t117 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1008 DGND DGND DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1009 Vxp.t85 casc_p.t259 a_1657_n21342.t7 AVDD.t203 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1010 bias_p bias_p AVDD.t92 AVDD.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1011 a_2458_6128.t182 a_2370_7428.t10 a_2458_6570.t4 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1012 a_1657_n21342.t91 a_1560_n22142.t85 AVDD.t171 AVDD.t159 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1013 a_32059_n4497.t2 casc_n.t147 a_32059_n4755.t11 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1014 a_2467_n30310.t83 casc_n.t148 Vop.t113 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1015 Vom.t35 casc_p.t260 a_2458_5328.t108 AVDD.t68 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1016 a_2467_n30310.t82 casc_n.t149 Vop.t112 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1017 a_1659_n4497.t58 casc_n.t150 Vxm.t55 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1018 a_2458_6128.t27 a_12760_n20342.t78 AVDD.t104 AVDD.t103 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1019 a_2458_5328.t7 Vinp.t34 Vxm.t3 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1020 a_32057_n14142.t3 bias_p.t77 a_32057_n15000.t0 AVDD.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1021 AVDD.t499 AVDD.t497 AVDD.t498 AVDD.t394 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1022 a_1657_n21342.t90 a_1560_n22142.t86 AVDD.t173 AVDD.t172 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1023 DGND Vom.t135 Vfold_bot_m.t44 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1024 DGND bias_var_n.t47 a_2467_n30310.t31 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1025 DGND DGND DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1026 Vop.t22 casc_p.t261 a_2458_6128.t151 AVDD.t148 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1027 a_2458_5328.t29 a_12760_n20342.t79 AVDD.t106 AVDD.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1028 Vxp.t12 Vinp.t35 Vfold_bot_m.t8 AVDD.t46 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1029 Vop.t21 casc_p.t262 a_2458_6128.t113 AVDD.t5 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1030 a_2458_6128.t191 bias_p.t78 AVDD.t759 AVDD.t148 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1031 level_shifter_up_5.xb_hv.t1 a_36259_n29829# DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1032 a_1659_n4497.t57 casc_n.t151 Vxm.t56 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1033 DGND level_shifter_up_7.x_hv.t5 a_32059_2049.t1 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1034 a_36699_n29829# hyst[0].t2 DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1035 Vxp.t84 casc_p.t263 a_1657_n21342.t39 AVDD.t163 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1036 DGND bias_n.t50 a_1659_n4497.t95 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1037 AVDD.t496 AVDD.t494 AVDD.t495 AVDD.t370 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1038 DGND DGND DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1039 DGND DGND DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1040 Vom.t34 casc_p.t264 a_2458_5328.t107 AVDD.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1041 casc_p.t30 casc_p.t28 casc_p.t29 AVDD.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1042 AVDD.t809 level_shifter_up_5.xb_hv.t6 a_32057_n9600.t8 AVDD.t808 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1043 a_1657_n21342.t89 a_1560_n22142.t87 AVDD.t174 AVDD.t161 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1044 Vom.t33 casc_p.t265 a_2458_5328.t106 AVDD.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1045 a_2458_5328.t13 Vinp.t36 Vxm.t8 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1046 a_32059_n4755.t20 a_35086_7130.t15 a_2458_6128.t196 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1047 a_2467_n30310.t81 casc_n.t152 Vop.t111 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1048 a_34648_11527# trim[2].t2 AVDD.t746 AVDD.t745 sky130_fd_pr__pfet_g5v0d10v5 ad=1.45e+11p pd=1.58e+06u as=0p ps=0u w=500000u l=2e+06u
X1049 a_32057_n14142.t2 bias_p.t79 a_32057_n15000.t8 AVDD.t48 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1050 a_2458_6128.t88 Vinm.t35 Vxm.t36 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1051 a_27936_n27260.t5 level_shifter_up_2.xb_hv.t9 res_p_bot.t9 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X1052 casc_p.t27 casc_p.t25 casc_p.t26 AVDD.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1053 a_32057_n8742.t4 bias_p.t80 a_32057_n9600.t1 AVDD.t147 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1054 a_32057_n17742.t4 a_1560_n22142.t88 AVDD.t175 AVDD.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1055 a_2458_5328.t30 a_12760_n20342.t80 AVDD.t107 AVDD.t68 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1056 a_25030_4566.t1 a_24364_11382.t1 DGND sky130_fd_pr__res_high_po_2p85 l=3.192e+07u
X1057 a_2458_5328.t14 Vinp.t37 Vxm.t9 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1058 a_2370_n28652.t1 level_shifter_up_3.x_hv.t5 a_23013_n25097.t1 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X1059 a_32057_n8742.t5 bias_p.t81 a_32057_n9600.t0 AVDD.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1060 a_23032_4566.t0 level_shifter_up_7.x_hv.t6 a_27926_9740.t6 AVDD.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X1061 DGND DGND DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1062 a_2467_n30310.t80 casc_n.t153 Vop.t110 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1063 a_1657_n21342.t88 a_1560_n22142.t89 AVDD.t176 AVDD.t168 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1064 a_2458_5328.t31 a_12760_n20342.t81 AVDD.t108 AVDD.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1065 casc_n.t15 casc_n.t13 casc_n.t14 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1066 a_2458_5328.t15 Vinp.t38 Vxm.t10 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1067 a_32057_n13616.t8 casc_p.t266 a_32057_n14142.t27 AVDD.t147 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1068 a_12859_n4755# bias_n.t51 a_12859_n4209# DGND sky130_fd_pr__nfet_g5v0d10v5 ad=1.16e+12p pd=9.16e+06u as=0p ps=0u w=2e+06u l=4e+06u
X1069 DGND bias_var_n.t48 Vfold_bot_m.t29 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1070 a_12857_n17742.t1 a_1560_n22142.t90 AVDD.t177 AVDD.t93 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1071 a_32057_n15000.t22 level_shifter_up_0.xb_hv.t14 AVDD.t364 AVDD.t363 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1072 a_2458_5328.t32 a_12760_n20342.t82 AVDD.t109 AVDD.t66 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1073 Vxp.t83 casc_p.t267 a_1657_n21342.t40 AVDD.t159 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1074 bias_p.t7 level_shifter_up_4.x_hv.t4 AVDD.t250 AVDD.t249 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X1075 Vxp.t9 Vinm.t36 a_2467_n30310.t6 AVDD.t46 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1076 DGND bias_n.t52 a_1659_n4497.t30 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1077 AVDD.t493 AVDD.t491 AVDD.t492 AVDD.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1078 a_2467_n29152.t1 a_2370_n28652.t10 a_2467_n30310.t18 AVDD.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1079 a_24345_n31913# a_23679_n25097# DGND sky130_fd_pr__res_high_po_2p85 l=3.192e+07u
X1080 a_12857_n14142.t0 a_12760_n20342.t83 AVDD.t110 AVDD.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1081 Vop.t20 casc_p.t268 a_2458_6128.t112 AVDD.t113 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1082 a_9060_4530.t0 a_12760_n20342.t84 AVDD.t112 AVDD.t111 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1083 DGND Vom.t136 Vfold_bot_m.t43 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1084 a_32059_n4755.t19 a_35086_7130.t16 a_2458_6128.t197 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1085 a_1657_n21342.t87 a_1560_n22142.t91 AVDD.t178 AVDD.t155 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1086 a_2458_6128.t26 a_12760_n20342.t85 AVDD.t114 AVDD.t113 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1087 a_34128_n30483# trim[4].t3 DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1088 a_32057_n17742.t3 a_1560_n22142.t92 AVDD.t179 AVDD.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1089 Vom_stg2.t2 Vop_stg2.t4 DGND.t442 DGND.t441 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X1090 a_32057_n14142.t1 bias_p.t82 a_32057_n15000.t7 AVDD.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1091 DGND Vom.t137 a_2467_n30310.t51 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1092 Vxp.t147 Vinp.t39 Vfold_bot_m.t116 AVDD.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1093 a_1657_n21342.t86 a_1560_n22142.t93 AVDD.t180 AVDD.t157 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1094 a_1657_n21342.t85 a_1560_n22142.t94 AVDD.t193 AVDD.t172 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1095 a_1657_n21342.t84 a_1560_n22142.t95 AVDD.t195 AVDD.t194 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1096 a_2458_5328.t33 a_12760_n20342.t86 AVDD.t115 AVDD.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1097 a_32059_n3351.t10 bias_n.t53 a_32059_n4497.t15 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1098 a_33659_n1551.t0 bias_n.t54 a_33659_n2697.t4 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1099 Vom.t32 casc_p.t269 a_2458_5328.t105 AVDD.t15 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1100 Vom.t31 casc_p.t270 a_2458_5328.t104 AVDD.t5 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1101 a_32057_n14142.t0 bias_p.t83 a_32057_n15000.t6 AVDD.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1102 DGND bias_var_n.t49 Vfold_bot_m.t25 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1103 DGND bias_var_n.t50 Vfold_bot_m.t26 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1104 level_shifter_up_3.x_hv.t0 a_31928_n30483# DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1105 DGND bias_n.t55 a_11259_n2697# DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1106 a_1659_n4497.t56 casc_n.t154 Vxm.t57 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1107 a_1659_n4497.t55 casc_n.t155 Vxm.t58 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1108 a_2370_7428.t6 level_shifter_up_8.x_hv.t3 a_23032_4566.t17 AVDD.t152 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X1109 a_2458_5328.t47 bias_p.t84 AVDD.t186 AVDD.t5 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1110 a_1657_n21342.t83 a_1560_n22142.t96 AVDD.t197 AVDD.t196 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1111 Vxp.t82 casc_p.t271 a_1657_n21342.t41 AVDD.t163 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1112 Vom.t30 casc_p.t272 a_2458_5328.t103 AVDD.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1113 a_2458_6128.t25 a_12760_n20342.t87 AVDD.t116 AVDD.t85 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1114 DGND DGND DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1115 a_1560_n22142.t5 casc_p.t273 a_12857_n14142.t5 AVDD.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1116 a_1657_n21342.t82 a_1560_n22142.t97 AVDD.t198 AVDD.t163 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1117 a_32057_n13616.t22 casc_p.t274 a_32057_n14142.t26 AVDD.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1118 DGND DGND DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1119 AVDD.t490 AVDD.t488 AVDD.t489 AVDD.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1120 a_2458_5328.t48 bias_p.t85 AVDD.t187 AVDD.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1121 Vxp.t81 casc_p.t275 a_1657_n21342.t42 AVDD.t159 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1122 a_33657_n22200.t0 level_shifter_up_1.xb_hv.t7 AVDD.t728 AVDD.t727 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1123 a_32057_n17742.t2 a_1560_n22142.t98 AVDD.t199 AVDD.t48 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1124 Vxp.t80 casc_p.t276 a_1657_n21342.t43 AVDD.t168 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1125 Vxp.t79 casc_p.t277 a_1657_n21342.t44 AVDD.t168 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1126 casc_p.t24 casc_p.t22 casc_p.t23 AVDD.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1127 a_12760_n20342.t2 casc_p.t278 a_9060_4530.t9 AVDD.t93 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1128 a_35086_7130.t0 a_34666_7130.t13 DVDD.t11 DVDD.t10 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1129 DGND DGND DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1130 AVDD.t487 AVDD.t485 AVDD.t486 AVDD.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1131 DGND DGND DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1132 Vop.t19 casc_p.t279 a_2458_6128.t111 AVDD.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1133 DGND DGND DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1134 AVDD.t484 AVDD.t482 AVDD.t483 AVDD.t381 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1135 Vfold_bot_m.t77 casc_n.t156 Vom.t116 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1136 Vfold_bot_m.t76 casc_n.t157 Vom.t115 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1137 a_2458_5328.t34 a_12760_n20342.t88 AVDD.t117 AVDD.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1138 a_14459_n4497# casc_n.t158 a_12760_n20342.t4 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1139 a_14459_n2697# casc_n.t159 a_1560_n22142.t7 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1140 AVDD.t481 AVDD.t479 AVDD.t480 AVDD.t401 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1141 a_32057_n13616.t21 casc_p.t280 a_32057_n14142.t25 AVDD.t147 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1142 Vfold_bot_m.t75 casc_n.t160 Vom.t114 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1143 a_2458_5328.t49 bias_p.t86 AVDD.t188 AVDD.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1144 DGND bias_n.t56 a_1659_n4497.t20 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1145 Vxp.t78 casc_p.t281 a_1657_n21342.t45 AVDD.t159 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1146 Vxp.t77 casc_p.t282 a_1657_n21342.t46 AVDD.t155 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1147 Vxp.t148 Vinp.t40 Vfold_bot_m.t117 AVDD.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1148 a_1657_n21342.t81 a_1560_n22142.t99 AVDD.t200 AVDD.t166 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1149 DGND bias_n.t57 a_1659_n4497.t21 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1150 a_32057_n13616.t13 casc_p.t283 a_32057_n8742.t7 AVDD.t48 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1151 a_32057_n13616.t20 casc_p.t284 a_32057_n14142.t24 AVDD.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1152 Vop.t18 casc_p.t285 a_2458_6128.t110 AVDD.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1153 a_11160_n9542.t11 a_11160_n9542.t10 a_11257_n8742.t1 AVDD.t93 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1154 a_32057_n13616.t12 casc_p.t286 a_32057_n8742.t6 AVDD.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1155 a_12857_n15942.t0 a_1560_n22142.t100 AVDD.t201 AVDD.t111 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1156 Vom.t29 casc_p.t287 a_2458_5328.t102 AVDD.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1157 Vop.t17 casc_p.t288 a_2458_6128.t109 AVDD.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1158 a_11160_n9542.t9 a_11160_n9542.t8 a_11257_n8742.t0 AVDD.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1159 Vxp.t76 casc_p.t289 a_1657_n21342.t47 AVDD.t157 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1160 DGND bias_n.t58 a_1659_n4497.t22 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1161 a_2458_5328.t195 Vinp.t41 Vxm.t102 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1162 Vom.t28 casc_p.t290 a_2458_5328.t101 AVDD.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1163 AVDD.t478 AVDD.t476 AVDD.t477 AVDD.t366 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1164 a_32683_n30483# a_31928_n30483# AVDD.t191 AVDD.t190 sky130_fd_pr__pfet_g5v0d10v5 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=500000u
X1165 Vxp.t75 casc_p.t291 a_1657_n21342.t48 AVDD.t203 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1166 a_1659_n4497.t54 casc_n.t161 Vxm.t51 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1167 a_1657_n21342.t80 a_1560_n22142.t101 AVDD.t202 AVDD.t194 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1168 a_34648_11527# trim[2].t3 DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1169 a_1657_n21342.t79 a_1560_n22142.t102 AVDD.t204 AVDD.t203 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1170 a_32057_n17742.t1 a_1560_n22142.t103 AVDD.t205 AVDD.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1171 a_2458_6128.t24 a_12760_n20342.t89 AVDD.t118 AVDD.t103 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1172 a_23013_n25097.t20 level_shifter_up_3.x_hv.t6 a_2370_n28652.t0 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X1173 casc_p.t21 casc_p.t19 casc_p.t20 AVDD.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1174 a_35403_11527# a_34648_11527# AVDD.t41 AVDD.t40 sky130_fd_pr__pfet_g5v0d10v5 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=500000u
X1175 a_1657_n21342.t78 a_1560_n22142.t104 AVDD.t206 AVDD.t196 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1176 a_32057_n13616.t25 casc_p.t292 a_32057_n14142.t23 AVDD.t48 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1177 Vom.t27 casc_p.t293 a_2458_5328.t100 AVDD.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1178 DGND Vom.t138 Vfold_bot_m.t42 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1179 a_2458_6128.t23 a_12760_n20342.t90 AVDD.t119 AVDD.t85 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1180 DGND bias_var_n.t51 a_2467_n30310.t28 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1181 a_32057_n13616.t24 casc_p.t294 a_32057_n14142.t22 AVDD.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1182 a_2458_5328.t82 a_12760_n20342.t91 AVDD.t312 AVDD.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1183 Vxp.t10 Vinm.t37 a_2467_n30310.t7 AVDD.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1184 Vxp.t11 Vinm.t38 a_2467_n30310.t8 AVDD.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1185 a_2370_n29452.t6 level_shifter_up_3.x_hv.t7 res_p_bot.t4 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X1186 a_32059_2049.t5 bias_n.t59 a_32059_903.t5 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1187 DGND bias_n.t60 a_1659_n4497.t9 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1188 Vxp.t74 casc_p.t295 a_1657_n21342.t18 AVDD.t168 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1189 a_2458_6128.t183 a_2370_7428.t11 a_2458_6570.t5 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1190 AVDD.t475 AVDD.t473 AVDD.t474 AVDD.t370 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1191 DGND bias_n.t61 a_1659_n4497.t10 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1192 a_1560_n22142.t2 casc_p.t296 a_12857_n15942.t5 AVDD.t93 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1193 Vop.t16 casc_p.t297 a_2458_6128.t108 AVDD.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1194 a_32059_2049.t4 bias_n.t62 a_32059_903.t4 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1195 DGND bias_n.t63 a_1659_n4497.t11 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1196 a_1657_n21342.t77 a_1560_n22142.t105 AVDD.t207 AVDD.t161 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1197 a_12857_n19542.t1 a_12760_n20342.t92 AVDD.t313 AVDD.t93 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1198 Vxp.t73 casc_p.t298 a_1657_n21342.t19 AVDD.t166 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1199 AVDD.t472 AVDD.t470 AVDD.t471 AVDD.t401 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1200 AVDD.t826 level_shifter_up_0.xb_hv.t15 a_32057_n15000.t21 AVDD.t825 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1201 a_2467_n30310.t79 casc_n.t162 Vop.t105 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1202 Vxp.t150 Vinm.t39 a_2467_n30310.t118 AVDD.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1203 casc_p.t18 casc_p.t16 casc_p.t17 AVDD.t111 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1204 a_1657_n21342.t76 a_1560_n22142.t106 AVDD.t209 AVDD.t208 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1205 Vxp.t72 casc_p.t299 a_1657_n21342.t20 AVDD.t155 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1206 casc_n.t12 casc_n.t10 casc_n.t11 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1207 a_2467_n29152.t11 casc_p.t300 a_32057_n17742.t17 AVDD.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1208 a_2458_6128.t22 a_12760_n20342.t93 AVDD.t314 AVDD.t125 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1209 a_1657_n21342.t75 a_1560_n22142.t107 AVDD.t210 AVDD.t155 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1210 a_1657_n21342.t74 a_1560_n22142.t108 AVDD.t211 AVDD.t157 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1211 DGND Vom.t139 a_2467_n30310.t50 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1212 AVDD.t469 AVDD.t467 AVDD.t468 AVDD.t46 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1213 DGND bias_var_n.t52 Vfold_bot_m.t27 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1214 a_2458_5328.t83 a_12760_n20342.t94 AVDD.t315 AVDD.t66 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1215 a_1657_n21342.t73 a_1560_n22142.t109 AVDD.t212 AVDD.t166 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1216 a_32057_n21342.t2 bias_p.t87 a_32057_n22200.t8 AVDD.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1217 Vxp.t71 casc_p.t301 a_1657_n21342.t21 AVDD.t157 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1218 Vxp.t70 casc_p.t302 a_1657_n21342.t22 AVDD.t194 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1219 AVDD.t466 AVDD.t464 AVDD.t465 AVDD.t381 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1220 a_36328_n30483# trim[3].t2 DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1221 a_23032_4566.t1 level_shifter_up_7.x_hv.t7 a_27926_9740.t5 AVDD.t57 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X1222 Vom.t26 casc_p.t303 a_2458_5328.t99 AVDD.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1223 a_1657_n21342.t72 a_1560_n22142.t110 AVDD.t213 AVDD.t157 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1224 a_32057_n13616.t23 casc_p.t304 a_32057_n14142.t21 AVDD.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1225 Vop.t15 casc_p.t305 a_2458_6128.t107 AVDD.t103 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1226 a_12857_n17742.t0 a_1560_n22142.t111 AVDD.t214 AVDD.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1227 Vom.t25 casc_p.t306 a_2458_5328.t98 AVDD.t15 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1228 Vxp.t69 casc_p.t307 a_1657_n21342.t23 AVDD.t196 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1229 AVDD.t463 AVDD.t461 AVDD.t462 AVDD.t374 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1230 Vxp.t68 casc_p.t308 a_1657_n21342.t24 AVDD.t194 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1231 a_32057_n17742.t0 a_1560_n22142.t112 AVDD.t858 AVDD.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1232 DGND DGND DGND sky130_fd_pr__res_high_po_2p85 l=3.192e+07u
X1233 AVDD.t724 level_shifter_up_4.xb_hv.t7 level_shifter_up_4.x_hv.t0 AVDD.t723 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1234 a_1659_n4497.t53 casc_n.t163 Vxm.t92 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1235 casc_p.t15 casc_p.t13 casc_p.t14 AVDD.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1236 a_11257_n8742.t6 a_11160_n9542.t14 AVDD.t151 AVDD.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1237 a_23032_4566.t16 level_shifter_up_8.x_hv.t4 a_2370_7428.t5 AVDD.t153 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X1238 a_2458_6128.t21 a_12760_n20342.t95 AVDD.t316 AVDD.t74 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1239 a_1657_n21342.t71 a_1560_n22142.t113 AVDD.t859 AVDD.t172 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1240 DGND bias_n.t64 a_37477_903# DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.16e+12p ps=9.16e+06u w=2e+06u l=4e+06u
X1241 a_32057_n13616.t19 casc_p.t309 a_32057_n14142.t20 AVDD.t48 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1242 Vfold_bot_m.t74 casc_n.t164 Vom.t113 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1243 AVDD.t460 AVDD.t458 AVDD.t459 AVDD.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1244 AVDD.t457 AVDD.t455 AVDD.t456 AVDD.t370 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1245 a_32059_n897.t7 casc_n.t165 a_2458_6570.t7 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1246 DGND DGND DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1247 a_2467_n30310.t78 casc_n.t166 Vop.t104 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1248 a_2458_5328.t84 a_12760_n20342.t96 AVDD.t317 AVDD.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1249 Vom.t24 casc_p.t310 a_2458_5328.t164 AVDD.t5 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1250 Vxp.t149 Vinp.t42 Vfold_bot_m.t118 AVDD.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1251 AVDD.t137 AVDD.t138 DGND sky130_fd_pr__res_high_po_2p85 l=3.192e+07u
X1252 Vxp.t67 casc_p.t311 a_1657_n21342.t25 AVDD.t161 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1253 AVDD.t454 AVDD.t452 AVDD.t453 AVDD.t394 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1254 Vxp.t66 casc_p.t312 a_1657_n21342.t26 AVDD.t163 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1255 DGND bias_n.t65 a_1659_n4497.t0 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1256 Vom.t23 casc_p.t313 a_2458_5328.t163 AVDD.t15 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1257 Vop.t14 casc_p.t314 a_2458_6128.t125 AVDD.t103 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1258 Vom.t22 casc_p.t315 a_2458_5328.t162 AVDD.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1259 Vom.t21 casc_p.t316 a_2458_5328.t161 AVDD.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1260 bias_var_n.t3 casc_p.t317 a_12857_n17742.t5 AVDD.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1261 Vop.t13 casc_p.t318 a_2458_6128.t124 AVDD.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1262 Vom.t20 casc_p.t319 a_2458_5328.t160 AVDD.t66 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1263 a_2458_5328.t50 bias_p.t88 AVDD.t189 AVDD.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1264 AVDD.t451 AVDD.t449 AVDD.t450 AVDD.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1265 Vxp.t65 casc_p.t320 a_1657_n21342.t27 AVDD.t166 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1266 DVDD.t3 a_29758_4670.t0 a_29758_4670.t1 DVDD.t2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1267 DGND bias_n.t4 bias_n.t5 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1268 a_2370_7428.t4 level_shifter_up_8.x_hv.t5 a_23032_4566.t15 AVDD.t154 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X1269 casc_p.t12 casc_p.t10 casc_p.t11 AVDD.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1270 a_1560_n22142.t3 casc_p.t321 a_12857_n14142.t4 AVDD.t111 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1271 a_1657_n21342.t70 a_1560_n22142.t114 AVDD.t860 AVDD.t166 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1272 Vom.t19 casc_p.t322 a_2458_5328.t159 AVDD.t66 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1273 a_1657_n21342.t69 a_1560_n22142.t115 AVDD.t861 AVDD.t208 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1274 a_11257_n21342# bias_p.t89 AVDD.t146 AVDD.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1275 Vxp.t151 Vinm.t40 a_2467_n30310.t119 AVDD.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1276 a_2458_5328.t10 a_2370_6628.t11 a_2458_6570.t2 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1277 a_2458_5328.t17 Vinp.t43 Vxm.t14 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1278 Vop.t12 casc_p.t323 a_2458_6128.t123 AVDD.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1279 DGND bias_n.t66 a_1659_n4497.t1 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1280 a_2458_5328.t85 a_12760_n20342.t97 AVDD.t318 AVDD.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1281 level_shifter_up_4.xb_hv.t1 level_shifter_up_4.x_hv.t5 AVDD.t742 AVDD.t741 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1282 a_2458_6128.t20 a_12760_n20342.t98 AVDD.t319 AVDD.t125 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1283 a_2467_n29152.t10 casc_p.t324 a_32057_n17742.t16 AVDD.t147 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1284 a_2458_5328.t86 a_12760_n20342.t99 AVDD.t320 AVDD.t68 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1285 a_12760_n20342.t1 casc_p.t325 a_9060_4530.t8 AVDD.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1286 a_2458_6128.t199 Vinm.t41 Vxm.t103 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1287 a_2458_6128.t85 Vinm.t42 Vxm.t35 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1288 a_32059_n3351.t9 bias_n.t67 a_32059_n4497.t14 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1289 DGND bias_n.t68 a_11259_n4497# DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1290 Vfold_bot_m.t73 casc_n.t167 Vom.t112 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1291 a_33657_n21342.t0 bias_p.t90 a_33657_n22200.t4 AVDD.t147 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1292 a_2458_5328.t18 Vinp.t44 Vxm.t15 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1293 Vxp.t64 casc_p.t326 a_1657_n21342.t157 AVDD.t159 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1294 Vxp.t63 casc_p.t327 a_1657_n21342.t158 AVDD.t194 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1295 AVDD.t448 AVDD.t446 AVDD.t447 AVDD.t381 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1296 DGND trim[5].t2 a_31928_n30483# DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1297 a_32057_n13616.t18 casc_p.t328 a_32057_n14142.t19 AVDD.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1298 Vop.t11 casc_p.t329 a_2458_6128.t122 AVDD.t103 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1299 a_32057_n13616.t17 casc_p.t330 a_32057_n14142.t18 AVDD.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1300 DGND.t526 level_shifter_up_4.xb_hv.t8 a_31098_4670.t4 DGND.t525 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1301 a_2458_5328.t19 Vinp.t45 Vxm.t16 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1302 a_1657_n21342.t68 a_1560_n22142.t116 AVDD.t862 AVDD.t159 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1303 DGND bias_n.t69 a_1659_n4497.t7 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1304 res_p_bot.t3 level_shifter_up_3.x_hv.t8 a_2370_n29452.t7 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X1305 a_2458_6128.t19 a_12760_n20342.t100 AVDD.t321 AVDD.t103 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1306 Vxp.t34 Vinm.t43 a_2467_n30310.t38 AVDD.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1307 Vxp.t62 casc_p.t331 a_1657_n21342.t159 AVDD.t196 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1308 Vxp.t61 casc_p.t332 a_1657_n21342.t160 AVDD.t172 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1309 a_1659_n4497.t52 casc_n.t168 Vxm.t93 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1310 a_2458_6128.t198 a_35086_7130.t17 a_32059_n4755.t18 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1311 Vom.t18 casc_p.t333 a_2458_5328.t158 AVDD.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1312 a_32059_n3351.t4 level_shifter_up_0.x_hv.t8 DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1313 AVDD.t445 AVDD.t443 AVDD.t444 AVDD.t370 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1314 AVDD.t442 AVDD.t440 AVDD.t441 AVDD.t374 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1315 a_2458_5328.t44 a_34666_7130.t14 a_32059_n4755.t1 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1316 a_2458_5328.t87 a_12760_n20342.t101 AVDD.t322 AVDD.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1317 a_32059_n4497.t1 casc_n.t169 a_32059_n4755.t10 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1318 a_2467_n30310.t77 casc_n.t170 Vop.t103 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1319 AVDD.t32 en.t1 a_32299_n29829# AVDD.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1.45e+11p ps=1.58e+06u w=500000u l=2e+06u
X1320 a_32059_n3351.t8 bias_n.t70 a_32059_n4497.t13 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1321 DGND Vom.t140 Vfold_bot_m.t41 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1322 AVDD.t439 AVDD.t437 AVDD.t438 AVDD.t370 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1323 DGND bias_var_n.t53 a_2467_n30310.t109 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1324 a_2467_n30310.t76 casc_n.t171 Vop.t102 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1325 Vxp.t60 casc_p.t334 a_1657_n21342.t161 AVDD.t161 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1326 DGND bias_n.t71 a_1659_n4497.t8 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1327 a_2458_5328.t20 Vinp.t46 Vxm.t17 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1328 DGND bias_var_n.t54 Vfold_bot_m.t112 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1329 a_1659_n4497.t51 casc_n.t172 Vxm.t46 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1330 DGND Vom.t141 a_2467_n30310.t49 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1331 a_1657_n21342.t67 a_1560_n22142.t117 AVDD.t863 AVDD.t161 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1332 a_32683_n30483# a_31928_n30483# DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X1333 a_1657_n21342.t66 a_1560_n22142.t118 AVDD.t864 AVDD.t161 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1334 DGND level_shifter_up_4.xb_hv.t9 bias_n.t3 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X1335 a_2458_6128.t18 a_12760_n20342.t102 AVDD.t323 AVDD.t85 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1336 DGND bias_var_n bias_var_n DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1337 a_2467_n29152.t9 casc_p.t335 a_32057_n17742.t15 AVDD.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1338 a_1657_n21342.t65 a_1560_n22142.t119 AVDD.t865 AVDD.t172 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1339 Vxp.t59 casc_p.t336 a_1657_n21342.t162 AVDD.t208 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1340 DGND DGND DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1341 DGND a_34499_n29829# level_shifter_up_0.x_hv.t0 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1342 a_32057_n21342.t1 bias_p.t91 a_32057_n22200.t7 AVDD.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1343 Vxp.t58 casc_p.t337 a_1657_n21342.t163 AVDD.t168 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1344 Vom.t17 casc_p.t338 a_2458_5328.t157 AVDD.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1345 Vxp.t35 Vinm.t44 a_2467_n30310.t39 AVDD.t46 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1346 DGND DGND DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1347 a_12857_n19016.t3 casc_p.t339 a_12857_n19542.t5 AVDD.t93 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1348 Vom.t16 casc_p.t340 a_2458_5328.t156 AVDD.t66 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1349 a_1657_n21342.t64 a_1560_n22142.t120 AVDD.t866 AVDD.t168 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1350 Vxp.t22 Vinp.t47 Vfold_bot_m.t22 AVDD.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1351 a_2467_n29152.t2 a_2370_n29452.t11 Vfold_bot_m.t19 AVDD.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1352 a_2458_5328.t88 a_12760_n20342.t103 AVDD.t324 AVDD.t66 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1353 AVDD.t436 AVDD.t434 AVDD.t435 AVDD.t381 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1354 DGND a_12857_n19016.t13 a_32059_n897.t2 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1355 casc_n.t9 casc_n.t7 casc_n.t8 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1356 a_32057_n13616.t37 a_34666_7130.t15 Vfold_bot_m.t119 AVDD.t344 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1357 AVDD.t433 AVDD.t431 AVDD.t432 AVDD.t401 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1358 a_2467_n30310.t75 casc_n.t173 Vop.t101 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1359 casc_n.t6 casc_n.t4 casc_n.t5 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1360 a_2458_5328.t89 a_12760_n20342.t104 AVDD.t325 AVDD.t68 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1361 a_12859_n2697# casc_n.t174 a_9060_4172.t2 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1362 a_1560_n22142.t9 casc_p.t341 a_12857_n15942.t4 AVDD.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1363 a_2458_6128.t76 bias_p.t92 AVDD.t149 AVDD.t148 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1364 DGND en.t2 a_32299_n29829# DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1365 a_2458_5328.t90 a_12760_n20342.t105 AVDD.t326 AVDD.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1366 AVDD.t430 AVDD.t428 AVDD.t429 AVDD.t401 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1367 DGND hyst[0].t3 a_36699_n29829# DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1368 a_2458_5328.t76 a_12760_n20342.t106 AVDD.t297 AVDD.t113 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1369 casc_p.t65 casc_p.t64 a_11257_n8742.t8 AVDD.t111 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1370 a_12857_n19542.t0 a_12760_n20342.t107 AVDD.t298 AVDD.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1371 Vxp.t57 casc_p.t342 a_1657_n21342.t164 AVDD.t155 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1372 Vfold_bot_m.t72 casc_n.t175 Vom.t111 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1373 a_23013_n25097.t18 casc_p.t343 a_32057_n21342.t10 AVDD.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1374 a_2467_n29152.t8 casc_p.t344 a_32057_n17742.t14 AVDD.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1375 a_2458_6128.t17 a_12760_n20342.t108 AVDD.t299 AVDD.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1376 a_32057_n9600.t7 level_shifter_up_5.xb_hv.t7 AVDD.t811 AVDD.t810 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1377 level_shifter_up_6.x_hv.t0 level_shifter_up_6.xb_hv AVDD.t340 AVDD.t339 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1378 a_32057_n21342.t0 bias_p.t93 a_32057_n22200.t6 AVDD.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1379 a_2467_n29152.t19 a_2370_n28652.t11 a_2467_n30310.t110 AVDD.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1380 Vxp.t56 casc_p.t345 a_1657_n21342.t165 AVDD.t157 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1381 Vxp.t55 casc_p.t346 a_1657_n21342.t166 AVDD.t172 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1382 a_2458_6128.t89 Vinm.t45 Vxm.t37 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1383 a_2458_6128.t90 Vinm.t46 Vxm.t38 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1384 DGND bias_n.t72 a_1659_n4497.t23 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1385 DGND.t530 Vom_stg2.t4 a_29758_4670.t4 DGND.t529 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1386 AVDD.t182 level_shifter_up_1.x_hv level_shifter_up_1.xb_hv.t0 AVDD.t181 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1387 Vom.t15 casc_p.t347 a_2458_5328.t155 AVDD.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1388 a_2458_6128.t16 a_12760_n20342.t109 AVDD.t300 AVDD.t74 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1389 DGND bias_n.t73 a_1659_n4497.t24 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1390 a_25696_11382.t14 level_shifter_up_8.x_hv.t6 a_2370_6628.t7 AVDD.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X1391 Vxp.t23 Vinp.t48 Vfold_bot_m.t23 AVDD.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1392 Vom.t14 casc_p.t348 a_2458_5328.t154 AVDD.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1393 AVDD.t828 level_shifter_up_0.xb_hv.t16 a_32057_n15000.t20 AVDD.t827 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1394 a_1657_n21342.t63 a_1560_n22142.t121 AVDD.t867 AVDD.t172 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1395 DGND DGND DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1396 a_2458_5328.t77 a_12760_n20342.t110 AVDD.t301 AVDD.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1397 DGND DGND DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1398 Vom.t13 casc_p.t349 a_2458_5328.t153 AVDD.t5 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1399 DGND bias_n.t74 a_1659_n4497.t25 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1400 AVDD.t427 AVDD.t425 AVDD.t426 AVDD.t374 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1401 a_2458_5328.t78 a_12760_n20342.t111 AVDD.t302 AVDD.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1402 a_2467_n30310.t74 casc_n.t176 Vop.t95 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1403 Vop.t10 casc_p.t350 a_2458_6128.t121 AVDD.t85 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1404 Vxp.t54 casc_p.t351 a_1657_n21342.t167 AVDD.t163 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1405 casc_p.t9 casc_p.t7 casc_p.t8 AVDD.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1406 Vom.t12 casc_p.t352 a_2458_5328.t152 AVDD.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1407 Vxp.t24 Vinp.t49 Vfold_bot_m.t24 AVDD.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1408 AVDD.t744 level_shifter_up_4.x_hv.t6 bias_p.t8 AVDD.t743 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X1409 a_2467_n29152.t7 casc_p.t353 a_32057_n17742.t13 AVDD.t48 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1410 a_2458_6128.t15 a_12760_n20342.t112 AVDD.t303 AVDD.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1411 DGND Vom.t142 a_2467_n30310.t48 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1412 a_2467_n30310.t73 casc_n.t177 Vop.t94 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1413 DGND bias_var_n.t56 Vfold_bot_m.t113 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1414 a_33657_n21342.t1 bias_p.t94 a_33657_n22200.t3 AVDD.t48 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1415 Vxp.t53 casc_p.t354 a_1657_n21342.t182 AVDD.t208 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1416 a_25030_4566.t0 a_25696_11382.t1 DGND sky130_fd_pr__res_high_po_2p85 l=3.192e+07u
X1417 a_1659_n4497.t50 casc_n.t178 Vxm.t47 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1418 Vom.t11 casc_p.t355 a_2458_5328.t125 AVDD.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1419 a_32057_n15000.t19 level_shifter_up_0.xb_hv.t17 AVDD.t830 AVDD.t829 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1420 AVDD.t424 AVDD.t422 AVDD.t423 AVDD.t401 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1421 Vom.t10 casc_p.t356 a_2458_5328.t124 AVDD.t68 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1422 DGND bias_n.t75 a_1659_n4497.t26 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1423 Vom.t9 casc_p.t357 a_2458_5328.t123 AVDD.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1424 DGND DGND DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1425 a_2458_5328.t79 a_12760_n20342.t113 AVDD.t304 AVDD.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1426 AVDD.t421 AVDD.t419 AVDD.t420 AVDD.t381 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1427 Vxp.t38 Vinm.t47 a_2467_n30310.t58 AVDD.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1428 Vxp.t52 casc_p.t358 a_1657_n21342.t183 AVDD.t166 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1429 a_2458_6128.t93 Vinm.t48 Vxm.t39 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1430 a_32448_11527# trim[1].t2 AVDD.t766 AVDD.t765 sky130_fd_pr__pfet_g5v0d10v5 ad=1.45e+11p pd=1.58e+06u as=0p ps=0u w=500000u l=2e+06u
X1431 AVDD.t418 AVDD.t416 AVDD.t417 AVDD.t366 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1432 bias_var_n.t2 casc_p.t359 a_12857_n17742.t4 AVDD.t111 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1433 DGND bias_n.t76 a_1659_n4497.t36 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1434 a_31928_n30483# trim[5].t3 DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1435 a_2458_6128.t77 bias_p.t95 AVDD.t150 AVDD.t148 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1436 AVDD.t415 AVDD.t413 AVDD.t414 AVDD.t111 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1437 Vfold_bot_m.t71 casc_n.t179 Vom.t110 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1438 DGND level_shifter_up_6.x_hv.t7 a_35259_2049# DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1439 a_2458_6128.t14 a_12760_n20342.t114 AVDD.t305 AVDD.t125 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1440 a_2458_6128.t13 a_12760_n20342.t115 AVDD.t306 AVDD.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1441 a_36859_903# casc_n.t180 a_25696_11382.t11 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=1.16e+12p pd=9.16e+06u as=0p ps=0u w=2e+06u l=1e+06u
X1442 DGND bias_n.t77 a_1659_n4497.t37 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1443 DGND DGND DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1444 casc_n.t0 ibias.t5 AVDD.t26 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1445 Vxp.t39 Vinm.t49 a_2467_n30310.t64 AVDD.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1446 a_2370_n29452.t1 level_shifter_up_3.x_hv.t9 res_p_bot.t2 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X1447 DGND bias_var_n.t57 Vfold_bot_m.t114 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1448 Vxp.t40 Vinm.t50 a_2467_n30310.t65 AVDD.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1449 DGND bias_n.t78 a_14459_n2697# DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1450 AVDD.t837 bias_stg2.t8 a_29757_7018.t5 AVDD.t760 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1451 Vxp.t51 casc_p.t360 a_1657_n21342.t184 AVDD.t194 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1452 a_2458_6128.t12 a_12760_n20342.t116 AVDD.t307 AVDD.t74 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1453 a_2467_n29152.t6 casc_p.t361 a_32057_n17742.t12 AVDD.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1454 a_2458_5328.t80 a_12760_n20342.t117 AVDD.t308 AVDD.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1455 Vop.t9 casc_p.t362 a_2458_6128.t120 AVDD.t103 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1456 a_1657_n21342.t62 a_1560_n22142.t122 AVDD.t868 AVDD.t194 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1457 DGND bias_n.t79 a_1659_n4497.t38 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1458 a_33657_n21342.t6 bias_p.t96 a_33657_n22200.t2 AVDD.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1459 a_32059_n3351.t1 level_shifter_up_0.x_hv.t9 DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1460 Vxp.t50 casc_p.t363 a_1657_n21342.t185 AVDD.t196 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1461 DGND a_32299_n29829# a_31859_n29829# DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X1462 Vop.t8 casc_p.t364 a_2458_6128.t119 AVDD.t85 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1463 a_1657_n21342.t61 a_1560_n22142.t123 AVDD.t869 AVDD.t196 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1464 a_2458_6128.t11 a_12760_n20342.t118 AVDD.t309 AVDD.t85 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1465 a_2467_n30310.t72 casc_n.t181 Vop.t93 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1466 a_2458_6128.t177 bias_p.t97 AVDD.t733 AVDD.t5 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1467 DGND DGND DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1468 DGND a_33203_11527# level_shifter_up_7.xb_hv DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X1469 a_2458_6128.t10 a_12760_n20342.t119 AVDD.t310 AVDD.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1470 a_2458_5328.t42 Vinp.t50 Vxm.t27 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1471 AVDD.t412 AVDD.t410 AVDD.t411 AVDD.t370 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1472 Vfold_bot_m.t70 casc_n.t182 Vom.t109 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1473 a_2467_n30310.t71 casc_n.t183 Vop.t92 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1474 a_32059_n897.t6 casc_n.t184 a_2458_6570.t6 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1475 Vfold_bot_m.t69 casc_n.t185 Vom.t108 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1476 a_2458_6128.t62 Vinm.t51 Vxm.t5 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1477 a_32059_n4755.t17 a_35086_7130.t18 a_2458_6128.t195 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1478 Vxp.t49 casc_p.t365 a_1657_n21342.t186 AVDD.t161 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1479 DGND bias_var_n.t58 a_2467_n30310.t13 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1480 a_2458_5328.t81 a_12760_n20342.t120 AVDD.t311 AVDD.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1481 casc_p.t6 casc_p.t4 casc_p.t5 AVDD.t93 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1482 a_1659_n4497.t49 casc_n.t186 Vxm.t48 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1483 AVDD.t409 AVDD.t407 AVDD.t408 AVDD.t401 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1484 a_2458_5328.t72 a_12760_n20342.t121 AVDD.t289 AVDD.t113 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1485 Vom.t8 casc_p.t366 a_2458_5328.t122 AVDD.t68 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1486 AVDD.t406 AVDD.t404 AVDD.t405 AVDD.t394 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1487 DGND bias_n.t80 a_1659_n4497.t31 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1488 AVDD.t403 AVDD.t400 AVDD.t402 AVDD.t401 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1489 a_31003_11527# a_30248_11527# DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=500000u
X1490 a_2370_6628.t6 level_shifter_up_8.x_hv.t7 a_25696_11382.t13 AVDD.t28 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X1491 a_32299_n29829# en.t3 DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1492 Vop.t7 casc_p.t367 a_2458_6128.t150 AVDD.t125 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1493 Vxp.t48 casc_p.t368 a_1657_n21342.t187 AVDD.t155 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1494 a_32057_n13616.t36 a_35086_7130.t19 a_2467_n30310.t111 AVDD.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1495 Vom.t7 casc_p.t369 a_2458_5328.t121 AVDD.t66 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1496 a_23013_n25097.t17 casc_p.t370 a_32057_n21342.t9 AVDD.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1497 a_35259_903# casc_n.t187 a_23032_4566.t9 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1498 DGND DGND DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1499 a_2458_6128.t178 bias_p.t98 AVDD.t734 AVDD.t148 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1500 a_2458_5328.t180 bias_p.t99 AVDD.t735 AVDD.t15 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1501 AVDD.t813 level_shifter_up_5.xb_hv.t8 a_32057_n9600.t6 AVDD.t812 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1502 DGND DGND DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1503 Vxp.t47 casc_p.t371 a_1657_n21342.t188 AVDD.t157 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1504 a_12859_n4497# casc_n.t188 a_12859_n4755# DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1505 a_34666_7130.t1 a_31098_4670.t8 DVDD.t9 DVDD.t8 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1506 a_27926_9740.t4 level_shifter_up_7.x_hv.t8 a_23032_4566.t2 AVDD.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X1507 a_12857_n19016.t2 casc_p.t372 a_12857_n19542.t4 AVDD.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1508 DGND Vom.t143 a_2467_n30310.t47 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1509 DGND Vom.t144 a_2467_n30310.t46 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1510 a_32059_n3351.t2 level_shifter_up_0.x_hv.t10 DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1511 a_32059_n4755.t25 a_34666_7130.t16 a_2458_5328.t198 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1512 AVDD.t399 AVDD.t397 AVDD.t398 AVDD.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1513 a_11259_2049# ibias.t6 bias_n.t0 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1514 a_1659_n4497.t48 casc_n.t189 Vxm.t49 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1515 a_2458_5328.t73 a_12760_n20342.t122 AVDD.t290 AVDD.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1516 a_2458_5328.t16 Vinp.t51 Vxm.t13 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1517 a_23013_n25097.t8 casc_p.t373 a_32057_n21342.t8 AVDD.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1518 DGND bias_n.t81 a_1659_n4497.t32 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1519 a_9060_4530.t5 Vinp.t52 a_9060_4172.t1 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1520 a_2458_6128.t63 Vinm.t52 Vxm.t6 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1521 a_32057_n15000.t18 level_shifter_up_0.xb_hv.t18 AVDD.t832 AVDD.t831 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1522 Vxp.t46 casc_p.t374 a_1657_n21342.t189 AVDD.t172 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1523 a_1659_n4497.t47 casc_n.t190 Vxm.t50 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1524 Vop.t6 casc_p.t375 a_2458_6128.t149 AVDD.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1525 res_p_bot.t14 casc_p.t376 a_11257_n21342# AVDD.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1526 AVDD.t396 AVDD.t393 AVDD.t395 AVDD.t394 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1527 level_shifter_up_2.x_hv level_shifter_up_2.xb_hv.t10 AVDD.t708 AVDD.t707 sky130_fd_pr__pfet_g5v0d10v5 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=500000u
X1528 Vom.t6 casc_p.t377 a_2458_5328.t120 AVDD.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1529 Vxp.t17 Vinp.t53 Vfold_bot_m.t9 AVDD.t46 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1530 AVDD.t30 level_shifter_up_8.x_hv.t8 level_shifter_up_8.xb_hv.t0 AVDD.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1531 Vxp.t45 casc_p.t378 a_1657_n21342.t190 AVDD.t163 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1532 Vxp.t18 Vinp.t54 Vfold_bot_m.t10 AVDD.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1533 level_shifter_up_5.xb_hv.t0 level_shifter_up_5.x_hv.t5 AVDD.t267 AVDD.t266 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1534 DGND bias_n.t82 a_1659_n4497.t33 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1535 a_2458_5328.t74 a_12760_n20342.t123 AVDD.t291 AVDD.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1536 Vxp.t5 Vinm.t53 a_2467_n30310.t2 AVDD.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1537 AVDD.t392 AVDD.t390 AVDD.t391 AVDD.t374 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1538 a_2458_6128.t9 a_12760_n20342.t124 AVDD.t292 AVDD.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1539 a_2370_6628.t2 level_shifter_up_8.xb_hv.t9 a_23032_4566.t4 AVDD.t722 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X1540 a_32059_n4497.t0 casc_n.t191 a_32059_n4755.t9 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1541 a_33659_n2697.t0 casc_n.t192 a_32059_n4755.t5 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1542 a_32448_11527# trim[1].t3 DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1543 Vfold_bot_m.t68 casc_n.t193 Vom.t107 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1544 Vfold_bot_m.t67 casc_n.t194 Vom.t94 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1545 DGND bias_n.t83 a_1659_n4497.t34 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1546 a_11259_n2697# casc_n.t195 bias_p.t9 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1547 DGND trim[3].t3 a_36328_n30483# DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1548 Vom.t5 casc_p.t379 a_2458_5328.t119 AVDD.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1549 a_32059_n4755.t26 a_34666_7130.t17 a_2458_5328.t199 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1550 a_33203_11527# a_32448_11527# AVDD.t55 AVDD.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=500000u
X1551 DGND a_37083_n30483# level_shifter_up_1.xb_hv DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X1552 a_2458_5328.t75 a_12760_n20342.t125 AVDD.t293 AVDD.t113 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1553 a_2458_6128.t179 bias_p.t100 AVDD.t736 AVDD.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1554 Vfold_bot_m.t66 casc_n.t196 Vom.t93 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1555 res_p_bot.t1 level_shifter_up_3.x_hv.t10 a_2370_n29452.t2 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X1556 a_2467_n30310.t70 casc_n.t197 Vop.t91 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1557 Vxp.t44 casc_p.t380 a_1657_n21342.t191 AVDD.t166 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1558 a_32057_n13616.t11 casc_p.t381 a_32057_n8742.t11 AVDD.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1559 Vop.t5 casc_p.t382 a_2458_6128.t148 AVDD.t125 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1560 Vxp.t43 casc_p.t383 a_1657_n21342.t0 AVDD.t208 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1561 Vop.t4 casc_p.t384 a_2458_6128.t147 AVDD.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1562 Vxp.t42 casc_p.t385 a_1657_n21342.t1 AVDD.t203 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1563 a_32059_2049.t0 level_shifter_up_7.x_hv.t9 DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1564 Vom.t4 casc_p.t386 a_2458_5328.t118 AVDD.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1565 Vop.t3 casc_p.t387 a_2458_6128.t146 AVDD.t125 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1566 DGND DGND DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1567 a_1657_n21342.t60 a_1560_n22142.t124 AVDD.t870 AVDD.t208 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1568 a_1657_n21342.t59 a_1560_n22142.t125 AVDD.t871 AVDD.t203 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1569 AVDD.t389 AVDD.t387 AVDD.t388 AVDD.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1570 DGND bias_n.t84 a_1659_n4497.t16 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1571 a_2458_5328.t194 Vinp.t55 Vxm.t101 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1572 DGND bias_var_n.t59 Vfold_bot_m.t11 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1573 a_2458_6128.t8 a_12760_n20342.t126 AVDD.t294 AVDD.t125 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1574 DGND DGND DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1575 DGND DGND DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1576 a_2458_5328.t181 bias_p.t101 AVDD.t737 AVDD.t15 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1577 AVDD.t386 AVDD.t384 AVDD.t385 AVDD.t381 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1578 DGND a_12857_n19016.t4 a_12857_n19016.t5 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1579 Vom.t3 casc_p.t388 a_2458_5328.t117 AVDD.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1580 a_37477_903# casc_n.t198 bias_stg2.t0 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1581 a_31098_4670.t3 level_shifter_up_4.xb_hv.t10 DGND.t534 DGND.t533 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1582 AVDD.t383 AVDD.t380 AVDD.t382 AVDD.t381 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1583 Vfold_bot_m.t63 a_34666_7130.t18 a_32057_n13616.t32 AVDD.t344 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1584 Vop.t2 casc_p.t389 a_2458_6128.t145 AVDD.t103 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1585 Vxp.t146 Vinp.t56 Vfold_bot_m.t115 AVDD.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1586 AVDD.t379 AVDD.t377 AVDD.t378 AVDD.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1587 Vfold_bot_m.t64 a_34666_7130.t19 a_32057_n13616.t33 AVDD.t344 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1588 DGND bias_n.t85 a_36859_903# DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1589 a_2458_6128.t7 a_12760_n20342.t127 AVDD.t295 AVDD.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1590 DGND bias_var_n.t60 a_2467_n30310.t14 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1591 DGND DGND DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1592 DGND bias_var_n.t61 Vfold_bot_m.t12 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1593 a_14459_n4755.t1 bias_n.t86 a_14459_n4209# DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1594 a_35259_2049# bias_n.t87 a_35259_903# DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1595 a_1659_n4497.t46 casc_n.t199 Vxm.t91 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1596 a_2458_6128.t70 Vinm.t54 Vxm.t19 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1597 Vop.t1 casc_p.t390 a_2458_6128.t144 AVDD.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1598 Vom.t2 casc_p.t391 a_2458_5328.t116 AVDD.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1599 AVDD.t376 AVDD.t373 AVDD.t375 AVDD.t374 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1600 DGND bias_var_n.t62 Vfold_bot_m.t57 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1601 a_2458_6128.t6 a_12760_n20342.t128 AVDD.t296 AVDD.t74 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1602 DVDD.t1 a_29758_4670.t6 a_31098_4670.t1 DVDD.t0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1603 AVDD.t372 AVDD.t369 AVDD.t371 AVDD.t370 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1604 Vxp.t41 casc_p.t392 a_1657_n21342.t2 AVDD.t161 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1605 a_2458_6128.t71 Vinm.t55 Vxm.t20 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1606 a_2458_6128.t72 Vinm.t56 Vxm.t21 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1607 Vop.t0 casc_p.t393 a_2458_6128.t94 AVDD.t85 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1608 DGND DGND DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1609 AVDD.t368 AVDD.t365 AVDD.t367 AVDD.t366 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1610 DGND DGND DGND DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=8e+06u l=1.5e+06u
X1611 a_2458_6128.t180 bias_p.t102 AVDD.t738 AVDD.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1612 Vfold_bot_m.t65 casc_n.t200 Vom.t92 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1613 a_2467_n30310.t69 casc_n.t201 Vop.t80 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1614 a_33659_n1551.t2 bias_n.t88 a_33659_n2697.t3 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1615 DGND bias_var_n.t63 a_2467_n30310.t61 DGND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1616 Vom.t1 casc_p.t394 a_2458_5328.t115 AVDD.t15 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1617 a_25696_11382.t12 level_shifter_up_8.x_hv.t9 a_2370_6628.t5 AVDD.t61 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X1618 Vom.t0 casc_p.t395 a_2458_5328.t114 AVDD.t66 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
R0 casc_n.n192 casc_n.t16 48.206
R1 casc_n.n0 casc_n.t34 48.206
R2 casc_n.n47 casc_n.t28 48.206
R3 casc_n.n50 casc_n.t19 48.206
R4 casc_n.n89 casc_n.t31 48.206
R5 casc_n.n86 casc_n.t25 48.206
R6 casc_n.n83 casc_n.t10 48.206
R7 casc_n.n80 casc_n.t4 48.206
R8 casc_n.n31 casc_n.t22 48.206
R9 casc_n.n28 casc_n.t13 48.206
R10 casc_n.n51 casc_n.t198 24.574
R11 casc_n.n148 casc_n.t92 24.574
R12 casc_n.n1 casc_n.t88 24.574
R13 casc_n.n179 casc_n.t56 24.573
R14 casc_n.n34 casc_n.t87 24.573
R15 casc_n.n91 casc_n.t145 24.573
R16 casc_n.n135 casc_n.t66 24.573
R17 casc_n.n105 casc_n.t7 24.106
R18 casc_n.n103 casc_n.t126 23.982
R19 casc_n.n147 casc_n.t46 23.982
R20 casc_n.n179 casc_n.t136 23.982
R21 casc_n.n180 casc_n.t107 23.982
R22 casc_n.n181 casc_n.t38 23.982
R23 casc_n.n182 casc_n.t178 23.982
R24 casc_n.n183 casc_n.t85 23.982
R25 casc_n.n184 casc_n.t68 23.982
R26 casc_n.n185 casc_n.t151 23.982
R27 casc_n.n186 casc_n.t123 23.982
R28 casc_n.n187 casc_n.t48 23.982
R29 casc_n.n188 casc_n.t190 23.982
R30 casc_n.n189 casc_n.t143 23.982
R31 casc_n.n34 casc_n.t103 23.982
R32 casc_n.n35 casc_n.t44 23.982
R33 casc_n.n36 casc_n.t96 23.982
R34 casc_n.n37 casc_n.t39 23.982
R35 casc_n.n38 casc_n.t54 23.982
R36 casc_n.n39 casc_n.t161 23.982
R37 casc_n.n40 casc_n.t168 23.982
R38 casc_n.n41 casc_n.t104 23.982
R39 casc_n.n42 casc_n.t163 23.982
R40 casc_n.n43 casc_n.t97 23.982
R41 casc_n.n44 casc_n.t110 23.982
R42 casc_n.n77 casc_n.t115 23.982
R43 casc_n.n76 casc_n.t167 23.982
R44 casc_n.n75 casc_n.t102 23.982
R45 casc_n.n74 casc_n.t124 23.982
R46 casc_n.n73 casc_n.t59 23.982
R47 casc_n.n72 casc_n.t116 23.982
R48 casc_n.n71 casc_n.t105 23.982
R49 casc_n.n70 casc_n.t127 23.982
R50 casc_n.n69 casc_n.t62 23.982
R51 casc_n.n68 casc_n.t74 23.982
R52 casc_n.n67 casc_n.t176 23.982
R53 casc_n.n66 casc_n.t69 23.982
R54 casc_n.n65 casc_n.t171 23.982
R55 casc_n.n64 casc_n.t181 23.982
R56 casc_n.n63 casc_n.t130 23.982
R57 casc_n.n62 casc_n.t177 23.982
R58 casc_n.n61 casc_n.t118 23.982
R59 casc_n.n60 casc_n.t137 23.982
R60 casc_n.n59 casc_n.t131 23.982
R61 casc_n.n58 casc_n.t146 23.982
R62 casc_n.n57 casc_n.t78 23.982
R63 casc_n.n56 casc_n.t140 23.982
R64 casc_n.n55 casc_n.t73 23.982
R65 casc_n.n54 casc_n.t83 23.982
R66 casc_n.n53 casc_n.t187 23.982
R67 casc_n.n52 casc_n.t79 23.982
R68 casc_n.n51 casc_n.t180 23.982
R69 casc_n.n91 casc_n.t47 23.982
R70 casc_n.n92 casc_n.t189 23.982
R71 casc_n.n93 casc_n.t122 23.982
R72 casc_n.n94 casc_n.t91 23.982
R73 casc_n.n95 casc_n.t172 23.982
R74 casc_n.n96 casc_n.t155 23.982
R75 casc_n.n97 casc_n.t61 23.982
R76 casc_n.n98 casc_n.t37 23.982
R77 casc_n.n99 casc_n.t135 23.982
R78 casc_n.n100 casc_n.t106 23.982
R79 casc_n.n101 casc_n.t51 23.982
R80 casc_n.n102 casc_n.t195 23.982
R81 casc_n.n134 casc_n.t95 23.982
R82 casc_n.n133 casc_n.t174 23.982
R83 casc_n.n132 casc_n.t159 23.982
R84 casc_n.n131 casc_n.t64 23.982
R85 casc_n.n130 casc_n.t41 23.982
R86 casc_n.n129 casc_n.t139 23.982
R87 casc_n.n128 casc_n.t112 23.982
R88 casc_n.n127 casc_n.t183 23.982
R89 casc_n.n126 casc_n.t164 23.982
R90 casc_n.n125 casc_n.t86 23.982
R91 casc_n.n124 casc_n.t149 23.982
R92 casc_n.n123 casc_n.t50 23.982
R93 casc_n.n122 casc_n.t194 23.982
R94 casc_n.n121 casc_n.t99 23.982
R95 casc_n.n120 casc_n.t81 23.982
R96 casc_n.n119 casc_n.t173 23.982
R97 casc_n.n118 casc_n.t157 23.982
R98 casc_n.n117 casc_n.t63 23.982
R99 casc_n.n116 casc_n.t40 23.982
R100 casc_n.n115 casc_n.t138 23.982
R101 casc_n.n114 casc_n.t109 23.982
R102 casc_n.n113 casc_n.t182 23.982
R103 casc_n.n112 casc_n.t71 23.982
R104 casc_n.n111 casc_n.t152 23.982
R105 casc_n.n110 casc_n.t125 23.982
R106 casc_n.n109 casc_n.t49 23.982
R107 casc_n.n108 casc_n.t192 23.982
R108 casc_n.n107 casc_n.t98 23.982
R109 casc_n.n106 casc_n.t80 23.982
R110 casc_n.n135 casc_n.t144 23.982
R111 casc_n.n136 casc_n.t117 23.982
R112 casc_n.n137 casc_n.t43 23.982
R113 casc_n.n138 casc_n.t186 23.982
R114 casc_n.n139 casc_n.t90 23.982
R115 casc_n.n140 casc_n.t75 23.982
R116 casc_n.n141 casc_n.t154 23.982
R117 casc_n.n142 casc_n.t132 23.982
R118 casc_n.n143 casc_n.t55 23.982
R119 casc_n.n144 casc_n.t199 23.982
R120 casc_n.n145 casc_n.t150 23.982
R121 casc_n.n146 casc_n.t121 23.982
R122 casc_n.n176 casc_n.t188 23.982
R123 casc_n.n175 casc_n.t94 23.982
R124 casc_n.n174 casc_n.t77 23.982
R125 casc_n.n173 casc_n.t158 23.982
R126 casc_n.n172 casc_n.t134 23.982
R127 casc_n.n171 casc_n.t58 23.982
R128 casc_n.n170 casc_n.t201 23.982
R129 casc_n.n169 casc_n.t111 23.982
R130 casc_n.n168 casc_n.t84 23.982
R131 casc_n.n167 casc_n.t179 23.982
R132 casc_n.n166 casc_n.t67 23.982
R133 casc_n.n165 casc_n.t148 23.982
R134 casc_n.n164 casc_n.t120 23.982
R135 casc_n.n163 casc_n.t193 23.982
R136 casc_n.n162 casc_n.t170 23.982
R137 casc_n.n161 casc_n.t93 23.982
R138 casc_n.n160 casc_n.t76 23.982
R139 casc_n.n159 casc_n.t156 23.982
R140 casc_n.n158 casc_n.t133 23.982
R141 casc_n.n157 casc_n.t57 23.982
R142 casc_n.n156 casc_n.t200 23.982
R143 casc_n.n155 casc_n.t108 23.982
R144 casc_n.n154 casc_n.t162 23.982
R145 casc_n.n153 casc_n.t70 23.982
R146 casc_n.n152 casc_n.t45 23.982
R147 casc_n.n151 casc_n.t147 23.982
R148 casc_n.n150 casc_n.t119 23.982
R149 casc_n.n149 casc_n.t191 23.982
R150 casc_n.n148 casc_n.t169 23.982
R151 casc_n.n25 casc_n.t129 23.982
R152 casc_n.n24 casc_n.t53 23.982
R153 casc_n.n23 casc_n.t197 23.982
R154 casc_n.n22 casc_n.t101 23.982
R155 casc_n.n21 casc_n.t82 23.982
R156 casc_n.n20 casc_n.t175 23.982
R157 casc_n.n19 casc_n.t60 23.982
R158 casc_n.n18 casc_n.t142 23.982
R159 casc_n.n17 casc_n.t114 23.982
R160 casc_n.n16 casc_n.t185 23.982
R161 casc_n.n15 casc_n.t166 23.982
R162 casc_n.n14 casc_n.t89 23.982
R163 casc_n.n13 casc_n.t72 23.982
R164 casc_n.n12 casc_n.t153 23.982
R165 casc_n.n11 casc_n.t128 23.982
R166 casc_n.n10 casc_n.t52 23.982
R167 casc_n.n9 casc_n.t196 23.982
R168 casc_n.n8 casc_n.t100 23.982
R169 casc_n.n7 casc_n.t160 23.982
R170 casc_n.n6 casc_n.t65 23.982
R171 casc_n.n5 casc_n.t42 23.982
R172 casc_n.n4 casc_n.t141 23.982
R173 casc_n.n3 casc_n.t113 23.982
R174 casc_n.n2 casc_n.t184 23.982
R175 casc_n.n1 casc_n.t165 23.982
R176 casc_n.n191 casc_n.t17 8.293
R177 casc_n.n191 casc_n.t18 8.292
R178 casc_n.n27 casc_n.t14 8.291
R179 casc_n.n194 casc_n.t35 8.291
R180 casc_n.n194 casc_n.t36 8.289
R181 casc_n.n27 casc_n.t15 8.289
R182 casc_n.n104 casc_n.t9 8.274
R183 casc_n.n104 casc_n.t8 8.274
R184 casc_n.n49 casc_n.t20 8.27
R185 casc_n.n49 casc_n.t21 8.27
R186 casc_n.n79 casc_n.t5 8.27
R187 casc_n.n79 casc_n.t6 8.27
R188 casc_n.n85 casc_n.t26 8.27
R189 casc_n.n85 casc_n.t27 8.27
R190 casc_n.n46 casc_n.t29 8.267
R191 casc_n.n46 casc_n.t30 8.267
R192 casc_n.n82 casc_n.t11 8.267
R193 casc_n.n82 casc_n.t12 8.267
R194 casc_n.n88 casc_n.t32 8.267
R195 casc_n.n88 casc_n.t33 8.267
R196 casc_n.n30 casc_n.t23 8.267
R197 casc_n.n30 casc_n.t24 8.267
R198 casc_n.n33 casc_n.t0 8.266
R199 casc_n.n33 casc_n.t3 8.266
R200 casc_n.n32 casc_n.t2 8.266
R201 casc_n.n32 casc_n.t1 8.266
R202 casc_n.n178 casc_n.n177 2.199
R203 casc_n.n0 casc_n.n178 2.177
R204 casc_n.n196 casc_n.n90 1.867
R205 casc_n.n43 casc_n.n42 0.942
R206 casc_n.n41 casc_n.n40 0.942
R207 casc_n.n39 casc_n.n38 0.942
R208 casc_n.n37 casc_n.n36 0.942
R209 casc_n.n35 casc_n.n34 0.942
R210 casc_n.n52 casc_n.n51 0.942
R211 casc_n.n54 casc_n.n53 0.942
R212 casc_n.n56 casc_n.n55 0.942
R213 casc_n.n58 casc_n.n57 0.942
R214 casc_n.n60 casc_n.n59 0.942
R215 casc_n.n62 casc_n.n61 0.942
R216 casc_n.n64 casc_n.n63 0.942
R217 casc_n.n66 casc_n.n65 0.942
R218 casc_n.n68 casc_n.n67 0.942
R219 casc_n.n70 casc_n.n69 0.942
R220 casc_n.n72 casc_n.n71 0.942
R221 casc_n.n74 casc_n.n73 0.942
R222 casc_n.n76 casc_n.n75 0.942
R223 casc_n.n102 casc_n.n101 0.942
R224 casc_n.n100 casc_n.n99 0.942
R225 casc_n.n98 casc_n.n97 0.942
R226 casc_n.n96 casc_n.n95 0.942
R227 casc_n.n94 casc_n.n93 0.942
R228 casc_n.n92 casc_n.n91 0.942
R229 casc_n.n107 casc_n.n106 0.942
R230 casc_n.n109 casc_n.n108 0.942
R231 casc_n.n111 casc_n.n110 0.942
R232 casc_n.n113 casc_n.n112 0.942
R233 casc_n.n115 casc_n.n114 0.942
R234 casc_n.n117 casc_n.n116 0.942
R235 casc_n.n119 casc_n.n118 0.942
R236 casc_n.n121 casc_n.n120 0.942
R237 casc_n.n123 casc_n.n122 0.942
R238 casc_n.n125 casc_n.n124 0.942
R239 casc_n.n127 casc_n.n126 0.942
R240 casc_n.n129 casc_n.n128 0.942
R241 casc_n.n131 casc_n.n130 0.942
R242 casc_n.n133 casc_n.n132 0.942
R243 casc_n.n146 casc_n.n145 0.942
R244 casc_n.n144 casc_n.n143 0.942
R245 casc_n.n142 casc_n.n141 0.942
R246 casc_n.n140 casc_n.n139 0.942
R247 casc_n.n138 casc_n.n137 0.942
R248 casc_n.n136 casc_n.n135 0.942
R249 casc_n.n149 casc_n.n148 0.942
R250 casc_n.n151 casc_n.n150 0.942
R251 casc_n.n153 casc_n.n152 0.942
R252 casc_n.n155 casc_n.n154 0.942
R253 casc_n.n157 casc_n.n156 0.942
R254 casc_n.n159 casc_n.n158 0.942
R255 casc_n.n161 casc_n.n160 0.942
R256 casc_n.n163 casc_n.n162 0.942
R257 casc_n.n165 casc_n.n164 0.942
R258 casc_n.n167 casc_n.n166 0.942
R259 casc_n.n169 casc_n.n168 0.942
R260 casc_n.n171 casc_n.n170 0.942
R261 casc_n.n173 casc_n.n172 0.942
R262 casc_n.n175 casc_n.n174 0.942
R263 casc_n.n2 casc_n.n1 0.942
R264 casc_n.n4 casc_n.n3 0.942
R265 casc_n.n6 casc_n.n5 0.942
R266 casc_n.n8 casc_n.n7 0.942
R267 casc_n.n10 casc_n.n9 0.942
R268 casc_n.n12 casc_n.n11 0.942
R269 casc_n.n14 casc_n.n13 0.942
R270 casc_n.n16 casc_n.n15 0.942
R271 casc_n.n18 casc_n.n17 0.942
R272 casc_n.n20 casc_n.n19 0.942
R273 casc_n.n22 casc_n.n21 0.942
R274 casc_n.n24 casc_n.n23 0.942
R275 casc_n.n188 casc_n.n187 0.942
R276 casc_n.n186 casc_n.n185 0.942
R277 casc_n.n184 casc_n.n183 0.942
R278 casc_n.n182 casc_n.n181 0.942
R279 casc_n.n180 casc_n.n179 0.942
R280 casc_n.n0 casc_n.n195 0.75
R281 casc_n.n45 casc_n.n44 0.697
R282 casc_n.n78 casc_n.n77 0.697
R283 casc_n.n26 casc_n.n25 0.697
R284 casc_n.n190 casc_n.n189 0.697
R285 casc_n.n32 casc_n.n31 0.689
R286 casc_n.n44 casc_n.n43 0.592
R287 casc_n.n42 casc_n.n41 0.592
R288 casc_n.n40 casc_n.n39 0.592
R289 casc_n.n38 casc_n.n37 0.592
R290 casc_n.n36 casc_n.n35 0.592
R291 casc_n.n53 casc_n.n52 0.592
R292 casc_n.n55 casc_n.n54 0.592
R293 casc_n.n57 casc_n.n56 0.592
R294 casc_n.n59 casc_n.n58 0.592
R295 casc_n.n61 casc_n.n60 0.592
R296 casc_n.n63 casc_n.n62 0.592
R297 casc_n.n65 casc_n.n64 0.592
R298 casc_n.n67 casc_n.n66 0.592
R299 casc_n.n69 casc_n.n68 0.592
R300 casc_n.n71 casc_n.n70 0.592
R301 casc_n.n73 casc_n.n72 0.592
R302 casc_n.n75 casc_n.n74 0.592
R303 casc_n.n77 casc_n.n76 0.592
R304 casc_n.n101 casc_n.n100 0.592
R305 casc_n.n99 casc_n.n98 0.592
R306 casc_n.n97 casc_n.n96 0.592
R307 casc_n.n95 casc_n.n94 0.592
R308 casc_n.n93 casc_n.n92 0.592
R309 casc_n.n108 casc_n.n107 0.592
R310 casc_n.n110 casc_n.n109 0.592
R311 casc_n.n112 casc_n.n111 0.592
R312 casc_n.n114 casc_n.n113 0.592
R313 casc_n.n116 casc_n.n115 0.592
R314 casc_n.n118 casc_n.n117 0.592
R315 casc_n.n120 casc_n.n119 0.592
R316 casc_n.n122 casc_n.n121 0.592
R317 casc_n.n124 casc_n.n123 0.592
R318 casc_n.n126 casc_n.n125 0.592
R319 casc_n.n128 casc_n.n127 0.592
R320 casc_n.n130 casc_n.n129 0.592
R321 casc_n.n132 casc_n.n131 0.592
R322 casc_n.n134 casc_n.n133 0.592
R323 casc_n.n145 casc_n.n144 0.592
R324 casc_n.n143 casc_n.n142 0.592
R325 casc_n.n141 casc_n.n140 0.592
R326 casc_n.n139 casc_n.n138 0.592
R327 casc_n.n137 casc_n.n136 0.592
R328 casc_n.n150 casc_n.n149 0.592
R329 casc_n.n152 casc_n.n151 0.592
R330 casc_n.n154 casc_n.n153 0.592
R331 casc_n.n156 casc_n.n155 0.592
R332 casc_n.n158 casc_n.n157 0.592
R333 casc_n.n160 casc_n.n159 0.592
R334 casc_n.n162 casc_n.n161 0.592
R335 casc_n.n164 casc_n.n163 0.592
R336 casc_n.n166 casc_n.n165 0.592
R337 casc_n.n168 casc_n.n167 0.592
R338 casc_n.n170 casc_n.n169 0.592
R339 casc_n.n172 casc_n.n171 0.592
R340 casc_n.n174 casc_n.n173 0.592
R341 casc_n.n176 casc_n.n175 0.592
R342 casc_n.n3 casc_n.n2 0.592
R343 casc_n.n5 casc_n.n4 0.592
R344 casc_n.n7 casc_n.n6 0.592
R345 casc_n.n9 casc_n.n8 0.592
R346 casc_n.n11 casc_n.n10 0.592
R347 casc_n.n13 casc_n.n12 0.592
R348 casc_n.n15 casc_n.n14 0.592
R349 casc_n.n17 casc_n.n16 0.592
R350 casc_n.n19 casc_n.n18 0.592
R351 casc_n.n21 casc_n.n20 0.592
R352 casc_n.n23 casc_n.n22 0.592
R353 casc_n.n25 casc_n.n24 0.592
R354 casc_n.n189 casc_n.n188 0.592
R355 casc_n.n187 casc_n.n186 0.592
R356 casc_n.n185 casc_n.n184 0.592
R357 casc_n.n183 casc_n.n182 0.592
R358 casc_n.n181 casc_n.n180 0.592
R359 casc_n.n103 casc_n.n102 0.591
R360 casc_n.n147 casc_n.n146 0.591
R361 casc_n.n178 casc_n.n134 0.579
R362 casc_n.n177 casc_n.n176 0.579
R363 casc_n.n106 casc_n.n105 0.467
R364 casc_n.n84 casc_n.n83 0.453
R365 casc_n casc_n.n196 0.421
R366 casc_n.n33 casc_n.n32 0.365
R367 casc_n.n178 casc_n.n103 0.348
R368 casc_n.n177 casc_n.n147 0.348
R369 casc_n.n90 casc_n.n89 0.335
R370 casc_n.n192 casc_n.n191 0.263
R371 casc_n.n27 casc_n.n26 0.261
R372 casc_n.n49 casc_n.n48 0.248
R373 casc_n.n80 casc_n.n79 0.248
R374 casc_n.n86 casc_n.n85 0.248
R375 casc_n.n46 casc_n.n45 0.246
R376 casc_n.n83 casc_n.n82 0.246
R377 casc_n.n89 casc_n.n88 0.246
R378 casc_n.n31 casc_n.n30 0.246
R379 casc_n.n47 casc_n.n46 0.244
R380 casc_n.n82 casc_n.n81 0.244
R381 casc_n.n88 casc_n.n87 0.244
R382 casc_n.n30 casc_n.n29 0.244
R383 casc_n.n79 casc_n.n78 0.242
R384 casc_n.n85 casc_n.n84 0.242
R385 casc_n.n50 casc_n.n49 0.24
R386 casc_n.n195 casc_n.n194 0.239
R387 casc_n.n28 casc_n.n27 0.228
R388 casc_n.n194 casc_n.n193 0.228
R389 casc_n.n191 casc_n.n190 0.226
R390 casc_n.n196 casc_n.n0 0.177
R391 casc_n.n105 casc_n.n104 0.12
R392 casc_n.n90 casc_n.n50 0.105
R393 casc_n.n48 casc_n.n47 0.103
R394 casc_n.n81 casc_n.n80 0.103
R395 casc_n.n87 casc_n.n86 0.103
R396 casc_n.n29 casc_n.n28 0.103
R397 casc_n.n193 casc_n.n192 0.103
R398 casc_n casc_n.n33 0.028
R399 Vxm.n6 Vxm.t52 8.857
R400 Vxm.n3 Vxm.t66 8.857
R401 Vxm.n9 Vxm.t61 8.857
R402 Vxm.n1 Vxm.t55 8.857
R403 Vxm.n0 Vxm.t88 8.266
R404 Vxm.n42 Vxm.t76 8.266
R405 Vxm.n43 Vxm.t57 8.266
R406 Vxm.n53 Vxm.t65 8.266
R407 Vxm.n54 Vxm.t80 8.266
R408 Vxm.n126 Vxm.t48 8.266
R409 Vxm.n128 Vxm.t70 8.266
R410 Vxm.n127 Vxm.t62 8.266
R411 Vxm.n116 Vxm.t53 8.266
R412 Vxm.n115 Vxm.t63 8.266
R413 Vxm.n122 Vxm.t79 8.266
R414 Vxm.n123 Vxm.t84 8.266
R415 Vxm.n139 Vxm.t71 8.266
R416 Vxm.n140 Vxm.t82 8.266
R417 Vxm.n138 Vxm.t69 8.266
R418 Vxm.n63 Vxm.t87 8.266
R419 Vxm.n62 Vxm.t51 8.266
R420 Vxm.n50 Vxm.t93 8.266
R421 Vxm.n40 Vxm.t90 8.266
R422 Vxm.n56 Vxm.t58 8.266
R423 Vxm.n57 Vxm.t46 8.266
R424 Vxm.n130 Vxm.t81 8.266
R425 Vxm.n132 Vxm.t74 8.266
R426 Vxm.n131 Vxm.t49 8.266
R427 Vxm.n114 Vxm.t59 8.266
R428 Vxm.n113 Vxm.t89 8.266
R429 Vxm.n135 Vxm.t60 8.266
R430 Vxm.n136 Vxm.t68 8.266
R431 Vxm.n134 Vxm.t47 8.266
R432 Vxm.n60 Vxm.t86 8.266
R433 Vxm.n59 Vxm.t64 8.266
R434 Vxm.n47 Vxm.t56 8.266
R435 Vxm.n46 Vxm.t75 8.266
R436 Vxm.n7 Vxm.t73 8.266
R437 Vxm.n6 Vxm.t50 8.266
R438 Vxm.n119 Vxm.t72 8.266
R439 Vxm.n118 Vxm.t54 8.266
R440 Vxm.n41 Vxm.t67 8.266
R441 Vxm.n4 Vxm.t77 8.266
R442 Vxm.n3 Vxm.t78 8.266
R443 Vxm.n49 Vxm.t85 8.266
R444 Vxm.n10 Vxm.t92 8.266
R445 Vxm.n9 Vxm.t83 8.266
R446 Vxm.n1 Vxm.t91 8.266
R447 Vxm.n112 Vxm.n68 3.303
R448 Vxm.n52 Vxm.n51 3.193
R449 Vxm.n142 Vxm.n141 3.193
R450 Vxm.n65 Vxm.n64 3.193
R451 Vxm.n125 Vxm.n124 3.193
R452 Vxm.n39 Vxm.n11 3.193
R453 Vxm.n39 Vxm.n38 2.974
R454 Vxm.n21 Vxm.n20 2.66
R455 Vxm.n106 Vxm.n94 2.66
R456 Vxm.n24 Vxm.n23 2.66
R457 Vxm.n107 Vxm.n90 2.66
R458 Vxm.n27 Vxm.n26 2.66
R459 Vxm.n108 Vxm.n86 2.66
R460 Vxm.n30 Vxm.n29 2.66
R461 Vxm.n109 Vxm.n82 2.66
R462 Vxm.n141 Vxm.n137 2.199
R463 Vxm.n133 Vxm.n129 2.199
R464 Vxm.n137 Vxm.n133 2.199
R465 Vxm.n64 Vxm.n61 2.199
R466 Vxm.n58 Vxm.n55 2.199
R467 Vxm.n61 Vxm.n58 2.199
R468 Vxm.n124 Vxm.n121 2.199
R469 Vxm.n121 Vxm.n120 2.199
R470 Vxm.n120 Vxm.n117 2.199
R471 Vxm.n45 Vxm.n44 2.199
R472 Vxm.n48 Vxm.n45 2.199
R473 Vxm.n51 Vxm.n48 2.199
R474 Vxm.n68 Vxm.n67 2.199
R475 Vxm.n67 Vxm.n66 2.199
R476 Vxm.n5 Vxm.n2 2.199
R477 Vxm.n8 Vxm.n5 2.199
R478 Vxm.n11 Vxm.n8 2.199
R479 Vxm.n17 Vxm.t15 2.071
R480 Vxm.n14 Vxm.t22 2.071
R481 Vxm.n13 Vxm.t20 2.071
R482 Vxm.n12 Vxm.t10 2.071
R483 Vxm.n100 Vxm.t100 2.071
R484 Vxm.n101 Vxm.t25 2.071
R485 Vxm.n102 Vxm.t97 2.071
R486 Vxm.n103 Vxm.t34 2.071
R487 Vxm.n104 Vxm.t38 2.071
R488 Vxm.n99 Vxm.t98 2.071
R489 Vxm.n98 Vxm.t94 2.071
R490 Vxm.n97 Vxm.t37 2.071
R491 Vxm.n96 Vxm.t30 2.071
R492 Vxm.n95 Vxm.t41 2.071
R493 Vxm.n15 Vxm.t29 2.071
R494 Vxm.n94 Vxm.t8 2.071
R495 Vxm.n93 Vxm.t19 2.071
R496 Vxm.n92 Vxm.t36 2.071
R497 Vxm.n91 Vxm.t35 2.071
R498 Vxm.n19 Vxm.t32 2.071
R499 Vxm.n20 Vxm.t43 2.071
R500 Vxm.n90 Vxm.t18 2.071
R501 Vxm.n89 Vxm.t31 2.071
R502 Vxm.n88 Vxm.t1 2.071
R503 Vxm.n87 Vxm.t26 2.071
R504 Vxm.n22 Vxm.t7 2.071
R505 Vxm.n23 Vxm.t39 2.071
R506 Vxm.n86 Vxm.t42 2.071
R507 Vxm.n85 Vxm.t17 2.071
R508 Vxm.n84 Vxm.t96 2.071
R509 Vxm.n83 Vxm.t3 2.071
R510 Vxm.n25 Vxm.t101 2.071
R511 Vxm.n26 Vxm.t12 2.071
R512 Vxm.n82 Vxm.t27 2.071
R513 Vxm.n81 Vxm.t28 2.071
R514 Vxm.n80 Vxm.t5 2.071
R515 Vxm.n79 Vxm.t4 2.071
R516 Vxm.n28 Vxm.t24 2.071
R517 Vxm.n29 Vxm.t102 2.071
R518 Vxm.n78 Vxm.t21 2.071
R519 Vxm.n77 Vxm.t23 2.071
R520 Vxm.n76 Vxm.t9 2.071
R521 Vxm.n75 Vxm.t99 2.071
R522 Vxm.n74 Vxm.t95 2.071
R523 Vxm.n31 Vxm.t16 2.071
R524 Vxm.n32 Vxm.t33 2.071
R525 Vxm.n33 Vxm.t40 2.071
R526 Vxm.n73 Vxm.t44 2.071
R527 Vxm.n72 Vxm.t14 2.071
R528 Vxm.n71 Vxm.t45 2.071
R529 Vxm.n70 Vxm.t103 2.071
R530 Vxm.n69 Vxm.t6 2.071
R531 Vxm.n35 Vxm.t11 2.071
R532 Vxm.n36 Vxm.t2 2.071
R533 Vxm.n37 Vxm.t13 2.071
R534 Vxm.n16 Vxm.t0 2.069
R535 Vxm.n16 Vxm.n15 1.246
R536 Vxm.n96 Vxm.n95 1.246
R537 Vxm.n97 Vxm.n96 1.246
R538 Vxm.n98 Vxm.n97 1.246
R539 Vxm.n99 Vxm.n98 1.246
R540 Vxm.n20 Vxm.n19 1.246
R541 Vxm.n92 Vxm.n91 1.246
R542 Vxm.n93 Vxm.n92 1.246
R543 Vxm.n94 Vxm.n93 1.246
R544 Vxm.n23 Vxm.n22 1.246
R545 Vxm.n88 Vxm.n87 1.246
R546 Vxm.n89 Vxm.n88 1.246
R547 Vxm.n90 Vxm.n89 1.246
R548 Vxm.n26 Vxm.n25 1.246
R549 Vxm.n84 Vxm.n83 1.246
R550 Vxm.n85 Vxm.n84 1.246
R551 Vxm.n86 Vxm.n85 1.246
R552 Vxm.n29 Vxm.n28 1.246
R553 Vxm.n80 Vxm.n79 1.246
R554 Vxm.n81 Vxm.n80 1.246
R555 Vxm.n82 Vxm.n81 1.246
R556 Vxm.n33 Vxm.n32 1.246
R557 Vxm.n32 Vxm.n31 1.246
R558 Vxm.n75 Vxm.n74 1.246
R559 Vxm.n76 Vxm.n75 1.246
R560 Vxm.n77 Vxm.n76 1.246
R561 Vxm.n78 Vxm.n77 1.246
R562 Vxm.n37 Vxm.n36 1.246
R563 Vxm.n36 Vxm.n35 1.246
R564 Vxm.n70 Vxm.n69 1.246
R565 Vxm.n71 Vxm.n70 1.246
R566 Vxm.n72 Vxm.n71 1.246
R567 Vxm.n73 Vxm.n72 1.246
R568 Vxm.n104 Vxm.n103 1.246
R569 Vxm.n103 Vxm.n102 1.246
R570 Vxm.n102 Vxm.n101 1.246
R571 Vxm.n101 Vxm.n100 1.246
R572 Vxm.n13 Vxm.n12 1.246
R573 Vxm.n14 Vxm.n13 1.246
R574 Vxm.n17 Vxm.n16 1.246
R575 Vxm.n105 Vxm.n99 1.124
R576 Vxm.n18 Vxm.n17 1.124
R577 Vxm.n34 Vxm.n33 0.936
R578 Vxm.n110 Vxm.n78 0.936
R579 Vxm.n38 Vxm.n37 0.936
R580 Vxm.n111 Vxm.n73 0.936
R581 Vxm.n105 Vxm.n104 0.936
R582 Vxm.n18 Vxm.n14 0.936
R583 Vxm.n8 Vxm.n6 0.597
R584 Vxm.n48 Vxm.n46 0.597
R585 Vxm.n61 Vxm.n59 0.597
R586 Vxm.n137 Vxm.n134 0.597
R587 Vxm.n133 Vxm.n130 0.597
R588 Vxm.n58 Vxm.n56 0.597
R589 Vxm.n5 Vxm.n3 0.597
R590 Vxm.n45 Vxm.n41 0.597
R591 Vxm.n11 Vxm.n9 0.597
R592 Vxm.n51 Vxm.n49 0.597
R593 Vxm.n64 Vxm.n62 0.597
R594 Vxm.n141 Vxm.n138 0.597
R595 Vxm.n129 Vxm.n126 0.597
R596 Vxm.n55 Vxm.n53 0.597
R597 Vxm.n44 Vxm.n42 0.597
R598 Vxm.n2 Vxm.n1 0.597
R599 Vxm.n114 Vxm.n113 0.591
R600 Vxm.n136 Vxm.n135 0.591
R601 Vxm.n119 Vxm.n118 0.591
R602 Vxm.n132 Vxm.n131 0.591
R603 Vxm.n140 Vxm.n139 0.591
R604 Vxm.n123 Vxm.n122 0.591
R605 Vxm.n116 Vxm.n115 0.591
R606 Vxm.n128 Vxm.n127 0.591
R607 Vxm.n112 Vxm.n111 0.401
R608 Vxm.n52 Vxm.n39 0.376
R609 Vxm.n65 Vxm.n52 0.376
R610 Vxm.n142 Vxm.n125 0.376
R611 Vxm.n121 Vxm.n114 0.351
R612 Vxm.n8 Vxm.n7 0.351
R613 Vxm.n48 Vxm.n47 0.351
R614 Vxm.n61 Vxm.n60 0.351
R615 Vxm.n137 Vxm.n136 0.351
R616 Vxm.n120 Vxm.n119 0.351
R617 Vxm.n133 Vxm.n132 0.351
R618 Vxm.n58 Vxm.n57 0.351
R619 Vxm.n45 Vxm.n40 0.351
R620 Vxm.n5 Vxm.n4 0.351
R621 Vxm.n11 Vxm.n10 0.351
R622 Vxm.n51 Vxm.n50 0.351
R623 Vxm.n64 Vxm.n63 0.351
R624 Vxm.n141 Vxm.n140 0.351
R625 Vxm.n124 Vxm.n123 0.351
R626 Vxm.n117 Vxm.n116 0.351
R627 Vxm.n129 Vxm.n128 0.351
R628 Vxm.n55 Vxm.n54 0.351
R629 Vxm.n44 Vxm.n43 0.351
R630 Vxm.n2 Vxm.n0 0.351
R631 Vxm.n125 Vxm.n112 0.265
R632 Vxm Vxm.n142 0.193
R633 Vxm.n106 Vxm.n105 0.188
R634 Vxm.n107 Vxm.n106 0.188
R635 Vxm.n108 Vxm.n107 0.188
R636 Vxm.n109 Vxm.n108 0.188
R637 Vxm.n110 Vxm.n109 0.188
R638 Vxm.n111 Vxm.n110 0.188
R639 Vxm.n21 Vxm.n18 0.188
R640 Vxm.n24 Vxm.n21 0.188
R641 Vxm.n27 Vxm.n24 0.188
R642 Vxm.n30 Vxm.n27 0.188
R643 Vxm.n34 Vxm.n30 0.188
R644 Vxm.n38 Vxm.n34 0.188
R645 Vxm Vxm.n65 0.182
R646 a_1659_n4497.n69 a_1659_n4497.t10 8.266
R647 a_1659_n4497.n12 a_1659_n4497.t63 8.266
R648 a_1659_n4497.n12 a_1659_n4497.t13 8.266
R649 a_1659_n4497.n13 a_1659_n4497.t84 8.266
R650 a_1659_n4497.n13 a_1659_n4497.t23 8.266
R651 a_1659_n4497.n14 a_1659_n4497.t64 8.266
R652 a_1659_n4497.n14 a_1659_n4497.t27 8.266
R653 a_1659_n4497.n19 a_1659_n4497.t56 8.266
R654 a_1659_n4497.n19 a_1659_n4497.t40 8.266
R655 a_1659_n4497.n18 a_1659_n4497.t79 8.266
R656 a_1659_n4497.n18 a_1659_n4497.t16 8.266
R657 a_1659_n4497.n16 a_1659_n4497.t76 8.266
R658 a_1659_n4497.n16 a_1659_n4497.t28 8.266
R659 a_1659_n4497.n15 a_1659_n4497.t49 8.266
R660 a_1659_n4497.n15 a_1659_n4497.t95 8.266
R661 a_1659_n4497.n41 a_1659_n4497.t90 8.266
R662 a_1659_n4497.n41 a_1659_n4497.t0 8.266
R663 a_1659_n4497.n40 a_1659_n4497.t67 8.266
R664 a_1659_n4497.n40 a_1659_n4497.t45 8.266
R665 a_1659_n4497.n38 a_1659_n4497.t60 8.266
R666 a_1659_n4497.n38 a_1659_n4497.t3 8.266
R667 a_1659_n4497.n37 a_1659_n4497.t81 8.266
R668 a_1659_n4497.n37 a_1659_n4497.t38 8.266
R669 a_1659_n4497.n46 a_1659_n4497.t17 8.266
R670 a_1659_n4497.n46 a_1659_n4497.t77 8.266
R671 a_1659_n4497.n47 a_1659_n4497.t72 8.266
R672 a_1659_n4497.n47 a_1659_n4497.t25 8.266
R673 a_1659_n4497.n43 a_1659_n4497.t89 8.266
R674 a_1659_n4497.n43 a_1659_n4497.t24 8.266
R675 a_1659_n4497.n44 a_1659_n4497.t74 8.266
R676 a_1659_n4497.n44 a_1659_n4497.t14 8.266
R677 a_1659_n4497.n23 a_1659_n4497.t91 8.266
R678 a_1659_n4497.n23 a_1659_n4497.t12 8.266
R679 a_1659_n4497.n24 a_1659_n4497.t85 8.266
R680 a_1659_n4497.n24 a_1659_n4497.t19 8.266
R681 a_1659_n4497.n26 a_1659_n4497.t54 8.266
R682 a_1659_n4497.n26 a_1659_n4497.t18 8.266
R683 a_1659_n4497.n27 a_1659_n4497.t52 8.266
R684 a_1659_n4497.n27 a_1659_n4497.t37 8.266
R685 a_1659_n4497.n22 a_1659_n4497.t71 8.266
R686 a_1659_n4497.n22 a_1659_n4497.t36 8.266
R687 a_1659_n4497.n21 a_1659_n4497.t53 8.266
R688 a_1659_n4497.n21 a_1659_n4497.t2 8.266
R689 a_1659_n4497.n29 a_1659_n4497.t87 8.266
R690 a_1659_n4497.n29 a_1659_n4497.t44 8.266
R691 a_1659_n4497.n30 a_1659_n4497.t65 8.266
R692 a_1659_n4497.n30 a_1659_n4497.t9 8.266
R693 a_1659_n4497.n32 a_1659_n4497.t57 8.266
R694 a_1659_n4497.n32 a_1659_n4497.t11 8.266
R695 a_1659_n4497.n31 a_1659_n4497.t80 8.266
R696 a_1659_n4497.n31 a_1659_n4497.t33 8.266
R697 a_1659_n4497.n35 a_1659_n4497.t78 8.266
R698 a_1659_n4497.n35 a_1659_n4497.t34 8.266
R699 a_1659_n4497.n34 a_1659_n4497.t50 8.266
R700 a_1659_n4497.n34 a_1659_n4497.t5 8.266
R701 a_1659_n4497.n53 a_1659_n4497.t92 8.266
R702 a_1659_n4497.n53 a_1659_n4497.t6 8.266
R703 a_1659_n4497.n52 a_1659_n4497.t69 8.266
R704 a_1659_n4497.n52 a_1659_n4497.t20 8.266
R705 a_1659_n4497.n58 a_1659_n4497.t88 8.266
R706 a_1659_n4497.n58 a_1659_n4497.t7 8.266
R707 a_1659_n4497.n57 a_1659_n4497.t59 8.266
R708 a_1659_n4497.n57 a_1659_n4497.t4 8.266
R709 a_1659_n4497.n60 a_1659_n4497.t48 8.266
R710 a_1659_n4497.n60 a_1659_n4497.t30 8.266
R711 a_1659_n4497.n61 a_1659_n4497.t66 8.266
R712 a_1659_n4497.n61 a_1659_n4497.t35 8.266
R713 a_1659_n4497.n63 a_1659_n4497.t75 8.266
R714 a_1659_n4497.n63 a_1659_n4497.t29 8.266
R715 a_1659_n4497.n64 a_1659_n4497.t51 8.266
R716 a_1659_n4497.n64 a_1659_n4497.t94 8.266
R717 a_1659_n4497.n66 a_1659_n4497.t55 8.266
R718 a_1659_n4497.n66 a_1659_n4497.t41 8.266
R719 a_1659_n4497.n67 a_1659_n4497.t82 8.266
R720 a_1659_n4497.n67 a_1659_n4497.t26 8.266
R721 a_1659_n4497.n50 a_1659_n4497.t62 8.266
R722 a_1659_n4497.n50 a_1659_n4497.t21 8.266
R723 a_1659_n4497.n49 a_1659_n4497.t83 8.266
R724 a_1659_n4497.n49 a_1659_n4497.t31 8.266
R725 a_1659_n4497.n4 a_1659_n4497.t47 8.266
R726 a_1659_n4497.n4 a_1659_n4497.t43 8.266
R727 a_1659_n4497.n3 a_1659_n4497.t61 8.266
R728 a_1659_n4497.n3 a_1659_n4497.t1 8.266
R729 a_1659_n4497.n6 a_1659_n4497.t73 8.266
R730 a_1659_n4497.n6 a_1659_n4497.t15 8.266
R731 a_1659_n4497.n5 a_1659_n4497.t68 8.266
R732 a_1659_n4497.n5 a_1659_n4497.t32 8.266
R733 a_1659_n4497.n1 a_1659_n4497.t46 8.266
R734 a_1659_n4497.n1 a_1659_n4497.t22 8.266
R735 a_1659_n4497.n0 a_1659_n4497.t58 8.266
R736 a_1659_n4497.n0 a_1659_n4497.t39 8.266
R737 a_1659_n4497.n10 a_1659_n4497.t70 8.266
R738 a_1659_n4497.n10 a_1659_n4497.t42 8.266
R739 a_1659_n4497.n9 a_1659_n4497.t86 8.266
R740 a_1659_n4497.n9 a_1659_n4497.t8 8.266
R741 a_1659_n4497.t93 a_1659_n4497.n69 8.266
R742 a_1659_n4497.n51 a_1659_n4497.n48 2.199
R743 a_1659_n4497.n54 a_1659_n4497.n45 2.199
R744 a_1659_n4497.n62 a_1659_n4497.n54 2.199
R745 a_1659_n4497.n62 a_1659_n4497.n42 2.199
R746 a_1659_n4497.n65 a_1659_n4497.n36 2.199
R747 a_1659_n4497.n33 a_1659_n4497.n28 2.199
R748 a_1659_n4497.n68 a_1659_n4497.n33 2.199
R749 a_1659_n4497.n68 a_1659_n4497.n20 2.199
R750 a_1659_n4497.n11 a_1659_n4497.n8 2.199
R751 a_1659_n4497.n8 a_1659_n4497.n7 2.199
R752 a_1659_n4497.n56 a_1659_n4497.n55 2.199
R753 a_1659_n4497.n11 a_1659_n4497.n2 2.199
R754 a_1659_n4497.n59 a_1659_n4497.n58 0.434
R755 a_1659_n4497.n68 a_1659_n4497.n67 0.434
R756 a_1659_n4497.n65 a_1659_n4497.n64 0.434
R757 a_1659_n4497.n62 a_1659_n4497.n61 0.434
R758 a_1659_n4497.n51 a_1659_n4497.n50 0.434
R759 a_1659_n4497.n54 a_1659_n4497.n53 0.434
R760 a_1659_n4497.n36 a_1659_n4497.n35 0.434
R761 a_1659_n4497.n33 a_1659_n4497.n32 0.434
R762 a_1659_n4497.n28 a_1659_n4497.n27 0.434
R763 a_1659_n4497.n25 a_1659_n4497.n24 0.434
R764 a_1659_n4497.n45 a_1659_n4497.n44 0.434
R765 a_1659_n4497.n48 a_1659_n4497.n47 0.434
R766 a_1659_n4497.n39 a_1659_n4497.n38 0.434
R767 a_1659_n4497.n42 a_1659_n4497.n41 0.434
R768 a_1659_n4497.n17 a_1659_n4497.n16 0.434
R769 a_1659_n4497.n20 a_1659_n4497.n19 0.434
R770 a_1659_n4497.n12 a_1659_n4497.n11 0.434
R771 a_1659_n4497.n58 a_1659_n4497.n57 0.365
R772 a_1659_n4497.n67 a_1659_n4497.n66 0.365
R773 a_1659_n4497.n64 a_1659_n4497.n63 0.365
R774 a_1659_n4497.n61 a_1659_n4497.n60 0.365
R775 a_1659_n4497.n50 a_1659_n4497.n49 0.365
R776 a_1659_n4497.n53 a_1659_n4497.n52 0.365
R777 a_1659_n4497.n35 a_1659_n4497.n34 0.365
R778 a_1659_n4497.n32 a_1659_n4497.n31 0.365
R779 a_1659_n4497.n30 a_1659_n4497.n29 0.365
R780 a_1659_n4497.n4 a_1659_n4497.n3 0.365
R781 a_1659_n4497.n6 a_1659_n4497.n5 0.365
R782 a_1659_n4497.n22 a_1659_n4497.n21 0.365
R783 a_1659_n4497.n27 a_1659_n4497.n26 0.365
R784 a_1659_n4497.n24 a_1659_n4497.n23 0.365
R785 a_1659_n4497.n44 a_1659_n4497.n43 0.365
R786 a_1659_n4497.n47 a_1659_n4497.n46 0.365
R787 a_1659_n4497.n38 a_1659_n4497.n37 0.365
R788 a_1659_n4497.n41 a_1659_n4497.n40 0.365
R789 a_1659_n4497.n16 a_1659_n4497.n15 0.365
R790 a_1659_n4497.n19 a_1659_n4497.n18 0.365
R791 a_1659_n4497.n14 a_1659_n4497.n13 0.365
R792 a_1659_n4497.n1 a_1659_n4497.n0 0.365
R793 a_1659_n4497.n10 a_1659_n4497.n9 0.365
R794 a_1659_n4497.n69 a_1659_n4497.n12 0.365
R795 a_1659_n4497.n57 a_1659_n4497.n56 0.253
R796 a_1659_n4497.n69 a_1659_n4497.n68 0.253
R797 a_1659_n4497.n66 a_1659_n4497.n65 0.253
R798 a_1659_n4497.n63 a_1659_n4497.n62 0.253
R799 a_1659_n4497.n60 a_1659_n4497.n59 0.253
R800 a_1659_n4497.n52 a_1659_n4497.n51 0.253
R801 a_1659_n4497.n33 a_1659_n4497.n30 0.253
R802 a_1659_n4497.n8 a_1659_n4497.n4 0.253
R803 a_1659_n4497.n7 a_1659_n4497.n6 0.253
R804 a_1659_n4497.n28 a_1659_n4497.n22 0.253
R805 a_1659_n4497.n26 a_1659_n4497.n25 0.253
R806 a_1659_n4497.n40 a_1659_n4497.n39 0.253
R807 a_1659_n4497.n18 a_1659_n4497.n17 0.253
R808 a_1659_n4497.n20 a_1659_n4497.n14 0.253
R809 a_1659_n4497.n2 a_1659_n4497.n1 0.253
R810 a_1659_n4497.n11 a_1659_n4497.n10 0.253
R811 DGND.n66 DGND.t525 292.915
R812 DGND.t523 DGND.t533 217.25
R813 DGND.t525 DGND.t473 217.25
R814 DGND.n87 DGND.n79 149.834
R815 DGND.n101 DGND.n100 149.834
R816 DGND.n16 DGND.t523 108.625
R817 DGND.n2 DGND.n1 93.745
R818 DGND.n109 DGND.n108 90.903
R819 DGND.n118 DGND.n115 90.352
R820 DGND.n65 DGND.n19 89.912
R821 DGND.n87 DGND.n86 53.082
R822 DGND.n65 DGND.n64 42.026
R823 DGND.n65 DGND.n44 42.026
R824 DGND.n12 DGND.t442 33.615
R825 DGND.n11 DGND.t528 33.599
R826 DGND.n39 DGND.n27 28.03
R827 DGND.n61 DGND.n56 28.03
R828 DGND.n63 DGND.n61 28.03
R829 DGND.n40 DGND.n39 28.03
R830 DGND.n26 DGND.n24 35.67
R831 DGND.n54 DGND.n50 27.22
R832 DGND.n33 DGND.n28 20.357
R833 DGND.n60 DGND.n57 19.54
R834 DGND.n39 DGND.n33 18.384
R835 DGND.n61 DGND.n60 18.384
R836 DGND.n4 DGND.t219 18.351
R837 DGND.n97 DGND.t676 18.3
R838 DGND.n4 DGND.t518 17.874
R839 DGND.n50 DGND.n49 16.371
R840 DGND.n69 DGND.n68 13.783
R841 DGND.n86 DGND.n85 11.717
R842 DGND.n6 DGND.t534 8.265
R843 DGND.n6 DGND.t524 8.265
R844 DGND.n5 DGND.t474 8.265
R845 DGND.n5 DGND.t526 8.265
R846 DGND.n39 DGND.n38 6.317
R847 DGND.n111 DGND.n110 5.737
R848 DGND.n95 DGND.n94 5.64
R849 DGND.n14 DGND.t23 5.633
R850 DGND.n10 DGND.t615 5.155
R851 DGND.n118 DGND.n117 4.603
R852 DGND.n10 DGND.t530 4.132
R853 DGND.n12 DGND.t146 4.132
R854 DGND.n90 DGND.n76 3.579
R855 DGND.n15 DGND.n14 3.1
R856 DGND.n119 DGND.n118 2.457
R857 DGND.n16 DGND.n6 2.363
R858 DGND.n16 DGND.n5 2.363
R859 DGND.n13 DGND.n12 1.851
R860 DGND.n64 DGND.n63 1.62
R861 DGND.n44 DGND.n40 1.62
R862 DGND.n13 DGND.n11 1.37
R863 DGND.n111 DGND.n109 1.324
R864 DGND.n74 DGND.n73 0.976
R865 DGND.n70 DGND.n17 0.822
R866 DGND.n70 DGND.n69 0.822
R867 DGND.n27 DGND.n26 0.81
R868 DGND.n56 DGND.n54 0.81
R869 DGND DGND.n128 0.431
R870 DGND.n85 DGND.n82 0.376
R871 DGND.n14 DGND.n13 0.349
R872 DGND.n71 DGND.n16 0.335
R873 DGND.n75 DGND.n72 0.141
R874 DGND.n128 DGND.n3 0.128
R875 DGND.n68 DGND.n65 0.112
R876 DGND.n117 DGND.n116 0.11
R877 DGND.n102 DGND.n101 0.109
R878 DGND.t517 DGND.n102 0.109
R879 DGND.n123 DGND.n122 0.109
R880 DGND.t675 DGND.n123 0.109
R881 DGND.n88 DGND.n87 0.109
R882 DGND.t218 DGND.n88 0.109
R883 DGND.n128 DGND.n127 0.09
R884 DGND.n120 DGND.n112 0.068
R885 DGND.n96 DGND.n93 0.068
R886 DGND.n97 DGND.n4 0.051
R887 DGND.n24 DGND.n23 0.046
R888 DGND.n23 DGND.n22 0.046
R889 DGND.n38 DGND.n35 0.046
R890 DGND.n35 DGND.n34 0.046
R891 DGND.n38 DGND.n37 0.046
R892 DGND.n37 DGND.n36 0.046
R893 DGND.n65 DGND.n46 0.046
R894 DGND.n46 DGND.n45 0.046
R895 DGND.n82 DGND.n81 0.042
R896 DGND.n81 DGND.n80 0.042
R897 DGND.n100 DGND.n99 0.042
R898 DGND.n99 DGND.n98 0.042
R899 DGND.n108 DGND.n107 0.042
R900 DGND.n107 DGND.n106 0.042
R901 DGND.n115 DGND.n114 0.042
R902 DGND.n114 DGND.n113 0.042
R903 DGND.n1 DGND.n0 0.042
R904 DGND.n79 DGND.n78 0.042
R905 DGND.n78 DGND.n77 0.042
R906 DGND.n49 DGND.n48 0.04
R907 DGND.n33 DGND.n30 0.04
R908 DGND.n30 DGND.n29 0.04
R909 DGND.n33 DGND.n32 0.04
R910 DGND.n32 DGND.n31 0.04
R911 DGND.n60 DGND.n58 0.04
R912 DGND.n60 DGND.n59 0.04
R913 DGND.n68 DGND.n66 0.04
R914 DGND.n68 DGND.n67 0.04
R915 DGND.n112 DGND.n105 0.037
R916 DGND.n93 DGND.n91 0.037
R917 DGND.n91 DGND.n75 0.037
R918 DGND.n72 DGND.n71 0.035
R919 DGND.n27 DGND.n21 0.025
R920 DGND.n55 DGND.t527 0.025
R921 DGND.n56 DGND.n55 0.025
R922 DGND.n63 DGND.n62 0.025
R923 DGND.n62 DGND.t441 0.025
R924 DGND.n40 DGND.n20 0.025
R925 DGND.n85 DGND.n84 0.023
R926 DGND.n84 DGND.n83 0.023
R927 DGND.n121 DGND.n120 0.022
R928 DGND.n97 DGND.n96 0.02
R929 DGND.n8 DGND.n7 0.019
R930 DGND.n71 DGND.n70 0.017
R931 DGND.n105 DGND.n97 0.017
R932 DGND.n93 DGND.n92 0.017
R933 DGND.n75 DGND.n74 0.017
R934 DGND.n112 DGND.n111 0.017
R935 DGND.n120 DGND.n119 0.017
R936 DGND.n96 DGND.n95 0.017
R937 DGND.n3 DGND.n2 0.017
R938 DGND.n127 DGND.n121 0.015
R939 DGND.n52 DGND.n51 0.014
R940 DGND.t529 DGND.n52 0.014
R941 DGND.n26 DGND.n25 0.014
R942 DGND.n53 DGND.t529 0.014
R943 DGND.n54 DGND.n53 0.014
R944 DGND.n64 DGND.n47 0.014
R945 DGND.n44 DGND.n43 0.014
R946 DGND.n43 DGND.t22 0.014
R947 DGND.n19 DGND.n18 0.014
R948 DGND.t22 DGND.n42 0.014
R949 DGND.n42 DGND.n41 0.014
R950 DGND.n16 DGND.n9 0.01
R951 DGND.n9 DGND.n8 0.01
R952 DGND.n16 DGND.n15 0.01
R953 DGND.n11 DGND.n10 0.008
R954 DGND.n125 DGND.n124 0.003
R955 DGND.n89 DGND.t218 0.003
R956 DGND.n103 DGND.t517 0.003
R957 DGND.n104 DGND.n103 0.003
R958 DGND.n90 DGND.n89 0.003
R959 DGND.n126 DGND.n125 0.003
R960 DGND.n124 DGND.t675 0.001
R961 DGND.n91 DGND.n90 0.001
R962 DGND.n127 DGND.n126 0.001
R963 DGND.n105 DGND.n104 0.001
R964 AVDD.n3587 AVDD.n3582 459.931
R965 AVDD.n3474 AVDD.n3473 459.931
R966 AVDD.n1208 AVDD.n1205 459.931
R967 AVDD.n1367 AVDD.n1364 459.931
R968 AVDD.n1483 AVDD.n1480 459.931
R969 AVDD.n1571 AVDD.n1568 459.931
R970 AVDD.n1664 AVDD.n1661 459.931
R971 AVDD.n1780 AVDD.n1777 459.931
R972 AVDD.n1925 AVDD.n1922 459.931
R973 AVDD.n1992 AVDD.n1989 459.931
R974 AVDD.n2196 AVDD.n2193 459.931
R975 AVDD.n2071 AVDD.n2068 459.931
R976 AVDD.n2297 AVDD.n2294 459.931
R977 AVDD.n2407 AVDD.n2404 459.931
R978 AVDD.n2477 AVDD.n2474 459.931
R979 AVDD.n2571 AVDD.n2568 459.931
R980 AVDD.n2722 AVDD.n2719 459.931
R981 AVDD.n2789 AVDD.n2786 459.931
R982 AVDD.n2885 AVDD.n2882 459.931
R983 AVDD.n2951 AVDD.n2948 459.931
R984 AVDD.n3066 AVDD.n3063 459.931
R985 AVDD.n3176 AVDD.n3173 459.931
R986 AVDD.n3285 AVDD.n3282 459.931
R987 AVDD.n3350 AVDD.n3347 459.931
R988 AVDD.n4715 AVDD.n4712 459.931
R989 AVDD.n4940 AVDD.n4937 459.931
R990 AVDD.n4721 AVDD.n4718 459.931
R991 AVDD.n4946 AVDD.n4943 459.931
R992 AVDD.n3291 AVDD.n3288 459.931
R993 AVDD.n3356 AVDD.n3353 459.931
R994 AVDD.n3072 AVDD.n3069 459.931
R995 AVDD.n3182 AVDD.n3179 459.931
R996 AVDD.n2891 AVDD.n2888 459.931
R997 AVDD.n2957 AVDD.n2954 459.931
R998 AVDD.n2728 AVDD.n2725 459.931
R999 AVDD.n2795 AVDD.n2792 459.931
R1000 AVDD.n2483 AVDD.n2480 459.931
R1001 AVDD.n2577 AVDD.n2574 459.931
R1002 AVDD.n2303 AVDD.n2300 459.931
R1003 AVDD.n2413 AVDD.n2410 459.931
R1004 AVDD.n2202 AVDD.n2199 459.931
R1005 AVDD.n2077 AVDD.n2074 459.931
R1006 AVDD.n1931 AVDD.n1928 459.931
R1007 AVDD.n1998 AVDD.n1995 459.931
R1008 AVDD.n1670 AVDD.n1667 459.931
R1009 AVDD.n1786 AVDD.n1783 459.931
R1010 AVDD.n1489 AVDD.n1486 459.931
R1011 AVDD.n1577 AVDD.n1574 459.931
R1012 AVDD.n1214 AVDD.n1211 459.931
R1013 AVDD.n1373 AVDD.n1370 459.931
R1014 AVDD.n1307 AVDD.n1304 459.931
R1015 AVDD.n1113 AVDD.n1110 459.931
R1016 AVDD.n946 AVDD.n943 459.931
R1017 AVDD.n1008 AVDD.n1005 459.931
R1018 AVDD.n765 AVDD.n762 459.931
R1019 AVDD.n827 AVDD.n824 459.931
R1020 AVDD.n2507 AVDD.n2504 459.931
R1021 AVDD.n2601 AVDD.n2598 459.931
R1022 AVDD.n2327 AVDD.n2324 459.931
R1023 AVDD.n2437 AVDD.n2434 459.931
R1024 AVDD.n2226 AVDD.n2223 459.931
R1025 AVDD.n2101 AVDD.n2098 459.931
R1026 AVDD.n1955 AVDD.n1952 459.931
R1027 AVDD.n2022 AVDD.n2019 459.931
R1028 AVDD.n1694 AVDD.n1691 459.931
R1029 AVDD.n1810 AVDD.n1807 459.931
R1030 AVDD.n1513 AVDD.n1510 459.931
R1031 AVDD.n1601 AVDD.n1598 459.931
R1032 AVDD.n1238 AVDD.n1235 459.931
R1033 AVDD.n1397 AVDD.n1394 459.931
R1034 AVDD.n1331 AVDD.n1328 459.931
R1035 AVDD.n1137 AVDD.n1134 459.931
R1036 AVDD.n970 AVDD.n967 459.931
R1037 AVDD.n1032 AVDD.n1029 459.931
R1038 AVDD.n789 AVDD.n786 459.931
R1039 AVDD.n851 AVDD.n848 459.931
R1040 AVDD.n4757 AVDD.n4754 459.931
R1041 AVDD.n4934 AVDD.n4931 459.931
R1042 AVDD.n3327 AVDD.n3324 459.931
R1043 AVDD.n3344 AVDD.n3341 459.931
R1044 AVDD.n3108 AVDD.n3105 459.931
R1045 AVDD.n3170 AVDD.n3167 459.931
R1046 AVDD.n2927 AVDD.n2924 459.931
R1047 AVDD.n2945 AVDD.n2942 459.931
R1048 AVDD.n2764 AVDD.n2761 459.931
R1049 AVDD.n2783 AVDD.n2780 459.931
R1050 AVDD.n2519 AVDD.n2516 459.931
R1051 AVDD.n2565 AVDD.n2562 459.931
R1052 AVDD.n2339 AVDD.n2336 459.931
R1053 AVDD.n2401 AVDD.n2398 459.931
R1054 AVDD.n2238 AVDD.n2235 459.931
R1055 AVDD.n2065 AVDD.n2062 459.931
R1056 AVDD.n1967 AVDD.n1964 459.931
R1057 AVDD.n1986 AVDD.n1983 459.931
R1058 AVDD.n1706 AVDD.n1703 459.931
R1059 AVDD.n1774 AVDD.n1771 459.931
R1060 AVDD.n1525 AVDD.n1522 459.931
R1061 AVDD.n1565 AVDD.n1562 459.931
R1062 AVDD.n1250 AVDD.n1247 459.931
R1063 AVDD.n1360 AVDD.n1357 459.931
R1064 AVDD.n1343 AVDD.n1340 459.931
R1065 AVDD.n1101 AVDD.n1098 459.931
R1066 AVDD.n982 AVDD.n979 459.931
R1067 AVDD.n996 AVDD.n993 459.931
R1068 AVDD.n801 AVDD.n798 459.931
R1069 AVDD.n815 AVDD.n812 459.931
R1070 AVDD.n4806 AVDD.n4803 459.931
R1071 AVDD.n4582 AVDD.n4581 459.931
R1072 AVDD.n4500 AVDD.n4485 459.931
R1073 AVDD.n3578 AVDD.n3577 459.931
R1074 AVDD.n4584 AVDD.n4559 459.931
R1075 AVDD.n4800 AVDD.n4797 459.931
R1076 AVDD.n3635 AVDD.n3630 459.931
R1077 AVDD.n4586 AVDD.n4585 459.931
R1078 AVDD.n4532 AVDD.n4531 459.931
R1079 AVDD.n4794 AVDD.n4791 459.931
R1080 AVDD.n3627 AVDD.n3622 459.931
R1081 AVDD.n4534 AVDD.n4533 459.931
R1082 AVDD.n4456 AVDD.n4455 459.931
R1083 AVDD.n4788 AVDD.n4785 459.931
R1084 AVDD.n3619 AVDD.n3614 459.931
R1085 AVDD.n4502 AVDD.n4457 459.931
R1086 AVDD.n4579 AVDD.n4578 459.931
R1087 AVDD.n4782 AVDD.n4779 459.931
R1088 AVDD.n3611 AVDD.n3606 459.931
R1089 AVDD.n4469 AVDD.n4468 459.931
R1090 AVDD.n3603 AVDD.n3598 459.931
R1091 AVDD.n3723 AVDD.n3722 459.931
R1092 AVDD.n3721 AVDD.n3720 459.931
R1093 AVDD.n4776 AVDD.n4773 459.931
R1094 AVDD.n771 AVDD.n768 459.931
R1095 AVDD.n833 AVDD.n830 459.931
R1096 AVDD.n952 AVDD.n949 459.931
R1097 AVDD.n1014 AVDD.n1011 459.931
R1098 AVDD.n1313 AVDD.n1310 459.931
R1099 AVDD.n1119 AVDD.n1116 459.931
R1100 AVDD.n1220 AVDD.n1217 459.931
R1101 AVDD.n1379 AVDD.n1376 459.931
R1102 AVDD.n1495 AVDD.n1492 459.931
R1103 AVDD.n1583 AVDD.n1580 459.931
R1104 AVDD.n1676 AVDD.n1673 459.931
R1105 AVDD.n1792 AVDD.n1789 459.931
R1106 AVDD.n1937 AVDD.n1934 459.931
R1107 AVDD.n2004 AVDD.n2001 459.931
R1108 AVDD.n2208 AVDD.n2205 459.931
R1109 AVDD.n2083 AVDD.n2080 459.931
R1110 AVDD.n2309 AVDD.n2306 459.931
R1111 AVDD.n2419 AVDD.n2416 459.931
R1112 AVDD.n2489 AVDD.n2486 459.931
R1113 AVDD.n2583 AVDD.n2580 459.931
R1114 AVDD.n2734 AVDD.n2731 459.931
R1115 AVDD.n2801 AVDD.n2798 459.931
R1116 AVDD.n2897 AVDD.n2894 459.931
R1117 AVDD.n2963 AVDD.n2960 459.931
R1118 AVDD.n3078 AVDD.n3075 459.931
R1119 AVDD.n3188 AVDD.n3185 459.931
R1120 AVDD.n3297 AVDD.n3294 459.931
R1121 AVDD.n3362 AVDD.n3359 459.931
R1122 AVDD.n4727 AVDD.n4724 459.931
R1123 AVDD.n4952 AVDD.n4949 459.931
R1124 AVDD.n777 AVDD.n774 459.931
R1125 AVDD.n839 AVDD.n836 459.931
R1126 AVDD.n958 AVDD.n955 459.931
R1127 AVDD.n1020 AVDD.n1017 459.931
R1128 AVDD.n1319 AVDD.n1316 459.931
R1129 AVDD.n1125 AVDD.n1122 459.931
R1130 AVDD.n1226 AVDD.n1223 459.931
R1131 AVDD.n1385 AVDD.n1382 459.931
R1132 AVDD.n1501 AVDD.n1498 459.931
R1133 AVDD.n1589 AVDD.n1586 459.931
R1134 AVDD.n1682 AVDD.n1679 459.931
R1135 AVDD.n1798 AVDD.n1795 459.931
R1136 AVDD.n1943 AVDD.n1940 459.931
R1137 AVDD.n2010 AVDD.n2007 459.931
R1138 AVDD.n2214 AVDD.n2211 459.931
R1139 AVDD.n2089 AVDD.n2086 459.931
R1140 AVDD.n2315 AVDD.n2312 459.931
R1141 AVDD.n2425 AVDD.n2422 459.931
R1142 AVDD.n2495 AVDD.n2492 459.931
R1143 AVDD.n2589 AVDD.n2586 459.931
R1144 AVDD.n2740 AVDD.n2737 459.931
R1145 AVDD.n2807 AVDD.n2804 459.931
R1146 AVDD.n2903 AVDD.n2900 459.931
R1147 AVDD.n2969 AVDD.n2966 459.931
R1148 AVDD.n3084 AVDD.n3081 459.931
R1149 AVDD.n3194 AVDD.n3191 459.931
R1150 AVDD.n3303 AVDD.n3300 459.931
R1151 AVDD.n3368 AVDD.n3365 459.931
R1152 AVDD.n4733 AVDD.n4730 459.931
R1153 AVDD.n4958 AVDD.n4955 459.931
R1154 AVDD.n783 AVDD.n780 459.931
R1155 AVDD.n845 AVDD.n842 459.931
R1156 AVDD.n964 AVDD.n961 459.931
R1157 AVDD.n1026 AVDD.n1023 459.931
R1158 AVDD.n1325 AVDD.n1322 459.931
R1159 AVDD.n1131 AVDD.n1128 459.931
R1160 AVDD.n1232 AVDD.n1229 459.931
R1161 AVDD.n1391 AVDD.n1388 459.931
R1162 AVDD.n1507 AVDD.n1504 459.931
R1163 AVDD.n1595 AVDD.n1592 459.931
R1164 AVDD.n1688 AVDD.n1685 459.931
R1165 AVDD.n1804 AVDD.n1801 459.931
R1166 AVDD.n1949 AVDD.n1946 459.931
R1167 AVDD.n2016 AVDD.n2013 459.931
R1168 AVDD.n2220 AVDD.n2217 459.931
R1169 AVDD.n2095 AVDD.n2092 459.931
R1170 AVDD.n2321 AVDD.n2318 459.931
R1171 AVDD.n2431 AVDD.n2428 459.931
R1172 AVDD.n2501 AVDD.n2498 459.931
R1173 AVDD.n2595 AVDD.n2592 459.931
R1174 AVDD.n2746 AVDD.n2743 459.931
R1175 AVDD.n2813 AVDD.n2810 459.931
R1176 AVDD.n2909 AVDD.n2906 459.931
R1177 AVDD.n2975 AVDD.n2972 459.931
R1178 AVDD.n3090 AVDD.n3087 459.931
R1179 AVDD.n3200 AVDD.n3197 459.931
R1180 AVDD.n3309 AVDD.n3306 459.931
R1181 AVDD.n3374 AVDD.n3371 459.931
R1182 AVDD.n4739 AVDD.n4736 459.931
R1183 AVDD.n4964 AVDD.n4961 459.931
R1184 AVDD.n2752 AVDD.n2749 459.931
R1185 AVDD.n2819 AVDD.n2816 459.931
R1186 AVDD.n2915 AVDD.n2912 459.931
R1187 AVDD.n2981 AVDD.n2978 459.931
R1188 AVDD.n3096 AVDD.n3093 459.931
R1189 AVDD.n3206 AVDD.n3203 459.931
R1190 AVDD.n3315 AVDD.n3312 459.931
R1191 AVDD.n3380 AVDD.n3377 459.931
R1192 AVDD.n4745 AVDD.n4742 459.931
R1193 AVDD.n4970 AVDD.n4967 459.931
R1194 AVDD.n795 AVDD.n792 459.931
R1195 AVDD.n857 AVDD.n854 459.931
R1196 AVDD.n976 AVDD.n973 459.931
R1197 AVDD.n1038 AVDD.n1035 459.931
R1198 AVDD.n1337 AVDD.n1334 459.931
R1199 AVDD.n1143 AVDD.n1140 459.931
R1200 AVDD.n1244 AVDD.n1241 459.931
R1201 AVDD.n1403 AVDD.n1400 459.931
R1202 AVDD.n1519 AVDD.n1516 459.931
R1203 AVDD.n1607 AVDD.n1604 459.931
R1204 AVDD.n1700 AVDD.n1697 459.931
R1205 AVDD.n1816 AVDD.n1813 459.931
R1206 AVDD.n1961 AVDD.n1958 459.931
R1207 AVDD.n2028 AVDD.n2025 459.931
R1208 AVDD.n2232 AVDD.n2229 459.931
R1209 AVDD.n2107 AVDD.n2104 459.931
R1210 AVDD.n2333 AVDD.n2330 459.931
R1211 AVDD.n2443 AVDD.n2440 459.931
R1212 AVDD.n2513 AVDD.n2510 459.931
R1213 AVDD.n2607 AVDD.n2604 459.931
R1214 AVDD.n2758 AVDD.n2755 459.931
R1215 AVDD.n2825 AVDD.n2822 459.931
R1216 AVDD.n2921 AVDD.n2918 459.931
R1217 AVDD.n2987 AVDD.n2984 459.931
R1218 AVDD.n3102 AVDD.n3099 459.931
R1219 AVDD.n3212 AVDD.n3209 459.931
R1220 AVDD.n3321 AVDD.n3318 459.931
R1221 AVDD.n3386 AVDD.n3383 459.931
R1222 AVDD.n4751 AVDD.n4748 459.931
R1223 AVDD.n4976 AVDD.n4973 459.931
R1224 AVDD.n3551 AVDD.n3550 459.931
R1225 AVDD.n4770 AVDD.n4767 459.931
R1226 AVDD.n3595 AVDD.n3590 459.931
R1227 AVDD.n3553 AVDD.n3552 459.931
R1228 AVDD.n4764 AVDD.n4761 459.931
R1229 AVDD.n3472 AVDD.n3471 459.931
R1230 AVDD.n1301 AVDD.n1298 459.931
R1231 AVDD.n1107 AVDD.n1104 459.931
R1232 AVDD.n940 AVDD.n937 459.931
R1233 AVDD.n1002 AVDD.n999 459.931
R1234 AVDD.n759 AVDD.n756 459.931
R1235 AVDD.n821 AVDD.n818 459.931
R1236 AVDD.n584 AVDD.n581 459.931
R1237 AVDD.n646 AVDD.n643 459.931
R1238 AVDD.n384 AVDD.n381 459.931
R1239 AVDD.n452 AVDD.n449 459.931
R1240 AVDD.n202 AVDD.n199 459.931
R1241 AVDD.n264 AVDD.n261 459.931
R1242 AVDD.n86 AVDD.n83 459.931
R1243 AVDD.n6516 AVDD.n6513 459.931
R1244 AVDD.n6453 AVDD.n6450 459.931
R1245 AVDD.n5964 AVDD.n5961 459.931
R1246 AVDD.n6008 AVDD.n6005 459.931
R1247 AVDD.n5762 AVDD.n5761 459.931
R1248 AVDD.n5760 AVDD.n5759 459.931
R1249 AVDD.n5766 AVDD.n5765 459.931
R1250 AVDD.n116 AVDD.n113 459.931
R1251 AVDD.n6546 AVDD.n6543 459.931
R1252 AVDD.n6483 AVDD.n6480 459.931
R1253 AVDD.n5994 AVDD.n5991 459.931
R1254 AVDD.n608 AVDD.n605 459.931
R1255 AVDD.n670 AVDD.n667 459.931
R1256 AVDD.n408 AVDD.n405 459.931
R1257 AVDD.n476 AVDD.n473 459.931
R1258 AVDD.n226 AVDD.n223 459.931
R1259 AVDD.n288 AVDD.n285 459.931
R1260 AVDD.n110 AVDD.n107 459.931
R1261 AVDD.n6540 AVDD.n6537 459.931
R1262 AVDD.n6477 AVDD.n6474 459.931
R1263 AVDD.n5988 AVDD.n5985 459.931
R1264 AVDD.n104 AVDD.n101 459.931
R1265 AVDD.n6534 AVDD.n6531 459.931
R1266 AVDD.n6471 AVDD.n6468 459.931
R1267 AVDD.n5982 AVDD.n5979 459.931
R1268 AVDD.n620 AVDD.n617 459.931
R1269 AVDD.n634 AVDD.n631 459.931
R1270 AVDD.n420 AVDD.n417 459.931
R1271 AVDD.n440 AVDD.n437 459.931
R1272 AVDD.n238 AVDD.n235 459.931
R1273 AVDD.n252 AVDD.n249 459.931
R1274 AVDD.n122 AVDD.n119 459.931
R1275 AVDD.n6504 AVDD.n6501 459.931
R1276 AVDD.n6459 AVDD.n6456 459.931
R1277 AVDD.n5970 AVDD.n5967 459.931
R1278 AVDD.n92 AVDD.n89 459.931
R1279 AVDD.n6522 AVDD.n6519 459.931
R1280 AVDD.n208 AVDD.n205 459.931
R1281 AVDD.n270 AVDD.n267 459.931
R1282 AVDD.n390 AVDD.n387 459.931
R1283 AVDD.n458 AVDD.n455 459.931
R1284 AVDD.n590 AVDD.n587 459.931
R1285 AVDD.n652 AVDD.n649 459.931
R1286 AVDD.n6465 AVDD.n6462 459.931
R1287 AVDD.n5976 AVDD.n5973 459.931
R1288 AVDD.n98 AVDD.n95 459.931
R1289 AVDD.n6528 AVDD.n6525 459.931
R1290 AVDD.n214 AVDD.n211 459.931
R1291 AVDD.n276 AVDD.n273 459.931
R1292 AVDD.n396 AVDD.n393 459.931
R1293 AVDD.n464 AVDD.n461 459.931
R1294 AVDD.n596 AVDD.n593 459.931
R1295 AVDD.n658 AVDD.n655 459.931
R1296 AVDD.n220 AVDD.n217 459.931
R1297 AVDD.n282 AVDD.n279 459.931
R1298 AVDD.n402 AVDD.n399 459.931
R1299 AVDD.n470 AVDD.n467 459.931
R1300 AVDD.n602 AVDD.n599 459.931
R1301 AVDD.n664 AVDD.n661 459.931
R1302 AVDD.n232 AVDD.n229 459.931
R1303 AVDD.n294 AVDD.n291 459.931
R1304 AVDD.n414 AVDD.n411 459.931
R1305 AVDD.n482 AVDD.n479 459.931
R1306 AVDD.n614 AVDD.n611 459.931
R1307 AVDD.n676 AVDD.n673 459.931
R1308 AVDD.n6489 AVDD.n6486 459.931
R1309 AVDD.n6000 AVDD.n5997 459.931
R1310 AVDD.n6050 AVDD.n6047 459.931
R1311 AVDD.n6274 AVDD.n6273 459.931
R1312 AVDD.n6272 AVDD.n6271 459.931
R1313 AVDD.n6276 AVDD.n6275 459.931
R1314 AVDD.n6044 AVDD.n6041 459.931
R1315 AVDD.n6251 AVDD.n6250 459.931
R1316 AVDD.n6249 AVDD.n6248 459.931
R1317 AVDD.n6253 AVDD.n6252 459.931
R1318 AVDD.n6038 AVDD.n6035 459.931
R1319 AVDD.n6228 AVDD.n6227 459.931
R1320 AVDD.n6226 AVDD.n6225 459.931
R1321 AVDD.n6230 AVDD.n6229 459.931
R1322 AVDD.n6032 AVDD.n6029 459.931
R1323 AVDD.n6205 AVDD.n6204 459.931
R1324 AVDD.n6203 AVDD.n6202 459.931
R1325 AVDD.n6207 AVDD.n6206 459.931
R1326 AVDD.n6026 AVDD.n6023 459.931
R1327 AVDD.n6161 AVDD.n6160 459.931
R1328 AVDD.n6159 AVDD.n6158 459.931
R1329 AVDD.n6185 AVDD.n6162 459.931
R1330 AVDD.n6020 AVDD.n6017 459.931
R1331 AVDD.n6139 AVDD.n6107 459.931
R1332 AVDD.n6106 AVDD.n5801 459.931
R1333 AVDD.n6141 AVDD.n6140 459.931
R1334 AVDD.n5783 AVDD.n5782 459.931
R1335 AVDD.n5779 AVDD.n5778 459.931
R1336 AVDD.n6014 AVDD.n6011 459.931
R1337 AVDD.n5781 AVDD.n5780 459.931
R1338 AVDD.n378 AVDD.n375 459.931
R1339 AVDD.n446 AVDD.n443 459.931
R1340 AVDD.n578 AVDD.n575 459.931
R1341 AVDD.n640 AVDD.n637 459.931
R1342 AVDD.n196 AVDD.n193 459.931
R1343 AVDD.n258 AVDD.n255 459.931
R1344 AVDD.n6447 AVDD.n6444 459.931
R1345 AVDD.n5958 AVDD.n5955 459.931
R1346 AVDD.n80 AVDD.n77 459.931
R1347 AVDD.n6510 AVDD.n6507 459.931
R1348 AVDD.n3821 AVDD.n3813 361.655
R1349 AVDD.n3821 AVDD.n3820 361.655
R1350 AVDD.n3819 AVDD.n3814 361.655
R1351 AVDD.n3819 AVDD.n3815 361.655
R1352 AVDD.n3920 AVDD.n3917 361.655
R1353 AVDD.n3854 AVDD.n3849 361.655
R1354 AVDD.n3868 AVDD.n3864 361.655
R1355 AVDD.n3853 AVDD.n3850 361.655
R1356 AVDD.n3869 AVDD.n3863 361.655
R1357 AVDD.n3936 AVDD.n3930 361.655
R1358 AVDD.n3921 AVDD.n3916 361.655
R1359 AVDD.n3935 AVDD.n3931 361.655
R1360 AVDD.n4135 AVDD.n4132 361.655
R1361 AVDD.n4069 AVDD.n4064 361.655
R1362 AVDD.n4083 AVDD.n4079 361.655
R1363 AVDD.n4068 AVDD.n4065 361.655
R1364 AVDD.n4084 AVDD.n4078 361.655
R1365 AVDD.n4236 AVDD.n4221 361.655
R1366 AVDD.n4236 AVDD.n4235 361.655
R1367 AVDD.n4234 AVDD.n4229 361.655
R1368 AVDD.n4234 AVDD.n4230 361.655
R1369 AVDD.n4151 AVDD.n4145 361.655
R1370 AVDD.n4136 AVDD.n4131 361.655
R1371 AVDD.n4150 AVDD.n4146 361.655
R1372 AVDD.n6085 AVDD.n5808 361.655
R1373 AVDD.n6085 AVDD.n5809 361.655
R1374 AVDD.n5807 AVDD.n5802 361.655
R1375 AVDD.n5807 AVDD.n5803 361.655
R1376 AVDD.n5904 AVDD.n5901 361.655
R1377 AVDD.n5905 AVDD.n5886 361.655
R1378 AVDD.n5924 AVDD.n5913 361.655
R1379 AVDD.n5923 AVDD.n5920 361.655
R1380 AVDD.n3775 AVDD.n3770 361.655
R1381 AVDD.n3774 AVDD.n3771 361.655
R1382 AVDD.n3743 AVDD.n3740 361.655
R1383 AVDD.n3744 AVDD.n3738 361.655
R1384 AVDD.n3803 AVDD.n3801 338.068
R1385 AVDD.n3868 AVDD.n3865 338.068
R1386 AVDD.n3935 AVDD.n3932 338.068
R1387 AVDD.n4083 AVDD.n4080 338.068
R1388 AVDD.n4251 AVDD.n4249 338.068
R1389 AVDD.n4150 AVDD.n4147 338.068
R1390 AVDD.n5840 AVDD.n5838 338.068
R1391 AVDD.n6054 AVDD.n6052 338.068
R1392 AVDD.n3743 AVDD.n3739 338.068
R1393 AVDD.n3960 AVDD.n3827 225.128
R1394 AVDD.n4177 AVDD.n4042 225.128
R1395 AVDD.n3829 AVDD.n3828 185
R1396 AVDD.n4404 AVDD.n4403 185
R1397 AVDD.n4386 AVDD.n4385 185
R1398 AVDD.n4044 AVDD.n4043 185
R1399 AVDD.n140 AVDD.n139 185
R1400 AVDD.n6500 AVDD.n6499 185
R1401 AVDD.n27 AVDD.n26 185
R1402 AVDD.n5758 AVDD.n5757 185
R1403 AVDD.n6375 AVDD.n6374 185
R1404 AVDD.n30 AVDD.n29 185
R1405 AVDD.n3897 AVDD.n3896 172.032
R1406 AVDD.n3963 AVDD.n3962 172.032
R1407 AVDD.n4112 AVDD.n4111 172.032
R1408 AVDD.n3966 AVDD.n3965 163.011
R1409 AVDD.n3833 AVDD.n3832 163.011
R1410 AVDD.n3900 AVDD.n3899 163.011
R1411 AVDD.n4048 AVDD.n4047 163.011
R1412 AVDD.n4115 AVDD.n4114 163.011
R1413 AVDD.n4335 AVDD.t36 152.832
R1414 AVDD.t712 AVDD.n4349 145.566
R1415 AVDD.n3894 AVDD.n3893 142.553
R1416 AVDD.n4109 AVDD.n4108 142.553
R1417 AVDD.n5836 AVDD.n5833 142.544
R1418 AVDD.n24 AVDD.n21 142.544
R1419 AVDD.n66 AVDD.n65 142.541
R1420 AVDD.n6492 AVDD.n6491 142.541
R1421 AVDD.n5900 AVDD.n5899 142.44
R1422 AVDD.n137 AVDD.n136 142.439
R1423 AVDD.n6495 AVDD.n6494 142.439
R1424 AVDD.n4625 AVDD.t701 138.83
R1425 AVDD.n4651 AVDD.t503 138.83
R1426 AVDD.n3054 AVDD.t397 138.83
R1427 AVDD.n2940 AVDD.t611 138.83
R1428 AVDD.n2868 AVDD.t671 138.83
R1429 AVDD.n2352 AVDD.t605 138.83
R1430 AVDD.n2172 AVDD.t491 138.83
R1431 AVDD.n1657 AVDD.t686 138.83
R1432 AVDD.n1538 AVDD.t566 138.83
R1433 AVDD.n1470 AVDD.t452 138.83
R1434 AVDD.n4656 AVDD.t548 138.83
R1435 AVDD.n5041 AVDD.t521 138.83
R1436 AVDD.n1629 AVDD.t545 138.83
R1437 AVDD.n1539 AVDD.t680 138.83
R1438 AVDD.n2375 AVDD.t596 138.83
R1439 AVDD.n2353 AVDD.t377 138.83
R1440 AVDD.n3009 AVDD.t467 138.83
R1441 AVDD.n3031 AVDD.t387 138.83
R1442 AVDD.n1708 AVDD.t485 138.83
R1443 AVDD.n3121 AVDD.t509 138.83
R1444 AVDD.n5019 AVDD.t632 138.83
R1445 AVDD.n4631 AVDD.t668 138.83
R1446 AVDD.n4636 AVDD.t515 138.83
R1447 AVDD.n4638 AVDD.t365 138.83
R1448 AVDD.n4642 AVDD.t416 138.83
R1449 AVDD.n4644 AVDD.t608 138.83
R1450 AVDD.n4647 AVDD.t476 138.83
R1451 AVDD.n4628 AVDD.t650 138.83
R1452 AVDD.n1632 AVDD.t404 138.83
R1453 AVDD.n1634 AVDD.t599 138.83
R1454 AVDD.n1636 AVDD.t638 138.83
R1455 AVDD.n1638 AVDD.t497 138.83
R1456 AVDD.n1640 AVDD.t683 138.83
R1457 AVDD.n1642 AVDD.t527 138.83
R1458 AVDD.n1644 AVDD.t393 138.83
R1459 AVDD.n1646 AVDD.t590 138.83
R1460 AVDD.n3948 AVDD.n3947 128.687
R1461 AVDD.n4163 AVDD.n4162 128.687
R1462 AVDD.n3962 AVDD.n3825 127.764
R1463 AVDD.n4179 AVDD.n4040 127.764
R1464 AVDD.n3 AVDD.n2 121.193
R1465 AVDD.n5852 AVDD.n5851 121.193
R1466 AVDD.n5826 AVDD.n5825 121.193
R1467 AVDD.n3892 AVDD.n3891 121.098
R1468 AVDD.n3795 AVDD.n3794 121.098
R1469 AVDD.n4107 AVDD.n4106 121.098
R1470 AVDD.n5 AVDD.n4 121.098
R1471 AVDD.n5854 AVDD.n5853 121.098
R1472 AVDD.n3960 AVDD.n3959 119.34
R1473 AVDD.n4177 AVDD.n4176 119.34
R1474 AVDD.n4281 AVDD.t33 116.344
R1475 AVDD.n5895 AVDD.n5894 113.839
R1476 AVDD.t38 AVDD.t722 113.368
R1477 AVDD.t748 AVDD.t747 113.368
R1478 AVDD.n3979 AVDD.n3978 107.2
R1479 AVDD.n3846 AVDD.n3845 107.2
R1480 AVDD.n3913 AVDD.n3912 107.2
R1481 AVDD.n4061 AVDD.n4060 107.2
R1482 AVDD.n4128 AVDD.n4127 107.2
R1483 AVDD.n3959 AVDD.t262 105.788
R1484 AVDD.n4176 AVDD.t765 105.788
R1485 AVDD.n3825 AVDD.n3824 101.581
R1486 AVDD.n4040 AVDD.n4039 101.581
R1487 AVDD.n3947 AVDD.n3946 101.515
R1488 AVDD.n4162 AVDD.n4161 101.515
R1489 AVDD.n5700 AVDD.n5699 96.007
R1490 AVDD.n1366 AVDD.n1365 92.965
R1491 AVDD.n6376 AVDD.n6370 92.665
R1492 AVDD.n195 AVDD.n194 92.611
R1493 AVDD.n257 AVDD.n256 92.611
R1494 AVDD.n377 AVDD.n376 92.611
R1495 AVDD.n445 AVDD.n444 92.611
R1496 AVDD.n577 AVDD.n576 92.611
R1497 AVDD.n639 AVDD.n638 92.611
R1498 AVDD.n758 AVDD.n757 92.611
R1499 AVDD.n820 AVDD.n819 92.611
R1500 AVDD.n939 AVDD.n938 92.611
R1501 AVDD.n1001 AVDD.n1000 92.611
R1502 AVDD.n1300 AVDD.n1299 92.611
R1503 AVDD.n1106 AVDD.n1105 92.611
R1504 AVDD.n1207 AVDD.n1206 92.611
R1505 AVDD.n1482 AVDD.n1481 92.611
R1506 AVDD.n1570 AVDD.n1569 92.611
R1507 AVDD.n1663 AVDD.n1662 92.611
R1508 AVDD.n1779 AVDD.n1778 92.611
R1509 AVDD.n1924 AVDD.n1923 92.611
R1510 AVDD.n1991 AVDD.n1990 92.611
R1511 AVDD.n2195 AVDD.n2194 92.611
R1512 AVDD.n2070 AVDD.n2069 92.611
R1513 AVDD.n2296 AVDD.n2295 92.611
R1514 AVDD.n2406 AVDD.n2405 92.611
R1515 AVDD.n2476 AVDD.n2475 92.611
R1516 AVDD.n2570 AVDD.n2569 92.611
R1517 AVDD.n2721 AVDD.n2720 92.611
R1518 AVDD.n2788 AVDD.n2787 92.611
R1519 AVDD.n2884 AVDD.n2883 92.611
R1520 AVDD.n2950 AVDD.n2949 92.611
R1521 AVDD.n3065 AVDD.n3064 92.611
R1522 AVDD.n3175 AVDD.n3174 92.611
R1523 AVDD.n3284 AVDD.n3283 92.611
R1524 AVDD.n3349 AVDD.n3348 92.611
R1525 AVDD.n4763 AVDD.n4762 92.611
R1526 AVDD.n4714 AVDD.n4713 92.611
R1527 AVDD.n4939 AVDD.n4938 92.611
R1528 AVDD.n5957 AVDD.n5956 92.611
R1529 AVDD.n6446 AVDD.n6445 92.611
R1530 AVDD.n6007 AVDD.n6006 92.611
R1531 AVDD.n6043 AVDD.n6042 92.611
R1532 AVDD.n6482 AVDD.n6481 92.611
R1533 AVDD.n5993 AVDD.n5992 92.611
R1534 AVDD.n115 AVDD.n114 92.611
R1535 AVDD.n6545 AVDD.n6544 92.611
R1536 AVDD.n231 AVDD.n230 92.611
R1537 AVDD.n293 AVDD.n292 92.611
R1538 AVDD.n413 AVDD.n412 92.611
R1539 AVDD.n481 AVDD.n480 92.611
R1540 AVDD.n613 AVDD.n612 92.611
R1541 AVDD.n675 AVDD.n674 92.611
R1542 AVDD.n794 AVDD.n793 92.611
R1543 AVDD.n856 AVDD.n855 92.611
R1544 AVDD.n975 AVDD.n974 92.611
R1545 AVDD.n1037 AVDD.n1036 92.611
R1546 AVDD.n1336 AVDD.n1335 92.611
R1547 AVDD.n1142 AVDD.n1141 92.611
R1548 AVDD.n1243 AVDD.n1242 92.611
R1549 AVDD.n1402 AVDD.n1401 92.611
R1550 AVDD.n1518 AVDD.n1517 92.611
R1551 AVDD.n1606 AVDD.n1605 92.611
R1552 AVDD.n1699 AVDD.n1698 92.611
R1553 AVDD.n1815 AVDD.n1814 92.611
R1554 AVDD.n1960 AVDD.n1959 92.611
R1555 AVDD.n2027 AVDD.n2026 92.611
R1556 AVDD.n2332 AVDD.n2331 92.611
R1557 AVDD.n2442 AVDD.n2441 92.611
R1558 AVDD.n2512 AVDD.n2511 92.611
R1559 AVDD.n2606 AVDD.n2605 92.611
R1560 AVDD.n2757 AVDD.n2756 92.611
R1561 AVDD.n2824 AVDD.n2823 92.611
R1562 AVDD.n2920 AVDD.n2919 92.611
R1563 AVDD.n2986 AVDD.n2985 92.611
R1564 AVDD.n3101 AVDD.n3100 92.611
R1565 AVDD.n3211 AVDD.n3210 92.611
R1566 AVDD.n3320 AVDD.n3319 92.611
R1567 AVDD.n3385 AVDD.n3384 92.611
R1568 AVDD.n4750 AVDD.n4749 92.611
R1569 AVDD.n4975 AVDD.n4974 92.611
R1570 AVDD.n4799 AVDD.n4798 92.611
R1571 AVDD.n4793 AVDD.n4792 92.611
R1572 AVDD.n4744 AVDD.n4743 92.611
R1573 AVDD.n4969 AVDD.n4968 92.611
R1574 AVDD.n3314 AVDD.n3313 92.611
R1575 AVDD.n3379 AVDD.n3378 92.611
R1576 AVDD.n3095 AVDD.n3094 92.611
R1577 AVDD.n3205 AVDD.n3204 92.611
R1578 AVDD.n2914 AVDD.n2913 92.611
R1579 AVDD.n2980 AVDD.n2979 92.611
R1580 AVDD.n2751 AVDD.n2750 92.611
R1581 AVDD.n2818 AVDD.n2817 92.611
R1582 AVDD.n2506 AVDD.n2505 92.611
R1583 AVDD.n2600 AVDD.n2599 92.611
R1584 AVDD.n2326 AVDD.n2325 92.611
R1585 AVDD.n2436 AVDD.n2435 92.611
R1586 AVDD.n2225 AVDD.n2224 92.611
R1587 AVDD.n2100 AVDD.n2099 92.611
R1588 AVDD.n1954 AVDD.n1953 92.611
R1589 AVDD.n2021 AVDD.n2020 92.611
R1590 AVDD.n1693 AVDD.n1692 92.611
R1591 AVDD.n1809 AVDD.n1808 92.611
R1592 AVDD.n1512 AVDD.n1511 92.611
R1593 AVDD.n1600 AVDD.n1599 92.611
R1594 AVDD.n1237 AVDD.n1236 92.611
R1595 AVDD.n1396 AVDD.n1395 92.611
R1596 AVDD.n1330 AVDD.n1329 92.611
R1597 AVDD.n1136 AVDD.n1135 92.611
R1598 AVDD.n969 AVDD.n968 92.611
R1599 AVDD.n1031 AVDD.n1030 92.611
R1600 AVDD.n788 AVDD.n787 92.611
R1601 AVDD.n850 AVDD.n849 92.611
R1602 AVDD.n607 AVDD.n606 92.611
R1603 AVDD.n669 AVDD.n668 92.611
R1604 AVDD.n407 AVDD.n406 92.611
R1605 AVDD.n475 AVDD.n474 92.611
R1606 AVDD.n225 AVDD.n224 92.611
R1607 AVDD.n287 AVDD.n286 92.611
R1608 AVDD.n109 AVDD.n108 92.611
R1609 AVDD.n6539 AVDD.n6538 92.611
R1610 AVDD.n6476 AVDD.n6475 92.611
R1611 AVDD.n5987 AVDD.n5986 92.611
R1612 AVDD.n6037 AVDD.n6036 92.611
R1613 AVDD.n4787 AVDD.n4786 92.611
R1614 AVDD.n4738 AVDD.n4737 92.611
R1615 AVDD.n4963 AVDD.n4962 92.611
R1616 AVDD.n3308 AVDD.n3307 92.611
R1617 AVDD.n3373 AVDD.n3372 92.611
R1618 AVDD.n3089 AVDD.n3088 92.611
R1619 AVDD.n3199 AVDD.n3198 92.611
R1620 AVDD.n2908 AVDD.n2907 92.611
R1621 AVDD.n2974 AVDD.n2973 92.611
R1622 AVDD.n2745 AVDD.n2744 92.611
R1623 AVDD.n2812 AVDD.n2811 92.611
R1624 AVDD.n2500 AVDD.n2499 92.611
R1625 AVDD.n2594 AVDD.n2593 92.611
R1626 AVDD.n2320 AVDD.n2319 92.611
R1627 AVDD.n2430 AVDD.n2429 92.611
R1628 AVDD.n2219 AVDD.n2218 92.611
R1629 AVDD.n2094 AVDD.n2093 92.611
R1630 AVDD.n1948 AVDD.n1947 92.611
R1631 AVDD.n2015 AVDD.n2014 92.611
R1632 AVDD.n1687 AVDD.n1686 92.611
R1633 AVDD.n1803 AVDD.n1802 92.611
R1634 AVDD.n1506 AVDD.n1505 92.611
R1635 AVDD.n1594 AVDD.n1593 92.611
R1636 AVDD.n1231 AVDD.n1230 92.611
R1637 AVDD.n1390 AVDD.n1389 92.611
R1638 AVDD.n1324 AVDD.n1323 92.611
R1639 AVDD.n1130 AVDD.n1129 92.611
R1640 AVDD.n963 AVDD.n962 92.611
R1641 AVDD.n1025 AVDD.n1024 92.611
R1642 AVDD.n782 AVDD.n781 92.611
R1643 AVDD.n844 AVDD.n843 92.611
R1644 AVDD.n601 AVDD.n600 92.611
R1645 AVDD.n663 AVDD.n662 92.611
R1646 AVDD.n401 AVDD.n400 92.611
R1647 AVDD.n469 AVDD.n468 92.611
R1648 AVDD.n219 AVDD.n218 92.611
R1649 AVDD.n281 AVDD.n280 92.611
R1650 AVDD.n103 AVDD.n102 92.611
R1651 AVDD.n6533 AVDD.n6532 92.611
R1652 AVDD.n6470 AVDD.n6469 92.611
R1653 AVDD.n5981 AVDD.n5980 92.611
R1654 AVDD.n6031 AVDD.n6030 92.611
R1655 AVDD.n4781 AVDD.n4780 92.611
R1656 AVDD.n4732 AVDD.n4731 92.611
R1657 AVDD.n4957 AVDD.n4956 92.611
R1658 AVDD.n3302 AVDD.n3301 92.611
R1659 AVDD.n3367 AVDD.n3366 92.611
R1660 AVDD.n3083 AVDD.n3082 92.611
R1661 AVDD.n3193 AVDD.n3192 92.611
R1662 AVDD.n2902 AVDD.n2901 92.611
R1663 AVDD.n2968 AVDD.n2967 92.611
R1664 AVDD.n2739 AVDD.n2738 92.611
R1665 AVDD.n2806 AVDD.n2805 92.611
R1666 AVDD.n2494 AVDD.n2493 92.611
R1667 AVDD.n2588 AVDD.n2587 92.611
R1668 AVDD.n2314 AVDD.n2313 92.611
R1669 AVDD.n2424 AVDD.n2423 92.611
R1670 AVDD.n2213 AVDD.n2212 92.611
R1671 AVDD.n2088 AVDD.n2087 92.611
R1672 AVDD.n1942 AVDD.n1941 92.611
R1673 AVDD.n2009 AVDD.n2008 92.611
R1674 AVDD.n1681 AVDD.n1680 92.611
R1675 AVDD.n1797 AVDD.n1796 92.611
R1676 AVDD.n1500 AVDD.n1499 92.611
R1677 AVDD.n1588 AVDD.n1587 92.611
R1678 AVDD.n1225 AVDD.n1224 92.611
R1679 AVDD.n1384 AVDD.n1383 92.611
R1680 AVDD.n1318 AVDD.n1317 92.611
R1681 AVDD.n1124 AVDD.n1123 92.611
R1682 AVDD.n957 AVDD.n956 92.611
R1683 AVDD.n1019 AVDD.n1018 92.611
R1684 AVDD.n776 AVDD.n775 92.611
R1685 AVDD.n838 AVDD.n837 92.611
R1686 AVDD.n595 AVDD.n594 92.611
R1687 AVDD.n657 AVDD.n656 92.611
R1688 AVDD.n395 AVDD.n394 92.611
R1689 AVDD.n463 AVDD.n462 92.611
R1690 AVDD.n213 AVDD.n212 92.611
R1691 AVDD.n275 AVDD.n274 92.611
R1692 AVDD.n97 AVDD.n96 92.611
R1693 AVDD.n6527 AVDD.n6526 92.611
R1694 AVDD.n6464 AVDD.n6463 92.611
R1695 AVDD.n5975 AVDD.n5974 92.611
R1696 AVDD.n6025 AVDD.n6024 92.611
R1697 AVDD.n4775 AVDD.n4774 92.611
R1698 AVDD.n4726 AVDD.n4725 92.611
R1699 AVDD.n4951 AVDD.n4950 92.611
R1700 AVDD.n3296 AVDD.n3295 92.611
R1701 AVDD.n3361 AVDD.n3360 92.611
R1702 AVDD.n3077 AVDD.n3076 92.611
R1703 AVDD.n3187 AVDD.n3186 92.611
R1704 AVDD.n2896 AVDD.n2895 92.611
R1705 AVDD.n2962 AVDD.n2961 92.611
R1706 AVDD.n2733 AVDD.n2732 92.611
R1707 AVDD.n2800 AVDD.n2799 92.611
R1708 AVDD.n2488 AVDD.n2487 92.611
R1709 AVDD.n2582 AVDD.n2581 92.611
R1710 AVDD.n2308 AVDD.n2307 92.611
R1711 AVDD.n2418 AVDD.n2417 92.611
R1712 AVDD.n2207 AVDD.n2206 92.611
R1713 AVDD.n2082 AVDD.n2081 92.611
R1714 AVDD.n1936 AVDD.n1935 92.611
R1715 AVDD.n2003 AVDD.n2002 92.611
R1716 AVDD.n1675 AVDD.n1674 92.611
R1717 AVDD.n1791 AVDD.n1790 92.611
R1718 AVDD.n1494 AVDD.n1493 92.611
R1719 AVDD.n1582 AVDD.n1581 92.611
R1720 AVDD.n1219 AVDD.n1218 92.611
R1721 AVDD.n1378 AVDD.n1377 92.611
R1722 AVDD.n1312 AVDD.n1311 92.611
R1723 AVDD.n1118 AVDD.n1117 92.611
R1724 AVDD.n951 AVDD.n950 92.611
R1725 AVDD.n1013 AVDD.n1012 92.611
R1726 AVDD.n770 AVDD.n769 92.611
R1727 AVDD.n832 AVDD.n831 92.611
R1728 AVDD.n589 AVDD.n588 92.611
R1729 AVDD.n651 AVDD.n650 92.611
R1730 AVDD.n389 AVDD.n388 92.611
R1731 AVDD.n457 AVDD.n456 92.611
R1732 AVDD.n207 AVDD.n206 92.611
R1733 AVDD.n269 AVDD.n268 92.611
R1734 AVDD.n91 AVDD.n90 92.611
R1735 AVDD.n6521 AVDD.n6520 92.611
R1736 AVDD.n6458 AVDD.n6457 92.611
R1737 AVDD.n5969 AVDD.n5968 92.611
R1738 AVDD.n6019 AVDD.n6018 92.611
R1739 AVDD.n4769 AVDD.n4768 92.611
R1740 AVDD.n4720 AVDD.n4719 92.611
R1741 AVDD.n4945 AVDD.n4944 92.611
R1742 AVDD.n3290 AVDD.n3289 92.611
R1743 AVDD.n3355 AVDD.n3354 92.611
R1744 AVDD.n3071 AVDD.n3070 92.611
R1745 AVDD.n3181 AVDD.n3180 92.611
R1746 AVDD.n2890 AVDD.n2889 92.611
R1747 AVDD.n2956 AVDD.n2955 92.611
R1748 AVDD.n2727 AVDD.n2726 92.611
R1749 AVDD.n2794 AVDD.n2793 92.611
R1750 AVDD.n2482 AVDD.n2481 92.611
R1751 AVDD.n2576 AVDD.n2575 92.611
R1752 AVDD.n2302 AVDD.n2301 92.611
R1753 AVDD.n2412 AVDD.n2411 92.611
R1754 AVDD.n2201 AVDD.n2200 92.611
R1755 AVDD.n2076 AVDD.n2075 92.611
R1756 AVDD.n1930 AVDD.n1929 92.611
R1757 AVDD.n1997 AVDD.n1996 92.611
R1758 AVDD.n1669 AVDD.n1668 92.611
R1759 AVDD.n1785 AVDD.n1784 92.611
R1760 AVDD.n1488 AVDD.n1487 92.611
R1761 AVDD.n1576 AVDD.n1575 92.611
R1762 AVDD.n1213 AVDD.n1212 92.611
R1763 AVDD.n1372 AVDD.n1371 92.611
R1764 AVDD.n1306 AVDD.n1305 92.611
R1765 AVDD.n1112 AVDD.n1111 92.611
R1766 AVDD.n945 AVDD.n944 92.611
R1767 AVDD.n1007 AVDD.n1006 92.611
R1768 AVDD.n764 AVDD.n763 92.611
R1769 AVDD.n826 AVDD.n825 92.611
R1770 AVDD.n583 AVDD.n582 92.611
R1771 AVDD.n645 AVDD.n644 92.611
R1772 AVDD.n383 AVDD.n382 92.611
R1773 AVDD.n451 AVDD.n450 92.611
R1774 AVDD.n201 AVDD.n200 92.611
R1775 AVDD.n263 AVDD.n262 92.611
R1776 AVDD.n85 AVDD.n84 92.611
R1777 AVDD.n6515 AVDD.n6514 92.611
R1778 AVDD.n6452 AVDD.n6451 92.611
R1779 AVDD.n5963 AVDD.n5962 92.611
R1780 AVDD.n6013 AVDD.n6012 92.611
R1781 AVDD.n2231 AVDD.n2230 92.611
R1782 AVDD.n2106 AVDD.n2105 92.611
R1783 AVDD.n6488 AVDD.n6487 92.611
R1784 AVDD.n5999 AVDD.n5998 92.611
R1785 AVDD.n121 AVDD.n120 92.611
R1786 AVDD.n6503 AVDD.n6502 92.611
R1787 AVDD.n237 AVDD.n236 92.611
R1788 AVDD.n251 AVDD.n250 92.611
R1789 AVDD.n419 AVDD.n418 92.611
R1790 AVDD.n439 AVDD.n438 92.611
R1791 AVDD.n619 AVDD.n618 92.611
R1792 AVDD.n633 AVDD.n632 92.611
R1793 AVDD.n800 AVDD.n799 92.611
R1794 AVDD.n814 AVDD.n813 92.611
R1795 AVDD.n981 AVDD.n980 92.611
R1796 AVDD.n995 AVDD.n994 92.611
R1797 AVDD.n1342 AVDD.n1341 92.611
R1798 AVDD.n1100 AVDD.n1099 92.611
R1799 AVDD.n1249 AVDD.n1248 92.611
R1800 AVDD.n1359 AVDD.n1358 92.611
R1801 AVDD.n1524 AVDD.n1523 92.611
R1802 AVDD.n1564 AVDD.n1563 92.611
R1803 AVDD.n1705 AVDD.n1704 92.611
R1804 AVDD.n1773 AVDD.n1772 92.611
R1805 AVDD.n1966 AVDD.n1965 92.611
R1806 AVDD.n1985 AVDD.n1984 92.611
R1807 AVDD.n2237 AVDD.n2236 92.611
R1808 AVDD.n2064 AVDD.n2063 92.611
R1809 AVDD.n2338 AVDD.n2337 92.611
R1810 AVDD.n2400 AVDD.n2399 92.611
R1811 AVDD.n2518 AVDD.n2517 92.611
R1812 AVDD.n2564 AVDD.n2563 92.611
R1813 AVDD.n2763 AVDD.n2762 92.611
R1814 AVDD.n2782 AVDD.n2781 92.611
R1815 AVDD.n2926 AVDD.n2925 92.611
R1816 AVDD.n2944 AVDD.n2943 92.611
R1817 AVDD.n3107 AVDD.n3106 92.611
R1818 AVDD.n3169 AVDD.n3168 92.611
R1819 AVDD.n3326 AVDD.n3325 92.611
R1820 AVDD.n3343 AVDD.n3342 92.611
R1821 AVDD.n4756 AVDD.n4755 92.611
R1822 AVDD.n4933 AVDD.n4932 92.611
R1823 AVDD.n4805 AVDD.n4804 92.611
R1824 AVDD.n6049 AVDD.n6048 92.611
R1825 AVDD.n6509 AVDD.n6508 92.611
R1826 AVDD.n79 AVDD.n78 92.611
R1827 AVDD.n3794 AVDD.n3793 82.551
R1828 AVDD.n3891 AVDD.n3890 82.551
R1829 AVDD.n3946 AVDD.n3945 82.551
R1830 AVDD.n4106 AVDD.n4105 82.551
R1831 AVDD.n4403 AVDD.n4402 82.551
R1832 AVDD.n4161 AVDD.n4160 82.551
R1833 AVDD.n5825 AVDD.n5824 80.586
R1834 AVDD.n5851 AVDD.n5850 80.586
R1835 AVDD.n2 AVDD.n1 80.586
R1836 AVDD.n5919 AVDD.n5918 79.572
R1837 AVDD.n23 AVDD.n22 79.572
R1838 AVDD.n6410 AVDD.n11 79.572
R1839 AVDD.n5835 AVDD.n5834 79.572
R1840 AVDD.n3879 AVDD.n3878 79.325
R1841 AVDD.n3784 AVDD.n3783 79.325
R1842 AVDD.n4094 AVDD.n4093 79.325
R1843 AVDD.n3896 AVDD.n3829 78.37
R1844 AVDD.n4111 AVDD.n4044 78.37
R1845 AVDD.n3818 AVDD.n3816 73.788
R1846 AVDD.n3818 AVDD.n3817 73.788
R1847 AVDD.n3867 AVDD.n3866 73.788
R1848 AVDD.n3852 AVDD.n3851 73.788
R1849 AVDD.n3934 AVDD.n3933 73.788
R1850 AVDD.n3919 AVDD.n3918 73.788
R1851 AVDD.n4082 AVDD.n4081 73.788
R1852 AVDD.n4067 AVDD.n4066 73.788
R1853 AVDD.n4233 AVDD.n4231 73.788
R1854 AVDD.n4233 AVDD.n4232 73.788
R1855 AVDD.n4149 AVDD.n4148 73.788
R1856 AVDD.n4134 AVDD.n4133 73.788
R1857 AVDD.n3773 AVDD.n3772 73.788
R1858 AVDD.n3742 AVDD.n3741 73.788
R1859 AVDD.n5806 AVDD.n5804 73.788
R1860 AVDD.n5806 AVDD.n5805 73.788
R1861 AVDD.n5903 AVDD.n5902 73.788
R1862 AVDD.n5922 AVDD.n5921 73.788
R1863 AVDD.n4348 AVDD.n4344 69.532
R1864 AVDD.n3893 AVDD.t142 69.302
R1865 AVDD.n4108 AVDD.t745 69.302
R1866 AVDD.t739 AVDD.n4036 69.302
R1867 AVDD.t52 AVDD.n5826 69.302
R1868 AVDD.t275 AVDD.n5852 69.302
R1869 AVDD.t31 AVDD.n3 69.302
R1870 AVDD.t731 AVDD.n3795 69.001
R1871 AVDD.t142 AVDD.n3892 69.001
R1872 AVDD.t745 AVDD.n4107 69.001
R1873 AVDD.t739 AVDD.n4037 69.001
R1874 AVDD.t275 AVDD.n5854 69.001
R1875 AVDD.t31 AVDD.n5 69.001
R1876 AVDD.n4350 AVDD.t712 68.164
R1877 AVDD.t57 AVDD.t58 67.249
R1878 AVDD.t154 AVDD.t153 67.249
R1879 AVDD.t4 AVDD.t152 67.249
R1880 AVDD.n5888 AVDD.n5887 66.321
R1881 AVDD.t709 AVDD.t721 64.269
R1882 AVDD.n1346 AVDD.n1345 61.804
R1883 AVDD.n134 AVDD.n133 57.682
R1884 AVDD.n4371 AVDD.t37 56.684
R1885 AVDD.n4371 AVDD.t38 56.684
R1886 AVDD.n4294 AVDD.t748 56.684
R1887 AVDD.n4294 AVDD.t39 56.684
R1888 level_shifter_up_5.VDD_HV AVDD.t53 56.029
R1889 AVDD.n3791 AVDD.t732 56.027
R1890 AVDD.n3830 AVDD.t143 56.027
R1891 AVDD.n3958 AVDD.t263 56.027
R1892 AVDD.n4045 AVDD.t746 56.027
R1893 AVDD.n4035 AVDD.t740 56.027
R1894 AVDD.n4175 AVDD.t766 56.027
R1895 AVDD.n6069 AVDD.t276 56.027
R1896 AVDD.n0 AVDD.t32 56.027
R1897 AVDD.n4296 AVDD.n4291 55.036
R1898 AVDD.t152 AVDD.n4379 54.48
R1899 AVDD.t709 AVDD.t61 48.947
R1900 AVDD.n4304 AVDD.n4268 48.202
R1901 AVDD.n4486 AVDD.t482 48.2
R1902 AVDD.n4491 AVDD.t569 48.2
R1903 AVDD.n4588 AVDD.t551 48.2
R1904 AVDD.n4536 AVDD.t373 48.2
R1905 AVDD.n4504 AVDD.t533 48.2
R1906 AVDD.n4428 AVDD.t698 48.2
R1907 AVDD.n3725 AVDD.t524 48.2
R1908 AVDD.n3555 AVDD.t665 48.2
R1909 AVDD.n3467 AVDD.t644 48.2
R1910 AVDD.n3469 AVDD.t512 48.2
R1911 AVDD.n5764 AVDD.t674 48.2
R1912 AVDD.n5763 AVDD.t369 48.2
R1913 AVDD.n5776 AVDD.t410 48.2
R1914 AVDD.n5793 AVDD.t704 48.2
R1915 AVDD.n5800 AVDD.t587 48.2
R1916 AVDD.n6143 AVDD.t542 48.2
R1917 AVDD.n6157 AVDD.t443 48.2
R1918 AVDD.n6187 AVDD.t407 48.2
R1919 AVDD.n6200 AVDD.t620 48.2
R1920 AVDD.n6209 AVDD.t578 48.2
R1921 AVDD.n6224 AVDD.t455 48.2
R1922 AVDD.n6232 AVDD.t422 48.2
R1923 AVDD.n4555 AVDD.t434 48.2
R1924 AVDD.n4527 AVDD.t575 48.2
R1925 AVDD.n4451 AVDD.t419 48.2
R1926 AVDD.n4423 AVDD.t557 48.2
R1927 AVDD.n3716 AVDD.t384 48.2
R1928 AVDD.n3546 AVDD.t530 48.2
R1929 AVDD.n6247 AVDD.t635 48.2
R1930 AVDD.n6255 AVDD.t602 48.2
R1931 AVDD.n6270 AVDD.t689 48.2
R1932 AVDD.n6278 AVDD.t536 48.2
R1933 AVDD.n4182 AVDD.n4179 46.644
R1934 AVDD.n1430 AVDD.n1428 46.545
R1935 AVDD.n1430 AVDD.n1429 46.545
R1936 AVDD.n1439 AVDD.n1438 46.545
R1937 AVDD.n1444 AVDD.n1443 46.545
R1938 AVDD.n1449 AVDD.n1448 46.545
R1939 AVDD.n1454 AVDD.n1453 46.545
R1940 AVDD.n1463 AVDD.n1462 45.228
R1941 AVDD.t749 AVDD.n4185 43.95
R1942 AVDD.n4409 AVDD.n3984 40.642
R1943 AVDD.n5665 AVDD.n5663 40.069
R1944 AVDD.n5665 AVDD.n5664 40.069
R1945 AVDD.n33 AVDD.n31 40.069
R1946 AVDD.n33 AVDD.n32 40.069
R1947 AVDD.n151 AVDD.n149 40.069
R1948 AVDD.n151 AVDD.n150 40.069
R1949 AVDD.n329 AVDD.n327 40.069
R1950 AVDD.n329 AVDD.n328 40.069
R1951 AVDD.n519 AVDD.n517 40.069
R1952 AVDD.n519 AVDD.n518 40.069
R1953 AVDD.n714 AVDD.n712 40.069
R1954 AVDD.n714 AVDD.n713 40.069
R1955 AVDD.n895 AVDD.n893 40.069
R1956 AVDD.n895 AVDD.n894 40.069
R1957 AVDD.n1066 AVDD.n1064 40.069
R1958 AVDD.n1066 AVDD.n1065 40.069
R1959 AVDD.n5591 AVDD.n5589 40.069
R1960 AVDD.n5591 AVDD.n5590 40.069
R1961 AVDD.n5540 AVDD.n5538 40.069
R1962 AVDD.n5540 AVDD.n5539 40.069
R1963 AVDD.n5495 AVDD.n5493 40.069
R1964 AVDD.n5495 AVDD.n5494 40.069
R1965 AVDD.n5444 AVDD.n5442 40.069
R1966 AVDD.n5444 AVDD.n5443 40.069
R1967 AVDD.n5391 AVDD.n5389 40.069
R1968 AVDD.n5391 AVDD.n5390 40.069
R1969 AVDD.n5345 AVDD.n5343 40.069
R1970 AVDD.n5345 AVDD.n5344 40.069
R1971 AVDD.n5294 AVDD.n5292 40.069
R1972 AVDD.n5294 AVDD.n5293 40.069
R1973 AVDD.n5244 AVDD.n5242 40.069
R1974 AVDD.n5244 AVDD.n5243 40.069
R1975 AVDD.n5196 AVDD.n5194 40.069
R1976 AVDD.n5196 AVDD.n5195 40.069
R1977 AVDD.n5145 AVDD.n5143 40.069
R1978 AVDD.n5145 AVDD.n5144 40.069
R1979 AVDD.n5094 AVDD.n5092 40.069
R1980 AVDD.n5094 AVDD.n5093 40.069
R1981 AVDD.n4902 AVDD.n4900 40.069
R1982 AVDD.n4902 AVDD.n4901 40.069
R1983 AVDD.n4690 AVDD.n4689 40.069
R1984 AVDD.n6356 AVDD.n6355 40.069
R1985 AVDD.n4203 AVDD.n4202 38.213
R1986 AVDD.n5915 AVDD.n5914 37.979
R1987 AVDD.t741 AVDD.n3756 37.472
R1988 AVDD.n3761 AVDD.n3758 36.297
R1989 AVDD.n4301 AVDD.t57 33.624
R1990 AVDD.n4301 AVDD.t711 33.624
R1991 AVDD.n4024 AVDD.t718 33.624
R1992 AVDD.n4378 AVDD.t154 33.624
R1993 AVDD.n4367 AVDD.n4358 32.376
R1994 AVDD.n4375 AVDD.n4330 32.23
R1995 AVDD.n4297 AVDD.n4283 31.722
R1996 AVDD.n4368 AVDD.n4352 31.722
R1997 AVDD.n4298 AVDD.n4276 31.623
R1998 AVDD.n4021 AVDD.n4006 31.623
R1999 AVDD.n3997 AVDD.n3992 31.623
R2000 AVDD.n4309 AVDD.n4265 31.623
R2001 AVDD.n4374 AVDD.n4338 31.623
R2002 AVDD.t709 AVDD.n4326 26.388
R2003 AVDD.n4018 AVDD.n4017 24.686
R2004 AVDD.n6359 AVDD.n5662 24.47
R2005 AVDD.n1276 AVDD.n1275 24.189
R2006 AVDD.n4376 AVDD.n4375 24
R2007 AVDD.n4374 AVDD.n4373 24
R2008 AVDD.n4373 AVDD.n4368 24
R2009 AVDD.n4297 AVDD.n4296 24
R2010 AVDD.n4303 AVDD.n4298 24
R2011 AVDD.t818 AVDD.n5919 21.638
R2012 AVDD.n1271 AVDD.n1270 21.107
R2013 AVDD.n4207 AVDD.t192 21.046
R2014 AVDD.n4266 AVDD.t56 20.855
R2015 AVDD.n3953 AVDD.n3952 20.329
R2016 AVDD.n4168 AVDD.n4167 20.329
R2017 AVDD.n4495 AVDD.n4494 20.22
R2018 AVDD.n3781 AVDD.n3780 20.034
R2019 AVDD.n3876 AVDD.n3875 20.034
R2020 AVDD.n3943 AVDD.n3942 20.034
R2021 AVDD.n4091 AVDD.n4090 20.034
R2022 AVDD.n4033 AVDD.n4032 20.034
R2023 AVDD.n4158 AVDD.n4157 20.034
R2024 AVDD.n6416 AVDD.n6415 20.034
R2025 AVDD.n5822 AVDD.n5821 20.034
R2026 AVDD.n5881 AVDD.n5880 20.034
R2027 AVDD.n135 AVDD.n134 20.023
R2028 AVDD.t185 AVDD.n4378 20.004
R2029 AVDD.n3789 AVDD.n3788 19.756
R2030 AVDD.n3884 AVDD.n3883 19.756
R2031 AVDD.n3954 AVDD.n3953 19.756
R2032 AVDD.n4099 AVDD.n4098 19.756
R2033 AVDD.n4396 AVDD.n4395 19.756
R2034 AVDD.n4169 AVDD.n4168 19.756
R2035 AVDD.n9 AVDD.n8 19.756
R2036 AVDD.n5811 AVDD.n5810 19.756
R2037 AVDD.n5856 AVDD.n5855 19.756
R2038 AVDD.n1276 AVDD.n1274 18.773
R2039 AVDD.n5650 AVDD.t5 18.648
R2040 AVDD.n5650 AVDD.t12 18.648
R2041 AVDD.n5642 AVDD.t15 18.648
R2042 AVDD.n5635 AVDD.t148 18.648
R2043 AVDD.n5635 AVDD.t10 18.648
R2044 AVDD.n1350 AVDD.n1349 17.803
R2045 AVDD.n4404 AVDD.n4401 17.126
R2046 AVDD.t806 AVDD.t760 16.92
R2047 AVDD.n4386 AVDD.n4384 16.92
R2048 AVDD.n4478 AVDD.n4477 16.832
R2049 AVDD.t49 AVDD.n132 16.654
R2050 AVDD.t12 AVDD.n248 16.654
R2051 AVDD.n5740 AVDD.t370 16.595
R2052 AVDD.t5 AVDD.n314 16.595
R2053 AVDD.t15 AVDD.n502 16.595
R2054 AVDD.n4304 AVDD.n4303 15.802
R2055 AVDD.n6389 AVDD.t828 15.794
R2056 AVDD.n6409 AVDD.n6408 15.657
R2057 AVDD.n14 AVDD.t715 15.396
R2058 AVDD.n6398 AVDD.t280 15.212
R2059 AVDD.n6366 AVDD.t728 15.137
R2060 AVDD.t31 AVDD.t812 15.129
R2061 AVDD.n138 AVDD.t49 15.129
R2062 AVDD.n1353 AVDD.n1352 15.072
R2063 AVDD.n17 AVDD.t726 15.063
R2064 AVDD.n6369 AVDD.t100 14.755
R2065 AVDD.n3872 AVDD.t834 14.684
R2066 AVDD.n3939 AVDD.t730 14.684
R2067 AVDD.n3800 AVDD.t191 14.684
R2068 AVDD.n4087 AVDD.t41 14.684
R2069 AVDD.n4154 AVDD.t55 14.684
R2070 AVDD.n4255 AVDD.t807 14.684
R2071 AVDD.n3737 AVDD.t839 14.684
R2072 AVDD.n5832 AVDD.t342 14.684
R2073 AVDD.n6058 AVDD.t96 14.684
R2074 AVDD.n3834 AVDD.t182 14.673
R2075 AVDD.n3857 AVDD.t768 14.673
R2076 AVDD.n3902 AVDD.t145 14.673
R2077 AVDD.n3924 AVDD.t708 14.673
R2078 AVDD.n3968 AVDD.t1 14.673
R2079 AVDD.n3812 AVDD.t764 14.673
R2080 AVDD.n4049 AVDD.t30 14.673
R2081 AVDD.n4072 AVDD.t720 14.673
R2082 AVDD.n4117 AVDD.t216 14.673
R2083 AVDD.n4139 AVDD.t271 14.673
R2084 AVDD.n4239 AVDD.t340 14.673
R2085 AVDD.n4038 AVDD.t750 14.673
R2086 AVDD.n3753 AVDD.t742 14.673
R2087 AVDD.n3778 AVDD.t724 14.673
R2088 AVDD.n6072 AVDD.t267 14.673
R2089 AVDD.n5849 AVDD.t354 14.673
R2090 AVDD.n5885 AVDD.t265 14.673
R2091 AVDD.n5927 AVDD.t819 14.673
R2092 AVDD.n4322 AVDD.t3 14.471
R2093 AVDD.n5254 AVDD.t660 14.438
R2094 AVDD.n5305 AVDD.t501 14.438
R2095 AVDD.n2050 AVDD.t450 14.432
R2096 AVDD.n2058 AVDD.t414 14.432
R2097 AVDD.n5817 AVDD.n5813 14.425
R2098 AVDD.n2465 AVDD.t573 14.27
R2099 AVDD.n2053 AVDD.t618 14.27
R2100 AVDD.n5251 AVDD.t489 14.254
R2101 AVDD.n2470 AVDD.t654 14.254
R2102 AVDD.n5876 AVDD.t287 14.25
R2103 AVDD.n5349 AVDD.t630 14.22
R2104 AVDD.n5408 AVDD.t696 14.201
R2105 AVDD.n5357 AVDD.t663 14.201
R2106 AVDD.n5297 AVDD.t459 14.14
R2107 AVDD.n4027 AVDD.t836 14.084
R2108 AVDD.n4207 AVDD.t835 14.079
R2109 AVDD.n5642 AVDD.n436 14.074
R2110 AVDD.n4389 AVDD.t710 13.849
R2111 AVDD.n4028 AVDD.t762 13.849
R2112 AVDD.n4198 AVDD.t837 13.849
R2113 AVDD.n12 AVDD.t22 13.849
R2114 AVDD.n316 AVDD.t274 13.849
R2115 AVDD.n315 AVDD.t51 13.849
R2116 AVDD.n508 AVDD.t272 13.849
R2117 AVDD.n505 AVDD.t759 13.849
R2118 AVDD.n703 AVDD.t19 13.849
R2119 AVDD.n702 AVDD.t132 13.849
R2120 AVDD.n884 AVDD.t114 13.849
R2121 AVDD.n883 AVDD.t258 13.849
R2122 AVDD.n5610 AVDD.t136 13.849
R2123 AVDD.n5609 AVDD.t251 13.849
R2124 AVDD.n1165 AVDD.t232 13.849
R2125 AVDD.n1164 AVDD.t126 13.849
R2126 AVDD.n5548 AVDD.t101 13.849
R2127 AVDD.n5547 AVDD.t82 13.849
R2128 AVDD.n1652 AVDD.t291 13.849
R2129 AVDD.n1651 AVDD.t231 13.849
R2130 AVDD.n5452 AVDD.t86 13.849
R2131 AVDD.n5451 AVDD.t301 13.849
R2132 AVDD.n5399 AVDD.t67 13.849
R2133 AVDD.n5398 AVDD.t451 13.849
R2134 AVDD.n2056 AVDD.t415 13.849
R2135 AVDD.n4909 AVDD.t769 13.849
R2136 AVDD.n4928 AVDD.t793 13.849
R2137 AVDD.n4929 AVDD.t866 13.849
R2138 AVDD.n5048 AVDD.t803 13.849
R2139 AVDD.n5049 AVDD.t869 13.849
R2140 AVDD.n5099 AVDD.t862 13.849
R2141 AVDD.n5100 AVDD.t776 13.849
R2142 AVDD.n5150 AVDD.t802 13.849
R2143 AVDD.n5151 AVDD.t868 13.849
R2144 AVDD.n2869 AVDD.t774 13.849
R2145 AVDD.n2870 AVDD.t870 13.849
R2146 AVDD.n2668 AVDD.t204 13.849
R2147 AVDD.n2669 AVDD.t273 13.849
R2148 AVDD.n2466 AVDD.t146 13.849
R2149 AVDD.n2467 AVDD.t574 13.849
R2150 AVDD.n2055 AVDD.t619 13.849
R2151 AVDD.n319 AVDD.t755 13.849
R2152 AVDD.n318 AVDD.t13 13.849
R2153 AVDD.n317 AVDD.t823 13.849
R2154 AVDD.n510 AVDD.t756 13.849
R2155 AVDD.n509 AVDD.t150 13.849
R2156 AVDD.n705 AVDD.t824 13.849
R2157 AVDD.n704 AVDD.t322 13.849
R2158 AVDD.n886 AVDD.t289 13.849
R2159 AVDD.n885 AVDD.t225 13.849
R2160 AVDD.n5612 AVDD.t299 13.849
R2161 AVDD.n5611 AVDD.t220 13.849
R2162 AVDD.n5599 AVDD.t230 13.849
R2163 AVDD.n5598 AVDD.t314 13.849
R2164 AVDD.n5558 AVDD.t300 13.849
R2165 AVDD.n5557 AVDD.t108 13.849
R2166 AVDD.n5507 AVDD.t242 13.849
R2167 AVDD.n5506 AVDD.t134 13.849
R2168 AVDD.n5462 AVDD.t116 13.849
R2169 AVDD.n5461 AVDD.t261 13.849
R2170 AVDD.n5411 AVDD.t102 13.849
R2171 AVDD.n5410 AVDD.t697 13.849
R2172 AVDD.n5355 AVDD.t664 13.849
R2173 AVDD.n5354 AVDD.t94 13.849
R2174 AVDD.n5312 AVDD.t92 13.849
R2175 AVDD.n5311 AVDD.t45 13.849
R2176 AVDD.n5261 AVDD.t44 13.849
R2177 AVDD.n5260 AVDD.t871 13.849
R2178 AVDD.n5211 AVDD.t788 13.849
R2179 AVDD.n5210 AVDD.t162 13.849
R2180 AVDD.n5163 AVDD.t845 13.849
R2181 AVDD.n5162 AVDD.t782 13.849
R2182 AVDD.n5112 AVDD.t173 13.849
R2183 AVDD.n5111 AVDD.t329 13.849
R2184 AVDD.n5061 AVDD.t846 13.849
R2185 AVDD.n5060 AVDD.t783 13.849
R2186 AVDD.n4827 AVDD.t331 13.849
R2187 AVDD.n4826 AVDD.t778 13.849
R2188 AVDD.n4599 AVDD.t785 13.849
R2189 AVDD.n3463 AVDD.t841 13.849
R2190 AVDD.n3454 AVDD.t328 13.849
R2191 AVDD.n3455 AVDD.t169 13.849
R2192 AVDD.n5058 AVDD.t336 13.849
R2193 AVDD.n5059 AVDD.t197 13.849
R2194 AVDD.n5109 AVDD.t160 13.849
R2195 AVDD.n5110 AVDD.t856 13.849
R2196 AVDD.n5160 AVDD.t335 13.849
R2197 AVDD.n5161 AVDD.t195 13.849
R2198 AVDD.n5208 AVDD.t848 13.849
R2199 AVDD.n5209 AVDD.t209 13.849
R2200 AVDD.n5207 AVDD.t780 13.849
R2201 AVDD.n5347 AVDD.t240 13.849
R2202 AVDD.n5393 AVDD.t257 13.849
R2203 AVDD.n5394 AVDD.t112 13.849
R2204 AVDD.n5446 AVDD.t131 13.849
R2205 AVDD.n5447 AVDD.t239 13.849
R2206 AVDD.n5497 AVDD.t106 13.849
R2207 AVDD.n5498 AVDD.t217 13.849
R2208 AVDD.n5542 AVDD.t235 13.849
R2209 AVDD.n5543 AVDD.t312 13.849
R2210 AVDD.n5593 AVDD.t243 13.849
R2211 AVDD.n5594 AVDD.t75 13.849
R2212 AVDD.n1062 AVDD.t223 13.849
R2213 AVDD.n1063 AVDD.t308 13.849
R2214 AVDD.n891 AVDD.t320 13.849
R2215 AVDD.n892 AVDD.t73 13.849
R2216 AVDD.n710 AVDD.t303 13.849
R2217 AVDD.n711 AVDD.t121 13.849
R2218 AVDD.n515 AVDD.t65 13.849
R2219 AVDD.n516 AVDD.t736 13.849
R2220 AVDD.n325 AVDD.t752 13.849
R2221 AVDD.n326 AVDD.t805 13.849
R2222 AVDD.n147 AVDD.t735 13.849
R2223 AVDD.n148 AVDD.t50 13.849
R2224 AVDD.n146 AVDD.t278 13.849
R2225 AVDD.n3462 AVDD.t167 13.849
R2226 AVDD.n3452 AVDD.t781 13.849
R2227 AVDD.n3453 AVDD.t338 13.849
R2228 AVDD.n5056 AVDD.t158 13.849
R2229 AVDD.n5057 AVDD.t855 13.849
R2230 AVDD.n5107 AVDD.t334 13.849
R2231 AVDD.n5108 AVDD.t193 13.849
R2232 AVDD.n5158 AVDD.t156 13.849
R2233 AVDD.n5159 AVDD.t853 13.849
R2234 AVDD.n5205 AVDD.t174 13.849
R2235 AVDD.n5206 AVDD.t795 13.849
R2236 AVDD.n5258 AVDD.t327 13.849
R2237 AVDD.n5259 AVDD.t347 13.849
R2238 AVDD.n5309 AVDD.t268 13.849
R2239 AVDD.n5310 AVDD.t110 13.849
R2240 AVDD.n2283 AVDD.t129 13.849
R2241 AVDD.n2284 AVDD.t238 13.849
R2242 AVDD.n5405 AVDD.t256 13.849
R2243 AVDD.n5406 AVDD.t109 13.849
R2244 AVDD.n5459 AVDD.t234 13.849
R2245 AVDD.n5460 AVDD.t119 13.849
R2246 AVDD.n5504 AVDD.t104 13.849
R2247 AVDD.n5505 AVDD.t246 13.849
R2248 AVDD.n5555 AVDD.t117 13.849
R2249 AVDD.n5556 AVDD.t307 13.849
R2250 AVDD.n5600 AVDD.t319 13.849
R2251 AVDD.n5601 AVDD.t71 13.849
R2252 AVDD.n5613 AVDD.t222 13.849
R2253 AVDD.n5614 AVDD.t306 13.849
R2254 AVDD.n887 AVDD.t63 13.849
R2255 AVDD.n888 AVDD.t293 13.849
R2256 AVDD.n706 AVDD.t302 13.849
R2257 AVDD.n707 AVDD.t753 13.849
R2258 AVDD.n511 AVDD.t734 13.849
R2259 AVDD.n512 AVDD.t8 13.849
R2260 AVDD.n320 AVDD.t751 13.849
R2261 AVDD.n321 AVDD.t350 13.849
R2262 AVDD.n322 AVDD.t6 13.849
R2263 AVDD.n3461 AVDD.t850 13.849
R2264 AVDD.n3450 AVDD.t330 13.849
R2265 AVDD.n3451 AVDD.t176 13.849
R2266 AVDD.n5054 AVDD.t844 13.849
R2267 AVDD.n5055 AVDD.t206 13.849
R2268 AVDD.n5105 AVDD.t171 13.849
R2269 AVDD.n5106 AVDD.t792 13.849
R2270 AVDD.n5156 AVDD.t842 13.849
R2271 AVDD.n5157 AVDD.t202 13.849
R2272 AVDD.n5203 AVDD.t857 13.849
R2273 AVDD.n5204 AVDD.t861 13.849
R2274 AVDD.n5255 AVDD.t784 13.849
R2275 AVDD.n5256 AVDD.t661 13.849
R2276 AVDD.n5307 AVDD.t502 13.849
R2277 AVDD.n5308 AVDD.t790 13.849
R2278 AVDD.n2281 AVDD.t840 13.849
R2279 AVDD.n2282 AVDD.t201 13.849
R2280 AVDD.n5403 AVDD.t165 13.849
R2281 AVDD.n5404 AVDD.t244 13.849
R2282 AVDD.n5457 AVDD.t115 13.849
R2283 AVDD.n5458 AVDD.t221 13.849
R2284 AVDD.n5502 AVDD.t241 13.849
R2285 AVDD.n5503 AVDD.t317 13.849
R2286 AVDD.n5553 AVDD.t219 13.849
R2287 AVDD.n5554 AVDD.t84 13.849
R2288 AVDD.n5602 AVDD.t229 13.849
R2289 AVDD.n5603 AVDD.t290 13.849
R2290 AVDD.n5615 AVDD.t325 13.849
R2291 AVDD.n5616 AVDD.t83 13.849
R2292 AVDD.n5622 AVDD.t310 13.849
R2293 AVDD.n5623 AVDD.t124 13.849
R2294 AVDD.n5629 AVDD.t78 13.849
R2295 AVDD.n5630 AVDD.t738 13.849
R2296 AVDD.n5636 AVDD.t754 13.849
R2297 AVDD.n5637 AVDD.t184 13.849
R2298 AVDD.n5643 AVDD.t737 13.849
R2299 AVDD.n5644 AVDD.t17 13.849
R2300 AVDD.n5651 AVDD.t183 13.849
R2301 AVDD.n5652 AVDD.t175 13.849
R2302 AVDD.n5653 AVDD.t843 13.849
R2303 AVDD.n5661 AVDD.t205 13.849
R2304 AVDD.n5660 AVDD.t170 13.849
R2305 AVDD.n5712 AVDD.t791 13.849
R2306 AVDD.n5711 AVDD.t199 13.849
R2307 AVDD.n4604 AVDD.t200 13.849
R2308 AVDD.n3448 AVDD.t164 13.849
R2309 AVDD.n3449 AVDD.t789 13.849
R2310 AVDD.n5052 AVDD.t180 13.849
R2311 AVDD.n5053 AVDD.t800 13.849
R2312 AVDD.n5103 AVDD.t852 13.849
R2313 AVDD.n5104 AVDD.t859 13.849
R2314 AVDD.n5154 AVDD.t178 13.849
R2315 AVDD.n5155 AVDD.t798 13.849
R2316 AVDD.n5201 AVDD.t207 13.849
R2317 AVDD.n5202 AVDD.t770 13.849
R2318 AVDD.n5249 AVDD.t337 13.849
R2319 AVDD.n5252 AVDD.t490 13.849
R2320 AVDD.n5302 AVDD.t655 13.849
R2321 AVDD.n5303 AVDD.t214 13.849
R2322 AVDD.n2279 AVDD.t177 13.849
R2323 AVDD.n2280 AVDD.t797 13.849
R2324 AVDD.n5401 AVDD.t849 13.849
R2325 AVDD.n5402 AVDD.t315 13.849
R2326 AVDD.n5455 AVDD.t245 13.849
R2327 AVDD.n5456 AVDD.t323 13.849
R2328 AVDD.n1655 AVDD.t118 13.849
R2329 AVDD.n1656 AVDD.t226 13.849
R2330 AVDD.n5551 AVDD.t318 13.849
R2331 AVDD.n5552 AVDD.t296 13.849
R2332 AVDD.n5604 AVDD.t305 13.849
R2333 AVDD.n5605 AVDD.t123 13.849
R2334 AVDD.n5617 AVDD.t69 13.849
R2335 AVDD.n5618 AVDD.t295 13.849
R2336 AVDD.n5624 AVDD.t120 13.849
R2337 AVDD.n5625 AVDD.t253 13.849
R2338 AVDD.n5631 AVDD.t292 13.849
R2339 AVDD.n5632 AVDD.t11 13.849
R2340 AVDD.n5638 AVDD.t277 13.849
R2341 AVDD.n5639 AVDD.t349 13.849
R2342 AVDD.n5645 AVDD.t757 13.849
R2343 AVDD.n5646 AVDD.t188 13.849
R2344 AVDD.n5654 AVDD.t348 13.849
R2345 AVDD.n5655 AVDD.t787 13.849
R2346 AVDD.n5656 AVDD.t179 13.849
R2347 AVDD.n5659 AVDD.t799 13.849
R2348 AVDD.n5658 AVDD.t851 13.849
R2349 AVDD.n6309 AVDD.t858 13.849
R2350 AVDD.n6308 AVDD.t794 13.849
R2351 AVDD.n3456 AVDD.t860 13.849
R2352 AVDD.n4904 AVDD.t198 13.849
R2353 AVDD.n4905 AVDD.t801 13.849
R2354 AVDD.n5096 AVDD.t213 13.849
R2355 AVDD.n5097 AVDD.t773 13.849
R2356 AVDD.n5147 AVDD.t796 13.849
R2357 AVDD.n5148 AVDD.t867 13.849
R2358 AVDD.n5198 AVDD.t210 13.849
R2359 AVDD.n5199 AVDD.t772 13.849
R2360 AVDD.n5246 AVDD.t863 13.849
R2361 AVDD.n5247 AVDD.t777 13.849
R2362 AVDD.n5298 AVDD.t854 13.849
R2363 AVDD.n5300 AVDD.t460 13.849
R2364 AVDD.n5351 AVDD.t631 13.849
R2365 AVDD.n5352 AVDD.t298 13.849
R2366 AVDD.n5395 AVDD.t313 13.849
R2367 AVDD.n5396 AVDD.t228 13.849
R2368 AVDD.n5448 AVDD.t218 13.849
R2369 AVDD.n5449 AVDD.t324 13.849
R2370 AVDD.n5499 AVDD.t224 13.849
R2371 AVDD.n5500 AVDD.t309 13.849
R2372 AVDD.n5544 AVDD.t321 13.849
R2373 AVDD.n5545 AVDD.t77 13.849
R2374 AVDD.n5595 AVDD.t304 13.849
R2375 AVDD.n5596 AVDD.t255 13.849
R2376 AVDD.n1060 AVDD.t294 13.849
R2377 AVDD.n1061 AVDD.t128 13.849
R2378 AVDD.n889 AVDD.t122 13.849
R2379 AVDD.n890 AVDD.t254 13.849
R2380 AVDD.n708 AVDD.t127 13.849
R2381 AVDD.n709 AVDD.t233 13.849
R2382 AVDD.n513 AVDD.t252 13.849
R2383 AVDD.n514 AVDD.t758 13.849
R2384 AVDD.n323 AVDD.t269 13.849
R2385 AVDD.n324 AVDD.t187 13.849
R2386 AVDD.n143 AVDD.t346 13.849
R2387 AVDD.n144 AVDD.t189 13.849
R2388 AVDD.n145 AVDD.t186 13.849
R2389 AVDD.n5647 AVDD.t733 13.849
R2390 AVDD.n5649 AVDD.t822 13.849
R2391 AVDD.n5648 AVDD.t16 13.849
R2392 AVDD.n5641 AVDD.t345 13.849
R2393 AVDD.n5640 AVDD.t149 13.849
R2394 AVDD.n5634 AVDD.t18 13.849
R2395 AVDD.n5633 AVDD.t79 13.849
R2396 AVDD.n5627 AVDD.t297 13.849
R2397 AVDD.n5626 AVDD.t259 13.849
R2398 AVDD.n5620 AVDD.t80 13.849
R2399 AVDD.n5619 AVDD.t107 13.849
R2400 AVDD.n5607 AVDD.t260 13.849
R2401 AVDD.n5606 AVDD.t227 13.849
R2402 AVDD.n5550 AVDD.t316 13.849
R2403 AVDD.n5549 AVDD.t133 13.849
R2404 AVDD.n1654 AVDD.t311 13.849
R2405 AVDD.n1653 AVDD.t236 13.849
R2406 AVDD.n5454 AVDD.t135 13.849
R2407 AVDD.n5453 AVDD.t326 13.849
R2408 AVDD.n5400 AVDD.t237 13.849
R2409 AVDD.n2672 AVDD.t151 13.849
R2410 AVDD.n2671 AVDD.t139 13.849
R2411 AVDD.n2670 AVDD.t771 13.849
R2412 AVDD.n2872 AVDD.t786 13.849
R2413 AVDD.n2871 AVDD.t864 13.849
R2414 AVDD.n5153 AVDD.t847 13.849
R2415 AVDD.n5152 AVDD.t775 13.849
R2416 AVDD.n5102 AVDD.t865 13.849
R2417 AVDD.n5101 AVDD.t332 13.849
R2418 AVDD.n5051 AVDD.t779 13.849
R2419 AVDD.n5050 AVDD.t211 13.849
R2420 AVDD.n3447 AVDD.t333 13.849
R2421 AVDD.n3446 AVDD.t804 13.849
R2422 AVDD.n4692 AVDD.t212 13.849
R2423 AVDD.n4215 AVDD.t761 13.848
R2424 AVDD.n3498 AVDD.t679 13.848
R2425 AVDD.n3498 AVDD.t463 13.848
R2426 AVDD.n4481 AVDD.t678 13.848
R2427 AVDD.n4481 AVDD.t462 13.848
R2428 AVDD.n4496 AVDD.t484 13.848
R2429 AVDD.n4493 AVDD.t483 13.848
R2430 AVDD.n4493 AVDD.t570 13.848
R2431 AVDD.n4496 AVDD.t571 13.848
R2432 AVDD.n4906 AVDD.t383 13.848
R2433 AVDD.n3483 AVDD.t382 13.848
R2434 AVDD.n3479 AVDD.t646 13.848
R2435 AVDD.n3487 AVDD.t645 13.848
R2436 AVDD.n3487 AVDD.t513 13.848
R2437 AVDD.n3479 AVDD.t514 13.848
R2438 AVDD.n3483 AVDD.t519 13.848
R2439 AVDD.n4906 AVDD.t520 13.848
R2440 AVDD.n5773 AVDD.t582 13.848
R2441 AVDD.n5773 AVDD.t540 13.848
R2442 AVDD.n6293 AVDD.t541 13.848
R2443 AVDD.n6293 AVDD.t583 13.848
R2444 AVDD.n5754 AVDD.t371 13.848
R2445 AVDD.n5754 AVDD.t675 13.848
R2446 AVDD.n5771 AVDD.t372 13.848
R2447 AVDD.n5771 AVDD.t676 13.848
R2448 AVDD.n5788 AVDD.t706 13.848
R2449 AVDD.n5788 AVDD.t412 13.848
R2450 AVDD.n5796 AVDD.t705 13.848
R2451 AVDD.n5796 AVDD.t411 13.848
R2452 AVDD.n5790 AVDD.t438 13.848
R2453 AVDD.n5790 AVDD.t402 13.848
R2454 AVDD.n6297 AVDD.t439 13.848
R2455 AVDD.n6297 AVDD.t403 13.848
R2456 AVDD.n5714 AVDD.t433 13.848
R2457 AVDD.n6147 AVDD.t474 13.848
R2458 AVDD.n6147 AVDD.t432 13.848
R2459 AVDD.n5714 AVDD.t475 13.848
R2460 AVDD.n6146 AVDD.t544 13.848
R2461 AVDD.n6146 AVDD.t589 13.848
R2462 AVDD.n6153 AVDD.t543 13.848
R2463 AVDD.n6153 AVDD.t588 13.848
R2464 AVDD.n5698 AVDD.t616 13.848
R2465 AVDD.n6191 AVDD.t648 13.848
R2466 AVDD.n6191 AVDD.t615 13.848
R2467 AVDD.n5698 AVDD.t649 13.848
R2468 AVDD.n6190 AVDD.t409 13.848
R2469 AVDD.n6190 AVDD.t445 13.848
R2470 AVDD.n6197 AVDD.t408 13.848
R2471 AVDD.n6197 AVDD.t444 13.848
R2472 AVDD.n6212 AVDD.t580 13.848
R2473 AVDD.n6212 AVDD.t622 13.848
R2474 AVDD.n6220 AVDD.t579 13.848
R2475 AVDD.n6220 AVDD.t621 13.848
R2476 AVDD.n6214 AVDD.t495 13.848
R2477 AVDD.n6214 AVDD.t471 13.848
R2478 AVDD.n5719 AVDD.t496 13.848
R2479 AVDD.n5719 AVDD.t472 13.848
R2480 AVDD.n6235 AVDD.t424 13.848
R2481 AVDD.n6235 AVDD.t457 13.848
R2482 AVDD.n6243 AVDD.t423 13.848
R2483 AVDD.n6243 AVDD.t456 13.848
R2484 AVDD.n6237 AVDD.t657 13.848
R2485 AVDD.n6237 AVDD.t627 13.848
R2486 AVDD.n5727 AVDD.t658 13.848
R2487 AVDD.n5727 AVDD.t628 13.848
R2488 AVDD.n3465 AVDD.t442 13.848
R2489 AVDD.n3465 AVDD.t643 13.848
R2490 AVDD.n4551 AVDD.t441 13.848
R2491 AVDD.n4551 AVDD.t642 13.848
R2492 AVDD.n4553 AVDD.t553 13.848
R2493 AVDD.n4553 AVDD.t436 13.848
R2494 AVDD.n4547 AVDD.t552 13.848
R2495 AVDD.n4547 AVDD.t435 13.848
R2496 AVDD.n4514 AVDD.t586 13.848
R2497 AVDD.n4514 AVDD.t466 13.848
R2498 AVDD.n4523 AVDD.t585 13.848
R2499 AVDD.n4523 AVDD.t465 13.848
R2500 AVDD.n4525 AVDD.t376 13.848
R2501 AVDD.n4525 AVDD.t577 13.848
R2502 AVDD.n4519 AVDD.t375 13.848
R2503 AVDD.n4519 AVDD.t576 13.848
R2504 AVDD.n4438 AVDD.t427 13.848
R2505 AVDD.n4438 AVDD.t625 13.848
R2506 AVDD.n4447 AVDD.t426 13.848
R2507 AVDD.n4447 AVDD.t624 13.848
R2508 AVDD.n4449 AVDD.t535 13.848
R2509 AVDD.n4449 AVDD.t421 13.848
R2510 AVDD.n4443 AVDD.t534 13.848
R2511 AVDD.n4443 AVDD.t420 13.848
R2512 AVDD.n3458 AVDD.t565 13.848
R2513 AVDD.n3458 AVDD.t448 13.848
R2514 AVDD.n4419 AVDD.t564 13.848
R2515 AVDD.n4419 AVDD.t447 13.848
R2516 AVDD.n4421 AVDD.t700 13.848
R2517 AVDD.n4421 AVDD.t559 13.848
R2518 AVDD.n4415 AVDD.t699 13.848
R2519 AVDD.n4415 AVDD.t558 13.848
R2520 AVDD.n3712 AVDD.t391 13.848
R2521 AVDD.n3712 AVDD.t594 13.848
R2522 AVDD.n3714 AVDD.t526 13.848
R2523 AVDD.n3714 AVDD.t386 13.848
R2524 AVDD.n3708 AVDD.t525 13.848
R2525 AVDD.n3708 AVDD.t385 13.848
R2526 AVDD.n4601 AVDD.t595 13.848
R2527 AVDD.n4601 AVDD.t392 13.848
R2528 AVDD.n3493 AVDD.t556 13.848
R2529 AVDD.n3493 AVDD.t694 13.848
R2530 AVDD.n3544 AVDD.t667 13.848
R2531 AVDD.n3544 AVDD.t532 13.848
R2532 AVDD.n3539 AVDD.t666 13.848
R2533 AVDD.n3539 AVDD.t531 13.848
R2534 AVDD.n3542 AVDD.t693 13.848
R2535 AVDD.n3542 AVDD.t555 13.848
R2536 AVDD.n6258 AVDD.t604 13.848
R2537 AVDD.n6258 AVDD.t637 13.848
R2538 AVDD.n6266 AVDD.t603 13.848
R2539 AVDD.n6266 AVDD.t636 13.848
R2540 AVDD.n6260 AVDD.t507 13.848
R2541 AVDD.n6260 AVDD.t480 13.848
R2542 AVDD.n5735 AVDD.t508 13.848
R2543 AVDD.n5735 AVDD.t481 13.848
R2544 AVDD.n6281 AVDD.t538 13.848
R2545 AVDD.n6281 AVDD.t691 13.848
R2546 AVDD.n6289 AVDD.t537 13.848
R2547 AVDD.n6289 AVDD.t690 13.848
R2548 AVDD.n6283 AVDD.t561 13.848
R2549 AVDD.n6283 AVDD.t429 13.848
R2550 AVDD.n5745 AVDD.t562 13.848
R2551 AVDD.n5745 AVDD.t430 13.848
R2552 AVDD.n6371 AVDD.t88 13.847
R2553 AVDD.n6371 AVDD.t98 13.847
R2554 AVDD.n6381 AVDD.t352 13.847
R2555 AVDD.n6381 AVDD.t60 13.847
R2556 AVDD.n6380 AVDD.t356 13.847
R2557 AVDD.n6380 AVDD.t809 13.847
R2558 AVDD.n6379 AVDD.t811 13.847
R2559 AVDD.n6379 AVDD.t813 13.847
R2560 AVDD.n6388 AVDD.t282 13.847
R2561 AVDD.n6388 AVDD.t360 13.847
R2562 AVDD.n6387 AVDD.t364 13.847
R2563 AVDD.n6387 AVDD.t826 13.847
R2564 AVDD.n6386 AVDD.t832 13.847
R2565 AVDD.n6386 AVDD.t286 13.847
R2566 AVDD.n6385 AVDD.t817 13.847
R2567 AVDD.n6385 AVDD.t284 13.847
R2568 AVDD.n6384 AVDD.t358 13.847
R2569 AVDD.n6384 AVDD.t362 13.847
R2570 AVDD.n6383 AVDD.t288 13.847
R2571 AVDD.n6383 AVDD.t821 13.847
R2572 AVDD.n6382 AVDD.t830 13.847
R2573 AVDD.n6382 AVDD.t815 13.847
R2574 AVDD.t185 AVDD.t4 13.62
R2575 AVDD.n5876 AVDD.t820 13.546
R2576 AVDD.n4409 AVDD.n4404 12.999
R2577 AVDD.t31 AVDD.t810 12.666
R2578 AVDD.n4310 AVDD.t27 12.343
R2579 AVDD.n5817 AVDD.n5816 12.314
R2580 AVDD.n5628 AVDD.t64 12.28
R2581 AVDD.n5628 AVDD.t113 12.28
R2582 AVDD.n5621 AVDD.t72 12.28
R2583 AVDD.n5608 AVDD.t68 12.28
R2584 AVDD.n5608 AVDD.t70 12.28
R2585 AVDD.n5450 AVDD.t105 12.28
R2586 AVDD.n5397 AVDD.t111 12.28
R2587 AVDD.n5353 AVDD.t93 12.28
R2588 AVDD.n5301 AVDD.t43 12.28
R2589 AVDD.n5248 AVDD.t203 12.28
R2590 AVDD.n5200 AVDD.t194 12.28
R2591 AVDD.n5149 AVDD.t155 12.28
R2592 AVDD.n5098 AVDD.t196 12.28
R2593 AVDD.n5047 AVDD.t168 12.28
R2594 AVDD.n4597 AVDD.t374 12.28
R2595 AVDD.t339 AVDD.n4228 12.174
R2596 AVDD.t806 AVDD.n4248 12.174
R2597 AVDD.n4483 AVDD.t461 12.05
R2598 AVDD.n4562 AVDD.t440 12.05
R2599 AVDD.n4566 AVDD.t584 12.05
R2600 AVDD.n4472 AVDD.t425 12.05
R2601 AVDD.n4466 AVDD.t563 12.05
R2602 AVDD.n4462 AVDD.t390 12.05
R2603 AVDD.n4570 AVDD.t692 12.05
R2604 AVDD.n4573 AVDD.t518 12.05
R2605 AVDD.n3980 AVDD.n3979 11.67
R2606 AVDD.n3810 AVDD.n3809 11.67
R2607 AVDD.n3847 AVDD.n3846 11.67
R2608 AVDD.n3861 AVDD.n3860 11.67
R2609 AVDD.n3914 AVDD.n3913 11.67
R2610 AVDD.n3928 AVDD.n3927 11.67
R2611 AVDD.n4062 AVDD.n4061 11.67
R2612 AVDD.n4076 AVDD.n4075 11.67
R2613 AVDD.n4129 AVDD.n4128 11.67
R2614 AVDD.n4241 AVDD.n4240 11.67
R2615 AVDD.n4192 AVDD.n4191 11.67
R2616 AVDD.n4143 AVDD.n4142 11.67
R2617 AVDD.n3768 AVDD.n3767 11.67
R2618 AVDD.n3748 AVDD.n3747 11.67
R2619 AVDD.n5847 AVDD.n5846 11.67
R2620 AVDD.n6081 AVDD.n6080 11.67
R2621 AVDD.n5909 AVDD.n5908 11.67
R2622 AVDD.n5929 AVDD.n5928 11.67
R2623 AVDD.n4412 AVDD.n4411 11.66
R2624 AVDD.n6315 AVDD.n6312 11.259
R2625 AVDD.n6411 AVDD.n6410 11.259
R2626 AVDD.t818 AVDD.n5917 11.083
R2627 AVDD.t113 AVDD.n811 10.967
R2628 AVDD.t72 AVDD.n992 10.967
R2629 AVDD.n4924 AVDD.t166 10.967
R2630 AVDD.t64 AVDD.n882 10.928
R2631 AVDD.t62 AVDD.n1058 10.928
R2632 AVDD.t68 AVDD.n1163 10.928
R2633 AVDD.n4822 AVDD.t163 10.928
R2634 AVDD.n4185 AVDD.n4182 10.729
R2635 AVDD.n3994 AVDD.n3993 10.215
R2636 AVDD.n1059 AVDD.t62 10.156
R2637 AVDD.n6557 AVDD.n6556 10.154
R2638 AVDD.n5812 AVDD.n5811 10.067
R2639 AVDD.n5857 AVDD.n5856 10.067
R2640 AVDD.n10 AVDD.n9 10.067
R2641 AVDD.n3782 AVDD.n3781 10.063
R2642 AVDD.n3877 AVDD.n3876 10.063
R2643 AVDD.n3944 AVDD.n3943 10.063
R2644 AVDD.n4092 AVDD.n4091 10.063
R2645 AVDD.n4034 AVDD.n4033 10.063
R2646 AVDD.n4159 AVDD.n4158 10.063
R2647 AVDD.t185 AVDD.n4386 9.904
R2648 AVDD.t10 AVDD.n630 9.632
R2649 AVDD.t264 AVDD.n5890 9.5
R2650 AVDD.n6405 AVDD.n6403 9.5
R2651 AVDD.n4407 AVDD.n4406 9.353
R2652 AVDD.n17 AVDD.n16 9.314
R2653 AVDD.n3790 AVDD.n3789 9.3
R2654 AVDD.n3885 AVDD.n3884 9.3
R2655 AVDD.n3955 AVDD.n3954 9.3
R2656 AVDD.n4100 AVDD.n4099 9.3
R2657 AVDD.n4397 AVDD.n4396 9.3
R2658 AVDD.n4170 AVDD.n4169 9.3
R2659 AVDD.n6368 AVDD.n6367 9.3
R2660 AVDD.n5823 AVDD.n5822 9.3
R2661 AVDD.n5882 AVDD.n5881 9.3
R2662 AVDD.n6417 AVDD.n6416 9.3
R2663 AVDD.t281 AVDD.t827 9.265
R2664 AVDD.t816 AVDD.t285 9.265
R2665 AVDD.t351 AVDD.t59 9.265
R2666 AVDD.n142 AVDD.n141 9.188
R2667 AVDD.t264 AVDD.t351 9.148
R2668 AVDD.n6303 AVDD.n5758 9.03
R2669 AVDD.t361 AVDD.t344 8.972
R2670 AVDD.n4406 AVDD.n4405 8.892
R2671 AVDD.n1648 AVDD.t81 8.804
R2672 AVDD.t140 AVDD.n433 8.737
R2673 AVDD.t2 AVDD.t159 8.727
R2674 AVDD.n4494 AVDD.t343 8.691
R2675 AVDD.t279 AVDD.t147 8.503
R2676 AVDD.t148 AVDD.n701 8.327
R2677 AVDD.n701 AVDD.n698 8.268
R2678 AVDD.n4494 AVDD.t26 8.267
R2679 AVDD.n1558 AVDD.t76 8.186
R2680 AVDD.t24 AVDD.t66 8.109
R2681 AVDD.n4026 AVDD.n4021 7.977
R2682 AVDD.t7 AVDD.t140 7.916
R2683 AVDD.n3687 AVDD.n3686 7.854
R2684 AVDD.n4414 AVDD 7.615
R2685 AVDD.t357 AVDD.t21 7.564
R2686 AVDD.n4375 AVDD.n4374 7.466
R2687 AVDD.n4298 AVDD.n4297 7.466
R2688 AVDD.n1766 AVDD.t85 7.414
R2689 AVDD.t394 AVDD.t74 7.337
R2690 AVDD.t168 AVDD.t47 7.337
R2691 AVDD.n28 AVDD.n27 7.33
R2692 AVDD.n562 AVDD.n561 7.196
R2693 AVDD.n5896 AVDD.n5895 7.168
R2694 AVDD.n140 AVDD.t714 7.154
R2695 AVDD.n4316 AVDD.n4315 7.001
R2696 AVDD.n6138 AVDD.t825 6.978
R2697 AVDD.n314 AVDD.n297 6.978
R2698 AVDD.n502 AVDD.n485 6.978
R2699 AVDD.n4359 AVDD.t713 6.923
R2700 AVDD.n504 AVDD.t250 6.923
R2701 AVDD.n504 AVDD.t744 6.923
R2702 AVDD.n503 AVDD.t141 6.923
R2703 AVDD.n503 AVDD.t248 6.923
R2704 AVDD.n6490 AVDD.n6441 6.919
R2705 AVDD.n132 AVDD.n123 6.919
R2706 AVDD.n248 AVDD.n239 6.919
R2707 AVDD.n4628 AVDD.n4627 6.879
R2708 AVDD.n4647 AVDD.n4646 6.879
R2709 AVDD.n4642 AVDD.n4640 6.879
R2710 AVDD.n4642 AVDD.n4641 6.879
R2711 AVDD.n4636 AVDD.n4634 6.879
R2712 AVDD.n4636 AVDD.n4635 6.879
R2713 AVDD.n4651 AVDD.n4649 6.879
R2714 AVDD.n4651 AVDD.n4650 6.879
R2715 AVDD.n4625 AVDD.n4624 6.879
R2716 AVDD.n1467 AVDD.t125 6.796
R2717 AVDD.n5038 AVDD.t157 6.796
R2718 AVDD.n4027 AVDD.n3998 6.736
R2719 AVDD.n569 AVDD.n568 6.724
R2720 AVDD.t34 AVDD.t103 6.719
R2721 AVDD.t366 AVDD.t381 6.719
R2722 AVDD.n4829 AVDD.n4828 6.546
R2723 AVDD.n4868 AVDD.n4867 6.546
R2724 AVDD.n369 AVDD.n368 6.4
R2725 AVDD.n2645 AVDD.n2644 6.318
R2726 AVDD.n687 AVDD.n686 6.298
R2727 AVDD.n369 AVDD.n367 6.291
R2728 AVDD.n4479 AVDD.n4478 6.272
R2729 AVDD.n4807 AVDD.n4758 6.178
R2730 AVDD.n4368 AVDD.n4367 6.164
R2731 AVDD.t285 AVDD.n6321 6.157
R2732 AVDD.n5356 AVDD.t662 6.033
R2733 AVDD.n5304 AVDD.t500 6.032
R2734 AVDD.n2057 AVDD.t413 6.029
R2735 AVDD.n5407 AVDD.t695 6.029
R2736 AVDD.n5348 AVDD.t629 6.028
R2737 AVDD.n5253 AVDD.t659 6.027
R2738 AVDD.n2051 AVDD.t572 6.027
R2739 AVDD.n2052 AVDD.t617 6.027
R2740 AVDD.n6124 AVDD.t539 6.026
R2741 AVDD.n6164 AVDD.t400 6.026
R2742 AVDD.n6096 AVDD.t470 6.026
R2743 AVDD.n6100 AVDD.t626 6.026
R2744 AVDD.n6177 AVDD.t479 6.026
R2745 AVDD.n6181 AVDD.t428 6.026
R2746 AVDD.n4461 AVDD.t593 6.026
R2747 AVDD.n4465 AVDD.t446 6.026
R2748 AVDD.n4471 AVDD.t623 6.026
R2749 AVDD.n4565 AVDD.t464 6.026
R2750 AVDD.n4561 AVDD.t641 6.026
R2751 AVDD.n4483 AVDD.t677 6.025
R2752 AVDD.n4575 AVDD.t380 6.025
R2753 AVDD.n6125 AVDD.t581 6.025
R2754 AVDD.n6165 AVDD.t437 6.025
R2755 AVDD.n6131 AVDD.t431 6.025
R2756 AVDD.n6172 AVDD.t614 6.025
R2757 AVDD.n6097 AVDD.t494 6.025
R2758 AVDD.n6101 AVDD.t656 6.025
R2759 AVDD.n4570 AVDD.t554 6.025
R2760 AVDD.n6178 AVDD.t506 6.025
R2761 AVDD.n6182 AVDD.t560 6.025
R2762 AVDD.n2469 AVDD.t653 6.025
R2763 AVDD.n5250 AVDD.t488 6.025
R2764 AVDD.n2049 AVDD.t449 6.025
R2765 AVDD.n6130 AVDD.t473 6.023
R2766 AVDD.n6171 AVDD.t647 6.023
R2767 AVDD.n5296 AVDD.t458 6.02
R2768 AVDD.t275 AVDD.t357 5.981
R2769 AVDD.t95 AVDD.t829 5.981
R2770 AVDD.t829 AVDD.n6051 5.922
R2771 AVDD.t341 AVDD.n5837 5.805
R2772 AVDD.t760 AVDD.n4245 5.571
R2773 AVDD.n4367 AVDD.n4366 5.567
R2774 AVDD.n4313 AVDD.t28 5.533
R2775 AVDD.t35 AVDD.t353 5.453
R2776 AVDD.n28 AVDD.n25 5.453
R2777 AVDD.n6405 AVDD.n6404 5.101
R2778 AVDD.n1465 AVDD.n1463 4.896
R2779 AVDD.n560 AVDD.t90 4.85
R2780 AVDD.n1269 AVDD.t138 4.85
R2781 AVDD.n1273 AVDD.t137 4.828
R2782 AVDD.n567 AVDD.t89 4.828
R2783 AVDD.t827 AVDD.n5702 4.75
R2784 AVDD.n5917 AVDD.t279 4.75
R2785 AVDD.n3648 AVDD.n3647 4.736
R2786 AVDD.t709 AVDD.t716 4.681
R2787 AVDD.n1460 AVDD.n1458 4.673
R2788 AVDD.n1456 AVDD.n1454 4.673
R2789 AVDD.n1451 AVDD.n1449 4.673
R2790 AVDD.n1446 AVDD.n1444 4.673
R2791 AVDD.n1441 AVDD.n1439 4.673
R2792 AVDD.n1436 AVDD.n1434 4.673
R2793 AVDD.n1432 AVDD.n1430 4.673
R2794 AVDD.n1426 AVDD.n1424 4.673
R2795 AVDD.n6324 AVDD.t816 4.632
R2796 AVDD.n6362 AVDD.t725 4.632
R2797 AVDD.t808 AVDD.n6422 4.632
R2798 AVDD.n6376 AVDD.t87 4.632
R2799 AVDD.t247 AVDD.n424 4.632
R2800 AVDD.n3639 AVDD.n3638 4.628
R2801 AVDD.n3574 AVDD.n3573 4.628
R2802 AVDD.n3642 AVDD.n3641 4.628
R2803 AVDD.n3571 AVDD.n3570 4.628
R2804 AVDD.n3645 AVDD.n3644 4.628
R2805 AVDD.n3568 AVDD.n3567 4.628
R2806 AVDD.n1058 AVDD.n1041 4.595
R2807 AVDD.n1163 AVDD.n1146 4.595
R2808 AVDD.n1421 AVDD.n1406 4.595
R2809 AVDD.n1625 AVDD.n1610 4.595
R2810 AVDD.n1834 AVDD.n1819 4.595
R2811 AVDD.n2046 AVDD.n2031 4.595
R2812 AVDD.n2125 AVDD.n2110 4.595
R2813 AVDD.n2461 AVDD.n2446 4.595
R2814 AVDD.n2625 AVDD.n2610 4.595
R2815 AVDD.n3005 AVDD.n2990 4.595
R2816 AVDD.n3404 AVDD.n3389 4.595
R2817 AVDD.n4822 AVDD.n4807 4.595
R2818 AVDD.n436 AVDD.t7 4.574
R2819 AVDD.n5898 AVDD.n5897 4.571
R2820 AVDD.n630 AVDD.n621 4.556
R2821 AVDD.n811 AVDD.n802 4.556
R2822 AVDD.n992 AVDD.n983 4.556
R2823 AVDD.n1344 AVDD.n1295 4.556
R2824 AVDD.n1406 AVDD.n1356 4.556
R2825 AVDD.n1260 AVDD.n1251 4.556
R2826 AVDD.n1535 AVDD.n1526 4.556
R2827 AVDD.n1977 AVDD.n1968 4.556
R2828 AVDD.n2349 AVDD.n2340 4.556
R2829 AVDD.n2774 AVDD.n2765 4.556
R2830 AVDD.n2937 AVDD.n2928 4.556
R2831 AVDD.n3118 AVDD.n3109 4.556
R2832 AVDD.n3337 AVDD.n3328 4.556
R2833 AVDD.n4758 AVDD.n4709 4.556
R2834 AVDD.n3650 AVDD.n3637 4.556
R2835 AVDD.n4207 AVDD.n4201 4.539
R2836 AVDD.n5704 AVDD.t281 4.515
R2837 AVDD.t359 AVDD.t35 4.398
R2838 AVDD.n6403 AVDD.t355 4.398
R2839 AVDD.n6002 AVDD.t814 4.354
R2840 AVDD.t709 AVDD.t185 4.333
R2841 AVDD.n6430 AVDD.n6429 4.275
R2842 AVDD.n4388 AVDD.n4324 4.237
R2843 AVDD.n6376 AVDD.t9 4.222
R2844 AVDD.n698 AVDD.t743 4.222
R2845 AVDD.n3705 AVDD.t366 4.209
R2846 AVDD.n3594 AVDD.n3591 4.151
R2847 AVDD.n3602 AVDD.n3599 4.151
R2848 AVDD.n3610 AVDD.n3607 4.151
R2849 AVDD.n3618 AVDD.n3615 4.151
R2850 AVDD.n3626 AVDD.n3623 4.151
R2851 AVDD.n3634 AVDD.n3631 4.151
R2852 AVDD.n3586 AVDD.n3583 4.093
R2853 AVDD.n1269 AVDD.n1268 3.981
R2854 AVDD.n882 AVDD.n865 3.977
R2855 AVDD.n6117 AVDD.t831 3.959
R2856 AVDD.n1351 AVDD.n1350 3.956
R2857 AVDD.n4027 AVDD.t717 3.83
R2858 AVDD.t812 AVDD.t99 3.753
R2859 AVDD.n5900 AVDD.n5896 3.696
R2860 AVDD.t814 AVDD.n5935 3.694
R2861 AVDD.n28 AVDD.n20 3.694
R2862 AVDD.n5657 AVDD.n142 3.669
R2863 AVDD.t820 AVDD.n5875 3.577
R2864 AVDD.n3669 AVDD.n3650 3.552
R2865 AVDD.n6321 AVDD.n6318 3.518
R2866 AVDD.n5657 AVDD.n138 3.518
R2867 AVDD.n4825 AVDD.n4658 3.475
R2868 AVDD.n3564 AVDD.t549 3.47
R2869 AVDD.n3672 AVDD.t550 3.47
R2870 AVDD.n3677 AVDD.t702 3.47
R2871 AVDD.n3677 AVDD.t703 3.47
R2872 AVDD.n3699 AVDD.t651 3.47
R2873 AVDD.n3699 AVDD.t652 3.47
R2874 AVDD.n3702 AVDD.t504 3.47
R2875 AVDD.n3702 AVDD.t505 3.47
R2876 AVDD.n3445 AVDD.t398 3.47
R2877 AVDD.n3445 AVDD.t399 3.47
R2878 AVDD.n3254 AVDD.t612 3.47
R2879 AVDD.n3254 AVDD.t613 3.47
R2880 AVDD.n2778 AVDD.t672 3.47
R2881 AVDD.n2778 AVDD.t673 3.47
R2882 AVDD.n2667 AVDD.t606 3.47
R2883 AVDD.n2667 AVDD.t607 3.47
R2884 AVDD.n2261 AVDD.t492 3.47
R2885 AVDD.n2261 AVDD.t493 3.47
R2886 AVDD.n1981 AVDD.t687 3.47
R2887 AVDD.n1981 AVDD.t688 3.47
R2888 AVDD.n1875 AVDD.t567 3.47
R2889 AVDD.n1875 AVDD.t568 3.47
R2890 AVDD.n1264 AVDD.t453 3.47
R2891 AVDD.n1264 AVDD.t454 3.47
R2892 AVDD.n4828 AVDD.t522 3.47
R2893 AVDD.n4867 AVDD.t523 3.47
R2894 AVDD.n1175 AVDD.t547 3.47
R2895 AVDD.n1175 AVDD.t546 3.47
R2896 AVDD.n1853 AVDD.t681 3.47
R2897 AVDD.n1853 AVDD.t682 3.47
R2898 AVDD.n2189 AVDD.t598 3.47
R2899 AVDD.n2189 AVDD.t597 3.47
R2900 AVDD.n2645 AVDD.t378 3.47
R2901 AVDD.n2645 AVDD.t379 3.47
R2902 AVDD.n2689 AVDD.t469 3.47
R2903 AVDD.n2689 AVDD.t468 3.47
R2904 AVDD.n3232 AVDD.t388 3.47
R2905 AVDD.n3232 AVDD.t389 3.47
R2906 AVDD.n1894 AVDD.t486 3.47
R2907 AVDD.n1894 AVDD.t487 3.47
R2908 AVDD.n3423 AVDD.t510 3.47
R2909 AVDD.n3423 AVDD.t511 3.47
R2910 AVDD.n4847 AVDD.t633 3.47
R2911 AVDD.n4847 AVDD.t634 3.47
R2912 AVDD.n3687 AVDD.t670 3.47
R2913 AVDD.n3687 AVDD.t669 3.47
R2914 AVDD.n3690 AVDD.t516 3.47
R2915 AVDD.n3690 AVDD.t517 3.47
R2916 AVDD.n3683 AVDD.t367 3.47
R2917 AVDD.n3683 AVDD.t368 3.47
R2918 AVDD.n3693 AVDD.t417 3.47
R2919 AVDD.n3693 AVDD.t418 3.47
R2920 AVDD.n3680 AVDD.t609 3.47
R2921 AVDD.n3680 AVDD.t610 3.47
R2922 AVDD.n3696 AVDD.t477 3.47
R2923 AVDD.n3696 AVDD.t478 3.47
R2924 AVDD.n1177 AVDD.t405 3.47
R2925 AVDD.n1177 AVDD.t406 3.47
R2926 AVDD.n1179 AVDD.t600 3.47
R2927 AVDD.n1179 AVDD.t601 3.47
R2928 AVDD.n1181 AVDD.t639 3.47
R2929 AVDD.n1181 AVDD.t640 3.47
R2930 AVDD.n1183 AVDD.t498 3.47
R2931 AVDD.n1183 AVDD.t499 3.47
R2932 AVDD.n1185 AVDD.t684 3.47
R2933 AVDD.n1185 AVDD.t685 3.47
R2934 AVDD.n1187 AVDD.t528 3.47
R2935 AVDD.n1187 AVDD.t529 3.47
R2936 AVDD.n1190 AVDD.t395 3.47
R2937 AVDD.n1190 AVDD.t396 3.47
R2938 AVDD.n1192 AVDD.t591 3.47
R2939 AVDD.n1192 AVDD.t592 3.47
R2940 AVDD.n4631 AVDD.n4630 3.349
R2941 AVDD.n6410 AVDD.n6409 3.166
R2942 AVDD.n5397 AVDD.n2278 3.025
R2943 AVDD.n5098 AVDD.n3339 3.025
R2944 AVDD.n5450 AVDD.n2048 3.02
R2945 AVDD.n5149 AVDD.n3271 3.02
R2946 AVDD.t825 AVDD.n6117 2.991
R2947 AVDD.n2464 AVDD.n2463 2.887
R2948 AVDD.n5301 AVDD.n2560 2.882
R2949 AVDD.t827 AVDD.t401 2.873
R2950 AVDD.n421 AVDD.t249 2.873
R2951 AVDD.n4656 AVDD.n4655 2.826
R2952 AVDD.n6358 AVDD.n6324 2.814
R2953 AVDD.n2940 AVDD.n2939 2.811
R2954 AVDD.n1465 AVDD.n1464 2.803
R2955 AVDD.n1630 AVDD.n1629 2.803
R2956 AVDD.n1540 AVDD.n1539 2.803
R2957 AVDD.n1748 AVDD.n1747 2.803
R2958 AVDD.n1709 AVDD.n1708 2.803
R2959 AVDD.n2129 AVDD.n2128 2.803
R2960 AVDD.n2151 AVDD.n2150 2.803
R2961 AVDD.n2376 AVDD.n2375 2.803
R2962 AVDD.n2354 AVDD.n2353 2.803
R2963 AVDD.n2522 AVDD.n2521 2.803
R2964 AVDD.n2830 AVDD.n2829 2.803
R2965 AVDD.n3010 AVDD.n3009 2.803
R2966 AVDD.n3032 AVDD.n3031 2.803
R2967 AVDD.n3144 AVDD.n3143 2.803
R2968 AVDD.n3122 AVDD.n3121 2.803
R2969 AVDD.n4981 AVDD.n4980 2.803
R2970 AVDD.n5020 AVDD.n5019 2.803
R2971 AVDD.n4606 AVDD.n4605 2.803
R2972 AVDD.n4632 AVDD.n4631 2.803
R2973 AVDD.n5248 AVDD.n2868 2.801
R2974 AVDD.t743 AVDD.n679 2.756
R2975 AVDD.n3662 AVDD.n3661 2.686
R2976 AVDD.n3660 AVDD.n3659 2.686
R2977 AVDD.n3658 AVDD.n3657 2.686
R2978 AVDD.n3656 AVDD.n3655 2.686
R2979 AVDD.n3654 AVDD.n3653 2.686
R2980 AVDD.n3652 AVDD.n3651 2.686
R2981 AVDD.n1633 AVDD.n1632 2.686
R2982 AVDD.n1635 AVDD.n1634 2.686
R2983 AVDD.n1637 AVDD.n1636 2.686
R2984 AVDD.n1639 AVDD.n1638 2.686
R2985 AVDD.n1641 AVDD.n1640 2.686
R2986 AVDD.n1643 AVDD.n1642 2.686
R2987 AVDD.n1645 AVDD.n1644 2.686
R2988 AVDD.n1647 AVDD.n1646 2.686
R2989 AVDD.n3666 AVDD.n3665 2.686
R2990 AVDD.n3664 AVDD.n3663 2.686
R2991 AVDD.n3668 AVDD.n3667 2.686
R2992 AVDD.n4308 AVDD.n4304 2.677
R2993 AVDD.n1460 AVDD.n1459 2.676
R2994 AVDD.n1456 AVDD.n1455 2.676
R2995 AVDD.n1451 AVDD.n1450 2.676
R2996 AVDD.n1446 AVDD.n1445 2.676
R2997 AVDD.n1441 AVDD.n1440 2.676
R2998 AVDD.n1436 AVDD.n1435 2.676
R2999 AVDD.n1432 AVDD.n1431 2.676
R3000 AVDD.n1426 AVDD.n1425 2.676
R3001 AVDD.n4321 AVDD.n4316 2.659
R3002 AVDD.t829 AVDD.n6002 2.595
R3003 AVDD.n3445 AVDD.n3406 2.565
R3004 AVDD.n1981 AVDD.n1979 2.489
R3005 AVDD.n4309 AVDD.n4308 2.481
R3006 AVDD.n3998 AVDD.n3997 2.481
R3007 AVDD.n5501 AVDD.n1875 2.479
R3008 AVDD.t351 AVDD.t727 2.462
R3009 AVDD.n5047 AVDD.n5046 2.393
R3010 AVDD.n1190 AVDD.n1189 2.288
R3011 AVDD.t363 AVDD.n6110 2.287
R3012 AVDD.t816 AVDD.n6315 2.287
R3013 AVDD.n6138 AVDD.t363 2.287
R3014 AVDD.n1175 AVDD.n1174 2.275
R3015 AVDD.n5621 AVDD.n1059 2.123
R3016 AVDD.n4009 AVDD.n4008 2.109
R3017 AVDD.n4324 AVDD.n4321 2.003
R3018 AVDD.n5597 AVDD.n1265 1.995
R3019 AVDD.t285 AVDD.t48 1.935
R3020 AVDD.n1628 AVDD.n1627 1.879
R3021 AVDD.n6431 AVDD.n6430 1.875
R3022 AVDD.n5501 AVDD.n1769 1.874
R3023 AVDD.n507 AVDD.n503 1.873
R3024 AVDD.n506 AVDD.n504 1.854
R3025 AVDD.n6358 AVDD.t283 1.817
R3026 AVDD.n30 AVDD.n28 1.817
R3027 AVDD.t810 AVDD.n6490 1.817
R3028 AVDD.n5657 AVDD.n140 1.817
R3029 AVDD.n1538 AVDD.n1537 1.804
R3030 AVDD.n5597 AVDD.n1470 1.794
R3031 AVDD.n424 AVDD.n421 1.759
R3032 AVDD.n4388 AVDD.n4309 1.737
R3033 AVDD.n5900 AVDD.n5898 1.71
R3034 AVDD.n5042 AVDD.n5041 1.703
R3035 AVDD.t21 AVDD.t361 1.7
R3036 AVDD.t812 AVDD.n6549 1.7
R3037 AVDD.n5900 AVDD.t20 1.641
R3038 AVDD.n6549 AVDD.n6500 1.641
R3039 AVDD.n6090 AVDD.t359 1.627
R3040 AVDD.n3672 AVDD.n3671 1.622
R3041 AVDD.n1356 AVDD.n1344 1.621
R3042 AVDD.n1362 AVDD.n1361 1.6
R3043 AVDD.n6394 AVDD.n6393 1.583
R3044 AVDD.n2667 AVDD.n2627 1.557
R3045 AVDD.n5248 AVDD.n2778 1.552
R3046 AVDD.t99 AVDD.n6567 1.524
R3047 AVDD.n2778 AVDD.n2776 1.481
R3048 AVDD.n5301 AVDD.n2667 1.471
R3049 AVDD.n3542 AVDD.n3541 1.458
R3050 AVDD.n4021 AVDD.n4020 1.453
R3051 AVDD.n3997 AVDD.n3996 1.436
R3052 AVDD.t147 AVDD.n5915 1.407
R3053 AVDD.n6376 AVDD.n6371 1.289
R3054 AVDD.n6399 AVDD.n6381 1.289
R3055 AVDD.n6400 AVDD.n6380 1.289
R3056 AVDD.n6406 AVDD.n6379 1.289
R3057 AVDD.n6389 AVDD.n6388 1.289
R3058 AVDD.n6390 AVDD.n6387 1.289
R3059 AVDD.n6391 AVDD.n6386 1.289
R3060 AVDD.n6392 AVDD.n6385 1.289
R3061 AVDD.n6395 AVDD.n6384 1.289
R3062 AVDD.n6396 AVDD.n6383 1.289
R3063 AVDD.n6397 AVDD.n6382 1.289
R3064 AVDD.n4027 AVDD.n4026 1.24
R3065 AVDD.n4401 AVDD.n4031 1.238
R3066 AVDD.n3565 AVDD.n3564 1.214
R3067 AVDD.n3675 AVDD.n3672 1.214
R3068 AVDD.n4349 AVDD.n4348 1.173
R3069 AVDD.t814 AVDD.n5952 1.172
R3070 AVDD.n4999 AVDD.n4979 1.158
R3071 AVDD.n6399 AVDD.n6398 1.133
R3072 AVDD.n3028 AVDD.t161 1.081
R3073 AVDD.t25 AVDD.n3215 1.081
R3074 AVDD.n13 AVDD.n12 1.07
R3075 AVDD.n6290 AVDD.n6289 1.057
R3076 AVDD.n6284 AVDD.n6281 1.057
R3077 AVDD.n6284 AVDD.n6283 1.057
R3078 AVDD.n5748 AVDD.n5745 1.057
R3079 AVDD.n6267 AVDD.n6266 1.049
R3080 AVDD.n6261 AVDD.n6258 1.049
R3081 AVDD.n6261 AVDD.n6260 1.049
R3082 AVDD.n5738 AVDD.n5735 1.049
R3083 AVDD.n6244 AVDD.n6243 1.049
R3084 AVDD.n6238 AVDD.n6235 1.049
R3085 AVDD.n6238 AVDD.n6237 1.049
R3086 AVDD.n5730 AVDD.n5727 1.049
R3087 AVDD.n6221 AVDD.n6220 1.049
R3088 AVDD.n6215 AVDD.n6212 1.049
R3089 AVDD.n6215 AVDD.n6214 1.049
R3090 AVDD.n5722 AVDD.n5719 1.049
R3091 AVDD.n6198 AVDD.n6197 1.049
R3092 AVDD.n6192 AVDD.n6190 1.049
R3093 AVDD.n6192 AVDD.n6191 1.049
R3094 AVDD.n6154 AVDD.n6153 1.049
R3095 AVDD.n6148 AVDD.n6146 1.049
R3096 AVDD.n6148 AVDD.n6147 1.049
R3097 AVDD.n5797 AVDD.n5796 1.049
R3098 AVDD.n5791 AVDD.n5788 1.049
R3099 AVDD.n5791 AVDD.n5790 1.049
R3100 AVDD.n6300 AVDD.n6297 1.049
R3101 AVDD.n5755 AVDD.n5754 1.049
R3102 AVDD.n5774 AVDD.n5771 1.049
R3103 AVDD.n5774 AVDD.n5773 1.049
R3104 AVDD.n4020 AVDD.n4009 1.028
R3105 AVDD.t23 AVDD.t14 1.004
R3106 AVDD.n2848 AVDD.n2828 1.004
R3107 AVDD.n2171 AVDD.n2149 0.987
R3108 AVDD.n2396 AVDD.n2374 0.987
R3109 AVDD.n3052 AVDD.n3030 0.987
R3110 AVDD.n3164 AVDD.n3142 0.987
R3111 AVDD.n6294 AVDD.n6293 0.963
R3112 AVDD.n4413 AVDD.n3779 0.951
R3113 AVDD.n2169 AVDD.t130 0.926
R3114 AVDD.n3482 AVDD.n3481 0.908
R3115 AVDD.n4550 AVDD.n4549 0.893
R3116 AVDD.n4522 AVDD.n4521 0.893
R3117 AVDD.n4446 AVDD.n4445 0.893
R3118 AVDD.n4418 AVDD.n4417 0.893
R3119 AVDD.n3711 AVDD.n3710 0.893
R3120 AVDD.n3008 AVDD.n3007 0.871
R3121 AVDD.n5149 AVDD.n3165 0.866
R3122 AVDD.n15 AVDD.n13 0.812
R3123 AVDD.n3790 AVDD.n3787 0.808
R3124 AVDD.n3885 AVDD.n3882 0.808
R3125 AVDD.n3955 AVDD.n3951 0.808
R3126 AVDD.n4100 AVDD.n4097 0.808
R3127 AVDD.n4398 AVDD.n4397 0.808
R3128 AVDD.n4170 AVDD.n4166 0.808
R3129 AVDD.n5823 AVDD.n5820 0.803
R3130 AVDD.n5882 AVDD.n5879 0.803
R3131 AVDD.n6417 AVDD.n6414 0.803
R3132 AVDD.n2352 AVDD.n2351 0.796
R3133 AVDD.n4409 AVDD.n4028 0.788
R3134 AVDD.n5397 AVDD.n2172 0.786
R3135 AVDD.t725 AVDD.n30 0.762
R3136 AVDD.t59 AVDD.n5900 0.762
R3137 AVDD.n6410 AVDD.n6406 0.737
R3138 AVDD.n3675 AVDD.n3674 0.732
R3139 AVDD.n1470 AVDD.n1469 0.695
R3140 AVDD.n1650 AVDD.n1628 0.695
R3141 AVDD.n1560 AVDD.n1538 0.695
R3142 AVDD.n1769 AVDD.n1768 0.695
R3143 AVDD.n2172 AVDD.n2171 0.695
R3144 AVDD.n2374 AVDD.n2352 0.695
R3145 AVDD.n3030 AVDD.n3008 0.695
R3146 AVDD.n3165 AVDD.n3164 0.695
R3147 AVDD.n5041 AVDD.n5040 0.695
R3148 AVDD.n3674 AVDD.n3673 0.689
R3149 AVDD.n2059 AVDD.n2058 0.657
R3150 AVDD.n5398 AVDD.n2050 0.657
R3151 AVDD.n4355 AVDD.n4354 0.656
R3152 AVDD.n4358 AVDD.n4357 0.656
R3153 AVDD.n4346 AVDD.n4345 0.656
R3154 AVDD.n4489 AVDD.n4487 0.65
R3155 AVDD.n4558 AVDD.n4556 0.65
R3156 AVDD.n4530 AVDD.n4528 0.65
R3157 AVDD.n4454 AVDD.n4452 0.65
R3158 AVDD.n4426 AVDD.n4424 0.65
R3159 AVDD.n3719 AVDD.n3717 0.65
R3160 AVDD.n3549 AVDD.n3547 0.65
R3161 AVDD.n3470 AVDD.n3468 0.65
R3162 AVDD.n3556 AVDD.n3554 0.642
R3163 AVDD.n3726 AVDD.n3724 0.642
R3164 AVDD.n4429 AVDD.n4427 0.642
R3165 AVDD.n4505 AVDD.n4503 0.642
R3166 AVDD.n4537 AVDD.n4535 0.642
R3167 AVDD.n4589 AVDD.n4587 0.642
R3168 AVDD.n3477 AVDD.n3475 0.642
R3169 AVDD.n4492 AVDD.n4490 0.641
R3170 AVDD.n6408 AVDD.n6407 0.639
R3171 AVDD.n4008 AVDD.n4007 0.63
R3172 AVDD.n1658 AVDD.n1657 0.624
R3173 AVDD.n865 AVDD.n860 0.617
R3174 AVDD.n4481 AVDD.n4480 0.615
R3175 AVDD.n4342 AVDD.n4340 0.611
R3176 AVDD.n4280 AVDD.n4278 0.611
R3177 AVDD.n4005 AVDD.n4004 0.61
R3178 AVDD.n3991 AVDD.n3990 0.61
R3179 AVDD.n4264 AVDD.n4263 0.61
R3180 AVDD.n4275 AVDD.n4274 0.61
R3181 AVDD.n4290 AVDD.n4289 0.61
R3182 AVDD.n4337 AVDD.n4336 0.61
R3183 AVDD.n4016 AVDD.n4015 0.61
R3184 AVDD.n4334 AVDD.n4333 0.61
R3185 AVDD.n4287 AVDD.n4286 0.61
R3186 AVDD.n4272 AVDD.n4271 0.61
R3187 AVDD.n4261 AVDD.n4260 0.61
R3188 AVDD.n4002 AVDD.n4001 0.61
R3189 AVDD.n4012 AVDD.n4011 0.61
R3190 AVDD.n3988 AVDD.n3987 0.61
R3191 AVDD.n4338 AVDD.n4337 0.61
R3192 AVDD.n4333 AVDD.n4332 0.61
R3193 AVDD.n4340 AVDD.n4339 0.61
R3194 AVDD.n4351 AVDD.n4350 0.61
R3195 AVDD.n4291 AVDD.n4290 0.61
R3196 AVDD.n4286 AVDD.n4285 0.61
R3197 AVDD.n4278 AVDD.n4277 0.61
R3198 AVDD.n4282 AVDD.n4281 0.61
R3199 AVDD.n4276 AVDD.n4275 0.61
R3200 AVDD.n4271 AVDD.n4270 0.61
R3201 AVDD.n4265 AVDD.n4264 0.61
R3202 AVDD.n4260 AVDD.n4259 0.61
R3203 AVDD.n4006 AVDD.n4005 0.61
R3204 AVDD.n4001 AVDD.n4000 0.61
R3205 AVDD.n4015 AVDD.n4014 0.61
R3206 AVDD.n4011 AVDD.n4010 0.61
R3207 AVDD.n3992 AVDD.n3991 0.61
R3208 AVDD.n3987 AVDD.n3986 0.61
R3209 AVDD.n5045 AVDD.n5044 0.609
R3210 AVDD.n4306 AVDD.n4305 0.606
R3211 AVDD.n4330 AVDD.n4329 0.606
R3212 AVDD.n4326 AVDD.n4325 0.606
R3213 AVDD.n2048 AVDD.n1982 0.6
R3214 AVDD.n1627 AVDD.n1561 0.599
R3215 AVDD.n1836 AVDD.n1770 0.599
R3216 AVDD.n2463 AVDD.n2397 0.599
R3217 AVDD.n2627 AVDD.n2561 0.599
R3218 AVDD.n3007 AVDD.n2941 0.599
R3219 AVDD.n3406 AVDD.n3340 0.599
R3220 AVDD.n3339 AVDD.n3273 0.595
R3221 AVDD.n1423 AVDD.n1267 0.594
R3222 AVDD.n1262 AVDD.n1196 0.594
R3223 AVDD.n1537 AVDD.n1471 0.594
R3224 AVDD.n1979 AVDD.n1913 0.594
R3225 AVDD.n2351 AVDD.n2285 0.594
R3226 AVDD.n2776 AVDD.n2710 0.594
R3227 AVDD.n2939 AVDD.n2873 0.594
R3228 AVDD.n5046 AVDD.n5045 0.586
R3229 AVDD.n6398 AVDD.n6397 0.584
R3230 AVDD.n3712 AVDD.n3711 0.58
R3231 AVDD.n4601 AVDD.n4600 0.58
R3232 AVDD.n4419 AVDD.n4418 0.58
R3233 AVDD.n3458 AVDD.n3457 0.58
R3234 AVDD.n4447 AVDD.n4446 0.58
R3235 AVDD.n4438 AVDD.n4436 0.58
R3236 AVDD.n4523 AVDD.n4522 0.58
R3237 AVDD.n4514 AVDD.n4512 0.58
R3238 AVDD.n4551 AVDD.n4550 0.58
R3239 AVDD.n3465 AVDD.n3464 0.58
R3240 AVDD.n3483 AVDD.n3482 0.58
R3241 AVDD.n6280 AVDD.n6279 0.567
R3242 AVDD.n1265 AVDD.n1264 0.564
R3243 AVDD.n5770 AVDD.n5769 0.563
R3244 AVDD.n5787 AVDD.n5786 0.563
R3245 AVDD.n6145 AVDD.n6144 0.563
R3246 AVDD.n6189 AVDD.n6188 0.563
R3247 AVDD.n6211 AVDD.n6210 0.563
R3248 AVDD.n6234 AVDD.n6233 0.563
R3249 AVDD.n6257 AVDD.n6256 0.563
R3250 AVDD.n2149 AVDD.n2127 0.559
R3251 AVDD.n6288 AVDD.n6287 0.559
R3252 AVDD.n6265 AVDD.n6264 0.555
R3253 AVDD.n6242 AVDD.n6241 0.555
R3254 AVDD.n6219 AVDD.n6218 0.555
R3255 AVDD.n6196 AVDD.n6195 0.555
R3256 AVDD.n6152 AVDD.n6151 0.555
R3257 AVDD.n5795 AVDD.n5794 0.555
R3258 AVDD.n5753 AVDD.n5752 0.555
R3259 AVDD.n5353 AVDD.n2396 0.554
R3260 AVDD.n4354 AVDD.n4353 0.551
R3261 AVDD.n1875 AVDD.n1836 0.549
R3262 AVDD.n5450 AVDD.n1981 0.544
R3263 AVDD.n2559 AVDD.n2542 0.544
R3264 AVDD.n6002 AVDD.n6001 0.542
R3265 AVDD.n1727 AVDD.n1707 0.54
R3266 AVDD.n1469 AVDD.n1423 0.539
R3267 AVDD.n5040 AVDD.n5018 0.539
R3268 AVDD.n2278 AVDD.n2261 0.535
R3269 AVDD.n5546 AVDD.n1560 0.534
R3270 AVDD.n5306 AVDD.n5305 0.528
R3271 AVDD.n5257 AVDD.n5254 0.528
R3272 AVDD.t59 AVDD.n5893 0.527
R3273 AVDD.n6441 AVDD.t808 0.527
R3274 AVDD.t810 AVDD.n6496 0.527
R3275 AVDD.t87 AVDD.n6375 0.527
R3276 AVDD.n433 AVDD.t247 0.527
R3277 AVDD.n1746 AVDD.n1729 0.524
R3278 AVDD.n6406 AVDD.n6405 0.519
R3279 AVDD.n4283 AVDD.n4282 0.512
R3280 AVDD.n4352 AVDD.n4351 0.512
R3281 AVDD.n6391 AVDD.n6390 0.512
R3282 AVDD.n6397 AVDD.n6396 0.512
R3283 AVDD.n6400 AVDD.n6399 0.509
R3284 AVDD.n6395 AVDD.n6394 0.509
R3285 AVDD.n6283 AVDD.n6282 0.505
R3286 AVDD.n5745 AVDD.n5744 0.505
R3287 AVDD.n6260 AVDD.n6259 0.501
R3288 AVDD.n5735 AVDD.n5734 0.501
R3289 AVDD.n6237 AVDD.n6236 0.501
R3290 AVDD.n5727 AVDD.n5726 0.501
R3291 AVDD.n6214 AVDD.n6213 0.501
R3292 AVDD.n5719 AVDD.n5718 0.501
R3293 AVDD.n5698 AVDD.n5697 0.501
R3294 AVDD.n5714 AVDD.n5713 0.501
R3295 AVDD.n5790 AVDD.n5789 0.501
R3296 AVDD.n6297 AVDD.n6296 0.501
R3297 AVDD.n5773 AVDD.n5772 0.501
R3298 AVDD.n6293 AVDD.n6292 0.501
R3299 AVDD.n6390 AVDD.n6389 0.496
R3300 AVDD.n6392 AVDD.n6391 0.496
R3301 AVDD.n6396 AVDD.n6395 0.496
R3302 AVDD.n3142 AVDD.n3120 0.483
R3303 AVDD.n4410 AVDD.n4409 0.482
R3304 AVDD.n4347 AVDD.n4346 0.48
R3305 AVDD.n4357 AVDD.n4356 0.48
R3306 AVDD.n148 AVDD.n147 0.475
R3307 AVDD.n326 AVDD.n325 0.475
R3308 AVDD.n516 AVDD.n515 0.475
R3309 AVDD.n711 AVDD.n710 0.475
R3310 AVDD.n892 AVDD.n891 0.475
R3311 AVDD.n1063 AVDD.n1062 0.475
R3312 AVDD.n5594 AVDD.n5593 0.475
R3313 AVDD.n5543 AVDD.n5542 0.475
R3314 AVDD.n5498 AVDD.n5497 0.475
R3315 AVDD.n5447 AVDD.n5446 0.475
R3316 AVDD.n5394 AVDD.n5393 0.475
R3317 AVDD.n5209 AVDD.n5208 0.475
R3318 AVDD.n5161 AVDD.n5160 0.475
R3319 AVDD.n5110 AVDD.n5109 0.475
R3320 AVDD.n5059 AVDD.n5058 0.475
R3321 AVDD.n3455 AVDD.n3454 0.475
R3322 AVDD.n321 AVDD.n320 0.475
R3323 AVDD.n512 AVDD.n511 0.475
R3324 AVDD.n707 AVDD.n706 0.475
R3325 AVDD.n888 AVDD.n887 0.475
R3326 AVDD.n5614 AVDD.n5613 0.475
R3327 AVDD.n5601 AVDD.n5600 0.475
R3328 AVDD.n5556 AVDD.n5555 0.475
R3329 AVDD.n5505 AVDD.n5504 0.475
R3330 AVDD.n5460 AVDD.n5459 0.475
R3331 AVDD.n5406 AVDD.n5405 0.475
R3332 AVDD.n2284 AVDD.n2283 0.475
R3333 AVDD.n5310 AVDD.n5309 0.475
R3334 AVDD.n5259 AVDD.n5258 0.475
R3335 AVDD.n5206 AVDD.n5205 0.475
R3336 AVDD.n5159 AVDD.n5158 0.475
R3337 AVDD.n5108 AVDD.n5107 0.475
R3338 AVDD.n5057 AVDD.n5056 0.475
R3339 AVDD.n3453 AVDD.n3452 0.475
R3340 AVDD.n144 AVDD.n143 0.475
R3341 AVDD.n324 AVDD.n323 0.475
R3342 AVDD.n514 AVDD.n513 0.475
R3343 AVDD.n709 AVDD.n708 0.475
R3344 AVDD.n890 AVDD.n889 0.475
R3345 AVDD.n1061 AVDD.n1060 0.475
R3346 AVDD.n5596 AVDD.n5595 0.475
R3347 AVDD.n5545 AVDD.n5544 0.475
R3348 AVDD.n5500 AVDD.n5499 0.475
R3349 AVDD.n5449 AVDD.n5448 0.475
R3350 AVDD.n5396 AVDD.n5395 0.475
R3351 AVDD.n5352 AVDD.n5351 0.475
R3352 AVDD.n5247 AVDD.n5246 0.475
R3353 AVDD.n5199 AVDD.n5198 0.475
R3354 AVDD.n5148 AVDD.n5147 0.475
R3355 AVDD.n5097 AVDD.n5096 0.475
R3356 AVDD.n4905 AVDD.n4904 0.475
R3357 AVDD.n3447 AVDD.n3446 0.475
R3358 AVDD.n5051 AVDD.n5050 0.475
R3359 AVDD.n5102 AVDD.n5101 0.475
R3360 AVDD.n5153 AVDD.n5152 0.475
R3361 AVDD.n2872 AVDD.n2871 0.475
R3362 AVDD.n2671 AVDD.n2670 0.475
R3363 AVDD.n5454 AVDD.n5453 0.475
R3364 AVDD.n1654 AVDD.n1653 0.475
R3365 AVDD.n5550 AVDD.n5549 0.475
R3366 AVDD.n5607 AVDD.n5606 0.475
R3367 AVDD.n5620 AVDD.n5619 0.475
R3368 AVDD.n5627 AVDD.n5626 0.475
R3369 AVDD.n5634 AVDD.n5633 0.475
R3370 AVDD.n5641 AVDD.n5640 0.475
R3371 AVDD.n5649 AVDD.n5648 0.475
R3372 AVDD.n3541 AVDD.n3540 0.473
R3373 AVDD.n1264 AVDD.n1262 0.473
R3374 AVDD.n5200 AVDD.n3052 0.473
R3375 AVDD.n2867 AVDD.n2850 0.468
R3376 AVDD.n5299 AVDD.n5298 0.468
R3377 AVDD.n1768 AVDD.n1746 0.463
R3378 AVDD.n2061 AVDD.n2060 0.463
R3379 AVDD.n5098 AVDD.n3445 0.463
R3380 AVDD.t42 AVDD.n2239 0.463
R3381 AVDD.n2372 AVDD.t91 0.463
R3382 AVDD.n4549 AVDD.n4548 0.462
R3383 AVDD.n4521 AVDD.n4520 0.462
R3384 AVDD.n4445 AVDD.n4444 0.462
R3385 AVDD.n4417 AVDD.n4416 0.462
R3386 AVDD.n3710 AVDD.n3709 0.462
R3387 AVDD.n3271 AVDD.n3254 0.459
R3388 AVDD.n6289 AVDD.n6288 0.457
R3389 AVDD.n5711 AVDD.n5710 0.454
R3390 AVDD.n6308 AVDD.n6307 0.454
R3391 AVDD.n6266 AVDD.n6265 0.454
R3392 AVDD.n6243 AVDD.n6242 0.454
R3393 AVDD.n6220 AVDD.n6219 0.454
R3394 AVDD.n6197 AVDD.n6196 0.454
R3395 AVDD.n6153 AVDD.n6152 0.454
R3396 AVDD.n5796 AVDD.n5795 0.454
R3397 AVDD.n5754 AVDD.n5753 0.454
R3398 AVDD.n2056 AVDD.n2055 0.453
R3399 AVDD.n2467 AVDD.n2466 0.453
R3400 AVDD.n2669 AVDD.n2668 0.453
R3401 AVDD.n2870 AVDD.n2869 0.453
R3402 AVDD.n5151 AVDD.n5150 0.453
R3403 AVDD.n5100 AVDD.n5099 0.453
R3404 AVDD.n5049 AVDD.n5048 0.453
R3405 AVDD.n4929 AVDD.n4928 0.453
R3406 AVDD.n5546 AVDD.n1650 0.453
R3407 AVDD.n5452 AVDD.n5451 0.453
R3408 AVDD.n1652 AVDD.n1651 0.453
R3409 AVDD.n5548 AVDD.n5547 0.453
R3410 AVDD.n1165 AVDD.n1164 0.453
R3411 AVDD.n5610 AVDD.n5609 0.453
R3412 AVDD.n884 AVDD.n883 0.453
R3413 AVDD.n703 AVDD.n702 0.453
R3414 AVDD.n316 AVDD.n315 0.453
R3415 AVDD.n5652 AVDD.n5651 0.453
R3416 AVDD.n5644 AVDD.n5643 0.453
R3417 AVDD.n5637 AVDD.n5636 0.453
R3418 AVDD.n5630 AVDD.n5629 0.453
R3419 AVDD.n5623 AVDD.n5622 0.453
R3420 AVDD.n5616 AVDD.n5615 0.453
R3421 AVDD.n5603 AVDD.n5602 0.453
R3422 AVDD.n5554 AVDD.n5553 0.453
R3423 AVDD.n5503 AVDD.n5502 0.453
R3424 AVDD.n5458 AVDD.n5457 0.453
R3425 AVDD.n5404 AVDD.n5403 0.453
R3426 AVDD.n2282 AVDD.n2281 0.453
R3427 AVDD.n5308 AVDD.n5307 0.453
R3428 AVDD.n5256 AVDD.n5255 0.453
R3429 AVDD.n5204 AVDD.n5203 0.453
R3430 AVDD.n5157 AVDD.n5156 0.453
R3431 AVDD.n5106 AVDD.n5105 0.453
R3432 AVDD.n5055 AVDD.n5054 0.453
R3433 AVDD.n3451 AVDD.n3450 0.453
R3434 AVDD.n5655 AVDD.n5654 0.453
R3435 AVDD.n5646 AVDD.n5645 0.453
R3436 AVDD.n5639 AVDD.n5638 0.453
R3437 AVDD.n5632 AVDD.n5631 0.453
R3438 AVDD.n5625 AVDD.n5624 0.453
R3439 AVDD.n5618 AVDD.n5617 0.453
R3440 AVDD.n5605 AVDD.n5604 0.453
R3441 AVDD.n5552 AVDD.n5551 0.453
R3442 AVDD.n1656 AVDD.n1655 0.453
R3443 AVDD.n5456 AVDD.n5455 0.453
R3444 AVDD.n5402 AVDD.n5401 0.453
R3445 AVDD.n2280 AVDD.n2279 0.453
R3446 AVDD.n5202 AVDD.n5201 0.453
R3447 AVDD.n5155 AVDD.n5154 0.453
R3448 AVDD.n5104 AVDD.n5103 0.453
R3449 AVDD.n5053 AVDD.n5052 0.453
R3450 AVDD.n3449 AVDD.n3448 0.453
R3451 AVDD.n4827 AVDD.n4826 0.453
R3452 AVDD.n5061 AVDD.n5060 0.453
R3453 AVDD.n5112 AVDD.n5111 0.453
R3454 AVDD.n5163 AVDD.n5162 0.453
R3455 AVDD.n5211 AVDD.n5210 0.453
R3456 AVDD.n5261 AVDD.n5260 0.453
R3457 AVDD.n5312 AVDD.n5311 0.453
R3458 AVDD.n5355 AVDD.n5354 0.453
R3459 AVDD.n5411 AVDD.n5410 0.453
R3460 AVDD.n5462 AVDD.n5461 0.453
R3461 AVDD.n5507 AVDD.n5506 0.453
R3462 AVDD.n5558 AVDD.n5557 0.453
R3463 AVDD.n5599 AVDD.n5598 0.453
R3464 AVDD.n5612 AVDD.n5611 0.453
R3465 AVDD.n886 AVDD.n885 0.453
R3466 AVDD.n705 AVDD.n704 0.453
R3467 AVDD.n510 AVDD.n509 0.453
R3468 AVDD.n318 AVDD.n317 0.453
R3469 AVDD.n5399 AVDD.n5398 0.452
R3470 AVDD.n5303 AVDD.n5302 0.452
R3471 AVDD.n5252 AVDD.n5249 0.452
R3472 AVDD.n3481 AVDD.n3480 0.45
R3473 AVDD.n4909 AVDD.n4908 0.449
R3474 AVDD.n3461 AVDD.n3460 0.449
R3475 AVDD.n4604 AVDD.n4603 0.449
R3476 AVDD.n4599 AVDD.n4598 0.449
R3477 AVDD.n6281 AVDD.n6280 0.449
R3478 AVDD.n5018 AVDD.n5001 0.448
R3479 AVDD.n6258 AVDD.n6257 0.446
R3480 AVDD.n6235 AVDD.n6234 0.446
R3481 AVDD.n6212 AVDD.n6211 0.446
R3482 AVDD.n6190 AVDD.n6189 0.446
R3483 AVDD.n6146 AVDD.n6145 0.446
R3484 AVDD.n5788 AVDD.n5787 0.446
R3485 AVDD.n5771 AVDD.n5770 0.446
R3486 AVDD.n2054 AVDD.n2053 0.422
R3487 AVDD.n2468 AVDD.n2465 0.422
R3488 AVDD.n6105 AVDD.n6090 0.416
R3489 AVDD.t9 AVDD.t97 0.41
R3490 AVDD.n4365 AVDD.n4364 0.406
R3491 AVDD.n4362 AVDD.n4361 0.406
R3492 AVDD.n4366 AVDD.n4365 0.406
R3493 AVDD.n4361 AVDD.n4360 0.406
R3494 AVDD.n4390 AVDD.n4389 0.402
R3495 AVDD.n5890 AVDD.n5889 0.388
R3496 AVDD.n2540 AVDD.n2520 0.386
R3497 AVDD.t46 AVDD.t208 0.386
R3498 AVDD.n3054 AVDD.n3053 0.382
R3499 AVDD.n5302 AVDD.n2470 0.372
R3500 AVDD.n5252 AVDD.n5251 0.372
R3501 AVDD.n6369 AVDD.n6368 0.365
R3502 AVDD.n5350 AVDD.n5349 0.361
R3503 AVDD.n5889 AVDD.n5888 0.326
R3504 AVDD.n621 AVDD.n572 0.308
R3505 AVDD.n1295 AVDD.n1278 0.308
R3506 AVDD.n3162 AVDD.t172 0.308
R3507 AVDD.n5358 AVDD.n5357 0.305
R3508 AVDD.n5409 AVDD.n5408 0.305
R3509 AVDD.n5829 AVDD.n5823 0.294
R3510 AVDD.n6061 AVDD.n5882 0.294
R3511 AVDD.n6418 AVDD.n6417 0.294
R3512 AVDD.n3797 AVDD.n3790 0.29
R3513 AVDD.n3886 AVDD.n3885 0.29
R3514 AVDD.n3956 AVDD.n3955 0.29
R3515 AVDD.n4101 AVDD.n4100 0.29
R3516 AVDD.n4397 AVDD.n4394 0.29
R3517 AVDD.n4171 AVDD.n4170 0.29
R3518 AVDD.n4220 AVDD.n4219 0.288
R3519 AVDD.n2052 AVDD.n2051 0.285
R3520 AVDD.n5299 AVDD.n5297 0.283
R3521 AVDD.n6377 AVDD.n6376 0.278
R3522 AVDD.n6359 AVDD.n6358 0.262
R3523 AVDD.n6359 AVDD.n5657 0.262
R3524 AVDD.n3273 AVDD.n3272 0.262
R3525 AVDD.n4482 AVDD.n4481 0.26
R3526 AVDD.n3484 AVDD.n3483 0.26
R3527 AVDD.n4552 AVDD.n4551 0.26
R3528 AVDD.n4524 AVDD.n4523 0.26
R3529 AVDD.n4448 AVDD.n4447 0.26
R3530 AVDD.n4420 AVDD.n4419 0.26
R3531 AVDD.n3713 AVDD.n3712 0.26
R3532 AVDD.n3543 AVDD.n3542 0.26
R3533 AVDD.n1274 AVDD.n1273 0.257
R3534 AVDD.n4479 AVDD.n4476 0.256
R3535 AVDD.n4497 AVDD.n4496 0.255
R3536 AVDD.n3485 AVDD.n3479 0.255
R3537 AVDD.n4554 AVDD.n4553 0.255
R3538 AVDD.n4526 AVDD.n4525 0.255
R3539 AVDD.n4450 AVDD.n4449 0.255
R3540 AVDD.n4422 AVDD.n4421 0.255
R3541 AVDD.n3715 AVDD.n3714 0.255
R3542 AVDD.n3545 AVDD.n3544 0.255
R3543 AVDD.n5738 AVDD.n5733 0.253
R3544 AVDD.n5730 AVDD.n5725 0.253
R3545 AVDD.n5722 AVDD.n5717 0.253
R3546 AVDD.n5748 AVDD.n5743 0.253
R3547 AVDD.n6300 AVDD.n6295 0.253
R3548 AVDD.n3488 AVDD.n3487 0.252
R3549 AVDD.n4592 AVDD.n4547 0.252
R3550 AVDD.n4540 AVDD.n4519 0.252
R3551 AVDD.n4508 AVDD.n4443 0.252
R3552 AVDD.n4432 AVDD.n4415 0.252
R3553 AVDD.n3729 AVDD.n3708 0.252
R3554 AVDD.n3559 AVDD.n3539 0.252
R3555 AVDD.n4495 AVDD.n4493 0.245
R3556 AVDD.n568 AVDD.n567 0.237
R3557 AVDD.n561 AVDD.n560 0.237
R3558 AVDD.n4028 AVDD.n4027 0.235
R3559 AVDD.n6378 AVDD.n6377 0.233
R3560 AVDD.n4207 AVDD.n4198 0.23
R3561 AVDD.n2868 AVDD.n2867 0.226
R3562 AVDD.n5200 AVDD.n2940 0.221
R3563 AVDD.n4348 AVDD.n4347 0.211
R3564 AVDD.n3120 AVDD.n3054 0.211
R3565 AVDD.n506 AVDD.n505 0.2
R3566 AVDD.n4413 AVDD.n4412 0.199
R3567 AVDD.n4597 AVDD.n4594 0.19
R3568 AVDD.n4597 AVDD.n3734 0.19
R3569 AVDD.n4597 AVDD.n4440 0.19
R3570 AVDD.n4597 AVDD.n4516 0.19
R3571 AVDD.n4597 AVDD.n4545 0.19
R3572 AVDD.n4597 AVDD.n3706 0.19
R3573 AVDD.n4597 AVDD.n3538 0.19
R3574 AVDD.n4597 AVDD.n3502 0.19
R3575 AVDD.n4824 AVDD.n4823 0.189
R3576 AVDD.n5750 AVDD.n5749 0.189
R3577 AVDD.n5742 AVDD.n5741 0.189
R3578 AVDD.n5732 AVDD.n5731 0.189
R3579 AVDD.n5724 AVDD.n5723 0.189
R3580 AVDD.n5708 AVDD.n5707 0.189
R3581 AVDD.n6305 AVDD.n6304 0.189
R3582 AVDD.n6302 AVDD.n6301 0.189
R3583 AVDD.n4926 AVDD.n4925 0.189
R3584 AVDD.n5747 AVDD.n5746 0.189
R3585 AVDD.n5737 AVDD.n5736 0.189
R3586 AVDD.n5729 AVDD.n5728 0.189
R3587 AVDD.n5721 AVDD.n5720 0.189
R3588 AVDD.n5706 AVDD.n5705 0.189
R3589 AVDD.n5716 AVDD.n5715 0.189
R3590 AVDD.n6299 AVDD.n6298 0.189
R3591 AVDD.n4207 AVDD.n4203 0.189
R3592 AVDD.n3996 AVDD.n3995 0.189
R3593 AVDD.n3995 AVDD.n3994 0.189
R3594 AVDD.n4020 AVDD.n4019 0.189
R3595 AVDD.n4019 AVDD.n4018 0.189
R3596 AVDD.n74 AVDD.n73 0.189
R3597 AVDD.n132 AVDD.n74 0.189
R3598 AVDD.n6558 AVDD.n6557 0.189
R3599 AVDD.n6567 AVDD.n6558 0.189
R3600 AVDD.n5952 AVDD.n5943 0.189
R3601 AVDD.n6432 AVDD.n6431 0.189
R3602 AVDD.n6441 AVDD.n6432 0.189
R3603 AVDD.n248 AVDD.n190 0.189
R3604 AVDD.n314 AVDD.n305 0.189
R3605 AVDD.n698 AVDD.n689 0.189
R3606 AVDD.n502 AVDD.n493 0.189
R3607 AVDD.n370 AVDD.n369 0.189
R3608 AVDD.n433 AVDD.n370 0.189
R3609 AVDD.n5875 AVDD.n5868 0.189
R3610 AVDD.t825 AVDD.n6118 0.189
R3611 AVDD.n5705 AVDD.n5704 0.189
R3612 AVDD.n5741 AVDD.n5740 0.189
R3613 AVDD.n5952 AVDD.n5951 0.189
R3614 AVDD.n698 AVDD.n681 0.189
R3615 AVDD.n433 AVDD.n362 0.189
R3616 AVDD.n502 AVDD.n487 0.189
R3617 AVDD.n248 AVDD.n184 0.189
R3618 AVDD.n314 AVDD.n299 0.189
R3619 AVDD.n698 AVDD.n683 0.189
R3620 AVDD.n433 AVDD.n364 0.189
R3621 AVDD.n502 AVDD.n489 0.189
R3622 AVDD.n248 AVDD.n186 0.189
R3623 AVDD.n314 AVDD.n301 0.189
R3624 AVDD.n698 AVDD.n693 0.189
R3625 AVDD.n433 AVDD.n428 0.189
R3626 AVDD.n502 AVDD.n497 0.189
R3627 AVDD.n248 AVDD.n243 0.189
R3628 AVDD.n314 AVDD.n309 0.189
R3629 AVDD.n132 AVDD.n127 0.189
R3630 AVDD.n6567 AVDD.n6562 0.189
R3631 AVDD.n6441 AVDD.n6436 0.189
R3632 AVDD.n5952 AVDD.n5947 0.189
R3633 AVDD.n698 AVDD.n685 0.189
R3634 AVDD.n433 AVDD.n366 0.189
R3635 AVDD.n502 AVDD.n491 0.189
R3636 AVDD.n248 AVDD.n188 0.189
R3637 AVDD.n314 AVDD.n303 0.189
R3638 AVDD.n132 AVDD.n72 0.189
R3639 AVDD.n6567 AVDD.n6555 0.189
R3640 AVDD.n6441 AVDD.n6428 0.189
R3641 AVDD.n5952 AVDD.n5941 0.189
R3642 AVDD.n6567 AVDD.n6566 0.189
R3643 AVDD.n132 AVDD.n131 0.189
R3644 AVDD.n314 AVDD.n313 0.189
R3645 AVDD.n248 AVDD.n247 0.189
R3646 AVDD.n502 AVDD.n501 0.189
R3647 AVDD.n433 AVDD.n432 0.189
R3648 AVDD.n698 AVDD.n697 0.189
R3649 AVDD.n6441 AVDD.n6426 0.189
R3650 AVDD.n5952 AVDD.n5939 0.189
R3651 AVDD.n132 AVDD.n70 0.189
R3652 AVDD.n6567 AVDD.n6553 0.189
R3653 AVDD.n6441 AVDD.n6438 0.189
R3654 AVDD.n5952 AVDD.n5949 0.189
R3655 AVDD.n132 AVDD.n129 0.189
R3656 AVDD.n6567 AVDD.n6564 0.189
R3657 AVDD.n248 AVDD.n245 0.189
R3658 AVDD.n314 AVDD.n311 0.189
R3659 AVDD.n433 AVDD.n430 0.189
R3660 AVDD.n502 AVDD.n499 0.189
R3661 AVDD.n698 AVDD.n695 0.189
R3662 AVDD.n6441 AVDD.n6424 0.189
R3663 AVDD.n5952 AVDD.n5937 0.189
R3664 AVDD.n132 AVDD.n68 0.189
R3665 AVDD.n6567 AVDD.n6551 0.189
R3666 AVDD.n6441 AVDD.n6440 0.189
R3667 AVDD.n5875 AVDD.n5874 0.189
R3668 AVDD.t825 AVDD.n6122 0.189
R3669 AVDD.n5875 AVDD.n5860 0.189
R3670 AVDD.t825 AVDD.n6111 0.189
R3671 AVDD.n5875 AVDD.n5872 0.189
R3672 AVDD.t825 AVDD.n6121 0.189
R3673 AVDD.n5875 AVDD.n5862 0.189
R3674 AVDD.t825 AVDD.n6112 0.189
R3675 AVDD.n5875 AVDD.n5870 0.189
R3676 AVDD.t825 AVDD.n6120 0.189
R3677 AVDD.n5875 AVDD.n5864 0.189
R3678 AVDD.t825 AVDD.n6114 0.189
R3679 AVDD.n5875 AVDD.n5866 0.189
R3680 AVDD.t825 AVDD.n6116 0.189
R3681 AVDD.n5740 AVDD.n5739 0.189
R3682 AVDD.n5704 AVDD.n5703 0.189
R3683 AVDD.n6441 AVDD.n6434 0.189
R3684 AVDD.n5952 AVDD.n5945 0.189
R3685 AVDD.n132 AVDD.n125 0.189
R3686 AVDD.n6567 AVDD.n6560 0.189
R3687 AVDD.n248 AVDD.n241 0.189
R3688 AVDD.n314 AVDD.n307 0.189
R3689 AVDD.n433 AVDD.n426 0.189
R3690 AVDD.n502 AVDD.n495 0.189
R3691 AVDD.n698 AVDD.n691 0.189
R3692 AVDD.n630 AVDD.n558 0.189
R3693 AVDD.n811 AVDD.n753 0.189
R3694 AVDD.n882 AVDD.n873 0.189
R3695 AVDD.n992 AVDD.n934 0.189
R3696 AVDD.n1058 AVDD.n1049 0.189
R3697 AVDD.n1295 AVDD.n1286 0.189
R3698 AVDD.n1163 AVDD.n1154 0.189
R3699 AVDD.n4822 AVDD.n4815 0.189
R3700 AVDD.n4709 AVDD.n4694 0.189
R3701 AVDD.n5016 AVDD.n5003 0.189
R3702 AVDD.n3337 AVDD.n3275 0.189
R3703 AVDD.n3404 AVDD.n3391 0.189
R3704 AVDD.n3118 AVDD.n3056 0.189
R3705 AVDD.n3269 AVDD.n3256 0.189
R3706 AVDD.n2937 AVDD.n2875 0.189
R3707 AVDD.n3005 AVDD.n2992 0.189
R3708 AVDD.n2774 AVDD.n2712 0.189
R3709 AVDD.n2865 AVDD.n2852 0.189
R3710 AVDD.n2557 AVDD.n2544 0.189
R3711 AVDD.n2625 AVDD.n2612 0.189
R3712 AVDD.n2349 AVDD.n2287 0.189
R3713 AVDD.n2461 AVDD.n2448 0.189
R3714 AVDD.n2276 AVDD.n2263 0.189
R3715 AVDD.n2125 AVDD.n2112 0.189
R3716 AVDD.n1977 AVDD.n1915 0.189
R3717 AVDD.n2046 AVDD.n2033 0.189
R3718 AVDD.n1744 AVDD.n1731 0.189
R3719 AVDD.n1834 AVDD.n1821 0.189
R3720 AVDD.n1535 AVDD.n1473 0.189
R3721 AVDD.n1625 AVDD.n1612 0.189
R3722 AVDD.n1260 AVDD.n1198 0.189
R3723 AVDD.n1421 AVDD.n1408 0.189
R3724 AVDD.n1295 AVDD.n1280 0.189
R3725 AVDD.n1163 AVDD.n1148 0.189
R3726 AVDD.n992 AVDD.n928 0.189
R3727 AVDD.n1058 AVDD.n1043 0.189
R3728 AVDD.n811 AVDD.n747 0.189
R3729 AVDD.n882 AVDD.n867 0.189
R3730 AVDD.n630 AVDD.n552 0.189
R3731 AVDD.n4709 AVDD.n4706 0.189
R3732 AVDD.n5016 AVDD.n5013 0.189
R3733 AVDD.n3337 AVDD.n3334 0.189
R3734 AVDD.n3404 AVDD.n3401 0.189
R3735 AVDD.n3118 AVDD.n3115 0.189
R3736 AVDD.n3269 AVDD.n3266 0.189
R3737 AVDD.n2937 AVDD.n2934 0.189
R3738 AVDD.n3005 AVDD.n3002 0.189
R3739 AVDD.n2774 AVDD.n2771 0.189
R3740 AVDD.n2865 AVDD.n2862 0.189
R3741 AVDD.n4709 AVDD.n4696 0.189
R3742 AVDD.n5016 AVDD.n5005 0.189
R3743 AVDD.n3337 AVDD.n3277 0.189
R3744 AVDD.n3404 AVDD.n3393 0.189
R3745 AVDD.n3118 AVDD.n3058 0.189
R3746 AVDD.n3269 AVDD.n3258 0.189
R3747 AVDD.n2937 AVDD.n2877 0.189
R3748 AVDD.n3005 AVDD.n2994 0.189
R3749 AVDD.n2774 AVDD.n2714 0.189
R3750 AVDD.n2865 AVDD.n2854 0.189
R3751 AVDD.n2557 AVDD.n2546 0.189
R3752 AVDD.n2625 AVDD.n2614 0.189
R3753 AVDD.n2349 AVDD.n2289 0.189
R3754 AVDD.n2461 AVDD.n2450 0.189
R3755 AVDD.n2276 AVDD.n2265 0.189
R3756 AVDD.n2125 AVDD.n2114 0.189
R3757 AVDD.n1977 AVDD.n1917 0.189
R3758 AVDD.n2046 AVDD.n2035 0.189
R3759 AVDD.n1744 AVDD.n1733 0.189
R3760 AVDD.n1834 AVDD.n1823 0.189
R3761 AVDD.n1535 AVDD.n1475 0.189
R3762 AVDD.n1625 AVDD.n1614 0.189
R3763 AVDD.n1260 AVDD.n1200 0.189
R3764 AVDD.n1421 AVDD.n1410 0.189
R3765 AVDD.n1295 AVDD.n1282 0.189
R3766 AVDD.n1163 AVDD.n1150 0.189
R3767 AVDD.n992 AVDD.n930 0.189
R3768 AVDD.n1058 AVDD.n1045 0.189
R3769 AVDD.n811 AVDD.n749 0.189
R3770 AVDD.n882 AVDD.n869 0.189
R3771 AVDD.n630 AVDD.n554 0.189
R3772 AVDD.n4709 AVDD.n4704 0.189
R3773 AVDD.n5016 AVDD.n5011 0.189
R3774 AVDD.n3337 AVDD.n3332 0.189
R3775 AVDD.n3404 AVDD.n3399 0.189
R3776 AVDD.n3118 AVDD.n3113 0.189
R3777 AVDD.n3269 AVDD.n3264 0.189
R3778 AVDD.n2937 AVDD.n2932 0.189
R3779 AVDD.n3005 AVDD.n3000 0.189
R3780 AVDD.n2774 AVDD.n2769 0.189
R3781 AVDD.n2865 AVDD.n2860 0.189
R3782 AVDD.n2557 AVDD.n2552 0.189
R3783 AVDD.n2625 AVDD.n2620 0.189
R3784 AVDD.n2349 AVDD.n2344 0.189
R3785 AVDD.n2461 AVDD.n2456 0.189
R3786 AVDD.n2276 AVDD.n2271 0.189
R3787 AVDD.n2125 AVDD.n2120 0.189
R3788 AVDD.n1977 AVDD.n1972 0.189
R3789 AVDD.n2046 AVDD.n2041 0.189
R3790 AVDD.n1744 AVDD.n1739 0.189
R3791 AVDD.n1834 AVDD.n1829 0.189
R3792 AVDD.n1535 AVDD.n1530 0.189
R3793 AVDD.n1625 AVDD.n1620 0.189
R3794 AVDD.n1260 AVDD.n1255 0.189
R3795 AVDD.n1421 AVDD.n1416 0.189
R3796 AVDD.n1295 AVDD.n1290 0.189
R3797 AVDD.n1163 AVDD.n1158 0.189
R3798 AVDD.n992 AVDD.n987 0.189
R3799 AVDD.n1058 AVDD.n1053 0.189
R3800 AVDD.n811 AVDD.n806 0.189
R3801 AVDD.n882 AVDD.n877 0.189
R3802 AVDD.n630 AVDD.n625 0.189
R3803 AVDD.n4709 AVDD.n4698 0.189
R3804 AVDD.n5016 AVDD.n5007 0.189
R3805 AVDD.n3337 AVDD.n3279 0.189
R3806 AVDD.n3404 AVDD.n3395 0.189
R3807 AVDD.n3118 AVDD.n3060 0.189
R3808 AVDD.n3269 AVDD.n3260 0.189
R3809 AVDD.n2937 AVDD.n2879 0.189
R3810 AVDD.n3005 AVDD.n2996 0.189
R3811 AVDD.n2774 AVDD.n2716 0.189
R3812 AVDD.n2865 AVDD.n2856 0.189
R3813 AVDD.n2557 AVDD.n2548 0.189
R3814 AVDD.n2625 AVDD.n2616 0.189
R3815 AVDD.n2349 AVDD.n2291 0.189
R3816 AVDD.n2461 AVDD.n2452 0.189
R3817 AVDD.n2276 AVDD.n2267 0.189
R3818 AVDD.n2125 AVDD.n2116 0.189
R3819 AVDD.n1977 AVDD.n1919 0.189
R3820 AVDD.n2046 AVDD.n2037 0.189
R3821 AVDD.n1744 AVDD.n1735 0.189
R3822 AVDD.n1834 AVDD.n1825 0.189
R3823 AVDD.n1535 AVDD.n1477 0.189
R3824 AVDD.n1625 AVDD.n1616 0.189
R3825 AVDD.n1260 AVDD.n1202 0.189
R3826 AVDD.n1421 AVDD.n1412 0.189
R3827 AVDD.n1295 AVDD.n1284 0.189
R3828 AVDD.n1163 AVDD.n1152 0.189
R3829 AVDD.n992 AVDD.n932 0.189
R3830 AVDD.n1058 AVDD.n1047 0.189
R3831 AVDD.n811 AVDD.n751 0.189
R3832 AVDD.n882 AVDD.n871 0.189
R3833 AVDD.n630 AVDD.n556 0.189
R3834 AVDD.n630 AVDD.n629 0.189
R3835 AVDD.n882 AVDD.n881 0.189
R3836 AVDD.n811 AVDD.n810 0.189
R3837 AVDD.n1058 AVDD.n1057 0.189
R3838 AVDD.n992 AVDD.n991 0.189
R3839 AVDD.n1163 AVDD.n1162 0.189
R3840 AVDD.n1295 AVDD.n1294 0.189
R3841 AVDD.n1421 AVDD.n1420 0.189
R3842 AVDD.n1260 AVDD.n1259 0.189
R3843 AVDD.n1625 AVDD.n1624 0.189
R3844 AVDD.n1535 AVDD.n1534 0.189
R3845 AVDD.n1834 AVDD.n1833 0.189
R3846 AVDD.n1744 AVDD.n1743 0.189
R3847 AVDD.n2046 AVDD.n2045 0.189
R3848 AVDD.n1977 AVDD.n1976 0.189
R3849 AVDD.n2125 AVDD.n2124 0.189
R3850 AVDD.n2276 AVDD.n2275 0.189
R3851 AVDD.n2461 AVDD.n2460 0.189
R3852 AVDD.n2349 AVDD.n2348 0.189
R3853 AVDD.n2625 AVDD.n2624 0.189
R3854 AVDD.n2557 AVDD.n2556 0.189
R3855 AVDD.n2865 AVDD.n2864 0.189
R3856 AVDD.n2774 AVDD.n2773 0.189
R3857 AVDD.n3005 AVDD.n3004 0.189
R3858 AVDD.n2937 AVDD.n2936 0.189
R3859 AVDD.n3269 AVDD.n3268 0.189
R3860 AVDD.n3118 AVDD.n3117 0.189
R3861 AVDD.n3404 AVDD.n3403 0.189
R3862 AVDD.n3337 AVDD.n3336 0.189
R3863 AVDD.n5016 AVDD.n5015 0.189
R3864 AVDD.n4709 AVDD.n4708 0.189
R3865 AVDD.n4822 AVDD.n4821 0.189
R3866 AVDD.n4924 AVDD.n4923 0.189
R3867 AVDD.n4822 AVDD.n4809 0.189
R3868 AVDD.n4924 AVDD.n4911 0.189
R3869 AVDD.n4822 AVDD.n4819 0.189
R3870 AVDD.n4924 AVDD.n4921 0.189
R3871 AVDD.n4822 AVDD.n4811 0.189
R3872 AVDD.n4924 AVDD.n4913 0.189
R3873 AVDD.n4822 AVDD.n4817 0.189
R3874 AVDD.n4924 AVDD.n4919 0.189
R3875 AVDD.n4822 AVDD.n4813 0.189
R3876 AVDD.n4924 AVDD.n4915 0.189
R3877 AVDD.n3706 AVDD.n3705 0.189
R3878 AVDD.n630 AVDD.n627 0.189
R3879 AVDD.n811 AVDD.n808 0.189
R3880 AVDD.n882 AVDD.n879 0.189
R3881 AVDD.n992 AVDD.n989 0.189
R3882 AVDD.n1058 AVDD.n1055 0.189
R3883 AVDD.n1295 AVDD.n1292 0.189
R3884 AVDD.n1163 AVDD.n1160 0.189
R3885 AVDD.n1260 AVDD.n1257 0.189
R3886 AVDD.n1421 AVDD.n1418 0.189
R3887 AVDD.n1535 AVDD.n1532 0.189
R3888 AVDD.n1625 AVDD.n1622 0.189
R3889 AVDD.n1744 AVDD.n1741 0.189
R3890 AVDD.n1834 AVDD.n1831 0.189
R3891 AVDD.n1977 AVDD.n1974 0.189
R3892 AVDD.n2046 AVDD.n2043 0.189
R3893 AVDD.n2276 AVDD.n2273 0.189
R3894 AVDD.n2125 AVDD.n2122 0.189
R3895 AVDD.n2349 AVDD.n2346 0.189
R3896 AVDD.n2461 AVDD.n2458 0.189
R3897 AVDD.n2557 AVDD.n2554 0.189
R3898 AVDD.n2625 AVDD.n2622 0.189
R3899 AVDD.n630 AVDD.n623 0.189
R3900 AVDD.n811 AVDD.n804 0.189
R3901 AVDD.n882 AVDD.n875 0.189
R3902 AVDD.n992 AVDD.n985 0.189
R3903 AVDD.n1058 AVDD.n1051 0.189
R3904 AVDD.n1295 AVDD.n1288 0.189
R3905 AVDD.n1163 AVDD.n1156 0.189
R3906 AVDD.n1260 AVDD.n1253 0.189
R3907 AVDD.n1421 AVDD.n1414 0.189
R3908 AVDD.n1535 AVDD.n1528 0.189
R3909 AVDD.n1625 AVDD.n1618 0.189
R3910 AVDD.n1744 AVDD.n1737 0.189
R3911 AVDD.n1834 AVDD.n1827 0.189
R3912 AVDD.n1977 AVDD.n1970 0.189
R3913 AVDD.n2046 AVDD.n2039 0.189
R3914 AVDD.n2276 AVDD.n2269 0.189
R3915 AVDD.n2125 AVDD.n2118 0.189
R3916 AVDD.n2349 AVDD.n2342 0.189
R3917 AVDD.n2461 AVDD.n2454 0.189
R3918 AVDD.n2557 AVDD.n2550 0.189
R3919 AVDD.n2625 AVDD.n2618 0.189
R3920 AVDD.n2774 AVDD.n2767 0.189
R3921 AVDD.n2865 AVDD.n2858 0.189
R3922 AVDD.n2937 AVDD.n2930 0.189
R3923 AVDD.n3005 AVDD.n2998 0.189
R3924 AVDD.n3118 AVDD.n3111 0.189
R3925 AVDD.n3269 AVDD.n3262 0.189
R3926 AVDD.n3337 AVDD.n3330 0.189
R3927 AVDD.n3404 AVDD.n3397 0.189
R3928 AVDD.n4709 AVDD.n4702 0.189
R3929 AVDD.n5016 AVDD.n5009 0.189
R3930 AVDD.n4924 AVDD.n4917 0.189
R3931 AVDD.n5018 AVDD.n5017 0.189
R3932 AVDD.n5017 AVDD.n5016 0.189
R3933 AVDD.n3338 AVDD.n3337 0.189
R3934 AVDD.n3406 AVDD.n3405 0.189
R3935 AVDD.n3405 AVDD.n3404 0.189
R3936 AVDD.n3120 AVDD.n3119 0.189
R3937 AVDD.n3119 AVDD.n3118 0.189
R3938 AVDD.n3270 AVDD.n3269 0.189
R3939 AVDD.n2939 AVDD.n2938 0.189
R3940 AVDD.n2938 AVDD.n2937 0.189
R3941 AVDD.n3007 AVDD.n3006 0.189
R3942 AVDD.n3006 AVDD.n3005 0.189
R3943 AVDD.n2776 AVDD.n2775 0.189
R3944 AVDD.n2775 AVDD.n2774 0.189
R3945 AVDD.n2867 AVDD.n2866 0.189
R3946 AVDD.n2866 AVDD.n2865 0.189
R3947 AVDD.n2559 AVDD.n2558 0.189
R3948 AVDD.n2558 AVDD.n2557 0.189
R3949 AVDD.n2627 AVDD.n2626 0.189
R3950 AVDD.n2626 AVDD.n2625 0.189
R3951 AVDD.n2351 AVDD.n2350 0.189
R3952 AVDD.n2350 AVDD.n2349 0.189
R3953 AVDD.n2463 AVDD.n2462 0.189
R3954 AVDD.n2462 AVDD.n2461 0.189
R3955 AVDD.n2277 AVDD.n2276 0.189
R3956 AVDD.n2127 AVDD.n2126 0.189
R3957 AVDD.n2126 AVDD.n2125 0.189
R3958 AVDD.n1979 AVDD.n1978 0.189
R3959 AVDD.n1978 AVDD.n1977 0.189
R3960 AVDD.n2047 AVDD.n2046 0.189
R3961 AVDD.n1746 AVDD.n1745 0.189
R3962 AVDD.n1745 AVDD.n1744 0.189
R3963 AVDD.n1836 AVDD.n1835 0.189
R3964 AVDD.n1835 AVDD.n1834 0.189
R3965 AVDD.n1537 AVDD.n1536 0.189
R3966 AVDD.n1536 AVDD.n1535 0.189
R3967 AVDD.n1627 AVDD.n1626 0.189
R3968 AVDD.n1626 AVDD.n1625 0.189
R3969 AVDD.n1262 AVDD.n1261 0.189
R3970 AVDD.n1261 AVDD.n1260 0.189
R3971 AVDD.n1423 AVDD.n1422 0.189
R3972 AVDD.n1422 AVDD.n1421 0.189
R3973 AVDD.n4700 AVDD.n4699 0.189
R3974 AVDD.n4709 AVDD.n4700 0.189
R3975 AVDD.n4823 AVDD.n4822 0.189
R3976 AVDD.n4925 AVDD.n4924 0.189
R3977 AVDD.n3650 AVDD.n3576 0.189
R3978 AVDD.n3640 AVDD.n3639 0.189
R3979 AVDD.n3650 AVDD.n3640 0.189
R3980 AVDD.n3575 AVDD.n3574 0.189
R3981 AVDD.n3650 AVDD.n3575 0.189
R3982 AVDD.n3643 AVDD.n3642 0.189
R3983 AVDD.n3650 AVDD.n3643 0.189
R3984 AVDD.n3572 AVDD.n3571 0.189
R3985 AVDD.n3650 AVDD.n3572 0.189
R3986 AVDD.n3646 AVDD.n3645 0.189
R3987 AVDD.n3650 AVDD.n3646 0.189
R3988 AVDD.n3569 AVDD.n3568 0.189
R3989 AVDD.n3650 AVDD.n3569 0.189
R3990 AVDD.n3649 AVDD.n3648 0.189
R3991 AVDD.n3650 AVDD.n3649 0.189
R3992 AVDD.n2278 AVDD.n2277 0.189
R3993 AVDD.n3339 AVDD.n3338 0.189
R3994 AVDD.n2048 AVDD.n2047 0.189
R3995 AVDD.n3271 AVDD.n3270 0.189
R3996 AVDD.n4356 AVDD.n4355 0.176
R3997 AVDD.t287 AVDD.n5858 0.175
R3998 AVDD.n689 AVDD.n688 0.164
R3999 AVDD.n1162 AVDD.n1161 0.159
R4000 AVDD.n1057 AVDD.n1056 0.159
R4001 AVDD.n881 AVDD.n880 0.159
R4002 AVDD.n691 AVDD.n690 0.159
R4003 AVDD.n695 AVDD.n694 0.159
R4004 AVDD.n697 AVDD.n696 0.159
R4005 AVDD.n501 AVDD.n500 0.159
R4006 AVDD.n313 AVDD.n312 0.159
R4007 AVDD.n6566 AVDD.n6565 0.159
R4008 AVDD.n685 AVDD.n684 0.159
R4009 AVDD.n693 AVDD.n692 0.159
R4010 AVDD.n683 AVDD.n682 0.159
R4011 AVDD.n681 AVDD.n680 0.159
R4012 AVDD.n5943 AVDD.n5942 0.159
R4013 AVDD.n305 AVDD.n304 0.159
R4014 AVDD.n493 AVDD.n492 0.159
R4015 AVDD.n5951 AVDD.n5950 0.159
R4016 AVDD.n487 AVDD.n486 0.159
R4017 AVDD.n299 AVDD.n298 0.159
R4018 AVDD.n489 AVDD.n488 0.159
R4019 AVDD.n301 AVDD.n300 0.159
R4020 AVDD.n497 AVDD.n496 0.159
R4021 AVDD.n309 AVDD.n308 0.159
R4022 AVDD.n6562 AVDD.n6561 0.159
R4023 AVDD.n5947 AVDD.n5946 0.159
R4024 AVDD.n491 AVDD.n490 0.159
R4025 AVDD.n303 AVDD.n302 0.159
R4026 AVDD.n6555 AVDD.n6554 0.159
R4027 AVDD.n5941 AVDD.n5940 0.159
R4028 AVDD.n5939 AVDD.n5938 0.159
R4029 AVDD.n6553 AVDD.n6552 0.159
R4030 AVDD.n5949 AVDD.n5948 0.159
R4031 AVDD.n6564 AVDD.n6563 0.159
R4032 AVDD.n311 AVDD.n310 0.159
R4033 AVDD.n499 AVDD.n498 0.159
R4034 AVDD.n5937 AVDD.n5936 0.159
R4035 AVDD.n6551 AVDD.n6550 0.159
R4036 AVDD.n6120 AVDD.n6119 0.159
R4037 AVDD.n6114 AVDD.n6113 0.159
R4038 AVDD.n6116 AVDD.n6115 0.159
R4039 AVDD.n5945 AVDD.n5944 0.159
R4040 AVDD.n6560 AVDD.n6559 0.159
R4041 AVDD.n307 AVDD.n306 0.159
R4042 AVDD.n495 AVDD.n494 0.159
R4043 AVDD.n873 AVDD.n872 0.159
R4044 AVDD.n1049 AVDD.n1048 0.159
R4045 AVDD.n1154 AVDD.n1153 0.159
R4046 AVDD.n4815 AVDD.n4814 0.159
R4047 AVDD.n5003 AVDD.n5002 0.159
R4048 AVDD.n3391 AVDD.n3390 0.159
R4049 AVDD.n3256 AVDD.n3255 0.159
R4050 AVDD.n2992 AVDD.n2991 0.159
R4051 AVDD.n2852 AVDD.n2851 0.159
R4052 AVDD.n2612 AVDD.n2611 0.159
R4053 AVDD.n2448 AVDD.n2447 0.159
R4054 AVDD.n2112 AVDD.n2111 0.159
R4055 AVDD.n2033 AVDD.n2032 0.159
R4056 AVDD.n1821 AVDD.n1820 0.159
R4057 AVDD.n1612 AVDD.n1611 0.159
R4058 AVDD.n1408 AVDD.n1407 0.159
R4059 AVDD.n1148 AVDD.n1147 0.159
R4060 AVDD.n1043 AVDD.n1042 0.159
R4061 AVDD.n867 AVDD.n866 0.159
R4062 AVDD.n5013 AVDD.n5012 0.159
R4063 AVDD.n3401 AVDD.n3400 0.159
R4064 AVDD.n3266 AVDD.n3265 0.159
R4065 AVDD.n3002 AVDD.n3001 0.159
R4066 AVDD.n2862 AVDD.n2861 0.159
R4067 AVDD.n5005 AVDD.n5004 0.159
R4068 AVDD.n3393 AVDD.n3392 0.159
R4069 AVDD.n3258 AVDD.n3257 0.159
R4070 AVDD.n2994 AVDD.n2993 0.159
R4071 AVDD.n2854 AVDD.n2853 0.159
R4072 AVDD.n2614 AVDD.n2613 0.159
R4073 AVDD.n2450 AVDD.n2449 0.159
R4074 AVDD.n2114 AVDD.n2113 0.159
R4075 AVDD.n2035 AVDD.n2034 0.159
R4076 AVDD.n1823 AVDD.n1822 0.159
R4077 AVDD.n1614 AVDD.n1613 0.159
R4078 AVDD.n1410 AVDD.n1409 0.159
R4079 AVDD.n1150 AVDD.n1149 0.159
R4080 AVDD.n1045 AVDD.n1044 0.159
R4081 AVDD.n869 AVDD.n868 0.159
R4082 AVDD.n5011 AVDD.n5010 0.159
R4083 AVDD.n3399 AVDD.n3398 0.159
R4084 AVDD.n3264 AVDD.n3263 0.159
R4085 AVDD.n3000 AVDD.n2999 0.159
R4086 AVDD.n2860 AVDD.n2859 0.159
R4087 AVDD.n2620 AVDD.n2619 0.159
R4088 AVDD.n2456 AVDD.n2455 0.159
R4089 AVDD.n2120 AVDD.n2119 0.159
R4090 AVDD.n2041 AVDD.n2040 0.159
R4091 AVDD.n1829 AVDD.n1828 0.159
R4092 AVDD.n1620 AVDD.n1619 0.159
R4093 AVDD.n1416 AVDD.n1415 0.159
R4094 AVDD.n1158 AVDD.n1157 0.159
R4095 AVDD.n1053 AVDD.n1052 0.159
R4096 AVDD.n877 AVDD.n876 0.159
R4097 AVDD.n5007 AVDD.n5006 0.159
R4098 AVDD.n3395 AVDD.n3394 0.159
R4099 AVDD.n3260 AVDD.n3259 0.159
R4100 AVDD.n2996 AVDD.n2995 0.159
R4101 AVDD.n2856 AVDD.n2855 0.159
R4102 AVDD.n2616 AVDD.n2615 0.159
R4103 AVDD.n2452 AVDD.n2451 0.159
R4104 AVDD.n2116 AVDD.n2115 0.159
R4105 AVDD.n2037 AVDD.n2036 0.159
R4106 AVDD.n1825 AVDD.n1824 0.159
R4107 AVDD.n1616 AVDD.n1615 0.159
R4108 AVDD.n1412 AVDD.n1411 0.159
R4109 AVDD.n1152 AVDD.n1151 0.159
R4110 AVDD.n1047 AVDD.n1046 0.159
R4111 AVDD.n871 AVDD.n870 0.159
R4112 AVDD.n1420 AVDD.n1419 0.159
R4113 AVDD.n1624 AVDD.n1623 0.159
R4114 AVDD.n1833 AVDD.n1832 0.159
R4115 AVDD.n2045 AVDD.n2044 0.159
R4116 AVDD.n2124 AVDD.n2123 0.159
R4117 AVDD.n2460 AVDD.n2459 0.159
R4118 AVDD.n2624 AVDD.n2623 0.159
R4119 AVDD.n2864 AVDD.n2863 0.159
R4120 AVDD.n3004 AVDD.n3003 0.159
R4121 AVDD.n3268 AVDD.n3267 0.159
R4122 AVDD.n3403 AVDD.n3402 0.159
R4123 AVDD.n5015 AVDD.n5014 0.159
R4124 AVDD.n4821 AVDD.n4820 0.159
R4125 AVDD.n4809 AVDD.n4808 0.159
R4126 AVDD.n4819 AVDD.n4818 0.159
R4127 AVDD.n4811 AVDD.n4810 0.159
R4128 AVDD.n4817 AVDD.n4816 0.159
R4129 AVDD.n4813 AVDD.n4812 0.159
R4130 AVDD.n879 AVDD.n878 0.159
R4131 AVDD.n1055 AVDD.n1054 0.159
R4132 AVDD.n1160 AVDD.n1159 0.159
R4133 AVDD.n1418 AVDD.n1417 0.159
R4134 AVDD.n1622 AVDD.n1621 0.159
R4135 AVDD.n1831 AVDD.n1830 0.159
R4136 AVDD.n2043 AVDD.n2042 0.159
R4137 AVDD.n2122 AVDD.n2121 0.159
R4138 AVDD.n2458 AVDD.n2457 0.159
R4139 AVDD.n2622 AVDD.n2621 0.159
R4140 AVDD.n875 AVDD.n874 0.159
R4141 AVDD.n1051 AVDD.n1050 0.159
R4142 AVDD.n1156 AVDD.n1155 0.159
R4143 AVDD.n1414 AVDD.n1413 0.159
R4144 AVDD.n1618 AVDD.n1617 0.159
R4145 AVDD.n1827 AVDD.n1826 0.159
R4146 AVDD.n2039 AVDD.n2038 0.159
R4147 AVDD.n2118 AVDD.n2117 0.159
R4148 AVDD.n2454 AVDD.n2453 0.159
R4149 AVDD.n2618 AVDD.n2617 0.159
R4150 AVDD.n2858 AVDD.n2857 0.159
R4151 AVDD.n2998 AVDD.n2997 0.159
R4152 AVDD.n3262 AVDD.n3261 0.159
R4153 AVDD.n3397 AVDD.n3396 0.159
R4154 AVDD.n5009 AVDD.n5008 0.159
R4155 AVDD.n4702 AVDD.n4701 0.159
R4156 AVDD.n3330 AVDD.n3329 0.159
R4157 AVDD.n3111 AVDD.n3110 0.159
R4158 AVDD.n2930 AVDD.n2929 0.159
R4159 AVDD.n2767 AVDD.n2766 0.159
R4160 AVDD.n2550 AVDD.n2549 0.159
R4161 AVDD.n2342 AVDD.n2341 0.159
R4162 AVDD.n2269 AVDD.n2268 0.159
R4163 AVDD.n1970 AVDD.n1969 0.159
R4164 AVDD.n1737 AVDD.n1736 0.159
R4165 AVDD.n1528 AVDD.n1527 0.159
R4166 AVDD.n1253 AVDD.n1252 0.159
R4167 AVDD.n1288 AVDD.n1287 0.159
R4168 AVDD.n985 AVDD.n984 0.159
R4169 AVDD.n804 AVDD.n803 0.159
R4170 AVDD.n2554 AVDD.n2553 0.159
R4171 AVDD.n2346 AVDD.n2345 0.159
R4172 AVDD.n2273 AVDD.n2272 0.159
R4173 AVDD.n1974 AVDD.n1973 0.159
R4174 AVDD.n1741 AVDD.n1740 0.159
R4175 AVDD.n1532 AVDD.n1531 0.159
R4176 AVDD.n1257 AVDD.n1256 0.159
R4177 AVDD.n1292 AVDD.n1291 0.159
R4178 AVDD.n989 AVDD.n988 0.159
R4179 AVDD.n808 AVDD.n807 0.159
R4180 AVDD.n1294 AVDD.n1293 0.159
R4181 AVDD.n991 AVDD.n990 0.159
R4182 AVDD.n810 AVDD.n809 0.159
R4183 AVDD.n751 AVDD.n750 0.159
R4184 AVDD.n932 AVDD.n931 0.159
R4185 AVDD.n1284 AVDD.n1283 0.159
R4186 AVDD.n1202 AVDD.n1201 0.159
R4187 AVDD.n1477 AVDD.n1476 0.159
R4188 AVDD.n1735 AVDD.n1734 0.159
R4189 AVDD.n1919 AVDD.n1918 0.159
R4190 AVDD.n2267 AVDD.n2266 0.159
R4191 AVDD.n2291 AVDD.n2290 0.159
R4192 AVDD.n2548 AVDD.n2547 0.159
R4193 AVDD.n2716 AVDD.n2715 0.159
R4194 AVDD.n2879 AVDD.n2878 0.159
R4195 AVDD.n3060 AVDD.n3059 0.159
R4196 AVDD.n3279 AVDD.n3278 0.159
R4197 AVDD.n4698 AVDD.n4697 0.159
R4198 AVDD.n806 AVDD.n805 0.159
R4199 AVDD.n987 AVDD.n986 0.159
R4200 AVDD.n1290 AVDD.n1289 0.159
R4201 AVDD.n1255 AVDD.n1254 0.159
R4202 AVDD.n1530 AVDD.n1529 0.159
R4203 AVDD.n1739 AVDD.n1738 0.159
R4204 AVDD.n1972 AVDD.n1971 0.159
R4205 AVDD.n2271 AVDD.n2270 0.159
R4206 AVDD.n2344 AVDD.n2343 0.159
R4207 AVDD.n2552 AVDD.n2551 0.159
R4208 AVDD.n2769 AVDD.n2768 0.159
R4209 AVDD.n2932 AVDD.n2931 0.159
R4210 AVDD.n3113 AVDD.n3112 0.159
R4211 AVDD.n3332 AVDD.n3331 0.159
R4212 AVDD.n4704 AVDD.n4703 0.159
R4213 AVDD.n749 AVDD.n748 0.159
R4214 AVDD.n930 AVDD.n929 0.159
R4215 AVDD.n1282 AVDD.n1281 0.159
R4216 AVDD.n1200 AVDD.n1199 0.159
R4217 AVDD.n1475 AVDD.n1474 0.159
R4218 AVDD.n1733 AVDD.n1732 0.159
R4219 AVDD.n1917 AVDD.n1916 0.159
R4220 AVDD.n2265 AVDD.n2264 0.159
R4221 AVDD.n2289 AVDD.n2288 0.159
R4222 AVDD.n2546 AVDD.n2545 0.159
R4223 AVDD.n2714 AVDD.n2713 0.159
R4224 AVDD.n2877 AVDD.n2876 0.159
R4225 AVDD.n3058 AVDD.n3057 0.159
R4226 AVDD.n3277 AVDD.n3276 0.159
R4227 AVDD.n4696 AVDD.n4695 0.159
R4228 AVDD.n2771 AVDD.n2770 0.159
R4229 AVDD.n2934 AVDD.n2933 0.159
R4230 AVDD.n3115 AVDD.n3114 0.159
R4231 AVDD.n3334 AVDD.n3333 0.159
R4232 AVDD.n4706 AVDD.n4705 0.159
R4233 AVDD.n747 AVDD.n746 0.159
R4234 AVDD.n928 AVDD.n927 0.159
R4235 AVDD.n1280 AVDD.n1279 0.159
R4236 AVDD.n1198 AVDD.n1197 0.159
R4237 AVDD.n1473 AVDD.n1472 0.159
R4238 AVDD.n1731 AVDD.n1730 0.159
R4239 AVDD.n1915 AVDD.n1914 0.159
R4240 AVDD.n2263 AVDD.n2262 0.159
R4241 AVDD.n2287 AVDD.n2286 0.159
R4242 AVDD.n2544 AVDD.n2543 0.159
R4243 AVDD.n2712 AVDD.n2711 0.159
R4244 AVDD.n2875 AVDD.n2874 0.159
R4245 AVDD.n3056 AVDD.n3055 0.159
R4246 AVDD.n3275 AVDD.n3274 0.159
R4247 AVDD.n4694 AVDD.n4693 0.159
R4248 AVDD.n1286 AVDD.n1285 0.159
R4249 AVDD.n934 AVDD.n933 0.159
R4250 AVDD.n753 AVDD.n752 0.159
R4251 AVDD.n426 AVDD.n425 0.159
R4252 AVDD.n241 AVDD.n240 0.159
R4253 AVDD.n125 AVDD.n124 0.159
R4254 AVDD.n6434 AVDD.n6433 0.159
R4255 AVDD.n68 AVDD.n67 0.159
R4256 AVDD.n6424 AVDD.n6423 0.159
R4257 AVDD.n627 AVDD.n626 0.159
R4258 AVDD.n430 AVDD.n429 0.159
R4259 AVDD.n245 AVDD.n244 0.159
R4260 AVDD.n129 AVDD.n128 0.159
R4261 AVDD.n6438 AVDD.n6437 0.159
R4262 AVDD.n70 AVDD.n69 0.159
R4263 AVDD.n6426 AVDD.n6425 0.159
R4264 AVDD.n629 AVDD.n628 0.159
R4265 AVDD.n432 AVDD.n431 0.159
R4266 AVDD.n247 AVDD.n246 0.159
R4267 AVDD.n131 AVDD.n130 0.159
R4268 AVDD.n6428 AVDD.n6427 0.159
R4269 AVDD.n72 AVDD.n71 0.159
R4270 AVDD.n188 AVDD.n187 0.159
R4271 AVDD.n366 AVDD.n365 0.159
R4272 AVDD.n6436 AVDD.n6435 0.159
R4273 AVDD.n127 AVDD.n126 0.159
R4274 AVDD.n243 AVDD.n242 0.159
R4275 AVDD.n428 AVDD.n427 0.159
R4276 AVDD.n186 AVDD.n185 0.159
R4277 AVDD.n364 AVDD.n363 0.159
R4278 AVDD.n184 AVDD.n183 0.159
R4279 AVDD.n362 AVDD.n361 0.159
R4280 AVDD.n5868 AVDD.n5867 0.159
R4281 AVDD.n190 AVDD.n189 0.159
R4282 AVDD.n6440 AVDD.n6439 0.159
R4283 AVDD.n5874 AVDD.n5873 0.159
R4284 AVDD.n5860 AVDD.n5859 0.159
R4285 AVDD.n5872 AVDD.n5871 0.159
R4286 AVDD.n5862 AVDD.n5861 0.159
R4287 AVDD.n5870 AVDD.n5869 0.159
R4288 AVDD.n5864 AVDD.n5863 0.159
R4289 AVDD.n5866 AVDD.n5865 0.159
R4290 AVDD.n558 AVDD.n557 0.159
R4291 AVDD.n552 AVDD.n551 0.159
R4292 AVDD.n554 AVDD.n553 0.159
R4293 AVDD.n625 AVDD.n624 0.159
R4294 AVDD.n556 AVDD.n555 0.159
R4295 AVDD.n1259 AVDD.n1258 0.159
R4296 AVDD.n1534 AVDD.n1533 0.159
R4297 AVDD.n1743 AVDD.n1742 0.159
R4298 AVDD.n1976 AVDD.n1975 0.159
R4299 AVDD.n2275 AVDD.n2274 0.159
R4300 AVDD.n2348 AVDD.n2347 0.159
R4301 AVDD.n2556 AVDD.n2555 0.159
R4302 AVDD.n2773 AVDD.n2772 0.159
R4303 AVDD.n2936 AVDD.n2935 0.159
R4304 AVDD.n3117 AVDD.n3116 0.159
R4305 AVDD.n3336 AVDD.n3335 0.159
R4306 AVDD.n4708 AVDD.n4707 0.159
R4307 AVDD.n4923 AVDD.n4922 0.159
R4308 AVDD.n4911 AVDD.n4910 0.159
R4309 AVDD.n4921 AVDD.n4920 0.159
R4310 AVDD.n4913 AVDD.n4912 0.159
R4311 AVDD.n4919 AVDD.n4918 0.159
R4312 AVDD.n4915 AVDD.n4914 0.159
R4313 AVDD.n623 AVDD.n622 0.159
R4314 AVDD.n4917 AVDD.n4916 0.159
R4315 AVDD.n4597 AVDD.n4596 0.154
R4316 AVDD.n4597 AVDD.n3707 0.154
R4317 AVDD.n4597 AVDD.n3735 0.154
R4318 AVDD.n4597 AVDD.n4442 0.154
R4319 AVDD.n4597 AVDD.n4518 0.154
R4320 AVDD.n4597 AVDD.n4546 0.154
R4321 AVDD.n4597 AVDD.n3495 0.154
R4322 AVDD.n507 AVDD.n506 0.153
R4323 AVDD.n5642 AVDD.n508 0.152
R4324 AVDD.n5650 AVDD.n146 0.152
R4325 AVDD.n5650 AVDD.n148 0.152
R4326 AVDD.n5642 AVDD.n326 0.152
R4327 AVDD.n5635 AVDD.n516 0.152
R4328 AVDD.n5628 AVDD.n711 0.152
R4329 AVDD.n5621 AVDD.n892 0.152
R4330 AVDD.n5608 AVDD.n1063 0.152
R4331 AVDD.n5597 AVDD.n5594 0.152
R4332 AVDD.n5546 AVDD.n5543 0.152
R4333 AVDD.n5501 AVDD.n5498 0.152
R4334 AVDD.n5450 AVDD.n5447 0.152
R4335 AVDD.n5397 AVDD.n5394 0.152
R4336 AVDD.n5353 AVDD.n5347 0.152
R4337 AVDD.n5248 AVDD.n5207 0.152
R4338 AVDD.n5248 AVDD.n5209 0.152
R4339 AVDD.n5200 AVDD.n5161 0.152
R4340 AVDD.n5149 AVDD.n5110 0.152
R4341 AVDD.n5098 AVDD.n5059 0.152
R4342 AVDD.n5047 AVDD.n3455 0.152
R4343 AVDD.n4825 AVDD.n3463 0.152
R4344 AVDD.n5650 AVDD.n322 0.152
R4345 AVDD.n5650 AVDD.n321 0.152
R4346 AVDD.n5642 AVDD.n512 0.152
R4347 AVDD.n5635 AVDD.n707 0.152
R4348 AVDD.n5628 AVDD.n888 0.152
R4349 AVDD.n5621 AVDD.n5614 0.152
R4350 AVDD.n5608 AVDD.n5601 0.152
R4351 AVDD.n5597 AVDD.n5556 0.152
R4352 AVDD.n5546 AVDD.n5505 0.152
R4353 AVDD.n5501 AVDD.n5460 0.152
R4354 AVDD.n5450 AVDD.n5406 0.152
R4355 AVDD.n5397 AVDD.n2284 0.152
R4356 AVDD.n5353 AVDD.n5310 0.152
R4357 AVDD.n5301 AVDD.n5259 0.152
R4358 AVDD.n5248 AVDD.n5206 0.152
R4359 AVDD.n5200 AVDD.n5159 0.152
R4360 AVDD.n5149 AVDD.n5108 0.152
R4361 AVDD.n5098 AVDD.n5057 0.152
R4362 AVDD.n5047 AVDD.n3453 0.152
R4363 AVDD.n4825 AVDD.n3462 0.152
R4364 AVDD.n5301 AVDD.n5300 0.152
R4365 AVDD.n5650 AVDD.n145 0.152
R4366 AVDD.n5650 AVDD.n144 0.152
R4367 AVDD.n5642 AVDD.n324 0.152
R4368 AVDD.n5635 AVDD.n514 0.152
R4369 AVDD.n5628 AVDD.n709 0.152
R4370 AVDD.n5621 AVDD.n890 0.152
R4371 AVDD.n5608 AVDD.n1061 0.152
R4372 AVDD.n5597 AVDD.n5596 0.152
R4373 AVDD.n5546 AVDD.n5545 0.152
R4374 AVDD.n5501 AVDD.n5500 0.152
R4375 AVDD.n5450 AVDD.n5449 0.152
R4376 AVDD.n5397 AVDD.n5396 0.152
R4377 AVDD.n5353 AVDD.n5352 0.152
R4378 AVDD.n5248 AVDD.n5247 0.152
R4379 AVDD.n5200 AVDD.n5199 0.152
R4380 AVDD.n5149 AVDD.n5148 0.152
R4381 AVDD.n5098 AVDD.n5097 0.152
R4382 AVDD.n5047 AVDD.n4905 0.152
R4383 AVDD.n4825 AVDD.n3456 0.152
R4384 AVDD.n4825 AVDD.n4692 0.152
R4385 AVDD.n5047 AVDD.n3447 0.152
R4386 AVDD.n5098 AVDD.n5051 0.152
R4387 AVDD.n5149 AVDD.n5102 0.152
R4388 AVDD.n5200 AVDD.n5153 0.152
R4389 AVDD.n5248 AVDD.n2872 0.152
R4390 AVDD.n5301 AVDD.n2671 0.152
R4391 AVDD.n5301 AVDD.n2672 0.152
R4392 AVDD.n5450 AVDD.n5400 0.152
R4393 AVDD.n5501 AVDD.n5454 0.152
R4394 AVDD.n5546 AVDD.n1654 0.152
R4395 AVDD.n5597 AVDD.n5550 0.152
R4396 AVDD.n5608 AVDD.n5607 0.152
R4397 AVDD.n5621 AVDD.n5620 0.152
R4398 AVDD.n5628 AVDD.n5627 0.152
R4399 AVDD.n5635 AVDD.n5634 0.152
R4400 AVDD.n5642 AVDD.n5641 0.152
R4401 AVDD.n5650 AVDD.n5649 0.152
R4402 AVDD.n5650 AVDD.n5647 0.152
R4403 AVDD.n2560 AVDD.n2559 0.151
R4404 AVDD.n5001 AVDD.n4930 0.151
R4405 AVDD.n4927 AVDD.n4909 0.147
R4406 AVDD.n5301 AVDD.n2669 0.147
R4407 AVDD.n5248 AVDD.n2870 0.147
R4408 AVDD.n5200 AVDD.n5151 0.147
R4409 AVDD.n5150 AVDD.n5149 0.147
R4410 AVDD.n5149 AVDD.n5100 0.147
R4411 AVDD.n5099 AVDD.n5098 0.147
R4412 AVDD.n5098 AVDD.n5049 0.147
R4413 AVDD.n5048 AVDD.n5047 0.147
R4414 AVDD.n5047 AVDD.n4929 0.147
R4415 AVDD.n4928 AVDD.n4927 0.147
R4416 AVDD.n5398 AVDD.n5397 0.147
R4417 AVDD.n5450 AVDD.n5399 0.147
R4418 AVDD.n5451 AVDD.n5450 0.147
R4419 AVDD.n5501 AVDD.n5452 0.147
R4420 AVDD.n5546 AVDD.n1652 0.147
R4421 AVDD.n5547 AVDD.n5546 0.147
R4422 AVDD.n5597 AVDD.n5548 0.147
R4423 AVDD.n5608 AVDD.n1165 0.147
R4424 AVDD.n5609 AVDD.n5608 0.147
R4425 AVDD.n5621 AVDD.n5610 0.147
R4426 AVDD.n5628 AVDD.n884 0.147
R4427 AVDD.n5635 AVDD.n703 0.147
R4428 AVDD.n5650 AVDD.n316 0.147
R4429 AVDD.n6358 AVDD.n5711 0.147
R4430 AVDD.n6358 AVDD.n5712 0.147
R4431 AVDD.n6359 AVDD.n5660 0.147
R4432 AVDD.n6359 AVDD.n5661 0.147
R4433 AVDD.n5657 AVDD.n5653 0.147
R4434 AVDD.n5657 AVDD.n5652 0.147
R4435 AVDD.n5651 AVDD.n5650 0.147
R4436 AVDD.n5650 AVDD.n5644 0.147
R4437 AVDD.n5643 AVDD.n5642 0.147
R4438 AVDD.n5642 AVDD.n5637 0.147
R4439 AVDD.n5636 AVDD.n5635 0.147
R4440 AVDD.n5635 AVDD.n5630 0.147
R4441 AVDD.n5629 AVDD.n5628 0.147
R4442 AVDD.n5628 AVDD.n5623 0.147
R4443 AVDD.n5622 AVDD.n5621 0.147
R4444 AVDD.n5621 AVDD.n5616 0.147
R4445 AVDD.n5608 AVDD.n5603 0.147
R4446 AVDD.n5597 AVDD.n5554 0.147
R4447 AVDD.n5546 AVDD.n5503 0.147
R4448 AVDD.n5502 AVDD.n5501 0.147
R4449 AVDD.n5501 AVDD.n5458 0.147
R4450 AVDD.n5450 AVDD.n5404 0.147
R4451 AVDD.n5397 AVDD.n2282 0.147
R4452 AVDD.n5353 AVDD.n5308 0.147
R4453 AVDD.n5248 AVDD.n5204 0.147
R4454 AVDD.n5200 AVDD.n5157 0.147
R4455 AVDD.n5149 AVDD.n5106 0.147
R4456 AVDD.n5098 AVDD.n5055 0.147
R4457 AVDD.n5047 AVDD.n3451 0.147
R4458 AVDD.n4825 AVDD.n3461 0.147
R4459 AVDD.n5302 AVDD.n5301 0.147
R4460 AVDD.n5301 AVDD.n5252 0.147
R4461 AVDD.n6358 AVDD.n6308 0.147
R4462 AVDD.n6358 AVDD.n6309 0.147
R4463 AVDD.n6359 AVDD.n5658 0.147
R4464 AVDD.n6359 AVDD.n5659 0.147
R4465 AVDD.n5657 AVDD.n5656 0.147
R4466 AVDD.n5657 AVDD.n5655 0.147
R4467 AVDD.n5650 AVDD.n5646 0.147
R4468 AVDD.n5642 AVDD.n5639 0.147
R4469 AVDD.n5635 AVDD.n5632 0.147
R4470 AVDD.n5628 AVDD.n5625 0.147
R4471 AVDD.n5621 AVDD.n5618 0.147
R4472 AVDD.n5608 AVDD.n5605 0.147
R4473 AVDD.n5597 AVDD.n5552 0.147
R4474 AVDD.n5546 AVDD.n1656 0.147
R4475 AVDD.n5501 AVDD.n5456 0.147
R4476 AVDD.n5450 AVDD.n5402 0.147
R4477 AVDD.n5397 AVDD.n2280 0.147
R4478 AVDD.n5353 AVDD.n5303 0.147
R4479 AVDD.n5249 AVDD.n5248 0.147
R4480 AVDD.n5248 AVDD.n5202 0.147
R4481 AVDD.n5201 AVDD.n5200 0.147
R4482 AVDD.n5200 AVDD.n5155 0.147
R4483 AVDD.n5149 AVDD.n5104 0.147
R4484 AVDD.n5098 AVDD.n5053 0.147
R4485 AVDD.n5047 AVDD.n3449 0.147
R4486 AVDD.n4825 AVDD.n4604 0.147
R4487 AVDD.n4825 AVDD.n4599 0.147
R4488 AVDD.n4826 AVDD.n4825 0.147
R4489 AVDD.n5047 AVDD.n4827 0.147
R4490 AVDD.n5098 AVDD.n5061 0.147
R4491 AVDD.n5149 AVDD.n5112 0.147
R4492 AVDD.n5200 AVDD.n5163 0.147
R4493 AVDD.n5248 AVDD.n5211 0.147
R4494 AVDD.n5301 AVDD.n5261 0.147
R4495 AVDD.n5353 AVDD.n5312 0.147
R4496 AVDD.n5354 AVDD.n5353 0.147
R4497 AVDD.n5450 AVDD.n5411 0.147
R4498 AVDD.n5501 AVDD.n5462 0.147
R4499 AVDD.n5546 AVDD.n5507 0.147
R4500 AVDD.n5597 AVDD.n5558 0.147
R4501 AVDD.n5598 AVDD.n5597 0.147
R4502 AVDD.n5608 AVDD.n5599 0.147
R4503 AVDD.n5621 AVDD.n5612 0.147
R4504 AVDD.n5628 AVDD.n886 0.147
R4505 AVDD.n5635 AVDD.n705 0.147
R4506 AVDD.n5642 AVDD.n510 0.147
R4507 AVDD.n5650 AVDD.n318 0.147
R4508 AVDD.n5650 AVDD.n319 0.147
R4509 AVDD.n5353 AVDD.n2468 0.146
R4510 AVDD.n5301 AVDD.n5257 0.146
R4511 AVDD.n5397 AVDD.n2059 0.144
R4512 AVDD.n5353 AVDD.n2464 0.141
R4513 AVDD.n3254 AVDD.n3166 0.141
R4514 AVDD.n5397 AVDD.n5358 0.139
R4515 AVDD.n5254 AVDD.n5253 0.136
R4516 AVDD.n2127 AVDD.n2061 0.136
R4517 AVDD.n5305 AVDD.n5304 0.131
R4518 AVDD.n2850 AVDD.n2779 0.131
R4519 AVDD.n6377 AVDD.n6369 0.13
R4520 AVDD.n6410 AVDD.n6378 0.126
R4521 AVDD.n2050 AVDD.n2049 0.119
R4522 AVDD.n6362 AVDD.n6359 0.117
R4523 AVDD.n6071 AVDD.n6069 0.116
R4524 AVDD.n5884 AVDD.n0 0.116
R4525 AVDD.n2058 AVDD.n2057 0.115
R4526 AVDD.n4483 AVDD.n4482 0.112
R4527 AVDD.n2470 AVDD.n2469 0.111
R4528 AVDD.n5251 AVDD.n5250 0.111
R4529 AVDD.n3901 level_shifter_up_1.VDD_HV 0.109
R4530 AVDD.n3967 level_shifter_up_2.VDD_HV 0.109
R4531 AVDD.n5408 AVDD.n5407 0.107
R4532 AVDD.n4116 AVDD 0.107
R4533 level_shifter_up_7.VDD_HV AVDD.n4174 0.107
R4534 AVDD.n508 AVDD.n507 0.104
R4535 AVDD.n5357 AVDD.n5356 0.103
R4536 AVDD.n2053 AVDD.n2052 0.102
R4537 AVDD.n6365 AVDD.n17 0.098
R4538 AVDD.n5297 AVDD.n5296 0.092
R4539 AVDD.n5047 AVDD.n5042 0.09
R4540 AVDD.n4315 AVDD.n4314 0.086
R4541 AVDD.n4314 AVDD.n4313 0.086
R4542 AVDD.n4311 AVDD.n4310 0.086
R4543 AVDD.n4267 AVDD.n4266 0.086
R4544 AVDD.n4223 AVDD.n4222 0.086
R4545 AVDD.n4228 AVDD.n4223 0.086
R4546 AVDD.n4228 AVDD.n4225 0.086
R4547 AVDD.n4228 AVDD.n4227 0.086
R4548 AVDD.n6366 AVDD.n6365 0.085
R4549 AVDD.n5349 AVDD.n5348 0.085
R4550 AVDD.n4312 AVDD.n4311 0.084
R4551 AVDD.n4411 AVDD.n4410 0.081
R4552 AVDD.n1267 AVDD.n1266 0.08
R4553 AVDD AVDD.n4413 0.079
R4554 AVDD.n5917 AVDD.n5916 0.079
R4555 AVDD.n4593 AVDD.n4592 0.074
R4556 AVDD.n4541 AVDD.n4540 0.074
R4557 AVDD.n4509 AVDD.n4508 0.074
R4558 AVDD.n3730 AVDD.n3729 0.074
R4559 AVDD.n3560 AVDD.n3559 0.074
R4560 AVDD.n3489 AVDD.n3488 0.074
R4561 AVDD.n4268 AVDD.n4267 0.073
R4562 AVDD.n4227 AVDD.n4226 0.073
R4563 AVDD.n4225 AVDD.n4224 0.072
R4564 AVDD.n3796 AVDD.t731 0.071
R4565 AVDD.t142 AVDD.n3887 0.071
R4566 AVDD.t262 AVDD.n3957 0.071
R4567 AVDD.t745 AVDD.n4102 0.071
R4568 AVDD.t765 AVDD.n4172 0.071
R4569 AVDD.n4554 AVDD.n4552 0.07
R4570 AVDD.n4526 AVDD.n4524 0.07
R4571 AVDD.n4450 AVDD.n4448 0.07
R4572 AVDD.n4422 AVDD.n4420 0.07
R4573 AVDD.n3715 AVDD.n3713 0.07
R4574 AVDD.n3545 AVDD.n3543 0.07
R4575 AVDD.n3485 AVDD.n3484 0.07
R4576 AVDD.n1729 AVDD.n1658 0.07
R4577 AVDD.n5828 AVDD.t52 0.07
R4578 AVDD.t275 AVDD.n6062 0.07
R4579 AVDD.t31 AVDD.n6419 0.07
R4580 AVDD.n5710 AVDD.n5709 0.07
R4581 AVDD.n6307 AVDD.n6306 0.07
R4582 AVDD.n4208 AVDD.n4197 0.063
R4583 AVDD.n4206 AVDD.n4205 0.063
R4584 AVDD.n3842 AVDD.n3840 0.063
R4585 AVDD.n3856 AVDD.n3848 0.063
R4586 AVDD.n3871 AVDD.n3862 0.063
R4587 AVDD.n3909 AVDD.n3907 0.063
R4588 AVDD.n3923 AVDD.n3915 0.063
R4589 AVDD.n3938 AVDD.n3929 0.063
R4590 AVDD.n3975 AVDD.n3973 0.063
R4591 AVDD.n3808 AVDD.n3806 0.063
R4592 AVDD.n4057 AVDD.n4055 0.063
R4593 AVDD.n4071 AVDD.n4063 0.063
R4594 AVDD.n4086 AVDD.n4077 0.063
R4595 AVDD.n4124 AVDD.n4122 0.063
R4596 AVDD.n4138 AVDD.n4130 0.063
R4597 AVDD.n4153 AVDD.n4144 0.063
R4598 AVDD.n4308 AVDD.n4307 0.063
R4599 AVDD.n4307 AVDD.n4306 0.063
R4600 AVDD.n4324 AVDD.n4323 0.063
R4601 AVDD.n4323 AVDD.n4322 0.063
R4602 AVDD.n4205 AVDD.n4204 0.063
R4603 AVDD.n4197 AVDD.n4196 0.063
R4604 AVDD.n2261 AVDD.n2259 0.06
R4605 AVDD.n3749 AVDD.n3746 0.06
R4606 AVDD.n3777 AVDD.n3769 0.06
R4607 AVDD.n3766 AVDD.n3764 0.06
R4608 AVDD.n5845 AVDD.n5843 0.06
R4609 AVDD.n6083 AVDD.n6082 0.06
R4610 AVDD.n6079 AVDD.n6077 0.06
R4611 AVDD.n6057 AVDD.n5932 0.06
R4612 AVDD.n5926 AVDD.n5912 0.06
R4613 AVDD.n5910 AVDD.n5907 0.06
R4614 AVDD.t739 level_shifter_up_6.VDD_HV 0.059
R4615 AVDD.n4195 AVDD.n4190 0.059
R4616 AVDD.n1277 AVDD.n1276 0.059
R4617 AVDD.n1278 AVDD.n1277 0.059
R4618 AVDD.n864 AVDD.n863 0.059
R4619 AVDD.n865 AVDD.n864 0.059
R4620 AVDD.n862 AVDD.n861 0.059
R4621 AVDD.n865 AVDD.n862 0.059
R4622 AVDD.n1272 AVDD.n1271 0.059
R4623 AVDD.n1278 AVDD.n1272 0.059
R4624 AVDD.n567 AVDD.n566 0.059
R4625 AVDD.n560 AVDD.n559 0.059
R4626 AVDD.n1270 AVDD.n1269 0.059
R4627 AVDD.n4597 AVDD.n4433 0.059
R4628 AVDD.n4195 AVDD.n4194 0.054
R4629 AVDD.n5044 AVDD.n5043 0.053
R4630 AVDD.n2542 AVDD.n2471 0.05
R4631 AVDD.n4220 AVDD.n4195 0.048
R4632 AVDD.t731 AVDD.n3791 0.047
R4633 AVDD.t142 AVDD.n3830 0.047
R4634 AVDD.t262 AVDD.n3958 0.047
R4635 AVDD.n4412 AVDD.n3981 0.047
R4636 AVDD.t745 AVDD.n4045 0.047
R4637 AVDD.t765 AVDD.n4175 0.047
R4638 AVDD.n5702 AVDD.n5701 0.047
R4639 AVDD.n6303 AVDD.n6294 0.047
R4640 AVDD.n4218 AVDD.n4216 0.043
R4641 AVDD.t52 level_shifter_up_5.VDD_HV 0.043
R4642 level_shifter_up_0.VDD_HV AVDD.t275 0.043
R4643 level_shifter_up_4.VDD_HV AVDD.t31 0.043
R4644 AVDD.n3500 AVDD.n3499 0.043
R4645 AVDD.n3536 AVDD.n3535 0.043
R4646 AVDD.n3848 AVDD.n3842 0.042
R4647 AVDD.n3862 AVDD.n3859 0.042
R4648 AVDD.n3915 AVDD.n3909 0.042
R4649 AVDD.n3929 AVDD.n3926 0.042
R4650 AVDD.n3981 AVDD.n3975 0.042
R4651 AVDD.n3811 AVDD.n3808 0.042
R4652 AVDD.n4063 AVDD.n4057 0.042
R4653 AVDD.n4077 AVDD.n4074 0.042
R4654 AVDD.n4130 AVDD.n4124 0.042
R4655 AVDD.n4144 AVDD.n4141 0.042
R4656 AVDD.n4543 AVDD.n4542 0.042
R4657 AVDD.n4511 AVDD.n4510 0.042
R4658 AVDD.n4435 AVDD.n4434 0.042
R4659 AVDD.n3732 AVDD.n3731 0.042
R4660 AVDD.n3562 AVDD.n3561 0.042
R4661 AVDD.n3491 AVDD.n3490 0.042
R4662 AVDD.n3834 AVDD.n3833 0.041
R4663 AVDD.n4049 AVDD.n4048 0.041
R4664 AVDD.n4433 AVDD.n4432 0.04
R4665 AVDD.n3787 AVDD.n3782 0.04
R4666 AVDD.n3882 AVDD.n3877 0.04
R4667 AVDD.n3951 AVDD.n3944 0.04
R4668 AVDD.n4097 AVDD.n4092 0.04
R4669 AVDD.n4398 AVDD.n4034 0.04
R4670 AVDD.n4166 AVDD.n4159 0.04
R4671 AVDD.n3751 AVDD.n3749 0.04
R4672 AVDD.n3769 AVDD.n3766 0.04
R4673 AVDD.n3753 AVDD.n3752 0.04
R4674 AVDD.n5820 AVDD.n5812 0.04
R4675 AVDD.n5848 AVDD.n5845 0.04
R4676 AVDD.n6082 AVDD.n6079 0.04
R4677 AVDD.n5879 AVDD.n5857 0.04
R4678 AVDD.n5932 AVDD.n5930 0.04
R4679 AVDD.n5912 AVDD.n5910 0.04
R4680 AVDD.n6414 AVDD.n10 0.04
R4681 AVDD.n5701 AVDD.n5700 0.04
R4682 AVDD.n3840 AVDD.n3834 0.039
R4683 AVDD.n3857 AVDD.n3856 0.039
R4684 AVDD.n3907 AVDD.n3902 0.039
R4685 AVDD.n3924 AVDD.n3923 0.039
R4686 AVDD.n3973 AVDD.n3968 0.039
R4687 AVDD.n3823 AVDD.n3812 0.039
R4688 AVDD.n4055 AVDD.n4049 0.039
R4689 AVDD.n4072 AVDD.n4071 0.039
R4690 AVDD.n4122 AVDD.n4117 0.039
R4691 AVDD.n4139 AVDD.n4138 0.039
R4692 AVDD.n4190 AVDD.n4038 0.039
R4693 AVDD.n3872 AVDD.n3871 0.038
R4694 AVDD.n3939 AVDD.n3938 0.038
R4695 AVDD.n3806 AVDD.n3800 0.038
R4696 AVDD.n4087 AVDD.n4086 0.038
R4697 AVDD.n4154 AVDD.n4153 0.038
R4698 AVDD.n4216 AVDD.n4214 0.037
R4699 AVDD.n3778 AVDD.n3777 0.037
R4700 AVDD.n3764 AVDD.n3753 0.037
R4701 AVDD.n6083 AVDD.n5849 0.037
R4702 AVDD.n6077 AVDD.n6072 0.037
R4703 AVDD.n5927 AVDD.n5926 0.037
R4704 AVDD.n5907 AVDD.n5885 0.037
R4705 AVDD.n4254 AVDD.n4244 0.036
R4706 AVDD.n3746 AVDD.n3737 0.036
R4707 AVDD.n5843 AVDD.n5832 0.036
R4708 AVDD.n6058 AVDD.n6057 0.036
R4709 level_shifter_up_6.VDD_HV AVDD.n4391 0.035
R4710 AVDD.n4498 AVDD.n4495 0.034
R4711 AVDD.n4498 AVDD.n4497 0.034
R4712 AVDD.n3486 AVDD.n3485 0.034
R4713 AVDD.n4591 AVDD.n4554 0.034
R4714 AVDD.n4539 AVDD.n4526 0.034
R4715 AVDD.n4507 AVDD.n4450 0.034
R4716 AVDD.n4431 AVDD.n4422 0.034
R4717 AVDD.n3728 AVDD.n3715 0.034
R4718 AVDD.n3558 AVDD.n3545 0.034
R4719 AVDD.n3488 AVDD.n3486 0.034
R4720 AVDD.n4592 AVDD.n4591 0.034
R4721 AVDD.n4540 AVDD.n4539 0.034
R4722 AVDD.n4508 AVDD.n4507 0.034
R4723 AVDD.n4432 AVDD.n4431 0.034
R4724 AVDD.n3729 AVDD.n3728 0.034
R4725 AVDD.n3559 AVDD.n3558 0.034
R4726 AVDD.n15 AVDD.n14 0.031
R4727 AVDD.n1355 AVDD.n1354 0.03
R4728 AVDD.n571 AVDD.n570 0.03
R4729 AVDD.n564 AVDD.n563 0.03
R4730 AVDD.n1348 AVDD.n1347 0.03
R4731 AVDD.n1354 AVDD.n1353 0.03
R4732 AVDD.n1347 AVDD.n1346 0.03
R4733 AVDD.n563 AVDD.n562 0.03
R4734 AVDD.n570 AVDD.n569 0.03
R4735 AVDD.n6368 AVDD.n6366 0.028
R4736 AVDD.n6378 AVDD.n15 0.026
R4737 AVDD.n688 AVDD.n687 0.026
R4738 AVDD.n3859 AVDD.n3857 0.024
R4739 AVDD.n3874 AVDD.n3872 0.024
R4740 AVDD.n3902 AVDD.n3901 0.024
R4741 AVDD.n3926 AVDD.n3924 0.024
R4742 AVDD.n3941 AVDD.n3939 0.024
R4743 AVDD.n3968 AVDD.n3967 0.024
R4744 AVDD.n3812 AVDD.n3811 0.024
R4745 AVDD.n3800 AVDD.n3799 0.024
R4746 AVDD.n4074 AVDD.n4072 0.024
R4747 AVDD.n4089 AVDD.n4087 0.024
R4748 AVDD.n4117 AVDD.n4116 0.024
R4749 AVDD.n4141 AVDD.n4139 0.024
R4750 AVDD.n4156 AVDD.n4154 0.024
R4751 AVDD.n4244 AVDD.n4242 0.024
R4752 AVDD.n4174 AVDD.n4038 0.024
R4753 AVDD.n3737 AVDD.n7 0.023
R4754 AVDD.n5832 AVDD.n5831 0.023
R4755 AVDD.n5849 AVDD.n5848 0.023
R4756 AVDD.n6072 AVDD.n6071 0.023
R4757 AVDD.n6060 AVDD.n6058 0.023
R4758 AVDD.n5930 AVDD.n5927 0.023
R4759 AVDD.n5885 AVDD.n5884 0.023
R4760 AVDD.n4239 AVDD.n4238 0.022
R4761 AVDD.n4255 AVDD.n4254 0.021
R4762 AVDD.n3836 AVDD.n3835 0.018
R4763 AVDD.t181 AVDD.n3836 0.018
R4764 AVDD.n3853 AVDD.n3852 0.018
R4765 AVDD.t767 AVDD.n3853 0.018
R4766 AVDD.n3868 AVDD.n3867 0.018
R4767 AVDD.t833 AVDD.n3868 0.018
R4768 AVDD.n3904 AVDD.n3903 0.018
R4769 AVDD.t144 AVDD.n3904 0.018
R4770 AVDD.n3970 AVDD.n3969 0.018
R4771 AVDD.t0 AVDD.n3970 0.018
R4772 AVDD.n3819 AVDD.n3818 0.018
R4773 AVDD.t763 AVDD.n3819 0.018
R4774 AVDD.n3803 AVDD.n3802 0.018
R4775 AVDD.t190 AVDD.n3803 0.018
R4776 AVDD.n3935 AVDD.n3934 0.018
R4777 AVDD.t729 AVDD.n3935 0.018
R4778 AVDD.n3920 AVDD.n3919 0.018
R4779 AVDD.t707 AVDD.n3920 0.018
R4780 AVDD.n4187 AVDD.n4186 0.018
R4781 AVDD.t749 AVDD.n4187 0.018
R4782 AVDD.n4234 AVDD.n4233 0.018
R4783 AVDD.t339 AVDD.n4234 0.018
R4784 AVDD.n4251 AVDD.n4250 0.018
R4785 AVDD.t806 AVDD.n4251 0.018
R4786 AVDD.n4051 AVDD.n4050 0.018
R4787 AVDD.t29 AVDD.n4051 0.018
R4788 AVDD.n4068 AVDD.n4067 0.018
R4789 AVDD.t719 AVDD.n4068 0.018
R4790 AVDD.n4083 AVDD.n4082 0.018
R4791 AVDD.t40 AVDD.n4083 0.018
R4792 AVDD.n4119 AVDD.n4118 0.018
R4793 AVDD.t215 AVDD.n4119 0.018
R4794 AVDD.n4150 AVDD.n4149 0.018
R4795 AVDD.t54 AVDD.n4150 0.018
R4796 AVDD.n4135 AVDD.n4134 0.018
R4797 AVDD.t270 AVDD.n4135 0.018
R4798 AVDD.t723 AVDD.n3774 0.018
R4799 AVDD.t838 AVDD.n3743 0.018
R4800 AVDD.n3760 AVDD.n3759 0.018
R4801 AVDD.n3774 AVDD.n3773 0.018
R4802 AVDD.n3743 AVDD.n3742 0.018
R4803 AVDD.t264 AVDD.n5904 0.018
R4804 AVDD.t818 AVDD.n5923 0.018
R4805 AVDD.t95 AVDD.n6054 0.018
R4806 AVDD.n5904 AVDD.n5903 0.018
R4807 AVDD.n5923 AVDD.n5922 0.018
R4808 AVDD.n6054 AVDD.n6053 0.018
R4809 AVDD.t266 AVDD.n6074 0.018
R4810 AVDD.t353 AVDD.n5807 0.018
R4811 AVDD.t341 AVDD.n5840 0.018
R4812 AVDD.n6074 AVDD.n6073 0.018
R4813 AVDD.n5807 AVDD.n5806 0.018
R4814 AVDD.n5840 AVDD.n5839 0.018
R4815 AVDD.n3761 AVDD.n3760 0.018
R4816 AVDD.n3859 AVDD.n3858 0.017
R4817 AVDD.n3848 AVDD.n3847 0.017
R4818 AVDD.n3842 AVDD.n3841 0.017
R4819 AVDD.n3862 AVDD.n3861 0.017
R4820 AVDD.n3874 AVDD.n3873 0.017
R4821 AVDD.n3926 AVDD.n3925 0.017
R4822 AVDD.n3901 AVDD.n3900 0.017
R4823 AVDD.n3909 AVDD.n3908 0.017
R4824 AVDD.n3915 AVDD.n3914 0.017
R4825 AVDD.n3929 AVDD.n3928 0.017
R4826 AVDD.n3941 AVDD.n3940 0.017
R4827 AVDD.n3808 AVDD.n3807 0.017
R4828 AVDD.n3811 AVDD.n3810 0.017
R4829 AVDD.n3967 AVDD.n3966 0.017
R4830 AVDD.n3975 AVDD.n3974 0.017
R4831 AVDD.n3981 AVDD.n3980 0.017
R4832 AVDD.n3799 AVDD.n3798 0.017
R4833 AVDD.n4074 AVDD.n4073 0.017
R4834 AVDD.n4063 AVDD.n4062 0.017
R4835 AVDD.n4057 AVDD.n4056 0.017
R4836 AVDD.n4077 AVDD.n4076 0.017
R4837 AVDD.n4089 AVDD.n4088 0.017
R4838 AVDD.n4141 AVDD.n4140 0.017
R4839 AVDD.n4116 AVDD.n4115 0.017
R4840 AVDD.n4124 AVDD.n4123 0.017
R4841 AVDD.n4130 AVDD.n4129 0.017
R4842 AVDD.n4242 AVDD.n4241 0.017
R4843 AVDD.n4244 AVDD.n4243 0.017
R4844 AVDD.n4257 AVDD.n4256 0.017
R4845 AVDD.n4144 AVDD.n4143 0.017
R4846 AVDD.n4156 AVDD.n4155 0.017
R4847 AVDD.n4174 AVDD.n4173 0.017
R4848 AVDD.n4194 AVDD.n4192 0.017
R4849 AVDD.n4194 AVDD.n4193 0.017
R4850 AVDD.n3766 AVDD.n3765 0.017
R4851 AVDD.n3751 AVDD.n3750 0.017
R4852 AVDD.n3769 AVDD.n3768 0.017
R4853 AVDD.n3749 AVDD.n3748 0.017
R4854 AVDD.n7 AVDD.n6 0.017
R4855 AVDD.n5845 AVDD.n5844 0.017
R4856 AVDD.n5831 AVDD.n5830 0.017
R4857 AVDD.n6071 AVDD.n6070 0.017
R4858 AVDD.n6079 AVDD.n6078 0.017
R4859 AVDD.n5848 AVDD.n5847 0.017
R4860 AVDD.n6082 AVDD.n6081 0.017
R4861 AVDD.n5932 AVDD.n5931 0.017
R4862 AVDD.n6060 AVDD.n6059 0.017
R4863 AVDD.n5884 AVDD.n5883 0.017
R4864 AVDD.n5910 AVDD.n5909 0.017
R4865 AVDD.n5930 AVDD.n5929 0.017
R4866 AVDD.n5912 AVDD.n5911 0.017
R4867 AVDD.n3886 AVDD.n3874 0.015
R4868 AVDD.n3956 AVDD.n3941 0.015
R4869 AVDD.n4412 AVDD.n3823 0.015
R4870 AVDD.n3799 AVDD.n3797 0.015
R4871 AVDD.n4101 AVDD.n4089 0.015
R4872 AVDD.n4171 AVDD.n4156 0.015
R4873 AVDD.n6418 AVDD.n7 0.015
R4874 AVDD.n5831 AVDD.n5829 0.015
R4875 AVDD.n6061 AVDD.n6060 0.015
R4876 AVDD.n4257 AVDD.n4255 0.014
R4877 AVDD.n3779 AVDD.n3778 0.014
R4878 AVDD.n3895 AVDD.n3894 0.014
R4879 AVDD.n3896 AVDD.n3895 0.014
R4880 AVDD.n3961 AVDD.n3960 0.014
R4881 AVDD.n3962 AVDD.n3961 0.014
R4882 AVDD.n4383 AVDD.n4382 0.014
R4883 AVDD.n4384 AVDD.n4383 0.014
R4884 AVDD.n4110 AVDD.n4109 0.014
R4885 AVDD.n4111 AVDD.n4110 0.014
R4886 AVDD.n4178 AVDD.n4177 0.014
R4887 AVDD.n4179 AVDD.n4178 0.014
R4888 AVDD.n6402 AVDD.n6401 0.014
R4889 AVDD.n6403 AVDD.n6402 0.014
R4890 AVDD.n6314 AVDD.n6313 0.014
R4891 AVDD.n6315 AVDD.n6314 0.014
R4892 AVDD.n4242 AVDD.n4239 0.013
R4893 AVDD.n4030 AVDD.n4029 0.013
R4894 AVDD.n4031 AVDD.n4030 0.013
R4895 AVDD.n4247 AVDD.n4246 0.013
R4896 AVDD.n4248 AVDD.n4247 0.013
R4897 AVDD.n4181 AVDD.n4180 0.013
R4898 AVDD.n4182 AVDD.n4181 0.013
R4899 AVDD.n6510 AVDD.n6509 0.013
R4900 AVDD.n6549 AVDD.n6510 0.013
R4901 AVDD.n80 AVDD.n79 0.013
R4902 AVDD.n123 AVDD.n80 0.013
R4903 AVDD.n5958 AVDD.n5957 0.013
R4904 AVDD.n6001 AVDD.n5958 0.013
R4905 AVDD.n6447 AVDD.n6446 0.013
R4906 AVDD.n6490 AVDD.n6447 0.013
R4907 AVDD.n258 AVDD.n257 0.013
R4908 AVDD.n297 AVDD.n258 0.013
R4909 AVDD.n196 AVDD.n195 0.013
R4910 AVDD.n239 AVDD.n196 0.013
R4911 AVDD.n640 AVDD.n639 0.013
R4912 AVDD.n679 AVDD.n640 0.013
R4913 AVDD.n446 AVDD.n445 0.013
R4914 AVDD.n485 AVDD.n446 0.013
R4915 AVDD.n378 AVDD.n377 0.013
R4916 AVDD.n421 AVDD.n378 0.013
R4917 AVDD.n5784 AVDD.n5779 0.013
R4918 AVDD.n5784 AVDD.n5781 0.013
R4919 AVDD.n6142 AVDD.n6106 0.013
R4920 AVDD.n6106 AVDD.n6105 0.013
R4921 AVDD.n6142 AVDD.n6139 0.013
R4922 AVDD.n6139 AVDD.n6138 0.013
R4923 AVDD.n6186 AVDD.n6159 0.013
R4924 AVDD.n6186 AVDD.n6161 0.013
R4925 AVDD.n6208 AVDD.n6203 0.013
R4926 AVDD.n6208 AVDD.n6205 0.013
R4927 AVDD.n6231 AVDD.n6226 0.013
R4928 AVDD.n6231 AVDD.n6228 0.013
R4929 AVDD.n6254 AVDD.n6249 0.013
R4930 AVDD.n6254 AVDD.n6251 0.013
R4931 AVDD.n6277 AVDD.n6272 0.013
R4932 AVDD.n6277 AVDD.n6274 0.013
R4933 AVDD.n676 AVDD.n675 0.013
R4934 AVDD.n679 AVDD.n676 0.013
R4935 AVDD.n482 AVDD.n481 0.013
R4936 AVDD.n485 AVDD.n482 0.013
R4937 AVDD.n414 AVDD.n413 0.013
R4938 AVDD.n421 AVDD.n414 0.013
R4939 AVDD.n294 AVDD.n293 0.013
R4940 AVDD.n297 AVDD.n294 0.013
R4941 AVDD.n232 AVDD.n231 0.013
R4942 AVDD.n239 AVDD.n232 0.013
R4943 AVDD.n664 AVDD.n663 0.013
R4944 AVDD.n679 AVDD.n664 0.013
R4945 AVDD.n470 AVDD.n469 0.013
R4946 AVDD.n485 AVDD.n470 0.013
R4947 AVDD.n402 AVDD.n401 0.013
R4948 AVDD.n421 AVDD.n402 0.013
R4949 AVDD.n282 AVDD.n281 0.013
R4950 AVDD.n297 AVDD.n282 0.013
R4951 AVDD.n220 AVDD.n219 0.013
R4952 AVDD.n239 AVDD.n220 0.013
R4953 AVDD.n658 AVDD.n657 0.013
R4954 AVDD.n679 AVDD.n658 0.013
R4955 AVDD.n464 AVDD.n463 0.013
R4956 AVDD.n485 AVDD.n464 0.013
R4957 AVDD.n396 AVDD.n395 0.013
R4958 AVDD.n421 AVDD.n396 0.013
R4959 AVDD.n276 AVDD.n275 0.013
R4960 AVDD.n297 AVDD.n276 0.013
R4961 AVDD.n214 AVDD.n213 0.013
R4962 AVDD.n239 AVDD.n214 0.013
R4963 AVDD.n6528 AVDD.n6527 0.013
R4964 AVDD.n6549 AVDD.n6528 0.013
R4965 AVDD.n98 AVDD.n97 0.013
R4966 AVDD.n123 AVDD.n98 0.013
R4967 AVDD.n5976 AVDD.n5975 0.013
R4968 AVDD.n6001 AVDD.n5976 0.013
R4969 AVDD.n6465 AVDD.n6464 0.013
R4970 AVDD.n6490 AVDD.n6465 0.013
R4971 AVDD.n652 AVDD.n651 0.013
R4972 AVDD.n679 AVDD.n652 0.013
R4973 AVDD.n458 AVDD.n457 0.013
R4974 AVDD.n485 AVDD.n458 0.013
R4975 AVDD.n390 AVDD.n389 0.013
R4976 AVDD.n421 AVDD.n390 0.013
R4977 AVDD.n270 AVDD.n269 0.013
R4978 AVDD.n297 AVDD.n270 0.013
R4979 AVDD.n208 AVDD.n207 0.013
R4980 AVDD.n239 AVDD.n208 0.013
R4981 AVDD.n6522 AVDD.n6521 0.013
R4982 AVDD.n6549 AVDD.n6522 0.013
R4983 AVDD.n92 AVDD.n91 0.013
R4984 AVDD.n123 AVDD.n92 0.013
R4985 AVDD.n5970 AVDD.n5969 0.013
R4986 AVDD.n6001 AVDD.n5970 0.013
R4987 AVDD.n6459 AVDD.n6458 0.013
R4988 AVDD.n6490 AVDD.n6459 0.013
R4989 AVDD.n6489 AVDD.n6488 0.013
R4990 AVDD.n6490 AVDD.n6489 0.013
R4991 AVDD.n6504 AVDD.n6503 0.013
R4992 AVDD.n6549 AVDD.n6504 0.013
R4993 AVDD.n122 AVDD.n121 0.013
R4994 AVDD.n123 AVDD.n122 0.013
R4995 AVDD.n252 AVDD.n251 0.013
R4996 AVDD.n297 AVDD.n252 0.013
R4997 AVDD.n238 AVDD.n237 0.013
R4998 AVDD.n239 AVDD.n238 0.013
R4999 AVDD.n440 AVDD.n439 0.013
R5000 AVDD.n485 AVDD.n440 0.013
R5001 AVDD.n420 AVDD.n419 0.013
R5002 AVDD.n421 AVDD.n420 0.013
R5003 AVDD.n634 AVDD.n633 0.013
R5004 AVDD.n679 AVDD.n634 0.013
R5005 AVDD.n5982 AVDD.n5981 0.013
R5006 AVDD.n6001 AVDD.n5982 0.013
R5007 AVDD.n6471 AVDD.n6470 0.013
R5008 AVDD.n6490 AVDD.n6471 0.013
R5009 AVDD.n6534 AVDD.n6533 0.013
R5010 AVDD.n6549 AVDD.n6534 0.013
R5011 AVDD.n104 AVDD.n103 0.013
R5012 AVDD.n123 AVDD.n104 0.013
R5013 AVDD.n5988 AVDD.n5987 0.013
R5014 AVDD.n6001 AVDD.n5988 0.013
R5015 AVDD.n6477 AVDD.n6476 0.013
R5016 AVDD.n6490 AVDD.n6477 0.013
R5017 AVDD.n6540 AVDD.n6539 0.013
R5018 AVDD.n6549 AVDD.n6540 0.013
R5019 AVDD.n110 AVDD.n109 0.013
R5020 AVDD.n123 AVDD.n110 0.013
R5021 AVDD.n288 AVDD.n287 0.013
R5022 AVDD.n297 AVDD.n288 0.013
R5023 AVDD.n226 AVDD.n225 0.013
R5024 AVDD.n239 AVDD.n226 0.013
R5025 AVDD.n476 AVDD.n475 0.013
R5026 AVDD.n485 AVDD.n476 0.013
R5027 AVDD.n408 AVDD.n407 0.013
R5028 AVDD.n421 AVDD.n408 0.013
R5029 AVDD.n670 AVDD.n669 0.013
R5030 AVDD.n679 AVDD.n670 0.013
R5031 AVDD.n5994 AVDD.n5993 0.013
R5032 AVDD.n6001 AVDD.n5994 0.013
R5033 AVDD.n6483 AVDD.n6482 0.013
R5034 AVDD.n6490 AVDD.n6483 0.013
R5035 AVDD.n6546 AVDD.n6545 0.013
R5036 AVDD.n6549 AVDD.n6546 0.013
R5037 AVDD.n116 AVDD.n115 0.013
R5038 AVDD.n123 AVDD.n116 0.013
R5039 AVDD.n6000 AVDD.n5999 0.013
R5040 AVDD.n6001 AVDD.n6000 0.013
R5041 AVDD.n6050 AVDD.n6049 0.013
R5042 AVDD.n6051 AVDD.n6050 0.013
R5043 AVDD.n6277 AVDD.n6276 0.013
R5044 AVDD.n6044 AVDD.n6043 0.013
R5045 AVDD.n6051 AVDD.n6044 0.013
R5046 AVDD.n6254 AVDD.n6253 0.013
R5047 AVDD.n6038 AVDD.n6037 0.013
R5048 AVDD.n6051 AVDD.n6038 0.013
R5049 AVDD.n6231 AVDD.n6230 0.013
R5050 AVDD.n6032 AVDD.n6031 0.013
R5051 AVDD.n6051 AVDD.n6032 0.013
R5052 AVDD.n6208 AVDD.n6207 0.013
R5053 AVDD.n6026 AVDD.n6025 0.013
R5054 AVDD.n6051 AVDD.n6026 0.013
R5055 AVDD.n6186 AVDD.n6185 0.013
R5056 AVDD.n6185 AVDD.n6184 0.013
R5057 AVDD.n6020 AVDD.n6019 0.013
R5058 AVDD.n6051 AVDD.n6020 0.013
R5059 AVDD.n6142 AVDD.n6141 0.013
R5060 AVDD.n6014 AVDD.n6013 0.013
R5061 AVDD.n6051 AVDD.n6014 0.013
R5062 AVDD.n5784 AVDD.n5783 0.013
R5063 AVDD.n5767 AVDD.n5762 0.013
R5064 AVDD.n5767 AVDD.n5760 0.013
R5065 AVDD.n6008 AVDD.n6007 0.013
R5066 AVDD.n6051 AVDD.n6008 0.013
R5067 AVDD.n5767 AVDD.n5766 0.013
R5068 AVDD.n5964 AVDD.n5963 0.013
R5069 AVDD.n6001 AVDD.n5964 0.013
R5070 AVDD.n6453 AVDD.n6452 0.013
R5071 AVDD.n6490 AVDD.n6453 0.013
R5072 AVDD.n6516 AVDD.n6515 0.013
R5073 AVDD.n6549 AVDD.n6516 0.013
R5074 AVDD.n86 AVDD.n85 0.013
R5075 AVDD.n123 AVDD.n86 0.013
R5076 AVDD.n264 AVDD.n263 0.013
R5077 AVDD.n297 AVDD.n264 0.013
R5078 AVDD.n202 AVDD.n201 0.013
R5079 AVDD.n239 AVDD.n202 0.013
R5080 AVDD.n452 AVDD.n451 0.013
R5081 AVDD.n485 AVDD.n452 0.013
R5082 AVDD.n384 AVDD.n383 0.013
R5083 AVDD.n421 AVDD.n384 0.013
R5084 AVDD.n646 AVDD.n645 0.013
R5085 AVDD.n679 AVDD.n646 0.013
R5086 AVDD.n578 AVDD.n577 0.013
R5087 AVDD.n621 AVDD.n578 0.013
R5088 AVDD.n821 AVDD.n820 0.013
R5089 AVDD.n860 AVDD.n821 0.013
R5090 AVDD.n759 AVDD.n758 0.013
R5091 AVDD.n802 AVDD.n759 0.013
R5092 AVDD.n1002 AVDD.n1001 0.013
R5093 AVDD.n1041 AVDD.n1002 0.013
R5094 AVDD.n940 AVDD.n939 0.013
R5095 AVDD.n983 AVDD.n940 0.013
R5096 AVDD.n1107 AVDD.n1106 0.013
R5097 AVDD.n1146 AVDD.n1107 0.013
R5098 AVDD.n1301 AVDD.n1300 0.013
R5099 AVDD.n1344 AVDD.n1301 0.013
R5100 AVDD.n4976 AVDD.n4975 0.013
R5101 AVDD.n4979 AVDD.n4976 0.013
R5102 AVDD.n4751 AVDD.n4750 0.013
R5103 AVDD.n4758 AVDD.n4751 0.013
R5104 AVDD.n3386 AVDD.n3385 0.013
R5105 AVDD.n3389 AVDD.n3386 0.013
R5106 AVDD.n3321 AVDD.n3320 0.013
R5107 AVDD.n3328 AVDD.n3321 0.013
R5108 AVDD.n3212 AVDD.n3211 0.013
R5109 AVDD.n3215 AVDD.n3212 0.013
R5110 AVDD.n3102 AVDD.n3101 0.013
R5111 AVDD.n3109 AVDD.n3102 0.013
R5112 AVDD.n2987 AVDD.n2986 0.013
R5113 AVDD.n2990 AVDD.n2987 0.013
R5114 AVDD.n2921 AVDD.n2920 0.013
R5115 AVDD.n2928 AVDD.n2921 0.013
R5116 AVDD.n2825 AVDD.n2824 0.013
R5117 AVDD.n2828 AVDD.n2825 0.013
R5118 AVDD.n2758 AVDD.n2757 0.013
R5119 AVDD.n2765 AVDD.n2758 0.013
R5120 AVDD.n2607 AVDD.n2606 0.013
R5121 AVDD.n2610 AVDD.n2607 0.013
R5122 AVDD.n2513 AVDD.n2512 0.013
R5123 AVDD.n2520 AVDD.n2513 0.013
R5124 AVDD.n2443 AVDD.n2442 0.013
R5125 AVDD.n2446 AVDD.n2443 0.013
R5126 AVDD.n2333 AVDD.n2332 0.013
R5127 AVDD.n2340 AVDD.n2333 0.013
R5128 AVDD.n2107 AVDD.n2106 0.013
R5129 AVDD.n2110 AVDD.n2107 0.013
R5130 AVDD.n2232 AVDD.n2231 0.013
R5131 AVDD.n2239 AVDD.n2232 0.013
R5132 AVDD.n2028 AVDD.n2027 0.013
R5133 AVDD.n2031 AVDD.n2028 0.013
R5134 AVDD.n1961 AVDD.n1960 0.013
R5135 AVDD.n1968 AVDD.n1961 0.013
R5136 AVDD.n1816 AVDD.n1815 0.013
R5137 AVDD.n1819 AVDD.n1816 0.013
R5138 AVDD.n1700 AVDD.n1699 0.013
R5139 AVDD.n1707 AVDD.n1700 0.013
R5140 AVDD.n1607 AVDD.n1606 0.013
R5141 AVDD.n1610 AVDD.n1607 0.013
R5142 AVDD.n1519 AVDD.n1518 0.013
R5143 AVDD.n1526 AVDD.n1519 0.013
R5144 AVDD.n1403 AVDD.n1402 0.013
R5145 AVDD.n1406 AVDD.n1403 0.013
R5146 AVDD.n1244 AVDD.n1243 0.013
R5147 AVDD.n1251 AVDD.n1244 0.013
R5148 AVDD.n1143 AVDD.n1142 0.013
R5149 AVDD.n1146 AVDD.n1143 0.013
R5150 AVDD.n1337 AVDD.n1336 0.013
R5151 AVDD.n1344 AVDD.n1337 0.013
R5152 AVDD.n1038 AVDD.n1037 0.013
R5153 AVDD.n1041 AVDD.n1038 0.013
R5154 AVDD.n976 AVDD.n975 0.013
R5155 AVDD.n983 AVDD.n976 0.013
R5156 AVDD.n857 AVDD.n856 0.013
R5157 AVDD.n860 AVDD.n857 0.013
R5158 AVDD.n795 AVDD.n794 0.013
R5159 AVDD.n802 AVDD.n795 0.013
R5160 AVDD.n614 AVDD.n613 0.013
R5161 AVDD.n621 AVDD.n614 0.013
R5162 AVDD.n4970 AVDD.n4969 0.013
R5163 AVDD.n4979 AVDD.n4970 0.013
R5164 AVDD.n4745 AVDD.n4744 0.013
R5165 AVDD.n4758 AVDD.n4745 0.013
R5166 AVDD.n3380 AVDD.n3379 0.013
R5167 AVDD.n3389 AVDD.n3380 0.013
R5168 AVDD.n3315 AVDD.n3314 0.013
R5169 AVDD.n3328 AVDD.n3315 0.013
R5170 AVDD.n3206 AVDD.n3205 0.013
R5171 AVDD.n3215 AVDD.n3206 0.013
R5172 AVDD.n3096 AVDD.n3095 0.013
R5173 AVDD.n3109 AVDD.n3096 0.013
R5174 AVDD.n2981 AVDD.n2980 0.013
R5175 AVDD.n2990 AVDD.n2981 0.013
R5176 AVDD.n2915 AVDD.n2914 0.013
R5177 AVDD.n2928 AVDD.n2915 0.013
R5178 AVDD.n2819 AVDD.n2818 0.013
R5179 AVDD.n2828 AVDD.n2819 0.013
R5180 AVDD.n2752 AVDD.n2751 0.013
R5181 AVDD.n2765 AVDD.n2752 0.013
R5182 AVDD.n4964 AVDD.n4963 0.013
R5183 AVDD.n4979 AVDD.n4964 0.013
R5184 AVDD.n4739 AVDD.n4738 0.013
R5185 AVDD.n4758 AVDD.n4739 0.013
R5186 AVDD.n3374 AVDD.n3373 0.013
R5187 AVDD.n3389 AVDD.n3374 0.013
R5188 AVDD.n3309 AVDD.n3308 0.013
R5189 AVDD.n3328 AVDD.n3309 0.013
R5190 AVDD.n3200 AVDD.n3199 0.013
R5191 AVDD.n3215 AVDD.n3200 0.013
R5192 AVDD.n3090 AVDD.n3089 0.013
R5193 AVDD.n3109 AVDD.n3090 0.013
R5194 AVDD.n2975 AVDD.n2974 0.013
R5195 AVDD.n2990 AVDD.n2975 0.013
R5196 AVDD.n2909 AVDD.n2908 0.013
R5197 AVDD.n2928 AVDD.n2909 0.013
R5198 AVDD.n2813 AVDD.n2812 0.013
R5199 AVDD.n2828 AVDD.n2813 0.013
R5200 AVDD.n2746 AVDD.n2745 0.013
R5201 AVDD.n2765 AVDD.n2746 0.013
R5202 AVDD.n2595 AVDD.n2594 0.013
R5203 AVDD.n2610 AVDD.n2595 0.013
R5204 AVDD.n2501 AVDD.n2500 0.013
R5205 AVDD.n2520 AVDD.n2501 0.013
R5206 AVDD.n2431 AVDD.n2430 0.013
R5207 AVDD.n2446 AVDD.n2431 0.013
R5208 AVDD.n2321 AVDD.n2320 0.013
R5209 AVDD.n2340 AVDD.n2321 0.013
R5210 AVDD.n2095 AVDD.n2094 0.013
R5211 AVDD.n2110 AVDD.n2095 0.013
R5212 AVDD.n2220 AVDD.n2219 0.013
R5213 AVDD.n2239 AVDD.n2220 0.013
R5214 AVDD.n2016 AVDD.n2015 0.013
R5215 AVDD.n2031 AVDD.n2016 0.013
R5216 AVDD.n1949 AVDD.n1948 0.013
R5217 AVDD.n1968 AVDD.n1949 0.013
R5218 AVDD.n1804 AVDD.n1803 0.013
R5219 AVDD.n1819 AVDD.n1804 0.013
R5220 AVDD.n1688 AVDD.n1687 0.013
R5221 AVDD.n1707 AVDD.n1688 0.013
R5222 AVDD.n1595 AVDD.n1594 0.013
R5223 AVDD.n1610 AVDD.n1595 0.013
R5224 AVDD.n1507 AVDD.n1506 0.013
R5225 AVDD.n1526 AVDD.n1507 0.013
R5226 AVDD.n1391 AVDD.n1390 0.013
R5227 AVDD.n1406 AVDD.n1391 0.013
R5228 AVDD.n1232 AVDD.n1231 0.013
R5229 AVDD.n1251 AVDD.n1232 0.013
R5230 AVDD.n1131 AVDD.n1130 0.013
R5231 AVDD.n1146 AVDD.n1131 0.013
R5232 AVDD.n1325 AVDD.n1324 0.013
R5233 AVDD.n1344 AVDD.n1325 0.013
R5234 AVDD.n1026 AVDD.n1025 0.013
R5235 AVDD.n1041 AVDD.n1026 0.013
R5236 AVDD.n964 AVDD.n963 0.013
R5237 AVDD.n983 AVDD.n964 0.013
R5238 AVDD.n845 AVDD.n844 0.013
R5239 AVDD.n860 AVDD.n845 0.013
R5240 AVDD.n783 AVDD.n782 0.013
R5241 AVDD.n802 AVDD.n783 0.013
R5242 AVDD.n602 AVDD.n601 0.013
R5243 AVDD.n621 AVDD.n602 0.013
R5244 AVDD.n4958 AVDD.n4957 0.013
R5245 AVDD.n4979 AVDD.n4958 0.013
R5246 AVDD.n4733 AVDD.n4732 0.013
R5247 AVDD.n4758 AVDD.n4733 0.013
R5248 AVDD.n3368 AVDD.n3367 0.013
R5249 AVDD.n3389 AVDD.n3368 0.013
R5250 AVDD.n3303 AVDD.n3302 0.013
R5251 AVDD.n3328 AVDD.n3303 0.013
R5252 AVDD.n3194 AVDD.n3193 0.013
R5253 AVDD.n3215 AVDD.n3194 0.013
R5254 AVDD.n3084 AVDD.n3083 0.013
R5255 AVDD.n3109 AVDD.n3084 0.013
R5256 AVDD.n2969 AVDD.n2968 0.013
R5257 AVDD.n2990 AVDD.n2969 0.013
R5258 AVDD.n2903 AVDD.n2902 0.013
R5259 AVDD.n2928 AVDD.n2903 0.013
R5260 AVDD.n2807 AVDD.n2806 0.013
R5261 AVDD.n2828 AVDD.n2807 0.013
R5262 AVDD.n2740 AVDD.n2739 0.013
R5263 AVDD.n2765 AVDD.n2740 0.013
R5264 AVDD.n2589 AVDD.n2588 0.013
R5265 AVDD.n2610 AVDD.n2589 0.013
R5266 AVDD.n2495 AVDD.n2494 0.013
R5267 AVDD.n2520 AVDD.n2495 0.013
R5268 AVDD.n2425 AVDD.n2424 0.013
R5269 AVDD.n2446 AVDD.n2425 0.013
R5270 AVDD.n2315 AVDD.n2314 0.013
R5271 AVDD.n2340 AVDD.n2315 0.013
R5272 AVDD.n2089 AVDD.n2088 0.013
R5273 AVDD.n2110 AVDD.n2089 0.013
R5274 AVDD.n2214 AVDD.n2213 0.013
R5275 AVDD.n2239 AVDD.n2214 0.013
R5276 AVDD.n2010 AVDD.n2009 0.013
R5277 AVDD.n2031 AVDD.n2010 0.013
R5278 AVDD.n1943 AVDD.n1942 0.013
R5279 AVDD.n1968 AVDD.n1943 0.013
R5280 AVDD.n1798 AVDD.n1797 0.013
R5281 AVDD.n1819 AVDD.n1798 0.013
R5282 AVDD.n1682 AVDD.n1681 0.013
R5283 AVDD.n1707 AVDD.n1682 0.013
R5284 AVDD.n1589 AVDD.n1588 0.013
R5285 AVDD.n1610 AVDD.n1589 0.013
R5286 AVDD.n1501 AVDD.n1500 0.013
R5287 AVDD.n1526 AVDD.n1501 0.013
R5288 AVDD.n1385 AVDD.n1384 0.013
R5289 AVDD.n1406 AVDD.n1385 0.013
R5290 AVDD.n1226 AVDD.n1225 0.013
R5291 AVDD.n1251 AVDD.n1226 0.013
R5292 AVDD.n1125 AVDD.n1124 0.013
R5293 AVDD.n1146 AVDD.n1125 0.013
R5294 AVDD.n1319 AVDD.n1318 0.013
R5295 AVDD.n1344 AVDD.n1319 0.013
R5296 AVDD.n1020 AVDD.n1019 0.013
R5297 AVDD.n1041 AVDD.n1020 0.013
R5298 AVDD.n958 AVDD.n957 0.013
R5299 AVDD.n983 AVDD.n958 0.013
R5300 AVDD.n839 AVDD.n838 0.013
R5301 AVDD.n860 AVDD.n839 0.013
R5302 AVDD.n777 AVDD.n776 0.013
R5303 AVDD.n802 AVDD.n777 0.013
R5304 AVDD.n596 AVDD.n595 0.013
R5305 AVDD.n621 AVDD.n596 0.013
R5306 AVDD.n4952 AVDD.n4951 0.013
R5307 AVDD.n4979 AVDD.n4952 0.013
R5308 AVDD.n4727 AVDD.n4726 0.013
R5309 AVDD.n4758 AVDD.n4727 0.013
R5310 AVDD.n3362 AVDD.n3361 0.013
R5311 AVDD.n3389 AVDD.n3362 0.013
R5312 AVDD.n3297 AVDD.n3296 0.013
R5313 AVDD.n3328 AVDD.n3297 0.013
R5314 AVDD.n3188 AVDD.n3187 0.013
R5315 AVDD.n3215 AVDD.n3188 0.013
R5316 AVDD.n3078 AVDD.n3077 0.013
R5317 AVDD.n3109 AVDD.n3078 0.013
R5318 AVDD.n2963 AVDD.n2962 0.013
R5319 AVDD.n2990 AVDD.n2963 0.013
R5320 AVDD.n2897 AVDD.n2896 0.013
R5321 AVDD.n2928 AVDD.n2897 0.013
R5322 AVDD.n2801 AVDD.n2800 0.013
R5323 AVDD.n2828 AVDD.n2801 0.013
R5324 AVDD.n2734 AVDD.n2733 0.013
R5325 AVDD.n2765 AVDD.n2734 0.013
R5326 AVDD.n2583 AVDD.n2582 0.013
R5327 AVDD.n2610 AVDD.n2583 0.013
R5328 AVDD.n2489 AVDD.n2488 0.013
R5329 AVDD.n2520 AVDD.n2489 0.013
R5330 AVDD.n2419 AVDD.n2418 0.013
R5331 AVDD.n2446 AVDD.n2419 0.013
R5332 AVDD.n2309 AVDD.n2308 0.013
R5333 AVDD.n2340 AVDD.n2309 0.013
R5334 AVDD.n2083 AVDD.n2082 0.013
R5335 AVDD.n2110 AVDD.n2083 0.013
R5336 AVDD.n2208 AVDD.n2207 0.013
R5337 AVDD.n2239 AVDD.n2208 0.013
R5338 AVDD.n2004 AVDD.n2003 0.013
R5339 AVDD.n2031 AVDD.n2004 0.013
R5340 AVDD.n1937 AVDD.n1936 0.013
R5341 AVDD.n1968 AVDD.n1937 0.013
R5342 AVDD.n1792 AVDD.n1791 0.013
R5343 AVDD.n1819 AVDD.n1792 0.013
R5344 AVDD.n1676 AVDD.n1675 0.013
R5345 AVDD.n1707 AVDD.n1676 0.013
R5346 AVDD.n1583 AVDD.n1582 0.013
R5347 AVDD.n1610 AVDD.n1583 0.013
R5348 AVDD.n1495 AVDD.n1494 0.013
R5349 AVDD.n1526 AVDD.n1495 0.013
R5350 AVDD.n1379 AVDD.n1378 0.013
R5351 AVDD.n1406 AVDD.n1379 0.013
R5352 AVDD.n1220 AVDD.n1219 0.013
R5353 AVDD.n1251 AVDD.n1220 0.013
R5354 AVDD.n1119 AVDD.n1118 0.013
R5355 AVDD.n1146 AVDD.n1119 0.013
R5356 AVDD.n1313 AVDD.n1312 0.013
R5357 AVDD.n1344 AVDD.n1313 0.013
R5358 AVDD.n1014 AVDD.n1013 0.013
R5359 AVDD.n1041 AVDD.n1014 0.013
R5360 AVDD.n952 AVDD.n951 0.013
R5361 AVDD.n983 AVDD.n952 0.013
R5362 AVDD.n833 AVDD.n832 0.013
R5363 AVDD.n860 AVDD.n833 0.013
R5364 AVDD.n771 AVDD.n770 0.013
R5365 AVDD.n802 AVDD.n771 0.013
R5366 AVDD.n590 AVDD.n589 0.013
R5367 AVDD.n621 AVDD.n590 0.013
R5368 AVDD.n4770 AVDD.n4769 0.013
R5369 AVDD.n4807 AVDD.n4770 0.013
R5370 AVDD.n3637 AVDD.n3578 0.013
R5371 AVDD.n620 AVDD.n619 0.013
R5372 AVDD.n621 AVDD.n620 0.013
R5373 AVDD.n815 AVDD.n814 0.013
R5374 AVDD.n860 AVDD.n815 0.013
R5375 AVDD.n801 AVDD.n800 0.013
R5376 AVDD.n802 AVDD.n801 0.013
R5377 AVDD.n996 AVDD.n995 0.013
R5378 AVDD.n1041 AVDD.n996 0.013
R5379 AVDD.n982 AVDD.n981 0.013
R5380 AVDD.n983 AVDD.n982 0.013
R5381 AVDD.n1101 AVDD.n1100 0.013
R5382 AVDD.n1146 AVDD.n1101 0.013
R5383 AVDD.n1343 AVDD.n1342 0.013
R5384 AVDD.n1344 AVDD.n1343 0.013
R5385 AVDD.n1360 AVDD.n1359 0.013
R5386 AVDD.n1406 AVDD.n1360 0.013
R5387 AVDD.n1250 AVDD.n1249 0.013
R5388 AVDD.n1251 AVDD.n1250 0.013
R5389 AVDD.n1565 AVDD.n1564 0.013
R5390 AVDD.n1610 AVDD.n1565 0.013
R5391 AVDD.n1525 AVDD.n1524 0.013
R5392 AVDD.n1526 AVDD.n1525 0.013
R5393 AVDD.n1774 AVDD.n1773 0.013
R5394 AVDD.n1819 AVDD.n1774 0.013
R5395 AVDD.n1706 AVDD.n1705 0.013
R5396 AVDD.n1707 AVDD.n1706 0.013
R5397 AVDD.n1986 AVDD.n1985 0.013
R5398 AVDD.n2031 AVDD.n1986 0.013
R5399 AVDD.n1967 AVDD.n1966 0.013
R5400 AVDD.n1968 AVDD.n1967 0.013
R5401 AVDD.n2065 AVDD.n2064 0.013
R5402 AVDD.n2110 AVDD.n2065 0.013
R5403 AVDD.n2238 AVDD.n2237 0.013
R5404 AVDD.n2239 AVDD.n2238 0.013
R5405 AVDD.n2401 AVDD.n2400 0.013
R5406 AVDD.n2446 AVDD.n2401 0.013
R5407 AVDD.n2339 AVDD.n2338 0.013
R5408 AVDD.n2340 AVDD.n2339 0.013
R5409 AVDD.n2565 AVDD.n2564 0.013
R5410 AVDD.n2610 AVDD.n2565 0.013
R5411 AVDD.n2519 AVDD.n2518 0.013
R5412 AVDD.n2520 AVDD.n2519 0.013
R5413 AVDD.n2783 AVDD.n2782 0.013
R5414 AVDD.n2828 AVDD.n2783 0.013
R5415 AVDD.n2764 AVDD.n2763 0.013
R5416 AVDD.n2765 AVDD.n2764 0.013
R5417 AVDD.n2945 AVDD.n2944 0.013
R5418 AVDD.n2990 AVDD.n2945 0.013
R5419 AVDD.n2927 AVDD.n2926 0.013
R5420 AVDD.n2928 AVDD.n2927 0.013
R5421 AVDD.n3170 AVDD.n3169 0.013
R5422 AVDD.n3215 AVDD.n3170 0.013
R5423 AVDD.n3108 AVDD.n3107 0.013
R5424 AVDD.n3109 AVDD.n3108 0.013
R5425 AVDD.n3344 AVDD.n3343 0.013
R5426 AVDD.n3389 AVDD.n3344 0.013
R5427 AVDD.n3327 AVDD.n3326 0.013
R5428 AVDD.n3328 AVDD.n3327 0.013
R5429 AVDD.n4934 AVDD.n4933 0.013
R5430 AVDD.n4979 AVDD.n4934 0.013
R5431 AVDD.n4757 AVDD.n4756 0.013
R5432 AVDD.n4758 AVDD.n4757 0.013
R5433 AVDD.n4806 AVDD.n4805 0.013
R5434 AVDD.n4807 AVDD.n4806 0.013
R5435 AVDD.n4800 AVDD.n4799 0.013
R5436 AVDD.n4807 AVDD.n4800 0.013
R5437 AVDD.n4590 AVDD.n4584 0.013
R5438 AVDD.n4584 AVDD.n4583 0.013
R5439 AVDD.n4590 AVDD.n4586 0.013
R5440 AVDD.n4794 AVDD.n4793 0.013
R5441 AVDD.n4807 AVDD.n4794 0.013
R5442 AVDD.n4538 AVDD.n4532 0.013
R5443 AVDD.n4538 AVDD.n4534 0.013
R5444 AVDD.n4788 AVDD.n4787 0.013
R5445 AVDD.n4807 AVDD.n4788 0.013
R5446 AVDD.n4506 AVDD.n4456 0.013
R5447 AVDD.n4506 AVDD.n4502 0.013
R5448 AVDD.n4502 AVDD.n4501 0.013
R5449 AVDD.n4782 AVDD.n4781 0.013
R5450 AVDD.n4807 AVDD.n4782 0.013
R5451 AVDD.n4583 AVDD.n4579 0.013
R5452 AVDD.n4501 AVDD.n4469 0.013
R5453 AVDD.n4776 AVDD.n4775 0.013
R5454 AVDD.n4807 AVDD.n4776 0.013
R5455 AVDD.n3727 AVDD.n3721 0.013
R5456 AVDD.n3727 AVDD.n3723 0.013
R5457 AVDD.n608 AVDD.n607 0.013
R5458 AVDD.n621 AVDD.n608 0.013
R5459 AVDD.n851 AVDD.n850 0.013
R5460 AVDD.n860 AVDD.n851 0.013
R5461 AVDD.n789 AVDD.n788 0.013
R5462 AVDD.n802 AVDD.n789 0.013
R5463 AVDD.n1032 AVDD.n1031 0.013
R5464 AVDD.n1041 AVDD.n1032 0.013
R5465 AVDD.n970 AVDD.n969 0.013
R5466 AVDD.n983 AVDD.n970 0.013
R5467 AVDD.n1137 AVDD.n1136 0.013
R5468 AVDD.n1146 AVDD.n1137 0.013
R5469 AVDD.n1331 AVDD.n1330 0.013
R5470 AVDD.n1344 AVDD.n1331 0.013
R5471 AVDD.n1397 AVDD.n1396 0.013
R5472 AVDD.n1406 AVDD.n1397 0.013
R5473 AVDD.n1238 AVDD.n1237 0.013
R5474 AVDD.n1251 AVDD.n1238 0.013
R5475 AVDD.n1601 AVDD.n1600 0.013
R5476 AVDD.n1610 AVDD.n1601 0.013
R5477 AVDD.n1513 AVDD.n1512 0.013
R5478 AVDD.n1526 AVDD.n1513 0.013
R5479 AVDD.n1810 AVDD.n1809 0.013
R5480 AVDD.n1819 AVDD.n1810 0.013
R5481 AVDD.n1694 AVDD.n1693 0.013
R5482 AVDD.n1707 AVDD.n1694 0.013
R5483 AVDD.n2022 AVDD.n2021 0.013
R5484 AVDD.n2031 AVDD.n2022 0.013
R5485 AVDD.n1955 AVDD.n1954 0.013
R5486 AVDD.n1968 AVDD.n1955 0.013
R5487 AVDD.n2101 AVDD.n2100 0.013
R5488 AVDD.n2110 AVDD.n2101 0.013
R5489 AVDD.n2226 AVDD.n2225 0.013
R5490 AVDD.n2239 AVDD.n2226 0.013
R5491 AVDD.n2437 AVDD.n2436 0.013
R5492 AVDD.n2446 AVDD.n2437 0.013
R5493 AVDD.n2327 AVDD.n2326 0.013
R5494 AVDD.n2340 AVDD.n2327 0.013
R5495 AVDD.n2601 AVDD.n2600 0.013
R5496 AVDD.n2610 AVDD.n2601 0.013
R5497 AVDD.n2507 AVDD.n2506 0.013
R5498 AVDD.n2520 AVDD.n2507 0.013
R5499 AVDD.n584 AVDD.n583 0.013
R5500 AVDD.n621 AVDD.n584 0.013
R5501 AVDD.n827 AVDD.n826 0.013
R5502 AVDD.n860 AVDD.n827 0.013
R5503 AVDD.n765 AVDD.n764 0.013
R5504 AVDD.n802 AVDD.n765 0.013
R5505 AVDD.n1008 AVDD.n1007 0.013
R5506 AVDD.n1041 AVDD.n1008 0.013
R5507 AVDD.n946 AVDD.n945 0.013
R5508 AVDD.n983 AVDD.n946 0.013
R5509 AVDD.n1113 AVDD.n1112 0.013
R5510 AVDD.n1146 AVDD.n1113 0.013
R5511 AVDD.n1307 AVDD.n1306 0.013
R5512 AVDD.n1344 AVDD.n1307 0.013
R5513 AVDD.n1373 AVDD.n1372 0.013
R5514 AVDD.n1406 AVDD.n1373 0.013
R5515 AVDD.n1214 AVDD.n1213 0.013
R5516 AVDD.n1251 AVDD.n1214 0.013
R5517 AVDD.n1577 AVDD.n1576 0.013
R5518 AVDD.n1610 AVDD.n1577 0.013
R5519 AVDD.n1489 AVDD.n1488 0.013
R5520 AVDD.n1526 AVDD.n1489 0.013
R5521 AVDD.n1786 AVDD.n1785 0.013
R5522 AVDD.n1819 AVDD.n1786 0.013
R5523 AVDD.n1670 AVDD.n1669 0.013
R5524 AVDD.n1707 AVDD.n1670 0.013
R5525 AVDD.n1998 AVDD.n1997 0.013
R5526 AVDD.n2031 AVDD.n1998 0.013
R5527 AVDD.n1931 AVDD.n1930 0.013
R5528 AVDD.n1968 AVDD.n1931 0.013
R5529 AVDD.n2077 AVDD.n2076 0.013
R5530 AVDD.n2110 AVDD.n2077 0.013
R5531 AVDD.n2202 AVDD.n2201 0.013
R5532 AVDD.n2239 AVDD.n2202 0.013
R5533 AVDD.n2413 AVDD.n2412 0.013
R5534 AVDD.n2446 AVDD.n2413 0.013
R5535 AVDD.n2303 AVDD.n2302 0.013
R5536 AVDD.n2340 AVDD.n2303 0.013
R5537 AVDD.n2577 AVDD.n2576 0.013
R5538 AVDD.n2610 AVDD.n2577 0.013
R5539 AVDD.n2483 AVDD.n2482 0.013
R5540 AVDD.n2520 AVDD.n2483 0.013
R5541 AVDD.n2795 AVDD.n2794 0.013
R5542 AVDD.n2828 AVDD.n2795 0.013
R5543 AVDD.n2728 AVDD.n2727 0.013
R5544 AVDD.n2765 AVDD.n2728 0.013
R5545 AVDD.n2957 AVDD.n2956 0.013
R5546 AVDD.n2990 AVDD.n2957 0.013
R5547 AVDD.n2891 AVDD.n2890 0.013
R5548 AVDD.n2928 AVDD.n2891 0.013
R5549 AVDD.n3182 AVDD.n3181 0.013
R5550 AVDD.n3215 AVDD.n3182 0.013
R5551 AVDD.n3072 AVDD.n3071 0.013
R5552 AVDD.n3109 AVDD.n3072 0.013
R5553 AVDD.n3356 AVDD.n3355 0.013
R5554 AVDD.n3389 AVDD.n3356 0.013
R5555 AVDD.n3291 AVDD.n3290 0.013
R5556 AVDD.n3328 AVDD.n3291 0.013
R5557 AVDD.n4946 AVDD.n4945 0.013
R5558 AVDD.n4979 AVDD.n4946 0.013
R5559 AVDD.n4721 AVDD.n4720 0.013
R5560 AVDD.n4758 AVDD.n4721 0.013
R5561 AVDD.n3557 AVDD.n3551 0.013
R5562 AVDD.n3557 AVDD.n3553 0.013
R5563 AVDD.n4764 AVDD.n4763 0.013
R5564 AVDD.n4807 AVDD.n4764 0.013
R5565 AVDD.n4940 AVDD.n4939 0.013
R5566 AVDD.n4979 AVDD.n4940 0.013
R5567 AVDD.n4715 AVDD.n4714 0.013
R5568 AVDD.n4758 AVDD.n4715 0.013
R5569 AVDD.n3350 AVDD.n3349 0.013
R5570 AVDD.n3389 AVDD.n3350 0.013
R5571 AVDD.n3285 AVDD.n3284 0.013
R5572 AVDD.n3328 AVDD.n3285 0.013
R5573 AVDD.n3176 AVDD.n3175 0.013
R5574 AVDD.n3215 AVDD.n3176 0.013
R5575 AVDD.n3066 AVDD.n3065 0.013
R5576 AVDD.n3109 AVDD.n3066 0.013
R5577 AVDD.n2951 AVDD.n2950 0.013
R5578 AVDD.n2990 AVDD.n2951 0.013
R5579 AVDD.n2885 AVDD.n2884 0.013
R5580 AVDD.n2928 AVDD.n2885 0.013
R5581 AVDD.n2789 AVDD.n2788 0.013
R5582 AVDD.n2828 AVDD.n2789 0.013
R5583 AVDD.n2722 AVDD.n2721 0.013
R5584 AVDD.n2765 AVDD.n2722 0.013
R5585 AVDD.n2571 AVDD.n2570 0.013
R5586 AVDD.n2610 AVDD.n2571 0.013
R5587 AVDD.n2477 AVDD.n2476 0.013
R5588 AVDD.n2520 AVDD.n2477 0.013
R5589 AVDD.n2407 AVDD.n2406 0.013
R5590 AVDD.n2446 AVDD.n2407 0.013
R5591 AVDD.n2297 AVDD.n2296 0.013
R5592 AVDD.n2340 AVDD.n2297 0.013
R5593 AVDD.n2071 AVDD.n2070 0.013
R5594 AVDD.n2110 AVDD.n2071 0.013
R5595 AVDD.n2196 AVDD.n2195 0.013
R5596 AVDD.n2239 AVDD.n2196 0.013
R5597 AVDD.n1992 AVDD.n1991 0.013
R5598 AVDD.n2031 AVDD.n1992 0.013
R5599 AVDD.n1925 AVDD.n1924 0.013
R5600 AVDD.n1968 AVDD.n1925 0.013
R5601 AVDD.n1780 AVDD.n1779 0.013
R5602 AVDD.n1819 AVDD.n1780 0.013
R5603 AVDD.n1664 AVDD.n1663 0.013
R5604 AVDD.n1707 AVDD.n1664 0.013
R5605 AVDD.n1571 AVDD.n1570 0.013
R5606 AVDD.n1610 AVDD.n1571 0.013
R5607 AVDD.n1483 AVDD.n1482 0.013
R5608 AVDD.n1526 AVDD.n1483 0.013
R5609 AVDD.n1367 AVDD.n1366 0.013
R5610 AVDD.n1406 AVDD.n1367 0.013
R5611 AVDD.n1208 AVDD.n1207 0.013
R5612 AVDD.n1251 AVDD.n1208 0.013
R5613 AVDD.n3478 AVDD.n3472 0.013
R5614 AVDD.n3478 AVDD.n3474 0.013
R5615 AVDD.n3587 AVDD.n3586 0.013
R5616 AVDD.n3637 AVDD.n3587 0.013
R5617 AVDD.n3595 AVDD.n3594 0.013
R5618 AVDD.n3637 AVDD.n3595 0.013
R5619 AVDD.n3603 AVDD.n3602 0.013
R5620 AVDD.n3637 AVDD.n3603 0.013
R5621 AVDD.n3611 AVDD.n3610 0.013
R5622 AVDD.n3637 AVDD.n3611 0.013
R5623 AVDD.n3619 AVDD.n3618 0.013
R5624 AVDD.n3637 AVDD.n3619 0.013
R5625 AVDD.n3627 AVDD.n3626 0.013
R5626 AVDD.n3637 AVDD.n3627 0.013
R5627 AVDD.n3635 AVDD.n3634 0.013
R5628 AVDD.n3637 AVDD.n3635 0.013
R5629 AVDD.n4583 AVDD.n4582 0.013
R5630 AVDD.n4500 AVDD.n4499 0.013
R5631 AVDD.n4501 AVDD.n4500 0.013
R5632 AVDD.n6362 AVDD.n6361 0.011
R5633 AVDD.n3791 level_shifter_up_3.VDD_HV 0.01
R5634 AVDD.n3830 level_shifter_up_1.VDD_HV 0.01
R5635 AVDD.n3958 level_shifter_up_2.VDD_HV 0.01
R5636 AVDD.n4045 AVDD 0.01
R5637 AVDD.n4175 level_shifter_up_7.VDD_HV 0.01
R5638 AVDD.n1751 AVDD.n1750 0.01
R5639 AVDD.n1766 AVDD.n1751 0.01
R5640 AVDD.n1543 AVDD.n1542 0.01
R5641 AVDD.n1558 AVDD.n1543 0.01
R5642 AVDD.n2132 AVDD.n2131 0.01
R5643 AVDD.n2147 AVDD.n2132 0.01
R5644 AVDD.n1712 AVDD.n1711 0.01
R5645 AVDD.n1727 AVDD.n1712 0.01
R5646 AVDD.n2379 AVDD.n2378 0.01
R5647 AVDD.n2394 AVDD.n2379 0.01
R5648 AVDD.n2154 AVDD.n2153 0.01
R5649 AVDD.n2169 AVDD.n2154 0.01
R5650 AVDD.n2525 AVDD.n2524 0.01
R5651 AVDD.n2540 AVDD.n2525 0.01
R5652 AVDD.n2357 AVDD.n2356 0.01
R5653 AVDD.n2372 AVDD.n2357 0.01
R5654 AVDD.n3013 AVDD.n3012 0.01
R5655 AVDD.n3028 AVDD.n3013 0.01
R5656 AVDD.n2833 AVDD.n2832 0.01
R5657 AVDD.n2848 AVDD.n2833 0.01
R5658 AVDD.n3147 AVDD.n3146 0.01
R5659 AVDD.n3162 AVDD.n3147 0.01
R5660 AVDD.n3035 AVDD.n3034 0.01
R5661 AVDD.n3050 AVDD.n3035 0.01
R5662 AVDD.n4984 AVDD.n4983 0.01
R5663 AVDD.n4999 AVDD.n4984 0.01
R5664 AVDD.n3125 AVDD.n3124 0.01
R5665 AVDD.n3140 AVDD.n3125 0.01
R5666 AVDD.n4609 AVDD.n4608 0.01
R5667 AVDD.n4658 AVDD.n4609 0.01
R5668 AVDD.n5023 AVDD.n5022 0.01
R5669 AVDD.n5038 AVDD.n5023 0.01
R5670 AVDD.n1753 AVDD.n1752 0.01
R5671 AVDD.n1766 AVDD.n1753 0.01
R5672 AVDD.n1545 AVDD.n1544 0.01
R5673 AVDD.n1558 AVDD.n1545 0.01
R5674 AVDD.n2134 AVDD.n2133 0.01
R5675 AVDD.n2147 AVDD.n2134 0.01
R5676 AVDD.n1714 AVDD.n1713 0.01
R5677 AVDD.n1727 AVDD.n1714 0.01
R5678 AVDD.n2381 AVDD.n2380 0.01
R5679 AVDD.n2394 AVDD.n2381 0.01
R5680 AVDD.n2156 AVDD.n2155 0.01
R5681 AVDD.n2169 AVDD.n2156 0.01
R5682 AVDD.n2527 AVDD.n2526 0.01
R5683 AVDD.n2540 AVDD.n2527 0.01
R5684 AVDD.n2359 AVDD.n2358 0.01
R5685 AVDD.n2372 AVDD.n2359 0.01
R5686 AVDD.n3015 AVDD.n3014 0.01
R5687 AVDD.n3028 AVDD.n3015 0.01
R5688 AVDD.n2835 AVDD.n2834 0.01
R5689 AVDD.n2848 AVDD.n2835 0.01
R5690 AVDD.n3149 AVDD.n3148 0.01
R5691 AVDD.n3162 AVDD.n3149 0.01
R5692 AVDD.n3037 AVDD.n3036 0.01
R5693 AVDD.n3050 AVDD.n3037 0.01
R5694 AVDD.n4986 AVDD.n4985 0.01
R5695 AVDD.n4999 AVDD.n4986 0.01
R5696 AVDD.n3127 AVDD.n3126 0.01
R5697 AVDD.n3140 AVDD.n3127 0.01
R5698 AVDD.n4611 AVDD.n4610 0.01
R5699 AVDD.n4658 AVDD.n4611 0.01
R5700 AVDD.n5025 AVDD.n5024 0.01
R5701 AVDD.n5038 AVDD.n5025 0.01
R5702 AVDD.n1755 AVDD.n1754 0.01
R5703 AVDD.n1766 AVDD.n1755 0.01
R5704 AVDD.n1547 AVDD.n1546 0.01
R5705 AVDD.n1558 AVDD.n1547 0.01
R5706 AVDD.n2136 AVDD.n2135 0.01
R5707 AVDD.n2147 AVDD.n2136 0.01
R5708 AVDD.n1716 AVDD.n1715 0.01
R5709 AVDD.n1727 AVDD.n1716 0.01
R5710 AVDD.n2383 AVDD.n2382 0.01
R5711 AVDD.n2394 AVDD.n2383 0.01
R5712 AVDD.n2158 AVDD.n2157 0.01
R5713 AVDD.n2169 AVDD.n2158 0.01
R5714 AVDD.n2529 AVDD.n2528 0.01
R5715 AVDD.n2540 AVDD.n2529 0.01
R5716 AVDD.n2361 AVDD.n2360 0.01
R5717 AVDD.n2372 AVDD.n2361 0.01
R5718 AVDD.n3017 AVDD.n3016 0.01
R5719 AVDD.n3028 AVDD.n3017 0.01
R5720 AVDD.n2837 AVDD.n2836 0.01
R5721 AVDD.n2848 AVDD.n2837 0.01
R5722 AVDD.n3151 AVDD.n3150 0.01
R5723 AVDD.n3162 AVDD.n3151 0.01
R5724 AVDD.n3039 AVDD.n3038 0.01
R5725 AVDD.n3050 AVDD.n3039 0.01
R5726 AVDD.n4988 AVDD.n4987 0.01
R5727 AVDD.n4999 AVDD.n4988 0.01
R5728 AVDD.n3129 AVDD.n3128 0.01
R5729 AVDD.n3140 AVDD.n3129 0.01
R5730 AVDD.n4613 AVDD.n4612 0.01
R5731 AVDD.n4658 AVDD.n4613 0.01
R5732 AVDD.n5027 AVDD.n5026 0.01
R5733 AVDD.n5038 AVDD.n5027 0.01
R5734 AVDD.n1757 AVDD.n1756 0.01
R5735 AVDD.n1766 AVDD.n1757 0.01
R5736 AVDD.n1549 AVDD.n1548 0.01
R5737 AVDD.n1558 AVDD.n1549 0.01
R5738 AVDD.n2138 AVDD.n2137 0.01
R5739 AVDD.n2147 AVDD.n2138 0.01
R5740 AVDD.n1718 AVDD.n1717 0.01
R5741 AVDD.n1727 AVDD.n1718 0.01
R5742 AVDD.n2385 AVDD.n2384 0.01
R5743 AVDD.n2394 AVDD.n2385 0.01
R5744 AVDD.n2160 AVDD.n2159 0.01
R5745 AVDD.n2169 AVDD.n2160 0.01
R5746 AVDD.n2531 AVDD.n2530 0.01
R5747 AVDD.n2540 AVDD.n2531 0.01
R5748 AVDD.n2363 AVDD.n2362 0.01
R5749 AVDD.n2372 AVDD.n2363 0.01
R5750 AVDD.n3019 AVDD.n3018 0.01
R5751 AVDD.n3028 AVDD.n3019 0.01
R5752 AVDD.n2839 AVDD.n2838 0.01
R5753 AVDD.n2848 AVDD.n2839 0.01
R5754 AVDD.n3153 AVDD.n3152 0.01
R5755 AVDD.n3162 AVDD.n3153 0.01
R5756 AVDD.n3041 AVDD.n3040 0.01
R5757 AVDD.n3050 AVDD.n3041 0.01
R5758 AVDD.n4990 AVDD.n4989 0.01
R5759 AVDD.n4999 AVDD.n4990 0.01
R5760 AVDD.n3131 AVDD.n3130 0.01
R5761 AVDD.n3140 AVDD.n3131 0.01
R5762 AVDD.n4615 AVDD.n4614 0.01
R5763 AVDD.n4658 AVDD.n4615 0.01
R5764 AVDD.n5029 AVDD.n5028 0.01
R5765 AVDD.n5038 AVDD.n5029 0.01
R5766 AVDD.n1759 AVDD.n1758 0.01
R5767 AVDD.n1766 AVDD.n1759 0.01
R5768 AVDD.n1551 AVDD.n1550 0.01
R5769 AVDD.n1558 AVDD.n1551 0.01
R5770 AVDD.n2140 AVDD.n2139 0.01
R5771 AVDD.n2147 AVDD.n2140 0.01
R5772 AVDD.n1720 AVDD.n1719 0.01
R5773 AVDD.n1727 AVDD.n1720 0.01
R5774 AVDD.n2387 AVDD.n2386 0.01
R5775 AVDD.n2394 AVDD.n2387 0.01
R5776 AVDD.n2162 AVDD.n2161 0.01
R5777 AVDD.n2169 AVDD.n2162 0.01
R5778 AVDD.n2533 AVDD.n2532 0.01
R5779 AVDD.n2540 AVDD.n2533 0.01
R5780 AVDD.n2365 AVDD.n2364 0.01
R5781 AVDD.n2372 AVDD.n2365 0.01
R5782 AVDD.n3021 AVDD.n3020 0.01
R5783 AVDD.n3028 AVDD.n3021 0.01
R5784 AVDD.n2841 AVDD.n2840 0.01
R5785 AVDD.n2848 AVDD.n2841 0.01
R5786 AVDD.n3155 AVDD.n3154 0.01
R5787 AVDD.n3162 AVDD.n3155 0.01
R5788 AVDD.n3043 AVDD.n3042 0.01
R5789 AVDD.n3050 AVDD.n3043 0.01
R5790 AVDD.n4992 AVDD.n4991 0.01
R5791 AVDD.n4999 AVDD.n4992 0.01
R5792 AVDD.n3133 AVDD.n3132 0.01
R5793 AVDD.n3140 AVDD.n3133 0.01
R5794 AVDD.n4617 AVDD.n4616 0.01
R5795 AVDD.n4658 AVDD.n4617 0.01
R5796 AVDD.n5031 AVDD.n5030 0.01
R5797 AVDD.n5038 AVDD.n5031 0.01
R5798 AVDD.n1761 AVDD.n1760 0.01
R5799 AVDD.n1766 AVDD.n1761 0.01
R5800 AVDD.n1553 AVDD.n1552 0.01
R5801 AVDD.n1558 AVDD.n1553 0.01
R5802 AVDD.n2142 AVDD.n2141 0.01
R5803 AVDD.n2147 AVDD.n2142 0.01
R5804 AVDD.n1722 AVDD.n1721 0.01
R5805 AVDD.n1727 AVDD.n1722 0.01
R5806 AVDD.n2389 AVDD.n2388 0.01
R5807 AVDD.n2394 AVDD.n2389 0.01
R5808 AVDD.n2164 AVDD.n2163 0.01
R5809 AVDD.n2169 AVDD.n2164 0.01
R5810 AVDD.n2535 AVDD.n2534 0.01
R5811 AVDD.n2540 AVDD.n2535 0.01
R5812 AVDD.n2367 AVDD.n2366 0.01
R5813 AVDD.n2372 AVDD.n2367 0.01
R5814 AVDD.n3023 AVDD.n3022 0.01
R5815 AVDD.n3028 AVDD.n3023 0.01
R5816 AVDD.n2843 AVDD.n2842 0.01
R5817 AVDD.n2848 AVDD.n2843 0.01
R5818 AVDD.n3157 AVDD.n3156 0.01
R5819 AVDD.n3162 AVDD.n3157 0.01
R5820 AVDD.n3045 AVDD.n3044 0.01
R5821 AVDD.n3050 AVDD.n3045 0.01
R5822 AVDD.n4994 AVDD.n4993 0.01
R5823 AVDD.n4999 AVDD.n4994 0.01
R5824 AVDD.n3135 AVDD.n3134 0.01
R5825 AVDD.n3140 AVDD.n3135 0.01
R5826 AVDD.n4619 AVDD.n4618 0.01
R5827 AVDD.n4658 AVDD.n4619 0.01
R5828 AVDD.n5033 AVDD.n5032 0.01
R5829 AVDD.n5038 AVDD.n5033 0.01
R5830 AVDD.n1763 AVDD.n1762 0.01
R5831 AVDD.n1766 AVDD.n1763 0.01
R5832 AVDD.n1555 AVDD.n1554 0.01
R5833 AVDD.n1558 AVDD.n1555 0.01
R5834 AVDD.n2144 AVDD.n2143 0.01
R5835 AVDD.n2147 AVDD.n2144 0.01
R5836 AVDD.n1724 AVDD.n1723 0.01
R5837 AVDD.n1727 AVDD.n1724 0.01
R5838 AVDD.n2391 AVDD.n2390 0.01
R5839 AVDD.n2394 AVDD.n2391 0.01
R5840 AVDD.n2166 AVDD.n2165 0.01
R5841 AVDD.n2169 AVDD.n2166 0.01
R5842 AVDD.n2537 AVDD.n2536 0.01
R5843 AVDD.n2540 AVDD.n2537 0.01
R5844 AVDD.n2369 AVDD.n2368 0.01
R5845 AVDD.n2372 AVDD.n2369 0.01
R5846 AVDD.n3025 AVDD.n3024 0.01
R5847 AVDD.n3028 AVDD.n3025 0.01
R5848 AVDD.n2845 AVDD.n2844 0.01
R5849 AVDD.n2848 AVDD.n2845 0.01
R5850 AVDD.n3159 AVDD.n3158 0.01
R5851 AVDD.n3162 AVDD.n3159 0.01
R5852 AVDD.n3047 AVDD.n3046 0.01
R5853 AVDD.n3050 AVDD.n3047 0.01
R5854 AVDD.n4996 AVDD.n4995 0.01
R5855 AVDD.n4999 AVDD.n4996 0.01
R5856 AVDD.n3137 AVDD.n3136 0.01
R5857 AVDD.n3140 AVDD.n3137 0.01
R5858 AVDD.n4621 AVDD.n4620 0.01
R5859 AVDD.n4658 AVDD.n4621 0.01
R5860 AVDD.n5035 AVDD.n5034 0.01
R5861 AVDD.n5038 AVDD.n5035 0.01
R5862 AVDD.n1765 AVDD.n1764 0.01
R5863 AVDD.n1766 AVDD.n1765 0.01
R5864 AVDD.n1557 AVDD.n1556 0.01
R5865 AVDD.n1558 AVDD.n1557 0.01
R5866 AVDD.n2146 AVDD.n2145 0.01
R5867 AVDD.n2147 AVDD.n2146 0.01
R5868 AVDD.n1726 AVDD.n1725 0.01
R5869 AVDD.n1727 AVDD.n1726 0.01
R5870 AVDD.n2393 AVDD.n2392 0.01
R5871 AVDD.n2394 AVDD.n2393 0.01
R5872 AVDD.n2168 AVDD.n2167 0.01
R5873 AVDD.n2169 AVDD.n2168 0.01
R5874 AVDD.n2539 AVDD.n2538 0.01
R5875 AVDD.n2540 AVDD.n2539 0.01
R5876 AVDD.n2371 AVDD.n2370 0.01
R5877 AVDD.n2372 AVDD.n2371 0.01
R5878 AVDD.n3027 AVDD.n3026 0.01
R5879 AVDD.n3028 AVDD.n3027 0.01
R5880 AVDD.n2847 AVDD.n2846 0.01
R5881 AVDD.n2848 AVDD.n2847 0.01
R5882 AVDD.n3161 AVDD.n3160 0.01
R5883 AVDD.n3162 AVDD.n3161 0.01
R5884 AVDD.n3049 AVDD.n3048 0.01
R5885 AVDD.n3050 AVDD.n3049 0.01
R5886 AVDD.n4998 AVDD.n4997 0.01
R5887 AVDD.n4999 AVDD.n4998 0.01
R5888 AVDD.n3139 AVDD.n3138 0.01
R5889 AVDD.n3140 AVDD.n3139 0.01
R5890 AVDD.n4623 AVDD.n4622 0.01
R5891 AVDD.n4658 AVDD.n4623 0.01
R5892 AVDD.n5037 AVDD.n5036 0.01
R5893 AVDD.n5038 AVDD.n5037 0.01
R5894 AVDD.n4656 AVDD.n4654 0.01
R5895 AVDD.n4654 AVDD.n4653 0.01
R5896 AVDD.n1631 AVDD.n1630 0.01
R5897 AVDD.n1648 AVDD.n1631 0.01
R5898 AVDD.n1461 AVDD.n1460 0.01
R5899 AVDD.n1467 AVDD.n1461 0.01
R5900 AVDD.n1648 AVDD.n1633 0.01
R5901 AVDD.n1457 AVDD.n1456 0.01
R5902 AVDD.n1467 AVDD.n1457 0.01
R5903 AVDD.n1648 AVDD.n1635 0.01
R5904 AVDD.n1452 AVDD.n1451 0.01
R5905 AVDD.n1467 AVDD.n1452 0.01
R5906 AVDD.n1648 AVDD.n1637 0.01
R5907 AVDD.n1447 AVDD.n1446 0.01
R5908 AVDD.n1467 AVDD.n1447 0.01
R5909 AVDD.n1648 AVDD.n1639 0.01
R5910 AVDD.n1442 AVDD.n1441 0.01
R5911 AVDD.n1467 AVDD.n1442 0.01
R5912 AVDD.n1648 AVDD.n1641 0.01
R5913 AVDD.n1437 AVDD.n1436 0.01
R5914 AVDD.n1467 AVDD.n1437 0.01
R5915 AVDD.n1648 AVDD.n1643 0.01
R5916 AVDD.n1433 AVDD.n1432 0.01
R5917 AVDD.n1467 AVDD.n1433 0.01
R5918 AVDD.n1648 AVDD.n1645 0.01
R5919 AVDD.n1650 AVDD.n1649 0.01
R5920 AVDD.n1649 AVDD.n1648 0.01
R5921 AVDD.n1469 AVDD.n1468 0.01
R5922 AVDD.n1468 AVDD.n1467 0.01
R5923 AVDD.n3669 AVDD.n3662 0.01
R5924 AVDD.n3669 AVDD.n3660 0.01
R5925 AVDD.n3669 AVDD.n3658 0.01
R5926 AVDD.n3669 AVDD.n3656 0.01
R5927 AVDD.n3669 AVDD.n3654 0.01
R5928 AVDD.n5021 AVDD.n5020 0.01
R5929 AVDD.n5038 AVDD.n5021 0.01
R5930 AVDD.n4982 AVDD.n4981 0.01
R5931 AVDD.n4999 AVDD.n4982 0.01
R5932 AVDD.n3669 AVDD.n3652 0.01
R5933 AVDD.n4633 AVDD.n4632 0.01
R5934 AVDD.n4653 AVDD.n4633 0.01
R5935 AVDD.n4607 AVDD.n4606 0.01
R5936 AVDD.n4658 AVDD.n4607 0.01
R5937 AVDD.n3011 AVDD.n3010 0.01
R5938 AVDD.n3028 AVDD.n3011 0.01
R5939 AVDD.n2377 AVDD.n2376 0.01
R5940 AVDD.n2394 AVDD.n2377 0.01
R5941 AVDD.n1749 AVDD.n1748 0.01
R5942 AVDD.n1766 AVDD.n1749 0.01
R5943 AVDD.n3033 AVDD.n3032 0.01
R5944 AVDD.n3050 AVDD.n3033 0.01
R5945 AVDD.n2355 AVDD.n2354 0.01
R5946 AVDD.n2372 AVDD.n2355 0.01
R5947 AVDD.n1710 AVDD.n1709 0.01
R5948 AVDD.n1727 AVDD.n1710 0.01
R5949 AVDD.n1541 AVDD.n1540 0.01
R5950 AVDD.n1558 AVDD.n1541 0.01
R5951 AVDD.n2130 AVDD.n2129 0.01
R5952 AVDD.n2147 AVDD.n2130 0.01
R5953 AVDD.n2152 AVDD.n2151 0.01
R5954 AVDD.n2169 AVDD.n2152 0.01
R5955 AVDD.n2523 AVDD.n2522 0.01
R5956 AVDD.n2540 AVDD.n2523 0.01
R5957 AVDD.n2831 AVDD.n2830 0.01
R5958 AVDD.n2848 AVDD.n2831 0.01
R5959 AVDD.n3145 AVDD.n3144 0.01
R5960 AVDD.n3162 AVDD.n3145 0.01
R5961 AVDD.n3123 AVDD.n3122 0.01
R5962 AVDD.n3140 AVDD.n3123 0.01
R5963 AVDD.n4637 AVDD.n4636 0.01
R5964 AVDD.n4653 AVDD.n4637 0.01
R5965 AVDD.n4639 AVDD.n4638 0.01
R5966 AVDD.n4653 AVDD.n4639 0.01
R5967 AVDD.n4643 AVDD.n4642 0.01
R5968 AVDD.n4653 AVDD.n4643 0.01
R5969 AVDD.n4645 AVDD.n4644 0.01
R5970 AVDD.n4653 AVDD.n4645 0.01
R5971 AVDD.n4648 AVDD.n4647 0.01
R5972 AVDD.n4653 AVDD.n4648 0.01
R5973 AVDD.n4629 AVDD.n4628 0.01
R5974 AVDD.n4653 AVDD.n4629 0.01
R5975 AVDD.n4657 AVDD.n4656 0.01
R5976 AVDD.n4658 AVDD.n4657 0.01
R5977 AVDD.n5040 AVDD.n5039 0.01
R5978 AVDD.n5039 AVDD.n5038 0.01
R5979 AVDD.n5001 AVDD.n5000 0.01
R5980 AVDD.n5000 AVDD.n4999 0.01
R5981 AVDD.n3142 AVDD.n3141 0.01
R5982 AVDD.n3141 AVDD.n3140 0.01
R5983 AVDD.n3164 AVDD.n3163 0.01
R5984 AVDD.n3163 AVDD.n3162 0.01
R5985 AVDD.n3052 AVDD.n3051 0.01
R5986 AVDD.n3051 AVDD.n3050 0.01
R5987 AVDD.n3030 AVDD.n3029 0.01
R5988 AVDD.n3029 AVDD.n3028 0.01
R5989 AVDD.n2850 AVDD.n2849 0.01
R5990 AVDD.n2849 AVDD.n2848 0.01
R5991 AVDD.n2542 AVDD.n2541 0.01
R5992 AVDD.n2541 AVDD.n2540 0.01
R5993 AVDD.n2374 AVDD.n2373 0.01
R5994 AVDD.n2373 AVDD.n2372 0.01
R5995 AVDD.n2396 AVDD.n2395 0.01
R5996 AVDD.n2395 AVDD.n2394 0.01
R5997 AVDD.n2171 AVDD.n2170 0.01
R5998 AVDD.n2170 AVDD.n2169 0.01
R5999 AVDD.n2149 AVDD.n2148 0.01
R6000 AVDD.n2148 AVDD.n2147 0.01
R6001 AVDD.n1729 AVDD.n1728 0.01
R6002 AVDD.n1728 AVDD.n1727 0.01
R6003 AVDD.n1768 AVDD.n1767 0.01
R6004 AVDD.n1767 AVDD.n1766 0.01
R6005 AVDD.n1560 AVDD.n1559 0.01
R6006 AVDD.n1559 AVDD.n1558 0.01
R6007 AVDD.n1427 AVDD.n1426 0.01
R6008 AVDD.n1467 AVDD.n1427 0.01
R6009 AVDD.n1648 AVDD.n1647 0.01
R6010 AVDD.n1466 AVDD.n1465 0.01
R6011 AVDD.n1467 AVDD.n1466 0.01
R6012 AVDD.n3669 AVDD.n3666 0.01
R6013 AVDD.n3669 AVDD.n3664 0.01
R6014 AVDD.n4652 AVDD.n4651 0.01
R6015 AVDD.n4653 AVDD.n4652 0.01
R6016 AVDD.n4626 AVDD.n4625 0.01
R6017 AVDD.n4653 AVDD.n4626 0.01
R6018 AVDD.n3669 AVDD.n3668 0.01
R6019 AVDD.n3671 AVDD.n3670 0.01
R6020 AVDD.n3670 AVDD.n3669 0.01
R6021 AVDD.t731 AVDD.n3792 0.009
R6022 AVDD.n6361 AVDD.n6360 0.009
R6023 AVDD.t52 AVDD.n5827 0.008
R6024 AVDD.n3537 AVDD.n3536 0.008
R6025 AVDD.n4544 AVDD.n4543 0.008
R6026 AVDD.n4515 AVDD.n4511 0.008
R6027 AVDD.n4439 AVDD.n4435 0.008
R6028 AVDD.n3733 AVDD.n3732 0.008
R6029 AVDD.n3563 AVDD.n3562 0.008
R6030 AVDD.n3494 AVDD.n3491 0.008
R6031 AVDD.n3501 AVDD.n3500 0.008
R6032 AVDD.n3889 AVDD.n3888 0.008
R6033 AVDD.t142 AVDD.n3889 0.008
R6034 AVDD.n3827 AVDD.n3826 0.008
R6035 AVDD.n4391 AVDD.n4257 0.008
R6036 AVDD.n4393 AVDD.n4392 0.008
R6037 AVDD.t739 AVDD.n4393 0.008
R6038 AVDD.n4104 AVDD.n4103 0.008
R6039 AVDD.t745 AVDD.n4104 0.008
R6040 AVDD.n4042 AVDD.n4041 0.008
R6041 AVDD.n4219 AVDD.n4218 0.008
R6042 AVDD.n5358 AVDD.n5355 0.008
R6043 AVDD.n3779 AVDD.n3751 0.008
R6044 AVDD.n6498 AVDD.n6497 0.008
R6045 AVDD.t31 AVDD.n6498 0.008
R6046 AVDD.n6068 AVDD.n6067 0.008
R6047 AVDD.t275 AVDD.n6068 0.008
R6048 AVDD.n5300 AVDD.n5299 0.007
R6049 AVDD.n3845 AVDD.n3844 0.007
R6050 AVDD.n3844 AVDD.n3843 0.007
R6051 AVDD.n3832 AVDD.n3831 0.007
R6052 AVDD.n3912 AVDD.n3911 0.007
R6053 AVDD.n3911 AVDD.n3910 0.007
R6054 AVDD.n3899 AVDD.n3898 0.007
R6055 AVDD.n3898 AVDD.n3897 0.007
R6056 AVDD.n3978 AVDD.n3977 0.007
R6057 AVDD.n3977 AVDD.n3976 0.007
R6058 AVDD.n3965 AVDD.n3964 0.007
R6059 AVDD.n3964 AVDD.n3963 0.007
R6060 AVDD.n4200 AVDD.n4199 0.007
R6061 AVDD.n4201 AVDD.n4200 0.007
R6062 AVDD.n4184 AVDD.n4183 0.007
R6063 AVDD.n4185 AVDD.n4184 0.007
R6064 AVDD.n4060 AVDD.n4059 0.007
R6065 AVDD.n4059 AVDD.n4058 0.007
R6066 AVDD.n4047 AVDD.n4046 0.007
R6067 AVDD.n4127 AVDD.n4126 0.007
R6068 AVDD.n4126 AVDD.n4125 0.007
R6069 AVDD.n4114 AVDD.n4113 0.007
R6070 AVDD.n4113 AVDD.n4112 0.007
R6071 AVDD.n3755 AVDD.n3754 0.007
R6072 AVDD.n3756 AVDD.n3755 0.007
R6073 AVDD.n3758 AVDD.n3757 0.007
R6074 AVDD.n19 AVDD.n18 0.007
R6075 AVDD.n20 AVDD.n19 0.007
R6076 AVDD.n5892 AVDD.n5891 0.007
R6077 AVDD.n5893 AVDD.n5892 0.007
R6078 AVDD.n6109 AVDD.n6108 0.007
R6079 AVDD.n6110 AVDD.n6109 0.007
R6080 AVDD.n6320 AVDD.n6319 0.007
R6081 AVDD.n6321 AVDD.n6320 0.007
R6082 AVDD.n4370 AVDD.n4369 0.006
R6083 AVDD.n4371 AVDD.n4370 0.006
R6084 AVDD.n4373 AVDD.n4372 0.006
R6085 AVDD.n4372 AVDD.n4371 0.006
R6086 AVDD.n4296 AVDD.n4295 0.006
R6087 AVDD.n4295 AVDD.n4294 0.006
R6088 AVDD.n4293 AVDD.n4292 0.006
R6089 AVDD.n4294 AVDD.n4293 0.006
R6090 AVDD.n4303 AVDD.n4302 0.006
R6091 AVDD.n4302 AVDD.n4301 0.006
R6092 AVDD.n4301 AVDD.n4300 0.006
R6093 AVDD.n4318 AVDD.n4317 0.006
R6094 AVDD.n4319 AVDD.n4318 0.006
R6095 AVDD.n4026 AVDD.n4025 0.006
R6096 AVDD.n4025 AVDD.n4024 0.006
R6097 AVDD.n4024 AVDD.n4023 0.006
R6098 AVDD.n4377 AVDD.n4376 0.006
R6099 AVDD.n4378 AVDD.n4377 0.006
R6100 AVDD.n4378 AVDD.n4328 0.006
R6101 AVDD.n4321 AVDD.n4320 0.006
R6102 AVDD.n4320 AVDD.n4319 0.006
R6103 AVDD.n3983 AVDD.n3982 0.006
R6104 AVDD.n6405 AVDD.n6400 0.006
R6105 AVDD.n6373 AVDD.n6372 0.006
R6106 AVDD.n6376 AVDD.n6373 0.006
R6107 AVDD.n372 AVDD.n371 0.006
R6108 AVDD.n424 AVDD.n372 0.006
R6109 AVDD.n423 AVDD.n422 0.006
R6110 AVDD.n424 AVDD.n423 0.006
R6111 AVDD.n4300 AVDD.n4299 0.006
R6112 AVDD.n4023 AVDD.n4022 0.006
R6113 AVDD.n4328 AVDD.n4327 0.006
R6114 AVDD.n5752 AVDD.n5751 0.005
R6115 AVDD.n5794 AVDD.n5793 0.005
R6116 AVDD.n6151 AVDD.n6150 0.005
R6117 AVDD.n6195 AVDD.n6194 0.005
R6118 AVDD.n6218 AVDD.n6217 0.005
R6119 AVDD.n6241 AVDD.n6240 0.005
R6120 AVDD.n6264 AVDD.n6263 0.005
R6121 AVDD.n6287 AVDD.n6286 0.005
R6122 AVDD.n6256 AVDD.n6255 0.005
R6123 AVDD.n6233 AVDD.n6232 0.005
R6124 AVDD.n6210 AVDD.n6209 0.005
R6125 AVDD.n6188 AVDD.n6187 0.005
R6126 AVDD.n6144 AVDD.n6143 0.005
R6127 AVDD.n5786 AVDD.n5785 0.005
R6128 AVDD.n5769 AVDD.n5768 0.005
R6129 AVDD.n6279 AVDD.n6278 0.005
R6130 AVDD.n4492 AVDD.n4491 0.005
R6131 AVDD.n3470 AVDD.n3469 0.005
R6132 AVDD.n3549 AVDD.n3548 0.005
R6133 AVDD.n3719 AVDD.n3718 0.005
R6134 AVDD.n4426 AVDD.n4425 0.005
R6135 AVDD.n4454 AVDD.n4453 0.005
R6136 AVDD.n4530 AVDD.n4529 0.005
R6137 AVDD.n4558 AVDD.n4557 0.005
R6138 AVDD.n4489 AVDD.n4488 0.005
R6139 AVDD.n4589 AVDD.n4588 0.005
R6140 AVDD.n4537 AVDD.n4536 0.005
R6141 AVDD.n4505 AVDD.n4504 0.005
R6142 AVDD.n4429 AVDD.n4428 0.005
R6143 AVDD.n3726 AVDD.n3725 0.005
R6144 AVDD.n3556 AVDD.n3555 0.005
R6145 AVDD.n3477 AVDD.n3476 0.005
R6146 AVDD.n5307 AVDD.n5306 0.005
R6147 AVDD.n4575 AVDD.n4572 0.005
R6148 AVDD.n6172 AVDD.n6171 0.005
R6149 AVDD.n6131 AVDD.n6130 0.005
R6150 AVDD.n3633 AVDD.n3632 0.005
R6151 AVDD.n3625 AVDD.n3624 0.005
R6152 AVDD.n3617 AVDD.n3616 0.005
R6153 AVDD.n3609 AVDD.n3608 0.005
R6154 AVDD.n3601 AVDD.n3600 0.005
R6155 AVDD.n3593 AVDD.n3592 0.005
R6156 AVDD.n3585 AVDD.n3584 0.005
R6157 AVDD.n4214 AVDD.n4212 0.005
R6158 AVDD.n3581 AVDD.n3580 0.005
R6159 AVDD.n3557 AVDD.n3546 0.005
R6160 AVDD.n3727 AVDD.n3716 0.005
R6161 AVDD.n4430 AVDD.n4423 0.005
R6162 AVDD.n4506 AVDD.n4451 0.005
R6163 AVDD.n4538 AVDD.n4527 0.005
R6164 AVDD.n4590 AVDD.n4555 0.005
R6165 AVDD.n6277 AVDD.n6270 0.005
R6166 AVDD.n6277 AVDD.n6269 0.005
R6167 AVDD.n6254 AVDD.n6247 0.005
R6168 AVDD.n6254 AVDD.n6246 0.005
R6169 AVDD.n6231 AVDD.n6224 0.005
R6170 AVDD.n6231 AVDD.n6223 0.005
R6171 AVDD.n6208 AVDD.n6201 0.005
R6172 AVDD.n6208 AVDD.n6200 0.005
R6173 AVDD.n6186 AVDD.n6157 0.005
R6174 AVDD.n6186 AVDD.n6156 0.005
R6175 AVDD.n6142 AVDD.n5800 0.005
R6176 AVDD.n6142 AVDD.n5799 0.005
R6177 AVDD.n5784 AVDD.n5777 0.005
R6178 AVDD.n5784 AVDD.n5776 0.005
R6179 AVDD.n5767 AVDD.n5763 0.005
R6180 AVDD.n5767 AVDD.n5764 0.005
R6181 AVDD.n4499 AVDD.n4486 0.005
R6182 AVDD.n3478 AVDD.n3467 0.005
R6183 AVDD.n3494 AVDD.n3493 0.005
R6184 AVDD.n4439 AVDD.n4438 0.005
R6185 AVDD.n4515 AVDD.n4514 0.005
R6186 AVDD.n3501 AVDD.n3498 0.005
R6187 AVDD.n76 AVDD.n75 0.005
R6188 AVDD.n123 AVDD.n76 0.005
R6189 AVDD.n6443 AVDD.n6442 0.005
R6190 AVDD.n6490 AVDD.n6443 0.005
R6191 AVDD.n5954 AVDD.n5953 0.005
R6192 AVDD.n6001 AVDD.n5954 0.005
R6193 AVDD.n6506 AVDD.n6505 0.005
R6194 AVDD.n6549 AVDD.n6506 0.005
R6195 AVDD.n192 AVDD.n191 0.005
R6196 AVDD.n239 AVDD.n192 0.005
R6197 AVDD.n254 AVDD.n253 0.005
R6198 AVDD.n297 AVDD.n254 0.005
R6199 AVDD.n700 AVDD.n699 0.005
R6200 AVDD.n701 AVDD.n700 0.005
R6201 AVDD.n435 AVDD.n434 0.005
R6202 AVDD.n436 AVDD.n435 0.005
R6203 AVDD.n374 AVDD.n373 0.005
R6204 AVDD.n421 AVDD.n374 0.005
R6205 AVDD.n442 AVDD.n441 0.005
R6206 AVDD.n485 AVDD.n442 0.005
R6207 AVDD.n636 AVDD.n635 0.005
R6208 AVDD.n679 AVDD.n636 0.005
R6209 AVDD.n6166 AVDD.n6165 0.005
R6210 AVDD.n6184 AVDD.n6166 0.005
R6211 AVDD.n6184 AVDD.n6174 0.005
R6212 AVDD.n6184 AVDD.n6175 0.005
R6213 AVDD.n6179 AVDD.n6178 0.005
R6214 AVDD.n6184 AVDD.n6179 0.005
R6215 AVDD.n6183 AVDD.n6182 0.005
R6216 AVDD.n6184 AVDD.n6183 0.005
R6217 AVDD.n672 AVDD.n671 0.005
R6218 AVDD.n679 AVDD.n672 0.005
R6219 AVDD.n410 AVDD.n409 0.005
R6220 AVDD.n421 AVDD.n410 0.005
R6221 AVDD.n478 AVDD.n477 0.005
R6222 AVDD.n485 AVDD.n478 0.005
R6223 AVDD.n228 AVDD.n227 0.005
R6224 AVDD.n239 AVDD.n228 0.005
R6225 AVDD.n290 AVDD.n289 0.005
R6226 AVDD.n297 AVDD.n290 0.005
R6227 AVDD.n660 AVDD.n659 0.005
R6228 AVDD.n679 AVDD.n660 0.005
R6229 AVDD.n398 AVDD.n397 0.005
R6230 AVDD.n421 AVDD.n398 0.005
R6231 AVDD.n466 AVDD.n465 0.005
R6232 AVDD.n485 AVDD.n466 0.005
R6233 AVDD.n216 AVDD.n215 0.005
R6234 AVDD.n239 AVDD.n216 0.005
R6235 AVDD.n278 AVDD.n277 0.005
R6236 AVDD.n297 AVDD.n278 0.005
R6237 AVDD.n654 AVDD.n653 0.005
R6238 AVDD.n679 AVDD.n654 0.005
R6239 AVDD.n392 AVDD.n391 0.005
R6240 AVDD.n421 AVDD.n392 0.005
R6241 AVDD.n460 AVDD.n459 0.005
R6242 AVDD.n485 AVDD.n460 0.005
R6243 AVDD.n210 AVDD.n209 0.005
R6244 AVDD.n239 AVDD.n210 0.005
R6245 AVDD.n272 AVDD.n271 0.005
R6246 AVDD.n297 AVDD.n272 0.005
R6247 AVDD.n94 AVDD.n93 0.005
R6248 AVDD.n123 AVDD.n94 0.005
R6249 AVDD.n6524 AVDD.n6523 0.005
R6250 AVDD.n6549 AVDD.n6524 0.005
R6251 AVDD.n6461 AVDD.n6460 0.005
R6252 AVDD.n6490 AVDD.n6461 0.005
R6253 AVDD.n5972 AVDD.n5971 0.005
R6254 AVDD.n6001 AVDD.n5972 0.005
R6255 AVDD.n648 AVDD.n647 0.005
R6256 AVDD.n679 AVDD.n648 0.005
R6257 AVDD.n386 AVDD.n385 0.005
R6258 AVDD.n421 AVDD.n386 0.005
R6259 AVDD.n454 AVDD.n453 0.005
R6260 AVDD.n485 AVDD.n454 0.005
R6261 AVDD.n204 AVDD.n203 0.005
R6262 AVDD.n239 AVDD.n204 0.005
R6263 AVDD.n266 AVDD.n265 0.005
R6264 AVDD.n297 AVDD.n266 0.005
R6265 AVDD.n88 AVDD.n87 0.005
R6266 AVDD.n123 AVDD.n88 0.005
R6267 AVDD.n6518 AVDD.n6517 0.005
R6268 AVDD.n6549 AVDD.n6518 0.005
R6269 AVDD.n6455 AVDD.n6454 0.005
R6270 AVDD.n6490 AVDD.n6455 0.005
R6271 AVDD.n5966 AVDD.n5965 0.005
R6272 AVDD.n6001 AVDD.n5966 0.005
R6273 AVDD.n6485 AVDD.n6484 0.005
R6274 AVDD.n6490 AVDD.n6485 0.005
R6275 AVDD.n5996 AVDD.n5995 0.005
R6276 AVDD.n6001 AVDD.n5996 0.005
R6277 AVDD.n118 AVDD.n117 0.005
R6278 AVDD.n123 AVDD.n118 0.005
R6279 AVDD.n6548 AVDD.n6547 0.005
R6280 AVDD.n6549 AVDD.n6548 0.005
R6281 AVDD.n234 AVDD.n233 0.005
R6282 AVDD.n239 AVDD.n234 0.005
R6283 AVDD.n296 AVDD.n295 0.005
R6284 AVDD.n297 AVDD.n296 0.005
R6285 AVDD.n416 AVDD.n415 0.005
R6286 AVDD.n421 AVDD.n416 0.005
R6287 AVDD.n484 AVDD.n483 0.005
R6288 AVDD.n485 AVDD.n484 0.005
R6289 AVDD.n678 AVDD.n677 0.005
R6290 AVDD.n679 AVDD.n678 0.005
R6291 AVDD.n6184 AVDD.n6168 0.005
R6292 AVDD.n6173 AVDD.n6172 0.005
R6293 AVDD.n6184 AVDD.n6173 0.005
R6294 AVDD.n6467 AVDD.n6466 0.005
R6295 AVDD.n6490 AVDD.n6467 0.005
R6296 AVDD.n5978 AVDD.n5977 0.005
R6297 AVDD.n6001 AVDD.n5978 0.005
R6298 AVDD.n100 AVDD.n99 0.005
R6299 AVDD.n123 AVDD.n100 0.005
R6300 AVDD.n6530 AVDD.n6529 0.005
R6301 AVDD.n6549 AVDD.n6530 0.005
R6302 AVDD.n6473 AVDD.n6472 0.005
R6303 AVDD.n6490 AVDD.n6473 0.005
R6304 AVDD.n5984 AVDD.n5983 0.005
R6305 AVDD.n6001 AVDD.n5984 0.005
R6306 AVDD.n106 AVDD.n105 0.005
R6307 AVDD.n123 AVDD.n106 0.005
R6308 AVDD.n6536 AVDD.n6535 0.005
R6309 AVDD.n6549 AVDD.n6536 0.005
R6310 AVDD.n222 AVDD.n221 0.005
R6311 AVDD.n239 AVDD.n222 0.005
R6312 AVDD.n284 AVDD.n283 0.005
R6313 AVDD.n297 AVDD.n284 0.005
R6314 AVDD.n404 AVDD.n403 0.005
R6315 AVDD.n421 AVDD.n404 0.005
R6316 AVDD.n472 AVDD.n471 0.005
R6317 AVDD.n485 AVDD.n472 0.005
R6318 AVDD.n666 AVDD.n665 0.005
R6319 AVDD.n679 AVDD.n666 0.005
R6320 AVDD.n6479 AVDD.n6478 0.005
R6321 AVDD.n6490 AVDD.n6479 0.005
R6322 AVDD.n5990 AVDD.n5989 0.005
R6323 AVDD.n6001 AVDD.n5990 0.005
R6324 AVDD.n112 AVDD.n111 0.005
R6325 AVDD.n123 AVDD.n112 0.005
R6326 AVDD.n6542 AVDD.n6541 0.005
R6327 AVDD.n6549 AVDD.n6542 0.005
R6328 AVDD.n6105 AVDD.n6104 0.005
R6329 AVDD.n6138 AVDD.n6137 0.005
R6330 AVDD.n6046 AVDD.n6045 0.005
R6331 AVDD.n6051 AVDD.n6046 0.005
R6332 AVDD.n6105 AVDD.n6103 0.005
R6333 AVDD.n6138 AVDD.n6136 0.005
R6334 AVDD.n6040 AVDD.n6039 0.005
R6335 AVDD.n6051 AVDD.n6040 0.005
R6336 AVDD.n6102 AVDD.n6101 0.005
R6337 AVDD.n6105 AVDD.n6102 0.005
R6338 AVDD.n6138 AVDD.n6135 0.005
R6339 AVDD.n6034 AVDD.n6033 0.005
R6340 AVDD.n6051 AVDD.n6034 0.005
R6341 AVDD.n6098 AVDD.n6097 0.005
R6342 AVDD.n6105 AVDD.n6098 0.005
R6343 AVDD.n6138 AVDD.n6134 0.005
R6344 AVDD.n6028 AVDD.n6027 0.005
R6345 AVDD.n6051 AVDD.n6028 0.005
R6346 AVDD.n6105 AVDD.n6094 0.005
R6347 AVDD.n6138 AVDD.n6133 0.005
R6348 AVDD.n6022 AVDD.n6021 0.005
R6349 AVDD.n6051 AVDD.n6022 0.005
R6350 AVDD.n6105 AVDD.n6093 0.005
R6351 AVDD.n6132 AVDD.n6131 0.005
R6352 AVDD.n6138 AVDD.n6132 0.005
R6353 AVDD.n6016 AVDD.n6015 0.005
R6354 AVDD.n6051 AVDD.n6016 0.005
R6355 AVDD.n6010 AVDD.n6009 0.005
R6356 AVDD.n6051 AVDD.n6010 0.005
R6357 AVDD.n6184 AVDD.n6167 0.005
R6358 AVDD.n6105 AVDD.n6091 0.005
R6359 AVDD.n6126 AVDD.n6125 0.005
R6360 AVDD.n6138 AVDD.n6126 0.005
R6361 AVDD.n6004 AVDD.n6003 0.005
R6362 AVDD.n6051 AVDD.n6004 0.005
R6363 AVDD.n6105 AVDD.n6092 0.005
R6364 AVDD.n6138 AVDD.n6127 0.005
R6365 AVDD.n6449 AVDD.n6448 0.005
R6366 AVDD.n6490 AVDD.n6449 0.005
R6367 AVDD.n5960 AVDD.n5959 0.005
R6368 AVDD.n6001 AVDD.n5960 0.005
R6369 AVDD.n82 AVDD.n81 0.005
R6370 AVDD.n123 AVDD.n82 0.005
R6371 AVDD.n6512 AVDD.n6511 0.005
R6372 AVDD.n6549 AVDD.n6512 0.005
R6373 AVDD.n198 AVDD.n197 0.005
R6374 AVDD.n239 AVDD.n198 0.005
R6375 AVDD.n260 AVDD.n259 0.005
R6376 AVDD.n297 AVDD.n260 0.005
R6377 AVDD.n380 AVDD.n379 0.005
R6378 AVDD.n421 AVDD.n380 0.005
R6379 AVDD.n448 AVDD.n447 0.005
R6380 AVDD.n485 AVDD.n448 0.005
R6381 AVDD.n642 AVDD.n641 0.005
R6382 AVDD.n679 AVDD.n642 0.005
R6383 AVDD.n574 AVDD.n573 0.005
R6384 AVDD.n621 AVDD.n574 0.005
R6385 AVDD.n755 AVDD.n754 0.005
R6386 AVDD.n802 AVDD.n755 0.005
R6387 AVDD.n817 AVDD.n816 0.005
R6388 AVDD.n860 AVDD.n817 0.005
R6389 AVDD.n936 AVDD.n935 0.005
R6390 AVDD.n983 AVDD.n936 0.005
R6391 AVDD.n998 AVDD.n997 0.005
R6392 AVDD.n1041 AVDD.n998 0.005
R6393 AVDD.n1297 AVDD.n1296 0.005
R6394 AVDD.n1344 AVDD.n1297 0.005
R6395 AVDD.n1103 AVDD.n1102 0.005
R6396 AVDD.n1146 AVDD.n1103 0.005
R6397 AVDD.n4571 AVDD.n4570 0.005
R6398 AVDD.n4583 AVDD.n4571 0.005
R6399 AVDD.n4501 AVDD.n4459 0.005
R6400 AVDD.n4747 AVDD.n4746 0.005
R6401 AVDD.n4758 AVDD.n4747 0.005
R6402 AVDD.n4972 AVDD.n4971 0.005
R6403 AVDD.n4979 AVDD.n4972 0.005
R6404 AVDD.n3317 AVDD.n3316 0.005
R6405 AVDD.n3328 AVDD.n3317 0.005
R6406 AVDD.n3382 AVDD.n3381 0.005
R6407 AVDD.n3389 AVDD.n3382 0.005
R6408 AVDD.n3098 AVDD.n3097 0.005
R6409 AVDD.n3109 AVDD.n3098 0.005
R6410 AVDD.n3208 AVDD.n3207 0.005
R6411 AVDD.n3215 AVDD.n3208 0.005
R6412 AVDD.n2917 AVDD.n2916 0.005
R6413 AVDD.n2928 AVDD.n2917 0.005
R6414 AVDD.n2983 AVDD.n2982 0.005
R6415 AVDD.n2990 AVDD.n2983 0.005
R6416 AVDD.n2754 AVDD.n2753 0.005
R6417 AVDD.n2765 AVDD.n2754 0.005
R6418 AVDD.n2821 AVDD.n2820 0.005
R6419 AVDD.n2828 AVDD.n2821 0.005
R6420 AVDD.n2509 AVDD.n2508 0.005
R6421 AVDD.n2520 AVDD.n2509 0.005
R6422 AVDD.n2603 AVDD.n2602 0.005
R6423 AVDD.n2610 AVDD.n2603 0.005
R6424 AVDD.n2329 AVDD.n2328 0.005
R6425 AVDD.n2340 AVDD.n2329 0.005
R6426 AVDD.n2439 AVDD.n2438 0.005
R6427 AVDD.n2446 AVDD.n2439 0.005
R6428 AVDD.n2228 AVDD.n2227 0.005
R6429 AVDD.n2239 AVDD.n2228 0.005
R6430 AVDD.n2103 AVDD.n2102 0.005
R6431 AVDD.n2110 AVDD.n2103 0.005
R6432 AVDD.n1957 AVDD.n1956 0.005
R6433 AVDD.n1968 AVDD.n1957 0.005
R6434 AVDD.n2024 AVDD.n2023 0.005
R6435 AVDD.n2031 AVDD.n2024 0.005
R6436 AVDD.n1696 AVDD.n1695 0.005
R6437 AVDD.n1707 AVDD.n1696 0.005
R6438 AVDD.n1812 AVDD.n1811 0.005
R6439 AVDD.n1819 AVDD.n1812 0.005
R6440 AVDD.n1515 AVDD.n1514 0.005
R6441 AVDD.n1526 AVDD.n1515 0.005
R6442 AVDD.n1603 AVDD.n1602 0.005
R6443 AVDD.n1610 AVDD.n1603 0.005
R6444 AVDD.n1240 AVDD.n1239 0.005
R6445 AVDD.n1251 AVDD.n1240 0.005
R6446 AVDD.n1399 AVDD.n1398 0.005
R6447 AVDD.n1406 AVDD.n1399 0.005
R6448 AVDD.n1333 AVDD.n1332 0.005
R6449 AVDD.n1344 AVDD.n1333 0.005
R6450 AVDD.n1139 AVDD.n1138 0.005
R6451 AVDD.n1146 AVDD.n1139 0.005
R6452 AVDD.n972 AVDD.n971 0.005
R6453 AVDD.n983 AVDD.n972 0.005
R6454 AVDD.n1034 AVDD.n1033 0.005
R6455 AVDD.n1041 AVDD.n1034 0.005
R6456 AVDD.n791 AVDD.n790 0.005
R6457 AVDD.n802 AVDD.n791 0.005
R6458 AVDD.n853 AVDD.n852 0.005
R6459 AVDD.n860 AVDD.n853 0.005
R6460 AVDD.n610 AVDD.n609 0.005
R6461 AVDD.n621 AVDD.n610 0.005
R6462 AVDD.n4741 AVDD.n4740 0.005
R6463 AVDD.n4758 AVDD.n4741 0.005
R6464 AVDD.n4966 AVDD.n4965 0.005
R6465 AVDD.n4979 AVDD.n4966 0.005
R6466 AVDD.n3311 AVDD.n3310 0.005
R6467 AVDD.n3328 AVDD.n3311 0.005
R6468 AVDD.n3376 AVDD.n3375 0.005
R6469 AVDD.n3389 AVDD.n3376 0.005
R6470 AVDD.n3092 AVDD.n3091 0.005
R6471 AVDD.n3109 AVDD.n3092 0.005
R6472 AVDD.n3202 AVDD.n3201 0.005
R6473 AVDD.n3215 AVDD.n3202 0.005
R6474 AVDD.n2911 AVDD.n2910 0.005
R6475 AVDD.n2928 AVDD.n2911 0.005
R6476 AVDD.n2977 AVDD.n2976 0.005
R6477 AVDD.n2990 AVDD.n2977 0.005
R6478 AVDD.n2748 AVDD.n2747 0.005
R6479 AVDD.n2765 AVDD.n2748 0.005
R6480 AVDD.n2815 AVDD.n2814 0.005
R6481 AVDD.n2828 AVDD.n2815 0.005
R6482 AVDD.n4735 AVDD.n4734 0.005
R6483 AVDD.n4758 AVDD.n4735 0.005
R6484 AVDD.n4960 AVDD.n4959 0.005
R6485 AVDD.n4979 AVDD.n4960 0.005
R6486 AVDD.n3305 AVDD.n3304 0.005
R6487 AVDD.n3328 AVDD.n3305 0.005
R6488 AVDD.n3370 AVDD.n3369 0.005
R6489 AVDD.n3389 AVDD.n3370 0.005
R6490 AVDD.n3086 AVDD.n3085 0.005
R6491 AVDD.n3109 AVDD.n3086 0.005
R6492 AVDD.n3196 AVDD.n3195 0.005
R6493 AVDD.n3215 AVDD.n3196 0.005
R6494 AVDD.n2905 AVDD.n2904 0.005
R6495 AVDD.n2928 AVDD.n2905 0.005
R6496 AVDD.n2971 AVDD.n2970 0.005
R6497 AVDD.n2990 AVDD.n2971 0.005
R6498 AVDD.n2742 AVDD.n2741 0.005
R6499 AVDD.n2765 AVDD.n2742 0.005
R6500 AVDD.n2809 AVDD.n2808 0.005
R6501 AVDD.n2828 AVDD.n2809 0.005
R6502 AVDD.n2497 AVDD.n2496 0.005
R6503 AVDD.n2520 AVDD.n2497 0.005
R6504 AVDD.n2591 AVDD.n2590 0.005
R6505 AVDD.n2610 AVDD.n2591 0.005
R6506 AVDD.n2317 AVDD.n2316 0.005
R6507 AVDD.n2340 AVDD.n2317 0.005
R6508 AVDD.n2427 AVDD.n2426 0.005
R6509 AVDD.n2446 AVDD.n2427 0.005
R6510 AVDD.n2216 AVDD.n2215 0.005
R6511 AVDD.n2239 AVDD.n2216 0.005
R6512 AVDD.n2091 AVDD.n2090 0.005
R6513 AVDD.n2110 AVDD.n2091 0.005
R6514 AVDD.n1945 AVDD.n1944 0.005
R6515 AVDD.n1968 AVDD.n1945 0.005
R6516 AVDD.n2012 AVDD.n2011 0.005
R6517 AVDD.n2031 AVDD.n2012 0.005
R6518 AVDD.n1684 AVDD.n1683 0.005
R6519 AVDD.n1707 AVDD.n1684 0.005
R6520 AVDD.n1800 AVDD.n1799 0.005
R6521 AVDD.n1819 AVDD.n1800 0.005
R6522 AVDD.n1503 AVDD.n1502 0.005
R6523 AVDD.n1526 AVDD.n1503 0.005
R6524 AVDD.n1591 AVDD.n1590 0.005
R6525 AVDD.n1610 AVDD.n1591 0.005
R6526 AVDD.n1228 AVDD.n1227 0.005
R6527 AVDD.n1251 AVDD.n1228 0.005
R6528 AVDD.n1387 AVDD.n1386 0.005
R6529 AVDD.n1406 AVDD.n1387 0.005
R6530 AVDD.n1321 AVDD.n1320 0.005
R6531 AVDD.n1344 AVDD.n1321 0.005
R6532 AVDD.n1127 AVDD.n1126 0.005
R6533 AVDD.n1146 AVDD.n1127 0.005
R6534 AVDD.n960 AVDD.n959 0.005
R6535 AVDD.n983 AVDD.n960 0.005
R6536 AVDD.n1022 AVDD.n1021 0.005
R6537 AVDD.n1041 AVDD.n1022 0.005
R6538 AVDD.n779 AVDD.n778 0.005
R6539 AVDD.n802 AVDD.n779 0.005
R6540 AVDD.n841 AVDD.n840 0.005
R6541 AVDD.n860 AVDD.n841 0.005
R6542 AVDD.n598 AVDD.n597 0.005
R6543 AVDD.n621 AVDD.n598 0.005
R6544 AVDD.n4729 AVDD.n4728 0.005
R6545 AVDD.n4758 AVDD.n4729 0.005
R6546 AVDD.n4954 AVDD.n4953 0.005
R6547 AVDD.n4979 AVDD.n4954 0.005
R6548 AVDD.n3299 AVDD.n3298 0.005
R6549 AVDD.n3328 AVDD.n3299 0.005
R6550 AVDD.n3364 AVDD.n3363 0.005
R6551 AVDD.n3389 AVDD.n3364 0.005
R6552 AVDD.n3080 AVDD.n3079 0.005
R6553 AVDD.n3109 AVDD.n3080 0.005
R6554 AVDD.n3190 AVDD.n3189 0.005
R6555 AVDD.n3215 AVDD.n3190 0.005
R6556 AVDD.n2899 AVDD.n2898 0.005
R6557 AVDD.n2928 AVDD.n2899 0.005
R6558 AVDD.n2965 AVDD.n2964 0.005
R6559 AVDD.n2990 AVDD.n2965 0.005
R6560 AVDD.n2736 AVDD.n2735 0.005
R6561 AVDD.n2765 AVDD.n2736 0.005
R6562 AVDD.n2803 AVDD.n2802 0.005
R6563 AVDD.n2828 AVDD.n2803 0.005
R6564 AVDD.n2491 AVDD.n2490 0.005
R6565 AVDD.n2520 AVDD.n2491 0.005
R6566 AVDD.n2585 AVDD.n2584 0.005
R6567 AVDD.n2610 AVDD.n2585 0.005
R6568 AVDD.n2311 AVDD.n2310 0.005
R6569 AVDD.n2340 AVDD.n2311 0.005
R6570 AVDD.n2421 AVDD.n2420 0.005
R6571 AVDD.n2446 AVDD.n2421 0.005
R6572 AVDD.n2210 AVDD.n2209 0.005
R6573 AVDD.n2239 AVDD.n2210 0.005
R6574 AVDD.n2085 AVDD.n2084 0.005
R6575 AVDD.n2110 AVDD.n2085 0.005
R6576 AVDD.n1939 AVDD.n1938 0.005
R6577 AVDD.n1968 AVDD.n1939 0.005
R6578 AVDD.n2006 AVDD.n2005 0.005
R6579 AVDD.n2031 AVDD.n2006 0.005
R6580 AVDD.n1678 AVDD.n1677 0.005
R6581 AVDD.n1707 AVDD.n1678 0.005
R6582 AVDD.n1794 AVDD.n1793 0.005
R6583 AVDD.n1819 AVDD.n1794 0.005
R6584 AVDD.n1497 AVDD.n1496 0.005
R6585 AVDD.n1526 AVDD.n1497 0.005
R6586 AVDD.n1585 AVDD.n1584 0.005
R6587 AVDD.n1610 AVDD.n1585 0.005
R6588 AVDD.n1222 AVDD.n1221 0.005
R6589 AVDD.n1251 AVDD.n1222 0.005
R6590 AVDD.n1381 AVDD.n1380 0.005
R6591 AVDD.n1406 AVDD.n1381 0.005
R6592 AVDD.n1315 AVDD.n1314 0.005
R6593 AVDD.n1344 AVDD.n1315 0.005
R6594 AVDD.n1121 AVDD.n1120 0.005
R6595 AVDD.n1146 AVDD.n1121 0.005
R6596 AVDD.n954 AVDD.n953 0.005
R6597 AVDD.n983 AVDD.n954 0.005
R6598 AVDD.n1016 AVDD.n1015 0.005
R6599 AVDD.n1041 AVDD.n1016 0.005
R6600 AVDD.n773 AVDD.n772 0.005
R6601 AVDD.n802 AVDD.n773 0.005
R6602 AVDD.n835 AVDD.n834 0.005
R6603 AVDD.n860 AVDD.n835 0.005
R6604 AVDD.n592 AVDD.n591 0.005
R6605 AVDD.n621 AVDD.n592 0.005
R6606 AVDD.n4723 AVDD.n4722 0.005
R6607 AVDD.n4758 AVDD.n4723 0.005
R6608 AVDD.n4948 AVDD.n4947 0.005
R6609 AVDD.n4979 AVDD.n4948 0.005
R6610 AVDD.n3293 AVDD.n3292 0.005
R6611 AVDD.n3328 AVDD.n3293 0.005
R6612 AVDD.n3358 AVDD.n3357 0.005
R6613 AVDD.n3389 AVDD.n3358 0.005
R6614 AVDD.n3074 AVDD.n3073 0.005
R6615 AVDD.n3109 AVDD.n3074 0.005
R6616 AVDD.n3184 AVDD.n3183 0.005
R6617 AVDD.n3215 AVDD.n3184 0.005
R6618 AVDD.n2893 AVDD.n2892 0.005
R6619 AVDD.n2928 AVDD.n2893 0.005
R6620 AVDD.n2959 AVDD.n2958 0.005
R6621 AVDD.n2990 AVDD.n2959 0.005
R6622 AVDD.n2730 AVDD.n2729 0.005
R6623 AVDD.n2765 AVDD.n2730 0.005
R6624 AVDD.n2797 AVDD.n2796 0.005
R6625 AVDD.n2828 AVDD.n2797 0.005
R6626 AVDD.n2485 AVDD.n2484 0.005
R6627 AVDD.n2520 AVDD.n2485 0.005
R6628 AVDD.n2579 AVDD.n2578 0.005
R6629 AVDD.n2610 AVDD.n2579 0.005
R6630 AVDD.n2305 AVDD.n2304 0.005
R6631 AVDD.n2340 AVDD.n2305 0.005
R6632 AVDD.n2415 AVDD.n2414 0.005
R6633 AVDD.n2446 AVDD.n2415 0.005
R6634 AVDD.n2204 AVDD.n2203 0.005
R6635 AVDD.n2239 AVDD.n2204 0.005
R6636 AVDD.n2079 AVDD.n2078 0.005
R6637 AVDD.n2110 AVDD.n2079 0.005
R6638 AVDD.n1933 AVDD.n1932 0.005
R6639 AVDD.n1968 AVDD.n1933 0.005
R6640 AVDD.n2000 AVDD.n1999 0.005
R6641 AVDD.n2031 AVDD.n2000 0.005
R6642 AVDD.n1672 AVDD.n1671 0.005
R6643 AVDD.n1707 AVDD.n1672 0.005
R6644 AVDD.n1788 AVDD.n1787 0.005
R6645 AVDD.n1819 AVDD.n1788 0.005
R6646 AVDD.n1491 AVDD.n1490 0.005
R6647 AVDD.n1526 AVDD.n1491 0.005
R6648 AVDD.n1579 AVDD.n1578 0.005
R6649 AVDD.n1610 AVDD.n1579 0.005
R6650 AVDD.n1216 AVDD.n1215 0.005
R6651 AVDD.n1251 AVDD.n1216 0.005
R6652 AVDD.n1375 AVDD.n1374 0.005
R6653 AVDD.n1406 AVDD.n1375 0.005
R6654 AVDD.n1309 AVDD.n1308 0.005
R6655 AVDD.n1344 AVDD.n1309 0.005
R6656 AVDD.n1115 AVDD.n1114 0.005
R6657 AVDD.n1146 AVDD.n1115 0.005
R6658 AVDD.n948 AVDD.n947 0.005
R6659 AVDD.n983 AVDD.n948 0.005
R6660 AVDD.n1010 AVDD.n1009 0.005
R6661 AVDD.n1041 AVDD.n1010 0.005
R6662 AVDD.n767 AVDD.n766 0.005
R6663 AVDD.n802 AVDD.n767 0.005
R6664 AVDD.n829 AVDD.n828 0.005
R6665 AVDD.n860 AVDD.n829 0.005
R6666 AVDD.n586 AVDD.n585 0.005
R6667 AVDD.n621 AVDD.n586 0.005
R6668 AVDD.n4766 AVDD.n4765 0.005
R6669 AVDD.n4807 AVDD.n4766 0.005
R6670 AVDD.n4583 AVDD.n4577 0.005
R6671 AVDD.n4583 AVDD.n4569 0.005
R6672 AVDD.n4467 AVDD.n4466 0.005
R6673 AVDD.n4501 AVDD.n4467 0.005
R6674 AVDD.n4583 AVDD.n4568 0.005
R6675 AVDD.n4473 AVDD.n4472 0.005
R6676 AVDD.n4501 AVDD.n4473 0.005
R6677 AVDD.n4567 AVDD.n4566 0.005
R6678 AVDD.n4583 AVDD.n4567 0.005
R6679 AVDD.n4501 AVDD.n4474 0.005
R6680 AVDD.n4563 AVDD.n4562 0.005
R6681 AVDD.n4583 AVDD.n4563 0.005
R6682 AVDD.n4501 AVDD.n4475 0.005
R6683 AVDD.n616 AVDD.n615 0.005
R6684 AVDD.n621 AVDD.n616 0.005
R6685 AVDD.n797 AVDD.n796 0.005
R6686 AVDD.n802 AVDD.n797 0.005
R6687 AVDD.n859 AVDD.n858 0.005
R6688 AVDD.n860 AVDD.n859 0.005
R6689 AVDD.n978 AVDD.n977 0.005
R6690 AVDD.n983 AVDD.n978 0.005
R6691 AVDD.n1040 AVDD.n1039 0.005
R6692 AVDD.n1041 AVDD.n1040 0.005
R6693 AVDD.n1339 AVDD.n1338 0.005
R6694 AVDD.n1344 AVDD.n1339 0.005
R6695 AVDD.n1145 AVDD.n1144 0.005
R6696 AVDD.n1146 AVDD.n1145 0.005
R6697 AVDD.n1246 AVDD.n1245 0.005
R6698 AVDD.n1251 AVDD.n1246 0.005
R6699 AVDD.n1405 AVDD.n1404 0.005
R6700 AVDD.n1406 AVDD.n1405 0.005
R6701 AVDD.n1521 AVDD.n1520 0.005
R6702 AVDD.n1526 AVDD.n1521 0.005
R6703 AVDD.n1609 AVDD.n1608 0.005
R6704 AVDD.n1610 AVDD.n1609 0.005
R6705 AVDD.n1702 AVDD.n1701 0.005
R6706 AVDD.n1707 AVDD.n1702 0.005
R6707 AVDD.n1818 AVDD.n1817 0.005
R6708 AVDD.n1819 AVDD.n1818 0.005
R6709 AVDD.n1963 AVDD.n1962 0.005
R6710 AVDD.n1968 AVDD.n1963 0.005
R6711 AVDD.n2030 AVDD.n2029 0.005
R6712 AVDD.n2031 AVDD.n2030 0.005
R6713 AVDD.n2234 AVDD.n2233 0.005
R6714 AVDD.n2239 AVDD.n2234 0.005
R6715 AVDD.n2109 AVDD.n2108 0.005
R6716 AVDD.n2110 AVDD.n2109 0.005
R6717 AVDD.n2335 AVDD.n2334 0.005
R6718 AVDD.n2340 AVDD.n2335 0.005
R6719 AVDD.n2445 AVDD.n2444 0.005
R6720 AVDD.n2446 AVDD.n2445 0.005
R6721 AVDD.n2515 AVDD.n2514 0.005
R6722 AVDD.n2520 AVDD.n2515 0.005
R6723 AVDD.n2609 AVDD.n2608 0.005
R6724 AVDD.n2610 AVDD.n2609 0.005
R6725 AVDD.n2760 AVDD.n2759 0.005
R6726 AVDD.n2765 AVDD.n2760 0.005
R6727 AVDD.n2827 AVDD.n2826 0.005
R6728 AVDD.n2828 AVDD.n2827 0.005
R6729 AVDD.n2923 AVDD.n2922 0.005
R6730 AVDD.n2928 AVDD.n2923 0.005
R6731 AVDD.n2989 AVDD.n2988 0.005
R6732 AVDD.n2990 AVDD.n2989 0.005
R6733 AVDD.n3104 AVDD.n3103 0.005
R6734 AVDD.n3109 AVDD.n3104 0.005
R6735 AVDD.n3214 AVDD.n3213 0.005
R6736 AVDD.n3215 AVDD.n3214 0.005
R6737 AVDD.n3323 AVDD.n3322 0.005
R6738 AVDD.n3328 AVDD.n3323 0.005
R6739 AVDD.n3388 AVDD.n3387 0.005
R6740 AVDD.n3389 AVDD.n3388 0.005
R6741 AVDD.n4753 AVDD.n4752 0.005
R6742 AVDD.n4758 AVDD.n4753 0.005
R6743 AVDD.n4978 AVDD.n4977 0.005
R6744 AVDD.n4979 AVDD.n4978 0.005
R6745 AVDD.n4802 AVDD.n4801 0.005
R6746 AVDD.n4807 AVDD.n4802 0.005
R6747 AVDD.n3637 AVDD.n3636 0.005
R6748 AVDD.n4796 AVDD.n4795 0.005
R6749 AVDD.n4807 AVDD.n4796 0.005
R6750 AVDD.n4790 AVDD.n4789 0.005
R6751 AVDD.n4807 AVDD.n4790 0.005
R6752 AVDD.n4784 AVDD.n4783 0.005
R6753 AVDD.n4807 AVDD.n4784 0.005
R6754 AVDD.n4778 AVDD.n4777 0.005
R6755 AVDD.n4807 AVDD.n4778 0.005
R6756 AVDD.n4772 AVDD.n4771 0.005
R6757 AVDD.n4807 AVDD.n4772 0.005
R6758 AVDD.n4463 AVDD.n4462 0.005
R6759 AVDD.n4501 AVDD.n4463 0.005
R6760 AVDD.n604 AVDD.n603 0.005
R6761 AVDD.n621 AVDD.n604 0.005
R6762 AVDD.n785 AVDD.n784 0.005
R6763 AVDD.n802 AVDD.n785 0.005
R6764 AVDD.n847 AVDD.n846 0.005
R6765 AVDD.n860 AVDD.n847 0.005
R6766 AVDD.n966 AVDD.n965 0.005
R6767 AVDD.n983 AVDD.n966 0.005
R6768 AVDD.n1028 AVDD.n1027 0.005
R6769 AVDD.n1041 AVDD.n1028 0.005
R6770 AVDD.n1327 AVDD.n1326 0.005
R6771 AVDD.n1344 AVDD.n1327 0.005
R6772 AVDD.n1133 AVDD.n1132 0.005
R6773 AVDD.n1146 AVDD.n1133 0.005
R6774 AVDD.n1234 AVDD.n1233 0.005
R6775 AVDD.n1251 AVDD.n1234 0.005
R6776 AVDD.n1393 AVDD.n1392 0.005
R6777 AVDD.n1406 AVDD.n1393 0.005
R6778 AVDD.n1509 AVDD.n1508 0.005
R6779 AVDD.n1526 AVDD.n1509 0.005
R6780 AVDD.n1597 AVDD.n1596 0.005
R6781 AVDD.n1610 AVDD.n1597 0.005
R6782 AVDD.n1690 AVDD.n1689 0.005
R6783 AVDD.n1707 AVDD.n1690 0.005
R6784 AVDD.n1806 AVDD.n1805 0.005
R6785 AVDD.n1819 AVDD.n1806 0.005
R6786 AVDD.n1951 AVDD.n1950 0.005
R6787 AVDD.n1968 AVDD.n1951 0.005
R6788 AVDD.n2018 AVDD.n2017 0.005
R6789 AVDD.n2031 AVDD.n2018 0.005
R6790 AVDD.n2222 AVDD.n2221 0.005
R6791 AVDD.n2239 AVDD.n2222 0.005
R6792 AVDD.n2097 AVDD.n2096 0.005
R6793 AVDD.n2110 AVDD.n2097 0.005
R6794 AVDD.n2323 AVDD.n2322 0.005
R6795 AVDD.n2340 AVDD.n2323 0.005
R6796 AVDD.n2433 AVDD.n2432 0.005
R6797 AVDD.n2446 AVDD.n2433 0.005
R6798 AVDD.n2503 AVDD.n2502 0.005
R6799 AVDD.n2520 AVDD.n2503 0.005
R6800 AVDD.n2597 AVDD.n2596 0.005
R6801 AVDD.n2610 AVDD.n2597 0.005
R6802 AVDD.n580 AVDD.n579 0.005
R6803 AVDD.n621 AVDD.n580 0.005
R6804 AVDD.n761 AVDD.n760 0.005
R6805 AVDD.n802 AVDD.n761 0.005
R6806 AVDD.n823 AVDD.n822 0.005
R6807 AVDD.n860 AVDD.n823 0.005
R6808 AVDD.n942 AVDD.n941 0.005
R6809 AVDD.n983 AVDD.n942 0.005
R6810 AVDD.n1004 AVDD.n1003 0.005
R6811 AVDD.n1041 AVDD.n1004 0.005
R6812 AVDD.n1303 AVDD.n1302 0.005
R6813 AVDD.n1344 AVDD.n1303 0.005
R6814 AVDD.n1109 AVDD.n1108 0.005
R6815 AVDD.n1146 AVDD.n1109 0.005
R6816 AVDD.n1210 AVDD.n1209 0.005
R6817 AVDD.n1251 AVDD.n1210 0.005
R6818 AVDD.n1369 AVDD.n1368 0.005
R6819 AVDD.n1406 AVDD.n1369 0.005
R6820 AVDD.n1485 AVDD.n1484 0.005
R6821 AVDD.n1526 AVDD.n1485 0.005
R6822 AVDD.n1573 AVDD.n1572 0.005
R6823 AVDD.n1610 AVDD.n1573 0.005
R6824 AVDD.n1666 AVDD.n1665 0.005
R6825 AVDD.n1707 AVDD.n1666 0.005
R6826 AVDD.n1782 AVDD.n1781 0.005
R6827 AVDD.n1819 AVDD.n1782 0.005
R6828 AVDD.n1927 AVDD.n1926 0.005
R6829 AVDD.n1968 AVDD.n1927 0.005
R6830 AVDD.n1994 AVDD.n1993 0.005
R6831 AVDD.n2031 AVDD.n1994 0.005
R6832 AVDD.n2198 AVDD.n2197 0.005
R6833 AVDD.n2239 AVDD.n2198 0.005
R6834 AVDD.n2073 AVDD.n2072 0.005
R6835 AVDD.n2110 AVDD.n2073 0.005
R6836 AVDD.n2299 AVDD.n2298 0.005
R6837 AVDD.n2340 AVDD.n2299 0.005
R6838 AVDD.n2409 AVDD.n2408 0.005
R6839 AVDD.n2446 AVDD.n2409 0.005
R6840 AVDD.n2479 AVDD.n2478 0.005
R6841 AVDD.n2520 AVDD.n2479 0.005
R6842 AVDD.n2573 AVDD.n2572 0.005
R6843 AVDD.n2610 AVDD.n2573 0.005
R6844 AVDD.n2724 AVDD.n2723 0.005
R6845 AVDD.n2765 AVDD.n2724 0.005
R6846 AVDD.n2791 AVDD.n2790 0.005
R6847 AVDD.n2828 AVDD.n2791 0.005
R6848 AVDD.n2887 AVDD.n2886 0.005
R6849 AVDD.n2928 AVDD.n2887 0.005
R6850 AVDD.n2953 AVDD.n2952 0.005
R6851 AVDD.n2990 AVDD.n2953 0.005
R6852 AVDD.n3068 AVDD.n3067 0.005
R6853 AVDD.n3109 AVDD.n3068 0.005
R6854 AVDD.n3178 AVDD.n3177 0.005
R6855 AVDD.n3215 AVDD.n3178 0.005
R6856 AVDD.n3287 AVDD.n3286 0.005
R6857 AVDD.n3328 AVDD.n3287 0.005
R6858 AVDD.n3352 AVDD.n3351 0.005
R6859 AVDD.n3389 AVDD.n3352 0.005
R6860 AVDD.n4717 AVDD.n4716 0.005
R6861 AVDD.n4758 AVDD.n4717 0.005
R6862 AVDD.n4942 AVDD.n4941 0.005
R6863 AVDD.n4979 AVDD.n4942 0.005
R6864 AVDD.n4760 AVDD.n4759 0.005
R6865 AVDD.n4807 AVDD.n4760 0.005
R6866 AVDD.n4711 AVDD.n4710 0.005
R6867 AVDD.n4758 AVDD.n4711 0.005
R6868 AVDD.n3281 AVDD.n3280 0.005
R6869 AVDD.n3328 AVDD.n3281 0.005
R6870 AVDD.n3346 AVDD.n3345 0.005
R6871 AVDD.n3389 AVDD.n3346 0.005
R6872 AVDD.n3062 AVDD.n3061 0.005
R6873 AVDD.n3109 AVDD.n3062 0.005
R6874 AVDD.n3172 AVDD.n3171 0.005
R6875 AVDD.n3215 AVDD.n3172 0.005
R6876 AVDD.n2881 AVDD.n2880 0.005
R6877 AVDD.n2928 AVDD.n2881 0.005
R6878 AVDD.n2947 AVDD.n2946 0.005
R6879 AVDD.n2990 AVDD.n2947 0.005
R6880 AVDD.n2718 AVDD.n2717 0.005
R6881 AVDD.n2765 AVDD.n2718 0.005
R6882 AVDD.n2785 AVDD.n2784 0.005
R6883 AVDD.n2828 AVDD.n2785 0.005
R6884 AVDD.n2473 AVDD.n2472 0.005
R6885 AVDD.n2520 AVDD.n2473 0.005
R6886 AVDD.n2567 AVDD.n2566 0.005
R6887 AVDD.n2610 AVDD.n2567 0.005
R6888 AVDD.n2293 AVDD.n2292 0.005
R6889 AVDD.n2340 AVDD.n2293 0.005
R6890 AVDD.n2403 AVDD.n2402 0.005
R6891 AVDD.n2446 AVDD.n2403 0.005
R6892 AVDD.n2192 AVDD.n2191 0.005
R6893 AVDD.n2239 AVDD.n2192 0.005
R6894 AVDD.n2067 AVDD.n2066 0.005
R6895 AVDD.n2110 AVDD.n2067 0.005
R6896 AVDD.n1921 AVDD.n1920 0.005
R6897 AVDD.n1968 AVDD.n1921 0.005
R6898 AVDD.n1988 AVDD.n1987 0.005
R6899 AVDD.n2031 AVDD.n1988 0.005
R6900 AVDD.n1660 AVDD.n1659 0.005
R6901 AVDD.n1707 AVDD.n1660 0.005
R6902 AVDD.n1776 AVDD.n1775 0.005
R6903 AVDD.n1819 AVDD.n1776 0.005
R6904 AVDD.n1479 AVDD.n1478 0.005
R6905 AVDD.n1526 AVDD.n1479 0.005
R6906 AVDD.n1567 AVDD.n1566 0.005
R6907 AVDD.n1610 AVDD.n1567 0.005
R6908 AVDD.n1204 AVDD.n1203 0.005
R6909 AVDD.n1251 AVDD.n1204 0.005
R6910 AVDD.n1363 AVDD.n1362 0.005
R6911 AVDD.n1406 AVDD.n1363 0.005
R6912 AVDD.n4936 AVDD.n4935 0.005
R6913 AVDD.n4979 AVDD.n4936 0.005
R6914 AVDD.n4576 AVDD.n4575 0.005
R6915 AVDD.n4583 AVDD.n4576 0.005
R6916 AVDD.n4501 AVDD.n4458 0.005
R6917 AVDD.n3637 AVDD.n3581 0.005
R6918 AVDD.n3589 AVDD.n3588 0.005
R6919 AVDD.n3637 AVDD.n3589 0.005
R6920 AVDD.n3597 AVDD.n3596 0.005
R6921 AVDD.n3637 AVDD.n3597 0.005
R6922 AVDD.n3605 AVDD.n3604 0.005
R6923 AVDD.n3637 AVDD.n3605 0.005
R6924 AVDD.n3613 AVDD.n3612 0.005
R6925 AVDD.n3637 AVDD.n3613 0.005
R6926 AVDD.n3621 AVDD.n3620 0.005
R6927 AVDD.n3637 AVDD.n3621 0.005
R6928 AVDD.n3629 AVDD.n3628 0.005
R6929 AVDD.n3637 AVDD.n3629 0.005
R6930 AVDD.n4484 AVDD.n4483 0.005
R6931 AVDD.n4501 AVDD.n4484 0.005
R6932 AVDD.n4583 AVDD.n4580 0.005
R6933 AVDD.n4212 AVDD.n4211 0.004
R6934 AVDD.n4344 AVDD.n4343 0.004
R6935 AVDD.n4218 AVDD.n4217 0.004
R6936 AVDD.n4411 AVDD.n3983 0.004
R6937 AVDD.n4908 AVDD.n4907 0.004
R6938 AVDD.n3460 AVDD.n3459 0.004
R6939 AVDD.n4603 AVDD.n4602 0.004
R6940 AVDD.n4598 AVDD.n3466 0.004
R6941 AVDD.n6087 AVDD.n6086 0.004
R6942 AVDD.t35 AVDD.n6087 0.004
R6943 AVDD.n6089 AVDD.n6088 0.004
R6944 AVDD.t35 AVDD.n6089 0.004
R6945 AVDD.n6064 AVDD.n6063 0.004
R6946 AVDD.t344 AVDD.n6064 0.004
R6947 AVDD.n6066 AVDD.n6065 0.004
R6948 AVDD.t344 AVDD.n6066 0.004
R6949 AVDD.n6421 AVDD.n6420 0.004
R6950 AVDD.n6422 AVDD.n6421 0.004
R6951 AVDD.n138 AVDD.n66 0.003
R6952 AVDD.n6496 AVDD.n6492 0.003
R6953 AVDD.n2059 AVDD.n2056 0.003
R6954 AVDD.n5351 AVDD.n5350 0.003
R6955 AVDD.n5410 AVDD.n5409 0.003
R6956 AVDD.n6394 AVDD.n6392 0.003
R6957 AVDD.n62 AVDD.n61 0.003
R6958 AVDD.n5657 AVDD.n62 0.003
R6959 AVDD.n64 AVDD.n63 0.003
R6960 AVDD.n5657 AVDD.n64 0.003
R6961 AVDD.n5670 AVDD.n5669 0.003
R6962 AVDD.n6359 AVDD.n5670 0.003
R6963 AVDD.n5668 AVDD.n5667 0.003
R6964 AVDD.n6359 AVDD.n5668 0.003
R6965 AVDD.n180 AVDD.n179 0.003
R6966 AVDD.n5650 AVDD.n180 0.003
R6967 AVDD.n182 AVDD.n181 0.003
R6968 AVDD.n5650 AVDD.n182 0.003
R6969 AVDD.n548 AVDD.n547 0.003
R6970 AVDD.n5635 AVDD.n548 0.003
R6971 AVDD.n550 AVDD.n549 0.003
R6972 AVDD.n5635 AVDD.n550 0.003
R6973 AVDD.n358 AVDD.n357 0.003
R6974 AVDD.n5642 AVDD.n358 0.003
R6975 AVDD.n360 AVDD.n359 0.003
R6976 AVDD.n5642 AVDD.n360 0.003
R6977 AVDD.n5666 AVDD.n5665 0.003
R6978 AVDD.n6359 AVDD.n5666 0.003
R6979 AVDD.n524 AVDD.n523 0.003
R6980 AVDD.n5635 AVDD.n524 0.003
R6981 AVDD.n526 AVDD.n525 0.003
R6982 AVDD.n5635 AVDD.n526 0.003
R6983 AVDD.n334 AVDD.n333 0.003
R6984 AVDD.n5642 AVDD.n334 0.003
R6985 AVDD.n336 AVDD.n335 0.003
R6986 AVDD.n5642 AVDD.n336 0.003
R6987 AVDD.n156 AVDD.n155 0.003
R6988 AVDD.n5650 AVDD.n156 0.003
R6989 AVDD.n158 AVDD.n157 0.003
R6990 AVDD.n5650 AVDD.n158 0.003
R6991 AVDD.n532 AVDD.n531 0.003
R6992 AVDD.n5635 AVDD.n532 0.003
R6993 AVDD.n534 AVDD.n533 0.003
R6994 AVDD.n5635 AVDD.n534 0.003
R6995 AVDD.n342 AVDD.n341 0.003
R6996 AVDD.n5642 AVDD.n342 0.003
R6997 AVDD.n344 AVDD.n343 0.003
R6998 AVDD.n5642 AVDD.n344 0.003
R6999 AVDD.n164 AVDD.n163 0.003
R7000 AVDD.n5650 AVDD.n164 0.003
R7001 AVDD.n166 AVDD.n165 0.003
R7002 AVDD.n5650 AVDD.n166 0.003
R7003 AVDD.n536 AVDD.n535 0.003
R7004 AVDD.n5635 AVDD.n536 0.003
R7005 AVDD.n538 AVDD.n537 0.003
R7006 AVDD.n5635 AVDD.n538 0.003
R7007 AVDD.n346 AVDD.n345 0.003
R7008 AVDD.n5642 AVDD.n346 0.003
R7009 AVDD.n348 AVDD.n347 0.003
R7010 AVDD.n5642 AVDD.n348 0.003
R7011 AVDD.n168 AVDD.n167 0.003
R7012 AVDD.n5650 AVDD.n168 0.003
R7013 AVDD.n170 AVDD.n169 0.003
R7014 AVDD.n5650 AVDD.n170 0.003
R7015 AVDD.n50 AVDD.n49 0.003
R7016 AVDD.n5657 AVDD.n50 0.003
R7017 AVDD.n52 AVDD.n51 0.003
R7018 AVDD.n5657 AVDD.n52 0.003
R7019 AVDD.n5682 AVDD.n5681 0.003
R7020 AVDD.n6359 AVDD.n5682 0.003
R7021 AVDD.n5680 AVDD.n5679 0.003
R7022 AVDD.n6359 AVDD.n5680 0.003
R7023 AVDD.n540 AVDD.n539 0.003
R7024 AVDD.n5635 AVDD.n540 0.003
R7025 AVDD.n542 AVDD.n541 0.003
R7026 AVDD.n5635 AVDD.n542 0.003
R7027 AVDD.n350 AVDD.n349 0.003
R7028 AVDD.n5642 AVDD.n350 0.003
R7029 AVDD.n352 AVDD.n351 0.003
R7030 AVDD.n5642 AVDD.n352 0.003
R7031 AVDD.n172 AVDD.n171 0.003
R7032 AVDD.n5650 AVDD.n172 0.003
R7033 AVDD.n174 AVDD.n173 0.003
R7034 AVDD.n5650 AVDD.n174 0.003
R7035 AVDD.n54 AVDD.n53 0.003
R7036 AVDD.n5657 AVDD.n54 0.003
R7037 AVDD.n56 AVDD.n55 0.003
R7038 AVDD.n5657 AVDD.n56 0.003
R7039 AVDD.n5678 AVDD.n5677 0.003
R7040 AVDD.n6359 AVDD.n5678 0.003
R7041 AVDD.n5676 AVDD.n5675 0.003
R7042 AVDD.n6359 AVDD.n5676 0.003
R7043 AVDD.n5696 AVDD.n5695 0.003
R7044 AVDD.n6359 AVDD.n5696 0.003
R7045 AVDD.n36 AVDD.n35 0.003
R7046 AVDD.n5657 AVDD.n36 0.003
R7047 AVDD.n34 AVDD.n33 0.003
R7048 AVDD.n5657 AVDD.n34 0.003
R7049 AVDD.n154 AVDD.n153 0.003
R7050 AVDD.n5650 AVDD.n154 0.003
R7051 AVDD.n152 AVDD.n151 0.003
R7052 AVDD.n5650 AVDD.n152 0.003
R7053 AVDD.n332 AVDD.n331 0.003
R7054 AVDD.n5642 AVDD.n332 0.003
R7055 AVDD.n330 AVDD.n329 0.003
R7056 AVDD.n5642 AVDD.n330 0.003
R7057 AVDD.n522 AVDD.n521 0.003
R7058 AVDD.n5635 AVDD.n522 0.003
R7059 AVDD.n520 AVDD.n519 0.003
R7060 AVDD.n5635 AVDD.n520 0.003
R7061 AVDD.n5686 AVDD.n5685 0.003
R7062 AVDD.n6359 AVDD.n5686 0.003
R7063 AVDD.n5684 AVDD.n5683 0.003
R7064 AVDD.n6359 AVDD.n5684 0.003
R7065 AVDD.n46 AVDD.n45 0.003
R7066 AVDD.n5657 AVDD.n46 0.003
R7067 AVDD.n48 AVDD.n47 0.003
R7068 AVDD.n5657 AVDD.n48 0.003
R7069 AVDD.n5690 AVDD.n5689 0.003
R7070 AVDD.n6359 AVDD.n5690 0.003
R7071 AVDD.n5688 AVDD.n5687 0.003
R7072 AVDD.n6359 AVDD.n5688 0.003
R7073 AVDD.n42 AVDD.n41 0.003
R7074 AVDD.n5657 AVDD.n42 0.003
R7075 AVDD.n44 AVDD.n43 0.003
R7076 AVDD.n5657 AVDD.n44 0.003
R7077 AVDD.n160 AVDD.n159 0.003
R7078 AVDD.n5650 AVDD.n160 0.003
R7079 AVDD.n162 AVDD.n161 0.003
R7080 AVDD.n5650 AVDD.n162 0.003
R7081 AVDD.n338 AVDD.n337 0.003
R7082 AVDD.n5642 AVDD.n338 0.003
R7083 AVDD.n340 AVDD.n339 0.003
R7084 AVDD.n5642 AVDD.n340 0.003
R7085 AVDD.n528 AVDD.n527 0.003
R7086 AVDD.n5635 AVDD.n528 0.003
R7087 AVDD.n530 AVDD.n529 0.003
R7088 AVDD.n5635 AVDD.n530 0.003
R7089 AVDD.n5694 AVDD.n5693 0.003
R7090 AVDD.n6359 AVDD.n5694 0.003
R7091 AVDD.n5692 AVDD.n5691 0.003
R7092 AVDD.n6359 AVDD.n5692 0.003
R7093 AVDD.n38 AVDD.n37 0.003
R7094 AVDD.n5657 AVDD.n38 0.003
R7095 AVDD.n40 AVDD.n39 0.003
R7096 AVDD.n5657 AVDD.n40 0.003
R7097 AVDD.n6291 AVDD.n6290 0.003
R7098 AVDD.n6303 AVDD.n6291 0.003
R7099 AVDD.n6357 AVDD.n6356 0.003
R7100 AVDD.n6358 AVDD.n6357 0.003
R7101 AVDD.n6354 AVDD.n6353 0.003
R7102 AVDD.n6358 AVDD.n6354 0.003
R7103 AVDD.n6285 AVDD.n6284 0.003
R7104 AVDD.n6303 AVDD.n6285 0.003
R7105 AVDD.n6268 AVDD.n6267 0.003
R7106 AVDD.n6303 AVDD.n6268 0.003
R7107 AVDD.n6352 AVDD.n6351 0.003
R7108 AVDD.n6358 AVDD.n6352 0.003
R7109 AVDD.n6350 AVDD.n6349 0.003
R7110 AVDD.n6358 AVDD.n6350 0.003
R7111 AVDD.n6262 AVDD.n6261 0.003
R7112 AVDD.n6303 AVDD.n6262 0.003
R7113 AVDD.n6245 AVDD.n6244 0.003
R7114 AVDD.n6303 AVDD.n6245 0.003
R7115 AVDD.n6348 AVDD.n6347 0.003
R7116 AVDD.n6358 AVDD.n6348 0.003
R7117 AVDD.n6346 AVDD.n6345 0.003
R7118 AVDD.n6358 AVDD.n6346 0.003
R7119 AVDD.n6239 AVDD.n6238 0.003
R7120 AVDD.n6303 AVDD.n6239 0.003
R7121 AVDD.n6222 AVDD.n6221 0.003
R7122 AVDD.n6303 AVDD.n6222 0.003
R7123 AVDD.n6344 AVDD.n6343 0.003
R7124 AVDD.n6358 AVDD.n6344 0.003
R7125 AVDD.n6342 AVDD.n6341 0.003
R7126 AVDD.n6358 AVDD.n6342 0.003
R7127 AVDD.n6216 AVDD.n6215 0.003
R7128 AVDD.n6303 AVDD.n6216 0.003
R7129 AVDD.n6199 AVDD.n6198 0.003
R7130 AVDD.n6303 AVDD.n6199 0.003
R7131 AVDD.n6340 AVDD.n6339 0.003
R7132 AVDD.n6358 AVDD.n6340 0.003
R7133 AVDD.n6338 AVDD.n6337 0.003
R7134 AVDD.n6358 AVDD.n6338 0.003
R7135 AVDD.n6193 AVDD.n6192 0.003
R7136 AVDD.n6303 AVDD.n6193 0.003
R7137 AVDD.n6155 AVDD.n6154 0.003
R7138 AVDD.n6303 AVDD.n6155 0.003
R7139 AVDD.n6336 AVDD.n6335 0.003
R7140 AVDD.n6358 AVDD.n6336 0.003
R7141 AVDD.n6334 AVDD.n6333 0.003
R7142 AVDD.n6358 AVDD.n6334 0.003
R7143 AVDD.n6149 AVDD.n6148 0.003
R7144 AVDD.n6303 AVDD.n6149 0.003
R7145 AVDD.n5798 AVDD.n5797 0.003
R7146 AVDD.n6303 AVDD.n5798 0.003
R7147 AVDD.n6332 AVDD.n6331 0.003
R7148 AVDD.n6358 AVDD.n6332 0.003
R7149 AVDD.n6330 AVDD.n6329 0.003
R7150 AVDD.n6358 AVDD.n6330 0.003
R7151 AVDD.n5792 AVDD.n5791 0.003
R7152 AVDD.n6303 AVDD.n5792 0.003
R7153 AVDD.n5756 AVDD.n5755 0.003
R7154 AVDD.n6303 AVDD.n5756 0.003
R7155 AVDD.n5775 AVDD.n5774 0.003
R7156 AVDD.n6303 AVDD.n5775 0.003
R7157 AVDD.n6328 AVDD.n6327 0.003
R7158 AVDD.n6358 AVDD.n6328 0.003
R7159 AVDD.n6326 AVDD.n6325 0.003
R7160 AVDD.n6358 AVDD.n6326 0.003
R7161 AVDD.n5674 AVDD.n5673 0.003
R7162 AVDD.n6359 AVDD.n5674 0.003
R7163 AVDD.n5672 AVDD.n5671 0.003
R7164 AVDD.n6359 AVDD.n5672 0.003
R7165 AVDD.n58 AVDD.n57 0.003
R7166 AVDD.n5657 AVDD.n58 0.003
R7167 AVDD.n60 AVDD.n59 0.003
R7168 AVDD.n5657 AVDD.n60 0.003
R7169 AVDD.n176 AVDD.n175 0.003
R7170 AVDD.n5650 AVDD.n176 0.003
R7171 AVDD.n178 AVDD.n177 0.003
R7172 AVDD.n5650 AVDD.n178 0.003
R7173 AVDD.n354 AVDD.n353 0.003
R7174 AVDD.n5642 AVDD.n354 0.003
R7175 AVDD.n356 AVDD.n355 0.003
R7176 AVDD.n5642 AVDD.n356 0.003
R7177 AVDD.n544 AVDD.n543 0.003
R7178 AVDD.n5635 AVDD.n544 0.003
R7179 AVDD.n546 AVDD.n545 0.003
R7180 AVDD.n5635 AVDD.n546 0.003
R7181 AVDD.n743 AVDD.n742 0.003
R7182 AVDD.n5628 AVDD.n743 0.003
R7183 AVDD.n745 AVDD.n744 0.003
R7184 AVDD.n5628 AVDD.n745 0.003
R7185 AVDD.n924 AVDD.n923 0.003
R7186 AVDD.n5621 AVDD.n924 0.003
R7187 AVDD.n926 AVDD.n925 0.003
R7188 AVDD.n5621 AVDD.n926 0.003
R7189 AVDD.n1095 AVDD.n1094 0.003
R7190 AVDD.n5608 AVDD.n1095 0.003
R7191 AVDD.n1097 AVDD.n1096 0.003
R7192 AVDD.n5608 AVDD.n1097 0.003
R7193 AVDD.n4662 AVDD.n4661 0.003
R7194 AVDD.n4825 AVDD.n4662 0.003
R7195 AVDD.n4897 AVDD.n4896 0.003
R7196 AVDD.n5047 AVDD.n4897 0.003
R7197 AVDD.n4895 AVDD.n4894 0.003
R7198 AVDD.n5047 AVDD.n4895 0.003
R7199 AVDD.n5089 AVDD.n5088 0.003
R7200 AVDD.n5098 AVDD.n5089 0.003
R7201 AVDD.n5087 AVDD.n5086 0.003
R7202 AVDD.n5098 AVDD.n5087 0.003
R7203 AVDD.n5140 AVDD.n5139 0.003
R7204 AVDD.n5149 AVDD.n5140 0.003
R7205 AVDD.n5138 AVDD.n5137 0.003
R7206 AVDD.n5149 AVDD.n5138 0.003
R7207 AVDD.n5191 AVDD.n5190 0.003
R7208 AVDD.n5200 AVDD.n5191 0.003
R7209 AVDD.n5189 AVDD.n5188 0.003
R7210 AVDD.n5200 AVDD.n5189 0.003
R7211 AVDD.n5239 AVDD.n5238 0.003
R7212 AVDD.n5248 AVDD.n5239 0.003
R7213 AVDD.n5237 AVDD.n5236 0.003
R7214 AVDD.n5248 AVDD.n5237 0.003
R7215 AVDD.n5289 AVDD.n5288 0.003
R7216 AVDD.n5301 AVDD.n5289 0.003
R7217 AVDD.n5287 AVDD.n5286 0.003
R7218 AVDD.n5301 AVDD.n5287 0.003
R7219 AVDD.n5340 AVDD.n5339 0.003
R7220 AVDD.n5353 AVDD.n5340 0.003
R7221 AVDD.n5338 AVDD.n5337 0.003
R7222 AVDD.n5353 AVDD.n5338 0.003
R7223 AVDD.n5386 AVDD.n5385 0.003
R7224 AVDD.n5397 AVDD.n5386 0.003
R7225 AVDD.n5384 AVDD.n5383 0.003
R7226 AVDD.n5397 AVDD.n5384 0.003
R7227 AVDD.n5439 AVDD.n5438 0.003
R7228 AVDD.n5450 AVDD.n5439 0.003
R7229 AVDD.n5437 AVDD.n5436 0.003
R7230 AVDD.n5450 AVDD.n5437 0.003
R7231 AVDD.n5490 AVDD.n5489 0.003
R7232 AVDD.n5501 AVDD.n5490 0.003
R7233 AVDD.n5488 AVDD.n5487 0.003
R7234 AVDD.n5501 AVDD.n5488 0.003
R7235 AVDD.n5535 AVDD.n5534 0.003
R7236 AVDD.n5546 AVDD.n5535 0.003
R7237 AVDD.n5533 AVDD.n5532 0.003
R7238 AVDD.n5546 AVDD.n5533 0.003
R7239 AVDD.n5586 AVDD.n5585 0.003
R7240 AVDD.n5597 AVDD.n5586 0.003
R7241 AVDD.n5584 AVDD.n5583 0.003
R7242 AVDD.n5597 AVDD.n5584 0.003
R7243 AVDD.n1071 AVDD.n1070 0.003
R7244 AVDD.n5608 AVDD.n1071 0.003
R7245 AVDD.n1073 AVDD.n1072 0.003
R7246 AVDD.n5608 AVDD.n1073 0.003
R7247 AVDD.n900 AVDD.n899 0.003
R7248 AVDD.n5621 AVDD.n900 0.003
R7249 AVDD.n902 AVDD.n901 0.003
R7250 AVDD.n5621 AVDD.n902 0.003
R7251 AVDD.n719 AVDD.n718 0.003
R7252 AVDD.n5628 AVDD.n719 0.003
R7253 AVDD.n721 AVDD.n720 0.003
R7254 AVDD.n5628 AVDD.n721 0.003
R7255 AVDD.n4893 AVDD.n4892 0.003
R7256 AVDD.n5047 AVDD.n4893 0.003
R7257 AVDD.n4891 AVDD.n4890 0.003
R7258 AVDD.n5047 AVDD.n4891 0.003
R7259 AVDD.n5085 AVDD.n5084 0.003
R7260 AVDD.n5098 AVDD.n5085 0.003
R7261 AVDD.n5083 AVDD.n5082 0.003
R7262 AVDD.n5098 AVDD.n5083 0.003
R7263 AVDD.n5136 AVDD.n5135 0.003
R7264 AVDD.n5149 AVDD.n5136 0.003
R7265 AVDD.n5134 AVDD.n5133 0.003
R7266 AVDD.n5149 AVDD.n5134 0.003
R7267 AVDD.n5187 AVDD.n5186 0.003
R7268 AVDD.n5200 AVDD.n5187 0.003
R7269 AVDD.n5185 AVDD.n5184 0.003
R7270 AVDD.n5200 AVDD.n5185 0.003
R7271 AVDD.n5235 AVDD.n5234 0.003
R7272 AVDD.n5248 AVDD.n5235 0.003
R7273 AVDD.n5233 AVDD.n5232 0.003
R7274 AVDD.n5248 AVDD.n5233 0.003
R7275 AVDD.n4889 AVDD.n4888 0.003
R7276 AVDD.n5047 AVDD.n4889 0.003
R7277 AVDD.n4887 AVDD.n4886 0.003
R7278 AVDD.n5047 AVDD.n4887 0.003
R7279 AVDD.n5081 AVDD.n5080 0.003
R7280 AVDD.n5098 AVDD.n5081 0.003
R7281 AVDD.n5079 AVDD.n5078 0.003
R7282 AVDD.n5098 AVDD.n5079 0.003
R7283 AVDD.n5132 AVDD.n5131 0.003
R7284 AVDD.n5149 AVDD.n5132 0.003
R7285 AVDD.n5130 AVDD.n5129 0.003
R7286 AVDD.n5149 AVDD.n5130 0.003
R7287 AVDD.n5183 AVDD.n5182 0.003
R7288 AVDD.n5200 AVDD.n5183 0.003
R7289 AVDD.n5181 AVDD.n5180 0.003
R7290 AVDD.n5200 AVDD.n5181 0.003
R7291 AVDD.n5231 AVDD.n5230 0.003
R7292 AVDD.n5248 AVDD.n5231 0.003
R7293 AVDD.n5229 AVDD.n5228 0.003
R7294 AVDD.n5248 AVDD.n5229 0.003
R7295 AVDD.n5281 AVDD.n5280 0.003
R7296 AVDD.n5301 AVDD.n5281 0.003
R7297 AVDD.n5279 AVDD.n5278 0.003
R7298 AVDD.n5301 AVDD.n5279 0.003
R7299 AVDD.n5332 AVDD.n5331 0.003
R7300 AVDD.n5353 AVDD.n5332 0.003
R7301 AVDD.n5330 AVDD.n5329 0.003
R7302 AVDD.n5353 AVDD.n5330 0.003
R7303 AVDD.n5378 AVDD.n5377 0.003
R7304 AVDD.n5397 AVDD.n5378 0.003
R7305 AVDD.n5376 AVDD.n5375 0.003
R7306 AVDD.n5397 AVDD.n5376 0.003
R7307 AVDD.n5431 AVDD.n5430 0.003
R7308 AVDD.n5450 AVDD.n5431 0.003
R7309 AVDD.n5429 AVDD.n5428 0.003
R7310 AVDD.n5450 AVDD.n5429 0.003
R7311 AVDD.n5482 AVDD.n5481 0.003
R7312 AVDD.n5501 AVDD.n5482 0.003
R7313 AVDD.n5480 AVDD.n5479 0.003
R7314 AVDD.n5501 AVDD.n5480 0.003
R7315 AVDD.n5527 AVDD.n5526 0.003
R7316 AVDD.n5546 AVDD.n5527 0.003
R7317 AVDD.n5525 AVDD.n5524 0.003
R7318 AVDD.n5546 AVDD.n5525 0.003
R7319 AVDD.n5578 AVDD.n5577 0.003
R7320 AVDD.n5597 AVDD.n5578 0.003
R7321 AVDD.n5576 AVDD.n5575 0.003
R7322 AVDD.n5597 AVDD.n5576 0.003
R7323 AVDD.n1079 AVDD.n1078 0.003
R7324 AVDD.n5608 AVDD.n1079 0.003
R7325 AVDD.n1081 AVDD.n1080 0.003
R7326 AVDD.n5608 AVDD.n1081 0.003
R7327 AVDD.n908 AVDD.n907 0.003
R7328 AVDD.n5621 AVDD.n908 0.003
R7329 AVDD.n910 AVDD.n909 0.003
R7330 AVDD.n5621 AVDD.n910 0.003
R7331 AVDD.n727 AVDD.n726 0.003
R7332 AVDD.n5628 AVDD.n727 0.003
R7333 AVDD.n729 AVDD.n728 0.003
R7334 AVDD.n5628 AVDD.n729 0.003
R7335 AVDD.n4885 AVDD.n4884 0.003
R7336 AVDD.n5047 AVDD.n4885 0.003
R7337 AVDD.n4883 AVDD.n4882 0.003
R7338 AVDD.n5047 AVDD.n4883 0.003
R7339 AVDD.n5077 AVDD.n5076 0.003
R7340 AVDD.n5098 AVDD.n5077 0.003
R7341 AVDD.n5075 AVDD.n5074 0.003
R7342 AVDD.n5098 AVDD.n5075 0.003
R7343 AVDD.n5128 AVDD.n5127 0.003
R7344 AVDD.n5149 AVDD.n5128 0.003
R7345 AVDD.n5126 AVDD.n5125 0.003
R7346 AVDD.n5149 AVDD.n5126 0.003
R7347 AVDD.n5179 AVDD.n5178 0.003
R7348 AVDD.n5200 AVDD.n5179 0.003
R7349 AVDD.n5177 AVDD.n5176 0.003
R7350 AVDD.n5200 AVDD.n5177 0.003
R7351 AVDD.n5227 AVDD.n5226 0.003
R7352 AVDD.n5248 AVDD.n5227 0.003
R7353 AVDD.n5225 AVDD.n5224 0.003
R7354 AVDD.n5248 AVDD.n5225 0.003
R7355 AVDD.n5277 AVDD.n5276 0.003
R7356 AVDD.n5301 AVDD.n5277 0.003
R7357 AVDD.n5275 AVDD.n5274 0.003
R7358 AVDD.n5301 AVDD.n5275 0.003
R7359 AVDD.n5328 AVDD.n5327 0.003
R7360 AVDD.n5353 AVDD.n5328 0.003
R7361 AVDD.n5326 AVDD.n5325 0.003
R7362 AVDD.n5353 AVDD.n5326 0.003
R7363 AVDD.n5374 AVDD.n5373 0.003
R7364 AVDD.n5397 AVDD.n5374 0.003
R7365 AVDD.n5372 AVDD.n5371 0.003
R7366 AVDD.n5397 AVDD.n5372 0.003
R7367 AVDD.n5427 AVDD.n5426 0.003
R7368 AVDD.n5450 AVDD.n5427 0.003
R7369 AVDD.n5425 AVDD.n5424 0.003
R7370 AVDD.n5450 AVDD.n5425 0.003
R7371 AVDD.n5478 AVDD.n5477 0.003
R7372 AVDD.n5501 AVDD.n5478 0.003
R7373 AVDD.n5476 AVDD.n5475 0.003
R7374 AVDD.n5501 AVDD.n5476 0.003
R7375 AVDD.n5523 AVDD.n5522 0.003
R7376 AVDD.n5546 AVDD.n5523 0.003
R7377 AVDD.n5521 AVDD.n5520 0.003
R7378 AVDD.n5546 AVDD.n5521 0.003
R7379 AVDD.n5574 AVDD.n5573 0.003
R7380 AVDD.n5597 AVDD.n5574 0.003
R7381 AVDD.n5572 AVDD.n5571 0.003
R7382 AVDD.n5597 AVDD.n5572 0.003
R7383 AVDD.n1083 AVDD.n1082 0.003
R7384 AVDD.n5608 AVDD.n1083 0.003
R7385 AVDD.n1085 AVDD.n1084 0.003
R7386 AVDD.n5608 AVDD.n1085 0.003
R7387 AVDD.n912 AVDD.n911 0.003
R7388 AVDD.n5621 AVDD.n912 0.003
R7389 AVDD.n914 AVDD.n913 0.003
R7390 AVDD.n5621 AVDD.n914 0.003
R7391 AVDD.n731 AVDD.n730 0.003
R7392 AVDD.n5628 AVDD.n731 0.003
R7393 AVDD.n733 AVDD.n732 0.003
R7394 AVDD.n5628 AVDD.n733 0.003
R7395 AVDD.n4881 AVDD.n4880 0.003
R7396 AVDD.n5047 AVDD.n4881 0.003
R7397 AVDD.n4879 AVDD.n4878 0.003
R7398 AVDD.n5047 AVDD.n4879 0.003
R7399 AVDD.n5073 AVDD.n5072 0.003
R7400 AVDD.n5098 AVDD.n5073 0.003
R7401 AVDD.n5071 AVDD.n5070 0.003
R7402 AVDD.n5098 AVDD.n5071 0.003
R7403 AVDD.n5124 AVDD.n5123 0.003
R7404 AVDD.n5149 AVDD.n5124 0.003
R7405 AVDD.n5122 AVDD.n5121 0.003
R7406 AVDD.n5149 AVDD.n5122 0.003
R7407 AVDD.n5175 AVDD.n5174 0.003
R7408 AVDD.n5200 AVDD.n5175 0.003
R7409 AVDD.n5173 AVDD.n5172 0.003
R7410 AVDD.n5200 AVDD.n5173 0.003
R7411 AVDD.n5223 AVDD.n5222 0.003
R7412 AVDD.n5248 AVDD.n5223 0.003
R7413 AVDD.n5221 AVDD.n5220 0.003
R7414 AVDD.n5248 AVDD.n5221 0.003
R7415 AVDD.n5273 AVDD.n5272 0.003
R7416 AVDD.n5301 AVDD.n5273 0.003
R7417 AVDD.n5271 AVDD.n5270 0.003
R7418 AVDD.n5301 AVDD.n5271 0.003
R7419 AVDD.n5324 AVDD.n5323 0.003
R7420 AVDD.n5353 AVDD.n5324 0.003
R7421 AVDD.n5322 AVDD.n5321 0.003
R7422 AVDD.n5353 AVDD.n5322 0.003
R7423 AVDD.n5370 AVDD.n5369 0.003
R7424 AVDD.n5397 AVDD.n5370 0.003
R7425 AVDD.n5368 AVDD.n5367 0.003
R7426 AVDD.n5397 AVDD.n5368 0.003
R7427 AVDD.n5423 AVDD.n5422 0.003
R7428 AVDD.n5450 AVDD.n5423 0.003
R7429 AVDD.n5421 AVDD.n5420 0.003
R7430 AVDD.n5450 AVDD.n5421 0.003
R7431 AVDD.n5474 AVDD.n5473 0.003
R7432 AVDD.n5501 AVDD.n5474 0.003
R7433 AVDD.n5472 AVDD.n5471 0.003
R7434 AVDD.n5501 AVDD.n5472 0.003
R7435 AVDD.n5519 AVDD.n5518 0.003
R7436 AVDD.n5546 AVDD.n5519 0.003
R7437 AVDD.n5517 AVDD.n5516 0.003
R7438 AVDD.n5546 AVDD.n5517 0.003
R7439 AVDD.n5570 AVDD.n5569 0.003
R7440 AVDD.n5597 AVDD.n5570 0.003
R7441 AVDD.n5568 AVDD.n5567 0.003
R7442 AVDD.n5597 AVDD.n5568 0.003
R7443 AVDD.n1087 AVDD.n1086 0.003
R7444 AVDD.n5608 AVDD.n1087 0.003
R7445 AVDD.n1089 AVDD.n1088 0.003
R7446 AVDD.n5608 AVDD.n1089 0.003
R7447 AVDD.n916 AVDD.n915 0.003
R7448 AVDD.n5621 AVDD.n916 0.003
R7449 AVDD.n918 AVDD.n917 0.003
R7450 AVDD.n5621 AVDD.n918 0.003
R7451 AVDD.n735 AVDD.n734 0.003
R7452 AVDD.n5628 AVDD.n735 0.003
R7453 AVDD.n737 AVDD.n736 0.003
R7454 AVDD.n5628 AVDD.n737 0.003
R7455 AVDD.n3526 AVDD.n3525 0.003
R7456 AVDD.n4597 AVDD.n3526 0.003
R7457 AVDD.n3528 AVDD.n3527 0.003
R7458 AVDD.n4597 AVDD.n3528 0.003
R7459 AVDD.n4666 AVDD.n4665 0.003
R7460 AVDD.n4825 AVDD.n4666 0.003
R7461 AVDD.n4668 AVDD.n4667 0.003
R7462 AVDD.n4825 AVDD.n4668 0.003
R7463 AVDD.n3534 AVDD.n3533 0.003
R7464 AVDD.n4597 AVDD.n3534 0.003
R7465 AVDD.n4660 AVDD.n4659 0.003
R7466 AVDD.n4825 AVDD.n4660 0.003
R7467 AVDD.n717 AVDD.n716 0.003
R7468 AVDD.n5628 AVDD.n717 0.003
R7469 AVDD.n715 AVDD.n714 0.003
R7470 AVDD.n5628 AVDD.n715 0.003
R7471 AVDD.n898 AVDD.n897 0.003
R7472 AVDD.n5621 AVDD.n898 0.003
R7473 AVDD.n896 AVDD.n895 0.003
R7474 AVDD.n5621 AVDD.n896 0.003
R7475 AVDD.n1069 AVDD.n1068 0.003
R7476 AVDD.n5608 AVDD.n1069 0.003
R7477 AVDD.n1067 AVDD.n1066 0.003
R7478 AVDD.n5608 AVDD.n1067 0.003
R7479 AVDD.n5588 AVDD.n5587 0.003
R7480 AVDD.n5597 AVDD.n5588 0.003
R7481 AVDD.n5592 AVDD.n5591 0.003
R7482 AVDD.n5597 AVDD.n5592 0.003
R7483 AVDD.n5537 AVDD.n5536 0.003
R7484 AVDD.n5546 AVDD.n5537 0.003
R7485 AVDD.n5541 AVDD.n5540 0.003
R7486 AVDD.n5546 AVDD.n5541 0.003
R7487 AVDD.n5492 AVDD.n5491 0.003
R7488 AVDD.n5501 AVDD.n5492 0.003
R7489 AVDD.n5496 AVDD.n5495 0.003
R7490 AVDD.n5501 AVDD.n5496 0.003
R7491 AVDD.n5441 AVDD.n5440 0.003
R7492 AVDD.n5450 AVDD.n5441 0.003
R7493 AVDD.n5445 AVDD.n5444 0.003
R7494 AVDD.n5450 AVDD.n5445 0.003
R7495 AVDD.n5388 AVDD.n5387 0.003
R7496 AVDD.n5397 AVDD.n5388 0.003
R7497 AVDD.n5392 AVDD.n5391 0.003
R7498 AVDD.n5397 AVDD.n5392 0.003
R7499 AVDD.n5342 AVDD.n5341 0.003
R7500 AVDD.n5353 AVDD.n5342 0.003
R7501 AVDD.n5346 AVDD.n5345 0.003
R7502 AVDD.n5353 AVDD.n5346 0.003
R7503 AVDD.n5291 AVDD.n5290 0.003
R7504 AVDD.n5301 AVDD.n5291 0.003
R7505 AVDD.n5295 AVDD.n5294 0.003
R7506 AVDD.n5301 AVDD.n5295 0.003
R7507 AVDD.n5241 AVDD.n5240 0.003
R7508 AVDD.n5248 AVDD.n5241 0.003
R7509 AVDD.n5245 AVDD.n5244 0.003
R7510 AVDD.n5248 AVDD.n5245 0.003
R7511 AVDD.n5193 AVDD.n5192 0.003
R7512 AVDD.n5200 AVDD.n5193 0.003
R7513 AVDD.n5197 AVDD.n5196 0.003
R7514 AVDD.n5200 AVDD.n5197 0.003
R7515 AVDD.n5142 AVDD.n5141 0.003
R7516 AVDD.n5149 AVDD.n5142 0.003
R7517 AVDD.n5146 AVDD.n5145 0.003
R7518 AVDD.n5149 AVDD.n5146 0.003
R7519 AVDD.n5091 AVDD.n5090 0.003
R7520 AVDD.n5098 AVDD.n5091 0.003
R7521 AVDD.n5095 AVDD.n5094 0.003
R7522 AVDD.n5098 AVDD.n5095 0.003
R7523 AVDD.n4899 AVDD.n4898 0.003
R7524 AVDD.n5047 AVDD.n4899 0.003
R7525 AVDD.n4903 AVDD.n4902 0.003
R7526 AVDD.n5047 AVDD.n4903 0.003
R7527 AVDD.n4691 AVDD.n4690 0.003
R7528 AVDD.n4825 AVDD.n4691 0.003
R7529 AVDD.n3508 AVDD.n3507 0.003
R7530 AVDD.n4597 AVDD.n3508 0.003
R7531 AVDD.n4688 AVDD.n4687 0.003
R7532 AVDD.n4825 AVDD.n4688 0.003
R7533 AVDD.n3510 AVDD.n3509 0.003
R7534 AVDD.n4597 AVDD.n3510 0.003
R7535 AVDD.n4686 AVDD.n4685 0.003
R7536 AVDD.n4825 AVDD.n4686 0.003
R7537 AVDD.n3512 AVDD.n3511 0.003
R7538 AVDD.n4597 AVDD.n3512 0.003
R7539 AVDD.n4684 AVDD.n4683 0.003
R7540 AVDD.n4825 AVDD.n4684 0.003
R7541 AVDD.n3514 AVDD.n3513 0.003
R7542 AVDD.n4597 AVDD.n3514 0.003
R7543 AVDD.n4682 AVDD.n4681 0.003
R7544 AVDD.n4825 AVDD.n4682 0.003
R7545 AVDD.n3516 AVDD.n3515 0.003
R7546 AVDD.n4597 AVDD.n3516 0.003
R7547 AVDD.n4680 AVDD.n4679 0.003
R7548 AVDD.n4825 AVDD.n4680 0.003
R7549 AVDD.n3518 AVDD.n3517 0.003
R7550 AVDD.n4597 AVDD.n3518 0.003
R7551 AVDD.n4678 AVDD.n4677 0.003
R7552 AVDD.n4825 AVDD.n4678 0.003
R7553 AVDD.n3520 AVDD.n3519 0.003
R7554 AVDD.n4597 AVDD.n3520 0.003
R7555 AVDD.n4676 AVDD.n4675 0.003
R7556 AVDD.n4825 AVDD.n4676 0.003
R7557 AVDD.n3522 AVDD.n3521 0.003
R7558 AVDD.n4597 AVDD.n3522 0.003
R7559 AVDD.n4674 AVDD.n4673 0.003
R7560 AVDD.n4825 AVDD.n4674 0.003
R7561 AVDD.n4672 AVDD.n4671 0.003
R7562 AVDD.n4825 AVDD.n4672 0.003
R7563 AVDD.n3524 AVDD.n3523 0.003
R7564 AVDD.n4597 AVDD.n3524 0.003
R7565 AVDD.n4670 AVDD.n4669 0.003
R7566 AVDD.n4825 AVDD.n4670 0.003
R7567 AVDD.n723 AVDD.n722 0.003
R7568 AVDD.n5628 AVDD.n723 0.003
R7569 AVDD.n725 AVDD.n724 0.003
R7570 AVDD.n5628 AVDD.n725 0.003
R7571 AVDD.n904 AVDD.n903 0.003
R7572 AVDD.n5621 AVDD.n904 0.003
R7573 AVDD.n906 AVDD.n905 0.003
R7574 AVDD.n5621 AVDD.n906 0.003
R7575 AVDD.n1075 AVDD.n1074 0.003
R7576 AVDD.n5608 AVDD.n1075 0.003
R7577 AVDD.n1077 AVDD.n1076 0.003
R7578 AVDD.n5608 AVDD.n1077 0.003
R7579 AVDD.n5582 AVDD.n5581 0.003
R7580 AVDD.n5597 AVDD.n5582 0.003
R7581 AVDD.n5580 AVDD.n5579 0.003
R7582 AVDD.n5597 AVDD.n5580 0.003
R7583 AVDD.n5531 AVDD.n5530 0.003
R7584 AVDD.n5546 AVDD.n5531 0.003
R7585 AVDD.n5529 AVDD.n5528 0.003
R7586 AVDD.n5546 AVDD.n5529 0.003
R7587 AVDD.n5486 AVDD.n5485 0.003
R7588 AVDD.n5501 AVDD.n5486 0.003
R7589 AVDD.n5484 AVDD.n5483 0.003
R7590 AVDD.n5501 AVDD.n5484 0.003
R7591 AVDD.n5435 AVDD.n5434 0.003
R7592 AVDD.n5450 AVDD.n5435 0.003
R7593 AVDD.n5433 AVDD.n5432 0.003
R7594 AVDD.n5450 AVDD.n5433 0.003
R7595 AVDD.n5382 AVDD.n5381 0.003
R7596 AVDD.n5397 AVDD.n5382 0.003
R7597 AVDD.n5380 AVDD.n5379 0.003
R7598 AVDD.n5397 AVDD.n5380 0.003
R7599 AVDD.n5336 AVDD.n5335 0.003
R7600 AVDD.n5353 AVDD.n5336 0.003
R7601 AVDD.n5334 AVDD.n5333 0.003
R7602 AVDD.n5353 AVDD.n5334 0.003
R7603 AVDD.n5285 AVDD.n5284 0.003
R7604 AVDD.n5301 AVDD.n5285 0.003
R7605 AVDD.n5283 AVDD.n5282 0.003
R7606 AVDD.n5301 AVDD.n5283 0.003
R7607 AVDD.n739 AVDD.n738 0.003
R7608 AVDD.n5628 AVDD.n739 0.003
R7609 AVDD.n741 AVDD.n740 0.003
R7610 AVDD.n5628 AVDD.n741 0.003
R7611 AVDD.n920 AVDD.n919 0.003
R7612 AVDD.n5621 AVDD.n920 0.003
R7613 AVDD.n922 AVDD.n921 0.003
R7614 AVDD.n5621 AVDD.n922 0.003
R7615 AVDD.n1091 AVDD.n1090 0.003
R7616 AVDD.n5608 AVDD.n1091 0.003
R7617 AVDD.n1093 AVDD.n1092 0.003
R7618 AVDD.n5608 AVDD.n1093 0.003
R7619 AVDD.n5566 AVDD.n5565 0.003
R7620 AVDD.n5597 AVDD.n5566 0.003
R7621 AVDD.n5564 AVDD.n5563 0.003
R7622 AVDD.n5597 AVDD.n5564 0.003
R7623 AVDD.n5515 AVDD.n5514 0.003
R7624 AVDD.n5546 AVDD.n5515 0.003
R7625 AVDD.n5513 AVDD.n5512 0.003
R7626 AVDD.n5546 AVDD.n5513 0.003
R7627 AVDD.n5470 AVDD.n5469 0.003
R7628 AVDD.n5501 AVDD.n5470 0.003
R7629 AVDD.n5468 AVDD.n5467 0.003
R7630 AVDD.n5501 AVDD.n5468 0.003
R7631 AVDD.n5419 AVDD.n5418 0.003
R7632 AVDD.n5450 AVDD.n5419 0.003
R7633 AVDD.n5417 AVDD.n5416 0.003
R7634 AVDD.n5450 AVDD.n5417 0.003
R7635 AVDD.n5366 AVDD.n5365 0.003
R7636 AVDD.n5397 AVDD.n5366 0.003
R7637 AVDD.n5364 AVDD.n5363 0.003
R7638 AVDD.n5397 AVDD.n5364 0.003
R7639 AVDD.n5320 AVDD.n5319 0.003
R7640 AVDD.n5353 AVDD.n5320 0.003
R7641 AVDD.n5318 AVDD.n5317 0.003
R7642 AVDD.n5353 AVDD.n5318 0.003
R7643 AVDD.n5269 AVDD.n5268 0.003
R7644 AVDD.n5301 AVDD.n5269 0.003
R7645 AVDD.n5267 AVDD.n5266 0.003
R7646 AVDD.n5301 AVDD.n5267 0.003
R7647 AVDD.n5219 AVDD.n5218 0.003
R7648 AVDD.n5248 AVDD.n5219 0.003
R7649 AVDD.n5217 AVDD.n5216 0.003
R7650 AVDD.n5248 AVDD.n5217 0.003
R7651 AVDD.n5171 AVDD.n5170 0.003
R7652 AVDD.n5200 AVDD.n5171 0.003
R7653 AVDD.n5169 AVDD.n5168 0.003
R7654 AVDD.n5200 AVDD.n5169 0.003
R7655 AVDD.n5120 AVDD.n5119 0.003
R7656 AVDD.n5149 AVDD.n5120 0.003
R7657 AVDD.n5118 AVDD.n5117 0.003
R7658 AVDD.n5149 AVDD.n5118 0.003
R7659 AVDD.n5069 AVDD.n5068 0.003
R7660 AVDD.n5098 AVDD.n5069 0.003
R7661 AVDD.n5067 AVDD.n5066 0.003
R7662 AVDD.n5098 AVDD.n5067 0.003
R7663 AVDD.n4877 AVDD.n4876 0.003
R7664 AVDD.n5047 AVDD.n4877 0.003
R7665 AVDD.n4875 AVDD.n4874 0.003
R7666 AVDD.n5047 AVDD.n4875 0.003
R7667 AVDD.n4664 AVDD.n4663 0.003
R7668 AVDD.n4825 AVDD.n4664 0.003
R7669 AVDD.n4873 AVDD.n4872 0.003
R7670 AVDD.n5047 AVDD.n4873 0.003
R7671 AVDD.n4871 AVDD.n4870 0.003
R7672 AVDD.n5047 AVDD.n4871 0.003
R7673 AVDD.n5065 AVDD.n5064 0.003
R7674 AVDD.n5098 AVDD.n5065 0.003
R7675 AVDD.n5063 AVDD.n5062 0.003
R7676 AVDD.n5098 AVDD.n5063 0.003
R7677 AVDD.n5116 AVDD.n5115 0.003
R7678 AVDD.n5149 AVDD.n5116 0.003
R7679 AVDD.n5114 AVDD.n5113 0.003
R7680 AVDD.n5149 AVDD.n5114 0.003
R7681 AVDD.n5167 AVDD.n5166 0.003
R7682 AVDD.n5200 AVDD.n5167 0.003
R7683 AVDD.n5165 AVDD.n5164 0.003
R7684 AVDD.n5200 AVDD.n5165 0.003
R7685 AVDD.n5215 AVDD.n5214 0.003
R7686 AVDD.n5248 AVDD.n5215 0.003
R7687 AVDD.n5213 AVDD.n5212 0.003
R7688 AVDD.n5248 AVDD.n5213 0.003
R7689 AVDD.n5265 AVDD.n5264 0.003
R7690 AVDD.n5301 AVDD.n5265 0.003
R7691 AVDD.n5263 AVDD.n5262 0.003
R7692 AVDD.n5301 AVDD.n5263 0.003
R7693 AVDD.n5316 AVDD.n5315 0.003
R7694 AVDD.n5353 AVDD.n5316 0.003
R7695 AVDD.n5314 AVDD.n5313 0.003
R7696 AVDD.n5353 AVDD.n5314 0.003
R7697 AVDD.n5362 AVDD.n5361 0.003
R7698 AVDD.n5397 AVDD.n5362 0.003
R7699 AVDD.n5360 AVDD.n5359 0.003
R7700 AVDD.n5397 AVDD.n5360 0.003
R7701 AVDD.n5415 AVDD.n5414 0.003
R7702 AVDD.n5450 AVDD.n5415 0.003
R7703 AVDD.n5413 AVDD.n5412 0.003
R7704 AVDD.n5450 AVDD.n5413 0.003
R7705 AVDD.n5466 AVDD.n5465 0.003
R7706 AVDD.n5501 AVDD.n5466 0.003
R7707 AVDD.n5464 AVDD.n5463 0.003
R7708 AVDD.n5501 AVDD.n5464 0.003
R7709 AVDD.n5511 AVDD.n5510 0.003
R7710 AVDD.n5546 AVDD.n5511 0.003
R7711 AVDD.n5509 AVDD.n5508 0.003
R7712 AVDD.n5546 AVDD.n5509 0.003
R7713 AVDD.n5562 AVDD.n5561 0.003
R7714 AVDD.n5597 AVDD.n5562 0.003
R7715 AVDD.n5560 AVDD.n5559 0.003
R7716 AVDD.n5597 AVDD.n5560 0.003
R7717 AVDD.n3530 AVDD.n3529 0.003
R7718 AVDD.n4597 AVDD.n3530 0.003
R7719 AVDD.n3532 AVDD.n3531 0.003
R7720 AVDD.n4597 AVDD.n3532 0.003
R7721 AVDD.n3504 AVDD.n3503 0.003
R7722 AVDD.n4597 AVDD.n3504 0.003
R7723 AVDD.n3506 AVDD.n3505 0.003
R7724 AVDD.n4597 AVDD.n3506 0.003
R7725 AVDD.n4480 AVDD.n4479 0.003
R7726 AVDD.n4315 AVDD.n4312 0.003
R7727 AVDD.n4381 AVDD.n4380 0.002
R7728 AVDD.n4394 AVDD.n4035 0.002
R7729 AVDD.n4408 AVDD.n4407 0.002
R7730 AVDD.n4409 AVDD.n4408 0.002
R7731 AVDD.n6069 level_shifter_up_0.VDD_HV 0.002
R7732 level_shifter_up_4.VDD_HV AVDD.n0 0.002
R7733 AVDD.n1850 AVDD.n1849 0.002
R7734 AVDD.t34 AVDD.n1850 0.002
R7735 AVDD.n1852 AVDD.n1851 0.002
R7736 AVDD.t34 AVDD.n1852 0.002
R7737 AVDD.n1889 AVDD.n1888 0.002
R7738 AVDD.t24 AVDD.n1889 0.002
R7739 AVDD.n1891 AVDD.n1890 0.002
R7740 AVDD.t24 AVDD.n1891 0.002
R7741 AVDD.n2186 AVDD.n2185 0.002
R7742 AVDD.t42 AVDD.n2186 0.002
R7743 AVDD.n2188 AVDD.n2187 0.002
R7744 AVDD.t42 AVDD.n2188 0.002
R7745 AVDD.n2641 AVDD.n2640 0.002
R7746 AVDD.t23 AVDD.n2641 0.002
R7747 AVDD.n2643 AVDD.n2642 0.002
R7748 AVDD.t23 AVDD.n2643 0.002
R7749 AVDD.n2686 AVDD.n2685 0.002
R7750 AVDD.t46 AVDD.n2686 0.002
R7751 AVDD.n2688 AVDD.n2687 0.002
R7752 AVDD.t46 AVDD.n2688 0.002
R7753 AVDD.n3229 AVDD.n3228 0.002
R7754 AVDD.t25 AVDD.n3229 0.002
R7755 AVDD.n3231 AVDD.n3230 0.002
R7756 AVDD.t25 AVDD.n3231 0.002
R7757 AVDD.n3420 AVDD.n3419 0.002
R7758 AVDD.t2 AVDD.n3420 0.002
R7759 AVDD.n3422 AVDD.n3421 0.002
R7760 AVDD.t2 AVDD.n3422 0.002
R7761 AVDD.n4844 AVDD.n4843 0.002
R7762 AVDD.t47 AVDD.n4844 0.002
R7763 AVDD.n4846 AVDD.n4845 0.002
R7764 AVDD.t47 AVDD.n4846 0.002
R7765 AVDD.n1860 AVDD.n1859 0.002
R7766 AVDD.t34 AVDD.n1860 0.002
R7767 AVDD.n1858 AVDD.n1857 0.002
R7768 AVDD.t34 AVDD.n1858 0.002
R7769 AVDD.n1899 AVDD.n1898 0.002
R7770 AVDD.t24 AVDD.n1899 0.002
R7771 AVDD.n1897 AVDD.n1896 0.002
R7772 AVDD.t24 AVDD.n1897 0.002
R7773 AVDD.n2245 AVDD.n2244 0.002
R7774 AVDD.t42 AVDD.n2245 0.002
R7775 AVDD.n2243 AVDD.n2242 0.002
R7776 AVDD.t42 AVDD.n2243 0.002
R7777 AVDD.n2652 AVDD.n2651 0.002
R7778 AVDD.t23 AVDD.n2652 0.002
R7779 AVDD.n2650 AVDD.n2649 0.002
R7780 AVDD.t23 AVDD.n2650 0.002
R7781 AVDD.n2696 AVDD.n2695 0.002
R7782 AVDD.t46 AVDD.n2696 0.002
R7783 AVDD.n2694 AVDD.n2693 0.002
R7784 AVDD.t46 AVDD.n2694 0.002
R7785 AVDD.n3239 AVDD.n3238 0.002
R7786 AVDD.t25 AVDD.n3239 0.002
R7787 AVDD.n3237 AVDD.n3236 0.002
R7788 AVDD.t25 AVDD.n3237 0.002
R7789 AVDD.n3430 AVDD.n3429 0.002
R7790 AVDD.t2 AVDD.n3430 0.002
R7791 AVDD.n3428 AVDD.n3427 0.002
R7792 AVDD.t2 AVDD.n3428 0.002
R7793 AVDD.n4854 AVDD.n4853 0.002
R7794 AVDD.t47 AVDD.n4854 0.002
R7795 AVDD.n4852 AVDD.n4851 0.002
R7796 AVDD.t47 AVDD.n4852 0.002
R7797 AVDD.n1846 AVDD.n1845 0.002
R7798 AVDD.t34 AVDD.n1846 0.002
R7799 AVDD.n1848 AVDD.n1847 0.002
R7800 AVDD.t34 AVDD.n1848 0.002
R7801 AVDD.n1885 AVDD.n1884 0.002
R7802 AVDD.t24 AVDD.n1885 0.002
R7803 AVDD.n1887 AVDD.n1886 0.002
R7804 AVDD.t24 AVDD.n1887 0.002
R7805 AVDD.n2182 AVDD.n2181 0.002
R7806 AVDD.t42 AVDD.n2182 0.002
R7807 AVDD.n2184 AVDD.n2183 0.002
R7808 AVDD.t42 AVDD.n2184 0.002
R7809 AVDD.n2637 AVDD.n2636 0.002
R7810 AVDD.t23 AVDD.n2637 0.002
R7811 AVDD.n2639 AVDD.n2638 0.002
R7812 AVDD.t23 AVDD.n2639 0.002
R7813 AVDD.n2682 AVDD.n2681 0.002
R7814 AVDD.t46 AVDD.n2682 0.002
R7815 AVDD.n2684 AVDD.n2683 0.002
R7816 AVDD.t46 AVDD.n2684 0.002
R7817 AVDD.n3225 AVDD.n3224 0.002
R7818 AVDD.t25 AVDD.n3225 0.002
R7819 AVDD.n3227 AVDD.n3226 0.002
R7820 AVDD.t25 AVDD.n3227 0.002
R7821 AVDD.n3416 AVDD.n3415 0.002
R7822 AVDD.t2 AVDD.n3416 0.002
R7823 AVDD.n3418 AVDD.n3417 0.002
R7824 AVDD.t2 AVDD.n3418 0.002
R7825 AVDD.n4840 AVDD.n4839 0.002
R7826 AVDD.t47 AVDD.n4840 0.002
R7827 AVDD.n4842 AVDD.n4841 0.002
R7828 AVDD.t47 AVDD.n4842 0.002
R7829 AVDD.n1864 AVDD.n1863 0.002
R7830 AVDD.t34 AVDD.n1864 0.002
R7831 AVDD.n1862 AVDD.n1861 0.002
R7832 AVDD.t34 AVDD.n1862 0.002
R7833 AVDD.n1903 AVDD.n1902 0.002
R7834 AVDD.t24 AVDD.n1903 0.002
R7835 AVDD.n1901 AVDD.n1900 0.002
R7836 AVDD.t24 AVDD.n1901 0.002
R7837 AVDD.n2249 AVDD.n2248 0.002
R7838 AVDD.t42 AVDD.n2249 0.002
R7839 AVDD.n2247 AVDD.n2246 0.002
R7840 AVDD.t42 AVDD.n2247 0.002
R7841 AVDD.n2656 AVDD.n2655 0.002
R7842 AVDD.t23 AVDD.n2656 0.002
R7843 AVDD.n2654 AVDD.n2653 0.002
R7844 AVDD.t23 AVDD.n2654 0.002
R7845 AVDD.n2700 AVDD.n2699 0.002
R7846 AVDD.t46 AVDD.n2700 0.002
R7847 AVDD.n2698 AVDD.n2697 0.002
R7848 AVDD.t46 AVDD.n2698 0.002
R7849 AVDD.n3243 AVDD.n3242 0.002
R7850 AVDD.t25 AVDD.n3243 0.002
R7851 AVDD.n3241 AVDD.n3240 0.002
R7852 AVDD.t25 AVDD.n3241 0.002
R7853 AVDD.n3434 AVDD.n3433 0.002
R7854 AVDD.t2 AVDD.n3434 0.002
R7855 AVDD.n3432 AVDD.n3431 0.002
R7856 AVDD.t2 AVDD.n3432 0.002
R7857 AVDD.n4858 AVDD.n4857 0.002
R7858 AVDD.t47 AVDD.n4858 0.002
R7859 AVDD.n4856 AVDD.n4855 0.002
R7860 AVDD.t47 AVDD.n4856 0.002
R7861 AVDD.n1842 AVDD.n1841 0.002
R7862 AVDD.t34 AVDD.n1842 0.002
R7863 AVDD.n1844 AVDD.n1843 0.002
R7864 AVDD.t34 AVDD.n1844 0.002
R7865 AVDD.n1881 AVDD.n1880 0.002
R7866 AVDD.t24 AVDD.n1881 0.002
R7867 AVDD.n1883 AVDD.n1882 0.002
R7868 AVDD.t24 AVDD.n1883 0.002
R7869 AVDD.n2178 AVDD.n2177 0.002
R7870 AVDD.t42 AVDD.n2178 0.002
R7871 AVDD.n2180 AVDD.n2179 0.002
R7872 AVDD.t42 AVDD.n2180 0.002
R7873 AVDD.n2633 AVDD.n2632 0.002
R7874 AVDD.t23 AVDD.n2633 0.002
R7875 AVDD.n2635 AVDD.n2634 0.002
R7876 AVDD.t23 AVDD.n2635 0.002
R7877 AVDD.n2678 AVDD.n2677 0.002
R7878 AVDD.t46 AVDD.n2678 0.002
R7879 AVDD.n2680 AVDD.n2679 0.002
R7880 AVDD.t46 AVDD.n2680 0.002
R7881 AVDD.n3221 AVDD.n3220 0.002
R7882 AVDD.t25 AVDD.n3221 0.002
R7883 AVDD.n3223 AVDD.n3222 0.002
R7884 AVDD.t25 AVDD.n3223 0.002
R7885 AVDD.n3412 AVDD.n3411 0.002
R7886 AVDD.t2 AVDD.n3412 0.002
R7887 AVDD.n3414 AVDD.n3413 0.002
R7888 AVDD.t2 AVDD.n3414 0.002
R7889 AVDD.n4836 AVDD.n4835 0.002
R7890 AVDD.t47 AVDD.n4836 0.002
R7891 AVDD.n4838 AVDD.n4837 0.002
R7892 AVDD.t47 AVDD.n4838 0.002
R7893 AVDD.n1868 AVDD.n1867 0.002
R7894 AVDD.t34 AVDD.n1868 0.002
R7895 AVDD.n1866 AVDD.n1865 0.002
R7896 AVDD.t34 AVDD.n1866 0.002
R7897 AVDD.n1907 AVDD.n1906 0.002
R7898 AVDD.t24 AVDD.n1907 0.002
R7899 AVDD.n1905 AVDD.n1904 0.002
R7900 AVDD.t24 AVDD.n1905 0.002
R7901 AVDD.n2253 AVDD.n2252 0.002
R7902 AVDD.t42 AVDD.n2253 0.002
R7903 AVDD.n2251 AVDD.n2250 0.002
R7904 AVDD.t42 AVDD.n2251 0.002
R7905 AVDD.n2660 AVDD.n2659 0.002
R7906 AVDD.t23 AVDD.n2660 0.002
R7907 AVDD.n2658 AVDD.n2657 0.002
R7908 AVDD.t23 AVDD.n2658 0.002
R7909 AVDD.n2704 AVDD.n2703 0.002
R7910 AVDD.t46 AVDD.n2704 0.002
R7911 AVDD.n2702 AVDD.n2701 0.002
R7912 AVDD.t46 AVDD.n2702 0.002
R7913 AVDD.n3247 AVDD.n3246 0.002
R7914 AVDD.t25 AVDD.n3247 0.002
R7915 AVDD.n3245 AVDD.n3244 0.002
R7916 AVDD.t25 AVDD.n3245 0.002
R7917 AVDD.n3438 AVDD.n3437 0.002
R7918 AVDD.t2 AVDD.n3438 0.002
R7919 AVDD.n3436 AVDD.n3435 0.002
R7920 AVDD.t2 AVDD.n3436 0.002
R7921 AVDD.n4862 AVDD.n4861 0.002
R7922 AVDD.t47 AVDD.n4862 0.002
R7923 AVDD.n4860 AVDD.n4859 0.002
R7924 AVDD.t47 AVDD.n4860 0.002
R7925 AVDD.n1838 AVDD.n1837 0.002
R7926 AVDD.t34 AVDD.n1838 0.002
R7927 AVDD.n1840 AVDD.n1839 0.002
R7928 AVDD.t34 AVDD.n1840 0.002
R7929 AVDD.n1877 AVDD.n1876 0.002
R7930 AVDD.t24 AVDD.n1877 0.002
R7931 AVDD.n1879 AVDD.n1878 0.002
R7932 AVDD.t24 AVDD.n1879 0.002
R7933 AVDD.n2174 AVDD.n2173 0.002
R7934 AVDD.t42 AVDD.n2174 0.002
R7935 AVDD.n2176 AVDD.n2175 0.002
R7936 AVDD.t42 AVDD.n2176 0.002
R7937 AVDD.n2629 AVDD.n2628 0.002
R7938 AVDD.t23 AVDD.n2629 0.002
R7939 AVDD.n2631 AVDD.n2630 0.002
R7940 AVDD.t23 AVDD.n2631 0.002
R7941 AVDD.n2674 AVDD.n2673 0.002
R7942 AVDD.t46 AVDD.n2674 0.002
R7943 AVDD.n2676 AVDD.n2675 0.002
R7944 AVDD.t46 AVDD.n2676 0.002
R7945 AVDD.n3217 AVDD.n3216 0.002
R7946 AVDD.t25 AVDD.n3217 0.002
R7947 AVDD.n3219 AVDD.n3218 0.002
R7948 AVDD.t25 AVDD.n3219 0.002
R7949 AVDD.n3408 AVDD.n3407 0.002
R7950 AVDD.t2 AVDD.n3408 0.002
R7951 AVDD.n3410 AVDD.n3409 0.002
R7952 AVDD.t2 AVDD.n3410 0.002
R7953 AVDD.n4832 AVDD.n4831 0.002
R7954 AVDD.t47 AVDD.n4832 0.002
R7955 AVDD.n4834 AVDD.n4833 0.002
R7956 AVDD.t47 AVDD.n4834 0.002
R7957 AVDD.n1872 AVDD.n1871 0.002
R7958 AVDD.t34 AVDD.n1872 0.002
R7959 AVDD.n1870 AVDD.n1869 0.002
R7960 AVDD.t34 AVDD.n1870 0.002
R7961 AVDD.n1911 AVDD.n1910 0.002
R7962 AVDD.t24 AVDD.n1911 0.002
R7963 AVDD.n1909 AVDD.n1908 0.002
R7964 AVDD.t24 AVDD.n1909 0.002
R7965 AVDD.n2257 AVDD.n2256 0.002
R7966 AVDD.t42 AVDD.n2257 0.002
R7967 AVDD.n2255 AVDD.n2254 0.002
R7968 AVDD.t42 AVDD.n2255 0.002
R7969 AVDD.n2664 AVDD.n2663 0.002
R7970 AVDD.t23 AVDD.n2664 0.002
R7971 AVDD.n2662 AVDD.n2661 0.002
R7972 AVDD.t23 AVDD.n2662 0.002
R7973 AVDD.n2708 AVDD.n2707 0.002
R7974 AVDD.t46 AVDD.n2708 0.002
R7975 AVDD.n2706 AVDD.n2705 0.002
R7976 AVDD.t46 AVDD.n2706 0.002
R7977 AVDD.n3251 AVDD.n3250 0.002
R7978 AVDD.t25 AVDD.n3251 0.002
R7979 AVDD.n3249 AVDD.n3248 0.002
R7980 AVDD.t25 AVDD.n3249 0.002
R7981 AVDD.n3442 AVDD.n3441 0.002
R7982 AVDD.t2 AVDD.n3442 0.002
R7983 AVDD.n3440 AVDD.n3439 0.002
R7984 AVDD.t2 AVDD.n3440 0.002
R7985 AVDD.n4866 AVDD.n4865 0.002
R7986 AVDD.t47 AVDD.n4866 0.002
R7987 AVDD.n4864 AVDD.n4863 0.002
R7988 AVDD.t47 AVDD.n4864 0.002
R7989 AVDD.n4830 AVDD.n4829 0.002
R7990 AVDD.t47 AVDD.n4830 0.002
R7991 AVDD.n3445 AVDD.n3443 0.002
R7992 AVDD.n3443 AVDD.t2 0.002
R7993 AVDD.n3254 AVDD.n3252 0.002
R7994 AVDD.n3252 AVDD.t25 0.002
R7995 AVDD.n2778 AVDD.n2709 0.002
R7996 AVDD.n2709 AVDD.t46 0.002
R7997 AVDD.n2667 AVDD.n2665 0.002
R7998 AVDD.n2665 AVDD.t23 0.002
R7999 AVDD.n2261 AVDD.n2258 0.002
R8000 AVDD.n2258 AVDD.t42 0.002
R8001 AVDD.n1981 AVDD.n1912 0.002
R8002 AVDD.n1912 AVDD.t24 0.002
R8003 AVDD.n1875 AVDD.n1873 0.002
R8004 AVDD.n1873 AVDD.t34 0.002
R8005 AVDD.n1264 AVDD.n1195 0.002
R8006 AVDD.n1195 AVDD.t394 0.002
R8007 AVDD.t394 AVDD.n1176 0.002
R8008 AVDD.t394 AVDD.n1172 0.002
R8009 AVDD.n1178 AVDD.n1177 0.002
R8010 AVDD.t394 AVDD.n1178 0.002
R8011 AVDD.n1180 AVDD.n1179 0.002
R8012 AVDD.t394 AVDD.n1180 0.002
R8013 AVDD.t394 AVDD.n1171 0.002
R8014 AVDD.t394 AVDD.n1170 0.002
R8015 AVDD.n1182 AVDD.n1181 0.002
R8016 AVDD.t394 AVDD.n1182 0.002
R8017 AVDD.n1184 AVDD.n1183 0.002
R8018 AVDD.t394 AVDD.n1184 0.002
R8019 AVDD.t394 AVDD.n1169 0.002
R8020 AVDD.t394 AVDD.n1168 0.002
R8021 AVDD.n1186 AVDD.n1185 0.002
R8022 AVDD.t394 AVDD.n1186 0.002
R8023 AVDD.n1188 AVDD.n1187 0.002
R8024 AVDD.t394 AVDD.n1188 0.002
R8025 AVDD.t394 AVDD.n1167 0.002
R8026 AVDD.t394 AVDD.n1166 0.002
R8027 AVDD.n1191 AVDD.n1190 0.002
R8028 AVDD.t394 AVDD.n1191 0.002
R8029 AVDD.n1264 AVDD.n1263 0.002
R8030 AVDD.t366 AVDD.n3698 0.002
R8031 AVDD.n3681 AVDD.n3680 0.002
R8032 AVDD.t366 AVDD.n3681 0.002
R8033 AVDD.t366 AVDD.n3695 0.002
R8034 AVDD.n3684 AVDD.n3683 0.002
R8035 AVDD.t366 AVDD.n3684 0.002
R8036 AVDD.t366 AVDD.n3692 0.002
R8037 AVDD.n3688 AVDD.n3687 0.002
R8038 AVDD.t366 AVDD.n3688 0.002
R8039 AVDD.t366 AVDD.n3689 0.002
R8040 AVDD.n3424 AVDD.n3423 0.002
R8041 AVDD.t2 AVDD.n3424 0.002
R8042 AVDD.n3233 AVDD.n3232 0.002
R8043 AVDD.t25 AVDD.n3233 0.002
R8044 AVDD.n2690 AVDD.n2689 0.002
R8045 AVDD.t46 AVDD.n2690 0.002
R8046 AVDD.n2646 AVDD.n2645 0.002
R8047 AVDD.t23 AVDD.n2646 0.002
R8048 AVDD.n2190 AVDD.n2189 0.002
R8049 AVDD.t42 AVDD.n2190 0.002
R8050 AVDD.n1176 AVDD.n1175 0.002
R8051 AVDD.n1854 AVDD.n1853 0.002
R8052 AVDD.t34 AVDD.n1854 0.002
R8053 AVDD.n1895 AVDD.n1894 0.002
R8054 AVDD.t24 AVDD.n1895 0.002
R8055 AVDD.n1856 AVDD.n1855 0.002
R8056 AVDD.t34 AVDD.n1856 0.002
R8057 AVDD.n1893 AVDD.n1892 0.002
R8058 AVDD.t24 AVDD.n1893 0.002
R8059 AVDD.n2241 AVDD.n2240 0.002
R8060 AVDD.t42 AVDD.n2241 0.002
R8061 AVDD.n2648 AVDD.n2647 0.002
R8062 AVDD.t23 AVDD.n2648 0.002
R8063 AVDD.n2692 AVDD.n2691 0.002
R8064 AVDD.t46 AVDD.n2692 0.002
R8065 AVDD.n3235 AVDD.n3234 0.002
R8066 AVDD.t25 AVDD.n3235 0.002
R8067 AVDD.n3426 AVDD.n3425 0.002
R8068 AVDD.t2 AVDD.n3426 0.002
R8069 AVDD.n4850 AVDD.n4849 0.002
R8070 AVDD.t47 AVDD.n4850 0.002
R8071 AVDD.n4848 AVDD.n4847 0.002
R8072 AVDD.t47 AVDD.n4848 0.002
R8073 AVDD.n3691 AVDD.n3690 0.002
R8074 AVDD.t366 AVDD.n3691 0.002
R8075 AVDD.t366 AVDD.n3685 0.002
R8076 AVDD.n3694 AVDD.n3693 0.002
R8077 AVDD.t366 AVDD.n3694 0.002
R8078 AVDD.t366 AVDD.n3682 0.002
R8079 AVDD.n3697 AVDD.n3696 0.002
R8080 AVDD.t366 AVDD.n3697 0.002
R8081 AVDD.t47 AVDD.n4869 0.002
R8082 AVDD.n4869 AVDD.n4868 0.002
R8083 AVDD.n3445 AVDD.n3444 0.002
R8084 AVDD.n3254 AVDD.n3253 0.002
R8085 AVDD.n2778 AVDD.n2777 0.002
R8086 AVDD.n2667 AVDD.n2666 0.002
R8087 AVDD.n2261 AVDD.n2260 0.002
R8088 AVDD.n1981 AVDD.n1980 0.002
R8089 AVDD.n1875 AVDD.n1874 0.002
R8090 AVDD.n1193 AVDD.n1192 0.002
R8091 AVDD.t394 AVDD.n1193 0.002
R8092 AVDD.t394 AVDD.n1194 0.002
R8093 AVDD.t394 AVDD.n1173 0.002
R8094 AVDD.t366 AVDD.n3704 0.002
R8095 AVDD.n3703 AVDD.n3702 0.002
R8096 AVDD.t366 AVDD.n3703 0.002
R8097 AVDD.t366 AVDD.n3701 0.002
R8098 AVDD.t366 AVDD.n3700 0.002
R8099 AVDD.n3700 AVDD.n3699 0.002
R8100 AVDD.n3678 AVDD.n3677 0.002
R8101 AVDD.t366 AVDD.n3678 0.002
R8102 AVDD.t366 AVDD.n3679 0.002
R8103 AVDD.t366 AVDD.n3566 0.002
R8104 AVDD.n3566 AVDD.n3565 0.002
R8105 AVDD.t366 AVDD.n3676 0.002
R8106 AVDD.n3676 AVDD.n3675 0.002
R8107 AVDD.n6317 AVDD.n6316 0.002
R8108 AVDD.n6318 AVDD.n6317 0.002
R8109 AVDD.n5815 AVDD.n5814 0.002
R8110 AVDD.n5816 AVDD.n5815 0.002
R8111 AVDD.n5934 AVDD.n5933 0.002
R8112 AVDD.n5935 AVDD.n5934 0.002
R8113 AVDD.n6311 AVDD.n6310 0.002
R8114 AVDD.n6312 AVDD.n6311 0.002
R8115 AVDD.n6323 AVDD.n6322 0.002
R8116 AVDD.n6324 AVDD.n6323 0.002
R8117 AVDD.n4209 AVDD.n4208 0.001
R8118 AVDD.n3838 AVDD.n3837 0.001
R8119 AVDD.n4053 AVDD.n4052 0.001
R8120 AVDD.n5710 AVDD.n5698 0.001
R8121 AVDD.n6307 AVDD.n5714 0.001
R8122 AVDD.t741 AVDD.n3761 0.001
R8123 AVDD.n4574 AVDD.n4573 0.001
R8124 AVDD.n6170 AVDD.n6169 0.001
R8125 AVDD.n6129 AVDD.n6128 0.001
R8126 AVDD.n4212 AVDD.n3983 0.001
R8127 AVDD.n3797 AVDD.n3796 0.001
R8128 AVDD.n3887 AVDD.n3886 0.001
R8129 AVDD.n3957 AVDD.n3956 0.001
R8130 AVDD.n4102 AVDD.n4101 0.001
R8131 AVDD.n4238 AVDD.n4220 0.001
R8132 AVDD.n4394 AVDD.t739 0.001
R8133 AVDD.n4391 AVDD.n4390 0.001
R8134 AVDD.n4172 AVDD.n4171 0.001
R8135 AVDD.n4216 AVDD.n4210 0.001
R8136 AVDD.n4216 AVDD.n4215 0.001
R8137 AVDD.n4214 AVDD.n4213 0.001
R8138 AVDD.n2055 AVDD.n2054 0.001
R8139 AVDD.n2468 AVDD.n2467 0.001
R8140 AVDD.n5257 AVDD.n5256 0.001
R8141 AVDD.n4597 AVDD.n4595 0.001
R8142 AVDD.n4597 AVDD.n4441 0.001
R8143 AVDD.n4597 AVDD.n4517 0.001
R8144 AVDD.n4598 AVDD.n4597 0.001
R8145 AVDD.n5829 AVDD.n5828 0.001
R8146 AVDD.n6062 AVDD.n6061 0.001
R8147 AVDD.n6419 AVDD.n6418 0.001
R8148 AVDD.n4597 AVDD.n3496 0.001
R8149 AVDD.n4597 AVDD.n3736 0.001
R8150 AVDD.n6131 AVDD.n6129 0.001
R8151 AVDD.n6172 AVDD.n6170 0.001
R8152 AVDD.n4575 AVDD.n4574 0.001
R8153 AVDD.n3839 AVDD.n3838 0.001
R8154 AVDD.n3854 AVDD.t767 0.001
R8155 AVDD.n3855 AVDD.n3854 0.001
R8156 AVDD.n3869 AVDD.t833 0.001
R8157 AVDD.n3870 AVDD.n3869 0.001
R8158 AVDD.n3905 AVDD.t144 0.001
R8159 AVDD.n3906 AVDD.n3905 0.001
R8160 AVDD.n3971 AVDD.t0 0.001
R8161 AVDD.n3821 AVDD.t763 0.001
R8162 AVDD.n3804 AVDD.t190 0.001
R8163 AVDD.n3922 AVDD.n3921 0.001
R8164 AVDD.n3921 AVDD.t707 0.001
R8165 AVDD.n3936 AVDD.t729 0.001
R8166 AVDD.n3937 AVDD.n3936 0.001
R8167 AVDD.n3972 AVDD.n3971 0.001
R8168 AVDD.n3822 AVDD.n3821 0.001
R8169 AVDD.n3805 AVDD.n3804 0.001
R8170 AVDD.n4188 AVDD.t749 0.001
R8171 AVDD.n4236 AVDD.t339 0.001
R8172 AVDD.n4237 AVDD.n4236 0.001
R8173 AVDD.n4252 AVDD.t806 0.001
R8174 AVDD.n4253 AVDD.n4252 0.001
R8175 AVDD.n4054 AVDD.n4053 0.001
R8176 AVDD.n4069 AVDD.t719 0.001
R8177 AVDD.n4070 AVDD.n4069 0.001
R8178 AVDD.n4084 AVDD.t40 0.001
R8179 AVDD.n4085 AVDD.n4084 0.001
R8180 AVDD.n4120 AVDD.t215 0.001
R8181 AVDD.n4121 AVDD.n4120 0.001
R8182 AVDD.n4137 AVDD.n4136 0.001
R8183 AVDD.n4136 AVDD.t270 0.001
R8184 AVDD.n4151 AVDD.t54 0.001
R8185 AVDD.n4152 AVDD.n4151 0.001
R8186 AVDD.n4189 AVDD.n4188 0.001
R8187 AVDD.n3745 AVDD.n3744 0.001
R8188 AVDD.n3744 AVDD.t838 0.001
R8189 AVDD.n3763 AVDD.n3762 0.001
R8190 AVDD.n3762 AVDD.t741 0.001
R8191 AVDD.n3776 AVDD.n3775 0.001
R8192 AVDD.n3775 AVDD.t723 0.001
R8193 AVDD.n6056 AVDD.n6055 0.001
R8194 AVDD.n6055 AVDD.t95 0.001
R8195 AVDD.n5906 AVDD.n5905 0.001
R8196 AVDD.n5905 AVDD.t264 0.001
R8197 AVDD.n5925 AVDD.n5924 0.001
R8198 AVDD.n5924 AVDD.t818 0.001
R8199 AVDD.n5842 AVDD.n5841 0.001
R8200 AVDD.n5841 AVDD.t341 0.001
R8201 AVDD.n6076 AVDD.n6075 0.001
R8202 AVDD.n6075 AVDD.t266 0.001
R8203 AVDD.n6085 AVDD.n6084 0.001
R8204 AVDD.t353 AVDD.n6085 0.001
R8205 AVDD.n3881 AVDD.n3880 0.001
R8206 AVDD.n3880 AVDD.n3879 0.001
R8207 AVDD.n3786 AVDD.n3785 0.001
R8208 AVDD.n3785 AVDD.n3784 0.001
R8209 AVDD.n3950 AVDD.n3949 0.001
R8210 AVDD.n3949 AVDD.n3948 0.001
R8211 AVDD.n4400 AVDD.n4399 0.001
R8212 AVDD.n4401 AVDD.n4400 0.001
R8213 AVDD.n4096 AVDD.n4095 0.001
R8214 AVDD.n4095 AVDD.n4094 0.001
R8215 AVDD.n4165 AVDD.n4164 0.001
R8216 AVDD.n4164 AVDD.n4163 0.001
R8217 AVDD.n6413 AVDD.n6412 0.001
R8218 AVDD.n6412 AVDD.n6411 0.001
R8219 AVDD.n5878 AVDD.n5877 0.001
R8220 AVDD.n5877 AVDD.n5876 0.001
R8221 AVDD.n5819 AVDD.n5818 0.001
R8222 AVDD.n5818 AVDD.n5817 0.001
R8223 AVDD.n5836 AVDD.n5835 0.001
R8224 AVDD.n5837 AVDD.n5836 0.001
R8225 AVDD.n24 AVDD.n23 0.001
R8226 AVDD.n25 AVDD.n24 0.001
R8227 AVDD.t185 AVDD.n4381 0.001
R8228 AVDD.n6364 AVDD.n6363 0.001
R8229 AVDD.n6363 AVDD.n6362 0.001
R8230 AVDD.n4342 AVDD.n4341 0.001
R8231 AVDD.n4350 AVDD.n4342 0.001
R8232 AVDD.n4280 AVDD.n4279 0.001
R8233 AVDD.n4281 AVDD.n4280 0.001
R8234 AVDD.n4561 AVDD.n4560 0.001
R8235 AVDD.n4565 AVDD.n4564 0.001
R8236 AVDD.n4471 AVDD.n4470 0.001
R8237 AVDD.n4465 AVDD.n4464 0.001
R8238 AVDD.n4461 AVDD.n4460 0.001
R8239 AVDD.n4462 AVDD.n4461 0.001
R8240 AVDD.n4466 AVDD.n4465 0.001
R8241 AVDD.n4472 AVDD.n4471 0.001
R8242 AVDD.n4566 AVDD.n4565 0.001
R8243 AVDD.n4562 AVDD.n4561 0.001
R8244 AVDD.n6181 AVDD.n6180 0.001
R8245 AVDD.n6182 AVDD.n6181 0.001
R8246 AVDD.n6177 AVDD.n6176 0.001
R8247 AVDD.n6178 AVDD.n6177 0.001
R8248 AVDD.n6100 AVDD.n6099 0.001
R8249 AVDD.n6101 AVDD.n6100 0.001
R8250 AVDD.n6096 AVDD.n6095 0.001
R8251 AVDD.n6097 AVDD.n6096 0.001
R8252 AVDD.n6164 AVDD.n6163 0.001
R8253 AVDD.n6165 AVDD.n6164 0.001
R8254 AVDD.n6124 AVDD.n6123 0.001
R8255 AVDD.n6125 AVDD.n6124 0.001
R8256 AVDD.n4388 AVDD.n4387 0.001
R8257 AVDD.n4387 AVDD.t709 0.001
R8258 AVDD.n4210 AVDD.n4209 0.001
R8259 AVDD.n4597 AVDD.n4593 0.001
R8260 AVDD.n4597 AVDD.n4541 0.001
R8261 AVDD.n4597 AVDD.n4509 0.001
R8262 AVDD.n4597 AVDD.n3730 0.001
R8263 AVDD.n4597 AVDD.n3560 0.001
R8264 AVDD.n4597 AVDD.n3489 0.001
R8265 AVDD.n4597 AVDD.n3501 0.001
R8266 AVDD.n4597 AVDD.n4544 0.001
R8267 AVDD.n4597 AVDD.n4515 0.001
R8268 AVDD.n4597 AVDD.n4439 0.001
R8269 AVDD.n4597 AVDD.n3733 0.001
R8270 AVDD.n4597 AVDD.n3563 0.001
R8271 AVDD.n4597 AVDD.n3494 0.001
R8272 AVDD.n4597 AVDD.n3537 0.001
R8273 AVDD.n4499 AVDD.n4498 0.001
R8274 AVDD.n3728 AVDD.n3727 0.001
R8275 AVDD.n4431 AVDD.n4430 0.001
R8276 AVDD.n4507 AVDD.n4506 0.001
R8277 AVDD.n4539 AVDD.n4538 0.001
R8278 AVDD.n4591 AVDD.n4590 0.001
R8279 AVDD.n3558 AVDD.n3557 0.001
R8280 AVDD.n3486 AVDD.n3478 0.001
R8281 AVDD.n3837 AVDD.t181 0.001
R8282 AVDD.n4052 AVDD.t29 0.001
R8283 AVDD.n3580 AVDD.n3579 0.001
R8284 AVDD.n3586 AVDD.n3585 0.001
R8285 AVDD.n3594 AVDD.n3593 0.001
R8286 AVDD.n3602 AVDD.n3601 0.001
R8287 AVDD.n3610 AVDD.n3609 0.001
R8288 AVDD.n3618 AVDD.n3617 0.001
R8289 AVDD.n3626 AVDD.n3625 0.001
R8290 AVDD.n3634 AVDD.n3633 0.001
R8291 AVDD.n3727 AVDD.n3726 0.001
R8292 AVDD.n4430 AVDD.n4429 0.001
R8293 AVDD.n4506 AVDD.n4505 0.001
R8294 AVDD.n4538 AVDD.n4537 0.001
R8295 AVDD.n4590 AVDD.n4589 0.001
R8296 AVDD.n3557 AVDD.n3556 0.001
R8297 AVDD.n3478 AVDD.n3477 0.001
R8298 AVDD.n3557 AVDD.n3549 0.001
R8299 AVDD.n3727 AVDD.n3719 0.001
R8300 AVDD.n4430 AVDD.n4426 0.001
R8301 AVDD.n4506 AVDD.n4454 0.001
R8302 AVDD.n4538 AVDD.n4530 0.001
R8303 AVDD.n4590 AVDD.n4558 0.001
R8304 AVDD.n3478 AVDD.n3470 0.001
R8305 AVDD.n4499 AVDD.n4489 0.001
R8306 AVDD.n4499 AVDD.n4492 0.001
R8307 AVDD.n6279 AVDD.n6277 0.001
R8308 AVDD.n6256 AVDD.n6254 0.001
R8309 AVDD.n6233 AVDD.n6231 0.001
R8310 AVDD.n6210 AVDD.n6208 0.001
R8311 AVDD.n6188 AVDD.n6186 0.001
R8312 AVDD.n6144 AVDD.n6142 0.001
R8313 AVDD.n5786 AVDD.n5784 0.001
R8314 AVDD.n5769 AVDD.n5767 0.001
R8315 AVDD.n4335 AVDD.n4334 0.001
R8316 AVDD.n4288 AVDD.n4287 0.001
R8317 AVDD.n4273 AVDD.n4272 0.001
R8318 AVDD.n4262 AVDD.n4261 0.001
R8319 AVDD.n4003 AVDD.n4002 0.001
R8320 AVDD.n4017 AVDD.n4012 0.001
R8321 AVDD.n3989 AVDD.n3988 0.001
R8322 AVDD.n4363 AVDD.n4362 0.001
R8323 AVDD.n4207 AVDD.n4206 0.001
R8324 AVDD.n6306 AVDD.n5716 0.001
R8325 AVDD.n5709 AVDD.n5706 0.001
R8326 AVDD.n5722 AVDD.n5721 0.001
R8327 AVDD.n5730 AVDD.n5729 0.001
R8328 AVDD.n5738 AVDD.n5737 0.001
R8329 AVDD.n5748 AVDD.n5747 0.001
R8330 AVDD.n6300 AVDD.n6299 0.001
R8331 AVDD.n4927 AVDD.n4926 0.001
R8332 AVDD.n4208 AVDD.n4207 0.001
R8333 AVDD.n1356 AVDD.n1348 0.001
R8334 AVDD.n572 AVDD.n564 0.001
R8335 AVDD.n3856 AVDD.n3855 0.001
R8336 AVDD.n3907 AVDD.n3906 0.001
R8337 AVDD.n3882 AVDD.n3881 0.001
R8338 AVDD.n3840 AVDD.n3839 0.001
R8339 AVDD.n3871 AVDD.n3870 0.001
R8340 AVDD.n3787 AVDD.n3786 0.001
R8341 AVDD.n3923 AVDD.n3922 0.001
R8342 AVDD.n3938 AVDD.n3937 0.001
R8343 AVDD.n3951 AVDD.n3950 0.001
R8344 AVDD.n3973 AVDD.n3972 0.001
R8345 AVDD.n3823 AVDD.n3822 0.001
R8346 AVDD.n3806 AVDD.n3805 0.001
R8347 AVDD.n4071 AVDD.n4070 0.001
R8348 AVDD.n4122 AVDD.n4121 0.001
R8349 AVDD.n4238 AVDD.n4237 0.001
R8350 AVDD.n4336 AVDD.n4335 0.001
R8351 AVDD.n4336 AVDD.n4331 0.001
R8352 AVDD.n4364 AVDD.n4363 0.001
R8353 AVDD.n4364 AVDD.n4359 0.001
R8354 AVDD.n4289 AVDD.n4288 0.001
R8355 AVDD.n4289 AVDD.n4284 0.001
R8356 AVDD.n4274 AVDD.n4273 0.001
R8357 AVDD.n4274 AVDD.n4269 0.001
R8358 AVDD.n4263 AVDD.n4262 0.001
R8359 AVDD.n4263 AVDD.n4258 0.001
R8360 AVDD.n4004 AVDD.n4003 0.001
R8361 AVDD.n4004 AVDD.n3999 0.001
R8362 AVDD.n4017 AVDD.n4016 0.001
R8363 AVDD.n4016 AVDD.n4013 0.001
R8364 AVDD.n3990 AVDD.n3989 0.001
R8365 AVDD.n3990 AVDD.n3985 0.001
R8366 AVDD.n4389 AVDD.n4388 0.001
R8367 AVDD.n4399 AVDD.n4398 0.001
R8368 AVDD.n4254 AVDD.n4253 0.001
R8369 AVDD.n4097 AVDD.n4096 0.001
R8370 AVDD.n4055 AVDD.n4054 0.001
R8371 AVDD.n4086 AVDD.n4085 0.001
R8372 AVDD.n4138 AVDD.n4137 0.001
R8373 AVDD.n4153 AVDD.n4152 0.001
R8374 AVDD.n4166 AVDD.n4165 0.001
R8375 AVDD.n4190 AVDD.n4189 0.001
R8376 AVDD.n3493 AVDD.n3492 0.001
R8377 AVDD.n4602 AVDD.n4601 0.001
R8378 AVDD.n3459 AVDD.n3458 0.001
R8379 AVDD.n4438 AVDD.n4437 0.001
R8380 AVDD.n4514 AVDD.n4513 0.001
R8381 AVDD.n3466 AVDD.n3465 0.001
R8382 AVDD.n3764 AVDD.n3763 0.001
R8383 AVDD.n6414 AVDD.n6413 0.001
R8384 AVDD.n3746 AVDD.n3745 0.001
R8385 AVDD.n3777 AVDD.n3776 0.001
R8386 AVDD.n5879 AVDD.n5878 0.001
R8387 AVDD.n6057 AVDD.n6056 0.001
R8388 AVDD.n5907 AVDD.n5906 0.001
R8389 AVDD.n5926 AVDD.n5925 0.001
R8390 AVDD.n5820 AVDD.n5819 0.001
R8391 AVDD.n5843 AVDD.n5842 0.001
R8392 AVDD.n6077 AVDD.n6076 0.001
R8393 AVDD.n6084 AVDD.n6083 0.001
R8394 AVDD.n137 AVDD.n135 0.001
R8395 AVDD.n138 AVDD.n137 0.001
R8396 AVDD.n6495 AVDD.n6493 0.001
R8397 AVDD.n6496 AVDD.n6495 0.001
R8398 AVDD.n6365 AVDD.n6364 0.001
R8399 AVDD.n6306 AVDD.n6305 0.001
R8400 AVDD.n6305 AVDD.n6303 0.001
R8401 AVDD.n5709 AVDD.n5708 0.001
R8402 AVDD.n5724 AVDD.n5722 0.001
R8403 AVDD.n6303 AVDD.n5724 0.001
R8404 AVDD.n5732 AVDD.n5730 0.001
R8405 AVDD.n6303 AVDD.n5732 0.001
R8406 AVDD.n5742 AVDD.n5738 0.001
R8407 AVDD.n6303 AVDD.n5742 0.001
R8408 AVDD.n5750 AVDD.n5748 0.001
R8409 AVDD.n6303 AVDD.n5750 0.001
R8410 AVDD.n6302 AVDD.n6300 0.001
R8411 AVDD.n6303 AVDD.n6302 0.001
R8412 AVDD.n1356 AVDD.n1355 0.001
R8413 AVDD.n1355 AVDD.n1351 0.001
R8414 AVDD.n572 AVDD.n571 0.001
R8415 AVDD.n571 AVDD.n565 0.001
R8416 AVDD.n4825 AVDD.n4824 0.001
R8417 AVDD.n4907 AVDD.n4906 0.001
R8418 AVDD.n3498 AVDD.n3497 0.001
R8419 AVDD.n4433 AVDD.n4414 0.001
R8420 a_1560_n22142.n60 a_1560_n22142.t6 14.771
R8421 a_1560_n22142.n61 a_1560_n22142.t5 14.771
R8422 a_1560_n22142.n320 a_1560_n22142.t9 14.286
R8423 a_1560_n22142.n331 a_1560_n22142.t1 14.27
R8424 a_1560_n22142.n60 a_1560_n22142.t0 13.849
R8425 a_1560_n22142.n61 a_1560_n22142.t3 13.849
R8426 a_1560_n22142.n332 a_1560_n22142.t4 13.849
R8427 a_1560_n22142.n321 a_1560_n22142.t2 13.849
R8428 a_1560_n22142.n335 a_1560_n22142.n334 13.623
R8429 a_1560_n22142.n3 a_1560_n22142.t100 12.05
R8430 a_1560_n22142.n3 a_1560_n22142.t81 12.05
R8431 a_1560_n22142.n2 a_1560_n22142.t50 12.05
R8432 a_1560_n22142.n2 a_1560_n22142.t31 12.05
R8433 a_1560_n22142.n18 a_1560_n22142.t111 12.05
R8434 a_1560_n22142.n18 a_1560_n22142.t90 12.05
R8435 a_1560_n22142.n39 a_1560_n22142.t16 12.05
R8436 a_1560_n22142.n39 a_1560_n22142.t108 12.05
R8437 a_1560_n22142.n40 a_1560_n22142.t14 12.05
R8438 a_1560_n22142.n40 a_1560_n22142.t72 12.05
R8439 a_1560_n22142.n41 a_1560_n22142.t83 12.05
R8440 a_1560_n22142.n41 a_1560_n22142.t19 12.05
R8441 a_1560_n22142.n46 a_1560_n22142.t21 12.05
R8442 a_1560_n22142.n46 a_1560_n22142.t77 12.05
R8443 a_1560_n22142.n53 a_1560_n22142.t89 12.05
R8444 a_1560_n22142.n53 a_1560_n22142.t26 12.05
R8445 a_1560_n22142.n54 a_1560_n22142.t42 12.05
R8446 a_1560_n22142.n54 a_1560_n22142.t93 12.05
R8447 a_1560_n22142.n59 a_1560_n22142.t54 12.05
R8448 a_1560_n22142.n59 a_1560_n22142.t110 12.05
R8449 a_1560_n22142.n50 a_1560_n22142.t99 12.05
R8450 a_1560_n22142.n50 a_1560_n22142.t80 12.05
R8451 a_1560_n22142.n52 a_1560_n22142.t32 12.05
R8452 a_1560_n22142.n52 a_1560_n22142.t13 12.05
R8453 a_1560_n22142.n51 a_1560_n22142.t82 12.05
R8454 a_1560_n22142.n51 a_1560_n22142.t70 12.05
R8455 a_1560_n22142.n44 a_1560_n22142.t23 12.05
R8456 a_1560_n22142.n44 a_1560_n22142.t11 12.05
R8457 a_1560_n22142.n42 a_1560_n22142.t109 12.05
R8458 a_1560_n22142.n42 a_1560_n22142.t57 12.05
R8459 a_1560_n22142.n20 a_1560_n22142.t75 12.05
R8460 a_1560_n22142.n20 a_1560_n22142.t60 12.05
R8461 a_1560_n22142.n21 a_1560_n22142.t41 12.05
R8462 a_1560_n22142.n21 a_1560_n22142.t125 12.05
R8463 a_1560_n22142.n24 a_1560_n22142.t106 12.05
R8464 a_1560_n22142.n24 a_1560_n22142.t69 12.05
R8465 a_1560_n22142.n25 a_1560_n22142.t48 12.05
R8466 a_1560_n22142.n25 a_1560_n22142.t10 12.05
R8467 a_1560_n22142.n26 a_1560_n22142.t115 12.05
R8468 a_1560_n22142.n26 a_1560_n22142.t73 12.05
R8469 a_1560_n22142.n19 a_1560_n22142.t59 12.05
R8470 a_1560_n22142.n19 a_1560_n22142.t20 12.05
R8471 a_1560_n22142.n13 a_1560_n22142.t66 12.05
R8472 a_1560_n22142.n13 a_1560_n22142.t36 12.05
R8473 a_1560_n22142.n10 a_1560_n22142.t124 12.05
R8474 a_1560_n22142.n10 a_1560_n22142.t102 12.05
R8475 a_1560_n22142.n5 a_1560_n22142.t112 12.05
R8476 a_1560_n22142.n5 a_1560_n22142.t47 12.05
R8477 a_1560_n22142.n4 a_1560_n22142.t44 12.05
R8478 a_1560_n22142.n4 a_1560_n22142.t98 12.05
R8479 a_1560_n22142.n7 a_1560_n22142.t40 12.05
R8480 a_1560_n22142.n7 a_1560_n22142.t92 12.05
R8481 a_1560_n22142.n6 a_1560_n22142.t88 12.05
R8482 a_1560_n22142.n6 a_1560_n22142.t25 12.05
R8483 a_1560_n22142.n9 a_1560_n22142.t52 12.05
R8484 a_1560_n22142.n9 a_1560_n22142.t33 12.05
R8485 a_1560_n22142.n8 a_1560_n22142.t103 12.05
R8486 a_1560_n22142.n8 a_1560_n22142.t84 12.05
R8487 a_1560_n22142.n11 a_1560_n22142.t122 12.05
R8488 a_1560_n22142.n11 a_1560_n22142.t63 12.05
R8489 a_1560_n22142.n14 a_1560_n22142.t61 12.05
R8490 a_1560_n22142.n14 a_1560_n22142.t117 12.05
R8491 a_1560_n22142.n27 a_1560_n22142.t51 12.05
R8492 a_1560_n22142.n27 a_1560_n22142.t105 12.05
R8493 a_1560_n22142.n30 a_1560_n22142.t101 12.05
R8494 a_1560_n22142.n30 a_1560_n22142.t39 12.05
R8495 a_1560_n22142.n29 a_1560_n22142.t35 12.05
R8496 a_1560_n22142.n29 a_1560_n22142.t87 12.05
R8497 a_1560_n22142.n28 a_1560_n22142.t95 12.05
R8498 a_1560_n22142.n28 a_1560_n22142.t30 12.05
R8499 a_1560_n22142.n15 a_1560_n22142.t123 12.05
R8500 a_1560_n22142.n15 a_1560_n22142.t116 12.05
R8501 a_1560_n22142.n57 a_1560_n22142.t62 12.05
R8502 a_1560_n22142.n57 a_1560_n22142.t49 12.05
R8503 a_1560_n22142.n48 a_1560_n22142.t53 12.05
R8504 a_1560_n22142.n48 a_1560_n22142.t34 12.05
R8505 a_1560_n22142.n49 a_1560_n22142.t104 12.05
R8506 a_1560_n22142.n49 a_1560_n22142.t85 12.05
R8507 a_1560_n22142.n45 a_1560_n22142.t37 12.05
R8508 a_1560_n22142.n45 a_1560_n22142.t17 12.05
R8509 a_1560_n22142.n32 a_1560_n22142.t119 12.05
R8510 a_1560_n22142.n32 a_1560_n22142.t64 12.05
R8511 a_1560_n22142.n33 a_1560_n22142.t86 12.05
R8512 a_1560_n22142.n33 a_1560_n22142.t71 12.05
R8513 a_1560_n22142.n34 a_1560_n22142.t38 12.05
R8514 a_1560_n22142.n34 a_1560_n22142.t18 12.05
R8515 a_1560_n22142.n35 a_1560_n22142.t94 12.05
R8516 a_1560_n22142.n35 a_1560_n22142.t76 12.05
R8517 a_1560_n22142.n47 a_1560_n22142.t45 12.05
R8518 a_1560_n22142.n47 a_1560_n22142.t24 12.05
R8519 a_1560_n22142.n31 a_1560_n22142.t113 12.05
R8520 a_1560_n22142.n31 a_1560_n22142.t91 12.05
R8521 a_1560_n22142.n56 a_1560_n22142.t121 12.05
R8522 a_1560_n22142.n56 a_1560_n22142.t107 12.05
R8523 a_1560_n22142.n12 a_1560_n22142.t65 12.05
R8524 a_1560_n22142.n12 a_1560_n22142.t55 12.05
R8525 a_1560_n22142.n38 a_1560_n22142.t96 12.05
R8526 a_1560_n22142.n38 a_1560_n22142.t78 12.05
R8527 a_1560_n22142.n37 a_1560_n22142.t28 12.05
R8528 a_1560_n22142.n37 a_1560_n22142.t12 12.05
R8529 a_1560_n22142.n36 a_1560_n22142.t68 12.05
R8530 a_1560_n22142.n36 a_1560_n22142.t15 12.05
R8531 a_1560_n22142.n23 a_1560_n22142.t27 12.05
R8532 a_1560_n22142.n23 a_1560_n22142.t79 12.05
R8533 a_1560_n22142.n22 a_1560_n22142.t29 12.05
R8534 a_1560_n22142.n22 a_1560_n22142.t118 12.05
R8535 a_1560_n22142.n43 a_1560_n22142.t74 12.05
R8536 a_1560_n22142.n43 a_1560_n22142.t67 12.05
R8537 a_1560_n22142.n17 a_1560_n22142.t58 12.05
R8538 a_1560_n22142.n17 a_1560_n22142.t46 12.05
R8539 a_1560_n22142.n58 a_1560_n22142.t114 12.05
R8540 a_1560_n22142.n58 a_1560_n22142.t97 12.05
R8541 a_1560_n22142.n16 a_1560_n22142.t120 12.05
R8542 a_1560_n22142.n16 a_1560_n22142.t56 12.05
R8543 a_1560_n22142.n55 a_1560_n22142.t43 12.05
R8544 a_1560_n22142.n55 a_1560_n22142.t22 12.05
R8545 a_1560_n22142.n315 a_1560_n22142.n1 10.648
R8546 a_1560_n22142.n325 a_1560_n22142.n323 9.3
R8547 a_1560_n22142.n325 a_1560_n22142.n324 9.3
R8548 a_1560_n22142.n329 a_1560_n22142.n327 9.3
R8549 a_1560_n22142.n329 a_1560_n22142.n328 9.3
R8550 a_1560_n22142.n243 a_1560_n22142.n241 9.3
R8551 a_1560_n22142.n243 a_1560_n22142.n242 9.3
R8552 a_1560_n22142.n137 a_1560_n22142.n135 9.3
R8553 a_1560_n22142.n137 a_1560_n22142.n136 9.3
R8554 a_1560_n22142.n133 a_1560_n22142.n131 9.3
R8555 a_1560_n22142.n133 a_1560_n22142.n132 9.3
R8556 a_1560_n22142.n129 a_1560_n22142.n127 9.3
R8557 a_1560_n22142.n129 a_1560_n22142.n128 9.3
R8558 a_1560_n22142.n105 a_1560_n22142.n103 9.3
R8559 a_1560_n22142.n105 a_1560_n22142.n104 9.3
R8560 a_1560_n22142.n73 a_1560_n22142.n71 9.3
R8561 a_1560_n22142.n73 a_1560_n22142.n72 9.3
R8562 a_1560_n22142.n69 a_1560_n22142.n67 9.3
R8563 a_1560_n22142.n69 a_1560_n22142.n68 9.3
R8564 a_1560_n22142.n86 a_1560_n22142.n84 9.3
R8565 a_1560_n22142.n86 a_1560_n22142.n85 9.3
R8566 a_1560_n22142.n77 a_1560_n22142.n75 9.3
R8567 a_1560_n22142.n77 a_1560_n22142.n76 9.3
R8568 a_1560_n22142.n81 a_1560_n22142.n79 9.3
R8569 a_1560_n22142.n81 a_1560_n22142.n80 9.3
R8570 a_1560_n22142.n114 a_1560_n22142.n112 9.3
R8571 a_1560_n22142.n114 a_1560_n22142.n113 9.3
R8572 a_1560_n22142.n122 a_1560_n22142.n120 9.3
R8573 a_1560_n22142.n122 a_1560_n22142.n121 9.3
R8574 a_1560_n22142.n230 a_1560_n22142.n228 9.3
R8575 a_1560_n22142.n230 a_1560_n22142.n229 9.3
R8576 a_1560_n22142.n226 a_1560_n22142.n224 9.3
R8577 a_1560_n22142.n226 a_1560_n22142.n225 9.3
R8578 a_1560_n22142.n212 a_1560_n22142.n210 9.3
R8579 a_1560_n22142.n212 a_1560_n22142.n211 9.3
R8580 a_1560_n22142.n208 a_1560_n22142.n206 9.3
R8581 a_1560_n22142.n208 a_1560_n22142.n207 9.3
R8582 a_1560_n22142.n204 a_1560_n22142.n202 9.3
R8583 a_1560_n22142.n204 a_1560_n22142.n203 9.3
R8584 a_1560_n22142.n238 a_1560_n22142.n236 9.3
R8585 a_1560_n22142.n238 a_1560_n22142.n237 9.3
R8586 a_1560_n22142.n273 a_1560_n22142.n271 9.3
R8587 a_1560_n22142.n273 a_1560_n22142.n272 9.3
R8588 a_1560_n22142.n287 a_1560_n22142.n285 9.3
R8589 a_1560_n22142.n287 a_1560_n22142.n286 9.3
R8590 a_1560_n22142.n310 a_1560_n22142.n308 9.3
R8591 a_1560_n22142.n310 a_1560_n22142.n309 9.3
R8592 a_1560_n22142.n314 a_1560_n22142.n312 9.3
R8593 a_1560_n22142.n314 a_1560_n22142.n313 9.3
R8594 a_1560_n22142.n301 a_1560_n22142.n299 9.3
R8595 a_1560_n22142.n301 a_1560_n22142.n300 9.3
R8596 a_1560_n22142.n305 a_1560_n22142.n303 9.3
R8597 a_1560_n22142.n305 a_1560_n22142.n304 9.3
R8598 a_1560_n22142.n293 a_1560_n22142.n291 9.3
R8599 a_1560_n22142.n293 a_1560_n22142.n292 9.3
R8600 a_1560_n22142.n297 a_1560_n22142.n295 9.3
R8601 a_1560_n22142.n297 a_1560_n22142.n296 9.3
R8602 a_1560_n22142.n282 a_1560_n22142.n280 9.3
R8603 a_1560_n22142.n282 a_1560_n22142.n281 9.3
R8604 a_1560_n22142.n268 a_1560_n22142.n266 9.3
R8605 a_1560_n22142.n268 a_1560_n22142.n267 9.3
R8606 a_1560_n22142.n199 a_1560_n22142.n197 9.3
R8607 a_1560_n22142.n199 a_1560_n22142.n198 9.3
R8608 a_1560_n22142.n185 a_1560_n22142.n183 9.3
R8609 a_1560_n22142.n185 a_1560_n22142.n184 9.3
R8610 a_1560_n22142.n189 a_1560_n22142.n187 9.3
R8611 a_1560_n22142.n189 a_1560_n22142.n188 9.3
R8612 a_1560_n22142.n193 a_1560_n22142.n191 9.3
R8613 a_1560_n22142.n193 a_1560_n22142.n192 9.3
R8614 a_1560_n22142.n260 a_1560_n22142.n258 9.3
R8615 a_1560_n22142.n260 a_1560_n22142.n259 9.3
R8616 a_1560_n22142.n96 a_1560_n22142.n94 9.3
R8617 a_1560_n22142.n96 a_1560_n22142.n95 9.3
R8618 a_1560_n22142.n92 a_1560_n22142.n90 9.3
R8619 a_1560_n22142.n92 a_1560_n22142.n91 9.3
R8620 a_1560_n22142.n110 a_1560_n22142.n108 9.3
R8621 a_1560_n22142.n110 a_1560_n22142.n109 9.3
R8622 a_1560_n22142.n172 a_1560_n22142.n170 9.3
R8623 a_1560_n22142.n172 a_1560_n22142.n171 9.3
R8624 a_1560_n22142.n168 a_1560_n22142.n166 9.3
R8625 a_1560_n22142.n168 a_1560_n22142.n167 9.3
R8626 a_1560_n22142.n164 a_1560_n22142.n162 9.3
R8627 a_1560_n22142.n164 a_1560_n22142.n163 9.3
R8628 a_1560_n22142.n160 a_1560_n22142.n158 9.3
R8629 a_1560_n22142.n160 a_1560_n22142.n159 9.3
R8630 a_1560_n22142.n101 a_1560_n22142.n99 9.3
R8631 a_1560_n22142.n101 a_1560_n22142.n100 9.3
R8632 a_1560_n22142.n180 a_1560_n22142.n178 9.3
R8633 a_1560_n22142.n180 a_1560_n22142.n179 9.3
R8634 a_1560_n22142.n277 a_1560_n22142.n275 9.3
R8635 a_1560_n22142.n277 a_1560_n22142.n276 9.3
R8636 a_1560_n22142.n144 a_1560_n22142.n142 9.3
R8637 a_1560_n22142.n144 a_1560_n22142.n143 9.3
R8638 a_1560_n22142.n148 a_1560_n22142.n146 9.3
R8639 a_1560_n22142.n148 a_1560_n22142.n147 9.3
R8640 a_1560_n22142.n152 a_1560_n22142.n150 9.3
R8641 a_1560_n22142.n152 a_1560_n22142.n151 9.3
R8642 a_1560_n22142.n216 a_1560_n22142.n214 9.3
R8643 a_1560_n22142.n216 a_1560_n22142.n215 9.3
R8644 a_1560_n22142.n220 a_1560_n22142.n218 9.3
R8645 a_1560_n22142.n220 a_1560_n22142.n219 9.3
R8646 a_1560_n22142.n118 a_1560_n22142.n116 9.3
R8647 a_1560_n22142.n118 a_1560_n22142.n117 9.3
R8648 a_1560_n22142.n248 a_1560_n22142.n246 9.3
R8649 a_1560_n22142.n248 a_1560_n22142.n247 9.3
R8650 a_1560_n22142.n253 a_1560_n22142.n251 9.3
R8651 a_1560_n22142.n253 a_1560_n22142.n252 9.3
R8652 a_1560_n22142.n65 a_1560_n22142.n63 9.3
R8653 a_1560_n22142.n65 a_1560_n22142.n64 9.3
R8654 a_1560_n22142.t8 a_1560_n22142.n335 8.857
R8655 a_1560_n22142.n335 a_1560_n22142.t7 8.268
R8656 a_1560_n22142.n334 a_1560_n22142.n333 2.236
R8657 a_1560_n22142.n244 a_1560_n22142.n58 1.326
R8658 a_1560_n22142.n264 a_1560_n22142.n56 1.326
R8659 a_1560_n22142.n33 a_1560_n22142.n173 1.322
R8660 a_1560_n22142.n34 a_1560_n22142.n174 1.322
R8661 a_1560_n22142.n35 a_1560_n22142.n175 1.322
R8662 a_1560_n22142.n47 a_1560_n22142.n176 1.322
R8663 a_1560_n22142.n181 a_1560_n22142.n31 1.322
R8664 a_1560_n22142.n278 a_1560_n22142.n12 1.322
R8665 a_1560_n22142.n37 a_1560_n22142.n153 1.322
R8666 a_1560_n22142.n38 a_1560_n22142.n154 1.322
R8667 a_1560_n22142.n45 a_1560_n22142.n155 1.322
R8668 a_1560_n22142.n97 a_1560_n22142.n48 1.322
R8669 a_1560_n22142.n263 a_1560_n22142.n57 1.322
R8670 a_1560_n22142.n262 a_1560_n22142.n15 1.322
R8671 a_1560_n22142.n23 a_1560_n22142.n221 1.322
R8672 a_1560_n22142.n29 a_1560_n22142.n194 1.322
R8673 a_1560_n22142.n30 a_1560_n22142.n195 1.322
R8674 a_1560_n22142.n200 a_1560_n22142.n27 1.322
R8675 a_1560_n22142.n269 a_1560_n22142.n14 1.322
R8676 a_1560_n22142.n283 a_1560_n22142.n11 1.322
R8677 a_1560_n22142.n21 a_1560_n22142.n231 1.322
R8678 a_1560_n22142.n24 a_1560_n22142.n232 1.322
R8679 a_1560_n22142.n25 a_1560_n22142.n233 1.322
R8680 a_1560_n22142.n26 a_1560_n22142.n234 1.322
R8681 a_1560_n22142.n239 a_1560_n22142.n19 1.322
R8682 a_1560_n22142.n317 a_1560_n22142.n13 1.322
R8683 a_1560_n22142.n316 a_1560_n22142.n10 1.322
R8684 a_1560_n22142.n43 a_1560_n22142.n123 1.322
R8685 a_1560_n22142.n44 a_1560_n22142.n124 1.322
R8686 a_1560_n22142.n52 a_1560_n22142.n82 1.322
R8687 a_1560_n22142.n87 a_1560_n22142.n50 1.322
R8688 a_1560_n22142.n249 a_1560_n22142.n17 1.322
R8689 a_1560_n22142.n40 a_1560_n22142.n138 1.322
R8690 a_1560_n22142.n41 a_1560_n22142.n139 1.322
R8691 a_1560_n22142.n88 a_1560_n22142.n54 1.322
R8692 a_1560_n22142.n256 a_1560_n22142.n59 1.322
R8693 a_1560_n22142.n255 a_1560_n22142.n16 1.322
R8694 a_1560_n22142.n319 a_1560_n22142.n18 1.267
R8695 a_1560_n22142.n330 a_1560_n22142.n2 1.267
R8696 a_1560_n22142.n1 a_1560_n22142.n5 1.245
R8697 a_1560_n22142.n306 a_1560_n22142.n7 1.245
R8698 a_1560_n22142.n0 a_1560_n22142.n9 1.245
R8699 a_1560_n22142.n320 a_1560_n22142.n55 0.961
R8700 a_1560_n22142.n331 a_1560_n22142.n3 0.961
R8701 a_1560_n22142.n333 a_1560_n22142.n332 0.849
R8702 a_1560_n22142.n334 a_1560_n22142.n61 0.834
R8703 a_1560_n22142.n319 a_1560_n22142.n239 0.834
R8704 a_1560_n22142.n318 a_1560_n22142.n317 0.834
R8705 a_1560_n22142.n3 a_1560_n22142.n322 0.752
R8706 a_1560_n22142.n2 a_1560_n22142.n326 0.752
R8707 a_1560_n22142.n18 a_1560_n22142.n240 0.752
R8708 a_1560_n22142.n39 a_1560_n22142.n134 0.752
R8709 a_1560_n22142.n40 a_1560_n22142.n130 0.752
R8710 a_1560_n22142.n41 a_1560_n22142.n126 0.752
R8711 a_1560_n22142.n46 a_1560_n22142.n102 0.752
R8712 a_1560_n22142.n53 a_1560_n22142.n70 0.752
R8713 a_1560_n22142.n54 a_1560_n22142.n66 0.752
R8714 a_1560_n22142.n50 a_1560_n22142.n83 0.752
R8715 a_1560_n22142.n52 a_1560_n22142.n74 0.752
R8716 a_1560_n22142.n51 a_1560_n22142.n78 0.752
R8717 a_1560_n22142.n44 a_1560_n22142.n111 0.752
R8718 a_1560_n22142.n42 a_1560_n22142.n119 0.752
R8719 a_1560_n22142.n20 a_1560_n22142.n227 0.752
R8720 a_1560_n22142.n21 a_1560_n22142.n223 0.752
R8721 a_1560_n22142.n24 a_1560_n22142.n209 0.752
R8722 a_1560_n22142.n25 a_1560_n22142.n205 0.752
R8723 a_1560_n22142.n26 a_1560_n22142.n201 0.752
R8724 a_1560_n22142.n19 a_1560_n22142.n235 0.752
R8725 a_1560_n22142.n13 a_1560_n22142.n270 0.752
R8726 a_1560_n22142.n10 a_1560_n22142.n284 0.752
R8727 a_1560_n22142.n5 a_1560_n22142.n307 0.752
R8728 a_1560_n22142.n4 a_1560_n22142.n311 0.752
R8729 a_1560_n22142.n7 a_1560_n22142.n298 0.752
R8730 a_1560_n22142.n6 a_1560_n22142.n302 0.752
R8731 a_1560_n22142.n9 a_1560_n22142.n290 0.752
R8732 a_1560_n22142.n8 a_1560_n22142.n294 0.752
R8733 a_1560_n22142.n11 a_1560_n22142.n279 0.752
R8734 a_1560_n22142.n14 a_1560_n22142.n265 0.752
R8735 a_1560_n22142.n27 a_1560_n22142.n196 0.752
R8736 a_1560_n22142.n30 a_1560_n22142.n182 0.752
R8737 a_1560_n22142.n29 a_1560_n22142.n186 0.752
R8738 a_1560_n22142.n28 a_1560_n22142.n190 0.752
R8739 a_1560_n22142.n15 a_1560_n22142.n257 0.752
R8740 a_1560_n22142.n48 a_1560_n22142.n93 0.752
R8741 a_1560_n22142.n49 a_1560_n22142.n89 0.752
R8742 a_1560_n22142.n45 a_1560_n22142.n107 0.752
R8743 a_1560_n22142.n32 a_1560_n22142.n169 0.752
R8744 a_1560_n22142.n33 a_1560_n22142.n165 0.752
R8745 a_1560_n22142.n34 a_1560_n22142.n161 0.752
R8746 a_1560_n22142.n35 a_1560_n22142.n157 0.752
R8747 a_1560_n22142.n47 a_1560_n22142.n98 0.752
R8748 a_1560_n22142.n31 a_1560_n22142.n177 0.752
R8749 a_1560_n22142.n12 a_1560_n22142.n274 0.752
R8750 a_1560_n22142.n38 a_1560_n22142.n141 0.752
R8751 a_1560_n22142.n37 a_1560_n22142.n145 0.752
R8752 a_1560_n22142.n36 a_1560_n22142.n149 0.752
R8753 a_1560_n22142.n23 a_1560_n22142.n213 0.752
R8754 a_1560_n22142.n22 a_1560_n22142.n217 0.752
R8755 a_1560_n22142.n43 a_1560_n22142.n115 0.752
R8756 a_1560_n22142.n17 a_1560_n22142.n245 0.752
R8757 a_1560_n22142.n16 a_1560_n22142.n250 0.752
R8758 a_1560_n22142.n55 a_1560_n22142.n62 0.752
R8759 a_1560_n22142.n59 a_1560_n22142.n255 0.556
R8760 a_1560_n22142.n57 a_1560_n22142.n262 0.556
R8761 a_1560_n22142.n173 a_1560_n22142.n32 0.552
R8762 a_1560_n22142.n174 a_1560_n22142.n33 0.552
R8763 a_1560_n22142.n175 a_1560_n22142.n34 0.552
R8764 a_1560_n22142.n176 a_1560_n22142.n35 0.552
R8765 a_1560_n22142.n181 a_1560_n22142.n47 0.552
R8766 a_1560_n22142.n153 a_1560_n22142.n36 0.552
R8767 a_1560_n22142.n154 a_1560_n22142.n37 0.552
R8768 a_1560_n22142.n155 a_1560_n22142.n38 0.552
R8769 a_1560_n22142.n156 a_1560_n22142.n45 0.552
R8770 a_1560_n22142.n97 a_1560_n22142.n49 0.552
R8771 a_1560_n22142.n15 a_1560_n22142.n261 0.552
R8772 a_1560_n22142.n221 a_1560_n22142.n22 0.552
R8773 a_1560_n22142.n222 a_1560_n22142.n23 0.552
R8774 a_1560_n22142.n194 a_1560_n22142.n28 0.552
R8775 a_1560_n22142.n195 a_1560_n22142.n29 0.552
R8776 a_1560_n22142.n200 a_1560_n22142.n30 0.552
R8777 a_1560_n22142.n231 a_1560_n22142.n20 0.552
R8778 a_1560_n22142.n232 a_1560_n22142.n21 0.552
R8779 a_1560_n22142.n233 a_1560_n22142.n24 0.552
R8780 a_1560_n22142.n234 a_1560_n22142.n25 0.552
R8781 a_1560_n22142.n239 a_1560_n22142.n26 0.552
R8782 a_1560_n22142.n13 a_1560_n22142.n316 0.552
R8783 a_1560_n22142.n10 a_1560_n22142.n315 0.552
R8784 a_1560_n22142.n123 a_1560_n22142.n42 0.552
R8785 a_1560_n22142.n124 a_1560_n22142.n43 0.552
R8786 a_1560_n22142.n125 a_1560_n22142.n44 0.552
R8787 a_1560_n22142.n82 a_1560_n22142.n51 0.552
R8788 a_1560_n22142.n87 a_1560_n22142.n52 0.552
R8789 a_1560_n22142.n138 a_1560_n22142.n39 0.552
R8790 a_1560_n22142.n139 a_1560_n22142.n40 0.552
R8791 a_1560_n22142.n140 a_1560_n22142.n41 0.552
R8792 a_1560_n22142.n106 a_1560_n22142.n46 0.552
R8793 a_1560_n22142.n88 a_1560_n22142.n53 0.552
R8794 a_1560_n22142.n16 a_1560_n22142.n254 0.552
R8795 a_1560_n22142.n333 a_1560_n22142.n321 0.521
R8796 a_1560_n22142.n334 a_1560_n22142.n60 0.506
R8797 a_1560_n22142.n55 a_1560_n22142.n319 0.496
R8798 a_1560_n22142.n3 a_1560_n22142.n330 0.496
R8799 a_1560_n22142.n18 a_1560_n22142.n318 0.489
R8800 a_1560_n22142.n1 a_1560_n22142.n4 0.485
R8801 a_1560_n22142.n306 a_1560_n22142.n6 0.485
R8802 a_1560_n22142.n0 a_1560_n22142.n8 0.485
R8803 a_1560_n22142.n0 a_1560_n22142.n306 0.442
R8804 a_1560_n22142.n1 a_1560_n22142.n0 0.441
R8805 a_1560_n22142.n332 a_1560_n22142.n331 0.437
R8806 a_1560_n22142.n321 a_1560_n22142.n320 0.421
R8807 a_1560_n22142.n176 a_1560_n22142.n156 0.417
R8808 a_1560_n22142.n156 a_1560_n22142.n106 0.417
R8809 a_1560_n22142.n155 a_1560_n22142.n140 0.417
R8810 a_1560_n22142.n140 a_1560_n22142.n125 0.417
R8811 a_1560_n22142.n232 a_1560_n22142.n222 0.417
R8812 a_1560_n22142.n315 a_1560_n22142.n289 0.417
R8813 a_1560_n22142.n289 a_1560_n22142.n288 0.417
R8814 a_1560_n22142.n316 a_1560_n22142.n283 0.417
R8815 a_1560_n22142.n283 a_1560_n22142.n278 0.417
R8816 a_1560_n22142.n255 a_1560_n22142.n249 0.417
R8817 a_1560_n22142.n239 a_1560_n22142.n200 0.417
R8818 a_1560_n22142.n200 a_1560_n22142.n181 0.417
R8819 a_1560_n22142.n181 a_1560_n22142.n97 0.417
R8820 a_1560_n22142.n97 a_1560_n22142.n88 0.417
R8821 a_1560_n22142.n88 a_1560_n22142.n87 0.417
R8822 a_1560_n22142.n317 a_1560_n22142.n269 0.417
R8823 a_1560_n22142.n269 a_1560_n22142.n264 0.417
R8824 a_1560_n22142.n264 a_1560_n22142.n263 0.417
R8825 a_1560_n22142.n263 a_1560_n22142.n256 0.417
R8826 a_1560_n22142.n256 a_1560_n22142.n244 0.417
R8827 a_1560_n22142.n9 a_1560_n22142.n293 0.285
R8828 a_1560_n22142.n8 a_1560_n22142.n297 0.285
R8829 a_1560_n22142.n7 a_1560_n22142.n301 0.285
R8830 a_1560_n22142.n6 a_1560_n22142.n305 0.285
R8831 a_1560_n22142.n5 a_1560_n22142.n310 0.285
R8832 a_1560_n22142.n4 a_1560_n22142.n314 0.285
R8833 a_1560_n22142.n55 a_1560_n22142.n65 0.281
R8834 a_1560_n22142.n54 a_1560_n22142.n69 0.281
R8835 a_1560_n22142.n53 a_1560_n22142.n73 0.281
R8836 a_1560_n22142.n52 a_1560_n22142.n77 0.281
R8837 a_1560_n22142.n51 a_1560_n22142.n81 0.281
R8838 a_1560_n22142.n50 a_1560_n22142.n86 0.281
R8839 a_1560_n22142.n49 a_1560_n22142.n92 0.281
R8840 a_1560_n22142.n48 a_1560_n22142.n96 0.281
R8841 a_1560_n22142.n47 a_1560_n22142.n101 0.281
R8842 a_1560_n22142.n46 a_1560_n22142.n105 0.281
R8843 a_1560_n22142.n45 a_1560_n22142.n110 0.281
R8844 a_1560_n22142.n44 a_1560_n22142.n114 0.281
R8845 a_1560_n22142.n43 a_1560_n22142.n118 0.281
R8846 a_1560_n22142.n42 a_1560_n22142.n122 0.281
R8847 a_1560_n22142.n41 a_1560_n22142.n129 0.281
R8848 a_1560_n22142.n40 a_1560_n22142.n133 0.281
R8849 a_1560_n22142.n39 a_1560_n22142.n137 0.281
R8850 a_1560_n22142.n38 a_1560_n22142.n144 0.281
R8851 a_1560_n22142.n37 a_1560_n22142.n148 0.281
R8852 a_1560_n22142.n36 a_1560_n22142.n152 0.281
R8853 a_1560_n22142.n35 a_1560_n22142.n160 0.281
R8854 a_1560_n22142.n34 a_1560_n22142.n164 0.281
R8855 a_1560_n22142.n33 a_1560_n22142.n168 0.281
R8856 a_1560_n22142.n32 a_1560_n22142.n172 0.281
R8857 a_1560_n22142.n31 a_1560_n22142.n180 0.281
R8858 a_1560_n22142.n30 a_1560_n22142.n185 0.281
R8859 a_1560_n22142.n29 a_1560_n22142.n189 0.281
R8860 a_1560_n22142.n28 a_1560_n22142.n193 0.281
R8861 a_1560_n22142.n27 a_1560_n22142.n199 0.281
R8862 a_1560_n22142.n26 a_1560_n22142.n204 0.281
R8863 a_1560_n22142.n25 a_1560_n22142.n208 0.281
R8864 a_1560_n22142.n24 a_1560_n22142.n212 0.281
R8865 a_1560_n22142.n23 a_1560_n22142.n216 0.281
R8866 a_1560_n22142.n22 a_1560_n22142.n220 0.281
R8867 a_1560_n22142.n21 a_1560_n22142.n226 0.281
R8868 a_1560_n22142.n20 a_1560_n22142.n230 0.281
R8869 a_1560_n22142.n19 a_1560_n22142.n238 0.281
R8870 a_1560_n22142.n18 a_1560_n22142.n243 0.281
R8871 a_1560_n22142.n17 a_1560_n22142.n248 0.281
R8872 a_1560_n22142.n16 a_1560_n22142.n253 0.281
R8873 a_1560_n22142.n15 a_1560_n22142.n260 0.281
R8874 a_1560_n22142.n14 a_1560_n22142.n268 0.281
R8875 a_1560_n22142.n13 a_1560_n22142.n273 0.281
R8876 a_1560_n22142.n12 a_1560_n22142.n277 0.281
R8877 a_1560_n22142.n11 a_1560_n22142.n282 0.281
R8878 a_1560_n22142.n10 a_1560_n22142.n287 0.281
R8879 a_1560_n22142.n3 a_1560_n22142.n325 0.281
R8880 a_1560_n22142.n2 a_1560_n22142.n329 0.281
R8881 a_1657_n21342.n95 a_1657_n21342.t100 13.851
R8882 a_1657_n21342.n116 a_1657_n21342.t135 13.851
R8883 a_1657_n21342.n77 a_1657_n21342.t88 13.851
R8884 a_1657_n21342.n40 a_1657_n21342.t69 13.851
R8885 a_1657_n21342.n41 a_1657_n21342.t80 13.851
R8886 a_1657_n21342.n68 a_1657_n21342.t126 13.851
R8887 a_1657_n21342.n80 a_1657_n21342.t78 13.851
R8888 a_1657_n21342.n113 a_1657_n21342.t81 13.851
R8889 a_1657_n21342.n71 a_1657_n21342.t127 13.851
R8890 a_1657_n21342.n74 a_1657_n21342.t121 13.851
R8891 a_1657_n21342.n14 a_1657_n21342.t115 13.851
R8892 a_1657_n21342.n36 a_1657_n21342.t122 13.851
R8893 a_1657_n21342.n33 a_1657_n21342.t71 13.851
R8894 a_1657_n21342.n50 a_1657_n21342.t128 13.851
R8895 a_1657_n21342.n57 a_1657_n21342.t139 13.851
R8896 a_1657_n21342.n54 a_1657_n21342.t90 13.851
R8897 a_1657_n21342.n92 a_1657_n21342.t138 13.851
R8898 a_1657_n21342.n98 a_1657_n21342.t150 13.851
R8899 a_1657_n21342.n110 a_1657_n21342.t70 13.851
R8900 a_1657_n21342.n24 a_1657_n21342.t120 13.851
R8901 a_1657_n21342.n27 a_1657_n21342.t112 13.851
R8902 a_1657_n21342.n30 a_1657_n21342.t63 13.851
R8903 a_1657_n21342.n9 a_1657_n21342.t108 13.851
R8904 a_1657_n21342.n10 a_1657_n21342.t113 13.851
R8905 a_1657_n21342.n61 a_1657_n21342.t76 13.851
R8906 a_1657_n21342.n65 a_1657_n21342.t84 13.851
R8907 a_1657_n21342.n62 a_1657_n21342.t130 13.851
R8908 a_1657_n21342.n107 a_1657_n21342.t83 13.851
R8909 a_1657_n21342.n104 a_1657_n21342.t92 13.851
R8910 a_1657_n21342.n101 a_1657_n21342.t142 13.851
R8911 a_1657_n21342.n83 a_1657_n21342.t73 13.851
R8912 a_1657_n21342.n86 a_1657_n21342.t148 13.851
R8913 a_1657_n21342.n89 a_1657_n21342.t106 13.851
R8914 a_1657_n21342.n51 a_1657_n21342.t65 13.851
R8915 a_1657_n21342.n44 a_1657_n21342.t137 13.851
R8916 a_1657_n21342.n47 a_1657_n21342.t99 13.851
R8917 a_1657_n21342.n1 a_1657_n21342.t60 13.851
R8918 a_1657_n21342.n5 a_1657_n21342.t62 13.851
R8919 a_1657_n21342.n2 a_1657_n21342.t109 13.851
R8920 a_1657_n21342.n21 a_1657_n21342.t61 13.851
R8921 a_1657_n21342.n18 a_1657_n21342.t64 13.851
R8922 a_1657_n21342.n15 a_1657_n21342.t116 13.851
R8923 a_1657_n21342.n125 a_1657_n21342.t93 13.851
R8924 a_1657_n21342.n128 a_1657_n21342.t143 13.851
R8925 a_1657_n21342.n131 a_1657_n21342.t131 13.851
R8926 a_1657_n21342.n134 a_1657_n21342.t85 13.851
R8927 a_1657_n21342.n137 a_1657_n21342.t133 13.851
R8928 a_1657_n21342.n140 a_1657_n21342.t124 13.851
R8929 a_1657_n21342.n141 a_1657_n21342.t7 13.849
R8930 a_1657_n21342.n140 a_1657_n21342.t182 13.849
R8931 a_1657_n21342.n138 a_1657_n21342.t89 13.849
R8932 a_1657_n21342.n138 a_1657_n21342.t52 13.849
R8933 a_1657_n21342.n137 a_1657_n21342.t158 13.849
R8934 a_1657_n21342.n135 a_1657_n21342.t98 13.849
R8935 a_1657_n21342.n135 a_1657_n21342.t11 13.849
R8936 a_1657_n21342.n134 a_1657_n21342.t56 13.849
R8937 a_1657_n21342.n132 a_1657_n21342.t147 13.849
R8938 a_1657_n21342.n132 a_1657_n21342.t45 13.849
R8939 a_1657_n21342.n131 a_1657_n21342.t159 13.849
R8940 a_1657_n21342.n129 a_1657_n21342.t97 13.849
R8941 a_1657_n21342.n129 a_1657_n21342.t12 13.849
R8942 a_1657_n21342.n128 a_1657_n21342.t18 13.849
R8943 a_1657_n21342.n126 a_1657_n21342.t104 13.849
R8944 a_1657_n21342.n126 a_1657_n21342.t179 13.849
R8945 a_1657_n21342.n125 a_1657_n21342.t16 13.849
R8946 a_1657_n21342.n15 a_1657_n21342.t191 13.849
R8947 a_1657_n21342.n16 a_1657_n21342.t125 13.849
R8948 a_1657_n21342.n16 a_1657_n21342.t167 13.849
R8949 a_1657_n21342.n18 a_1657_n21342.t174 13.849
R8950 a_1657_n21342.n19 a_1657_n21342.t118 13.849
R8951 a_1657_n21342.n19 a_1657_n21342.t188 13.849
R8952 a_1657_n21342.n21 a_1657_n21342.t4 13.849
R8953 a_1657_n21342.n22 a_1657_n21342.t68 13.849
R8954 a_1657_n21342.n22 a_1657_n21342.t169 13.849
R8955 a_1657_n21342.n2 a_1657_n21342.t156 13.849
R8956 a_1657_n21342.n3 a_1657_n21342.t119 13.849
R8957 a_1657_n21342.n3 a_1657_n21342.t187 13.849
R8958 a_1657_n21342.n5 a_1657_n21342.t3 13.849
R8959 a_1657_n21342.n6 a_1657_n21342.t111 13.849
R8960 a_1657_n21342.n6 a_1657_n21342.t2 13.849
R8961 a_1657_n21342.n45 a_1657_n21342.t66 13.849
R8962 a_1657_n21342.n45 a_1657_n21342.t172 13.849
R8963 a_1657_n21342.n44 a_1657_n21342.t24 13.849
R8964 a_1657_n21342.n52 a_1657_n21342.t110 13.849
R8965 a_1657_n21342.n52 a_1657_n21342.t155 13.849
R8966 a_1657_n21342.n51 a_1657_n21342.t173 13.849
R8967 a_1657_n21342.n90 a_1657_n21342.t149 13.849
R8968 a_1657_n21342.n90 a_1657_n21342.t42 13.849
R8969 a_1657_n21342.n89 a_1657_n21342.t177 13.849
R8970 a_1657_n21342.n87 a_1657_n21342.t74 13.849
R8971 a_1657_n21342.n87 a_1657_n21342.t36 13.849
R8972 a_1657_n21342.n86 a_1657_n21342.t44 13.849
R8973 a_1657_n21342.n84 a_1657_n21342.t117 13.849
R8974 a_1657_n21342.n84 a_1657_n21342.t190 13.849
R8975 a_1657_n21342.n83 a_1657_n21342.t37 13.849
R8976 a_1657_n21342.n101 a_1657_n21342.t19 13.849
R8977 a_1657_n21342.n102 a_1657_n21342.t153 13.849
R8978 a_1657_n21342.n102 a_1657_n21342.t39 13.849
R8979 a_1657_n21342.n104 a_1657_n21342.t17 13.849
R8980 a_1657_n21342.n105 a_1657_n21342.t145 13.849
R8981 a_1657_n21342.n105 a_1657_n21342.t47 13.849
R8982 a_1657_n21342.n107 a_1657_n21342.t58 13.849
R8983 a_1657_n21342.n108 a_1657_n21342.t96 13.849
R8984 a_1657_n21342.n108 a_1657_n21342.t13 13.849
R8985 a_1657_n21342.n62 a_1657_n21342.t160 13.849
R8986 a_1657_n21342.n63 a_1657_n21342.t146 13.849
R8987 a_1657_n21342.n63 a_1657_n21342.t46 13.849
R8988 a_1657_n21342.n31 a_1657_n21342.t75 13.849
R8989 a_1657_n21342.n31 a_1657_n21342.t164 13.849
R8990 a_1657_n21342.n30 a_1657_n21342.t189 13.849
R8991 a_1657_n21342.n28 a_1657_n21342.t123 13.849
R8992 a_1657_n21342.n28 a_1657_n21342.t29 13.849
R8993 a_1657_n21342.n27 a_1657_n21342.t171 13.849
R8994 a_1657_n21342.n25 a_1657_n21342.t72 13.849
R8995 a_1657_n21342.n25 a_1657_n21342.t165 13.849
R8996 a_1657_n21342.n24 a_1657_n21342.t35 13.849
R8997 a_1657_n21342.n96 a_1657_n21342.t107 13.849
R8998 a_1657_n21342.n96 a_1657_n21342.t176 13.849
R8999 a_1657_n21342.n95 a_1657_n21342.t9 13.849
R9000 a_1657_n21342.n98 a_1657_n21342.t43 13.849
R9001 a_1657_n21342.n99 a_1657_n21342.t102 13.849
R9002 a_1657_n21342.n99 a_1657_n21342.t181 13.849
R9003 a_1657_n21342.n92 a_1657_n21342.t23 13.849
R9004 a_1657_n21342.n93 a_1657_n21342.t152 13.849
R9005 a_1657_n21342.n93 a_1657_n21342.t40 13.849
R9006 a_1657_n21342.n75 a_1657_n21342.t134 13.849
R9007 a_1657_n21342.n75 a_1657_n21342.t157 13.849
R9008 a_1657_n21342.n74 a_1657_n21342.t185 13.849
R9009 a_1657_n21342.n78 a_1657_n21342.t140 13.849
R9010 a_1657_n21342.n78 a_1657_n21342.t21 13.849
R9011 a_1657_n21342.n77 a_1657_n21342.t53 13.849
R9012 a_1657_n21342.n117 a_1657_n21342.t151 13.849
R9013 a_1657_n21342.n117 a_1657_n21342.t41 13.849
R9014 a_1657_n21342.n116 a_1657_n21342.t27 13.849
R9015 a_1657_n21342.n80 a_1657_n21342.t32 13.849
R9016 a_1657_n21342.n81 a_1657_n21342.t91 13.849
R9017 a_1657_n21342.n81 a_1657_n21342.t49 13.849
R9018 a_1657_n21342.n68 a_1657_n21342.t166 13.849
R9019 a_1657_n21342.n69 a_1657_n21342.t141 13.849
R9020 a_1657_n21342.n69 a_1657_n21342.t20 13.849
R9021 a_1657_n21342.n41 a_1657_n21342.t30 13.849
R9022 a_1657_n21342.n42 a_1657_n21342.t129 13.849
R9023 a_1657_n21342.n42 a_1657_n21342.t161 13.849
R9024 a_1657_n21342.n40 a_1657_n21342.t168 13.849
R9025 a_1657_n21342.n39 a_1657_n21342.t101 13.849
R9026 a_1657_n21342.n39 a_1657_n21342.t8 13.849
R9027 a_1657_n21342.n72 a_1657_n21342.t86 13.849
R9028 a_1657_n21342.n72 a_1657_n21342.t55 13.849
R9029 a_1657_n21342.n71 a_1657_n21342.t163 13.849
R9030 a_1657_n21342.n114 a_1657_n21342.t94 13.849
R9031 a_1657_n21342.n114 a_1657_n21342.t15 13.849
R9032 a_1657_n21342.n113 a_1657_n21342.t28 13.849
R9033 a_1657_n21342.n33 a_1657_n21342.t38 13.849
R9034 a_1657_n21342.n34 a_1657_n21342.t87 13.849
R9035 a_1657_n21342.n34 a_1657_n21342.t54 13.849
R9036 a_1657_n21342.n36 a_1657_n21342.t184 13.849
R9037 a_1657_n21342.n37 a_1657_n21342.t77 13.849
R9038 a_1657_n21342.n37 a_1657_n21342.t33 13.849
R9039 a_1657_n21342.n14 a_1657_n21342.t0 13.849
R9040 a_1657_n21342.n13 a_1657_n21342.t144 13.849
R9041 a_1657_n21342.n13 a_1657_n21342.t48 13.849
R9042 a_1657_n21342.n54 a_1657_n21342.t50 13.849
R9043 a_1657_n21342.n55 a_1657_n21342.t103 13.849
R9044 a_1657_n21342.n55 a_1657_n21342.t180 13.849
R9045 a_1657_n21342.n57 a_1657_n21342.t22 13.849
R9046 a_1657_n21342.n58 a_1657_n21342.t95 13.849
R9047 a_1657_n21342.n58 a_1657_n21342.t14 13.849
R9048 a_1657_n21342.n50 a_1657_n21342.t162 13.849
R9049 a_1657_n21342.n49 a_1657_n21342.t59 13.849
R9050 a_1657_n21342.n49 a_1657_n21342.t5 13.849
R9051 a_1657_n21342.n111 a_1657_n21342.t82 13.849
R9052 a_1657_n21342.n111 a_1657_n21342.t26 13.849
R9053 a_1657_n21342.n110 a_1657_n21342.t183 13.849
R9054 a_1657_n21342.n10 a_1657_n21342.t170 13.849
R9055 a_1657_n21342.n11 a_1657_n21342.t67 13.849
R9056 a_1657_n21342.n11 a_1657_n21342.t186 13.849
R9057 a_1657_n21342.n9 a_1657_n21342.t175 13.849
R9058 a_1657_n21342.n8 a_1657_n21342.t132 13.849
R9059 a_1657_n21342.n8 a_1657_n21342.t51 13.849
R9060 a_1657_n21342.n65 a_1657_n21342.t57 13.849
R9061 a_1657_n21342.n66 a_1657_n21342.t136 13.849
R9062 a_1657_n21342.n66 a_1657_n21342.t25 13.849
R9063 a_1657_n21342.n61 a_1657_n21342.t34 13.849
R9064 a_1657_n21342.n60 a_1657_n21342.t105 13.849
R9065 a_1657_n21342.n60 a_1657_n21342.t178 13.849
R9066 a_1657_n21342.n47 a_1657_n21342.t10 13.849
R9067 a_1657_n21342.n46 a_1657_n21342.t114 13.849
R9068 a_1657_n21342.n46 a_1657_n21342.t1 13.849
R9069 a_1657_n21342.n1 a_1657_n21342.t6 13.849
R9070 a_1657_n21342.n0 a_1657_n21342.t79 13.849
R9071 a_1657_n21342.n0 a_1657_n21342.t31 13.849
R9072 a_1657_n21342.t154 a_1657_n21342.n141 13.849
R9073 a_1657_n21342.n94 a_1657_n21342.n91 2.199
R9074 a_1657_n21342.n106 a_1657_n21342.n100 2.199
R9075 a_1657_n21342.n29 a_1657_n21342.n23 2.199
R9076 a_1657_n21342.n82 a_1657_n21342.n76 2.199
R9077 a_1657_n21342.n133 a_1657_n21342.n82 2.199
R9078 a_1657_n21342.n133 a_1657_n21342.n109 2.199
R9079 a_1657_n21342.n109 a_1657_n21342.n94 2.199
R9080 a_1657_n21342.n56 a_1657_n21342.n53 2.199
R9081 a_1657_n21342.n127 a_1657_n21342.n118 2.199
R9082 a_1657_n21342.n118 a_1657_n21342.n115 2.199
R9083 a_1657_n21342.n115 a_1657_n21342.n112 2.199
R9084 a_1657_n21342.n35 a_1657_n21342.n32 2.199
R9085 a_1657_n21342.n136 a_1657_n21342.n70 2.199
R9086 a_1657_n21342.n124 a_1657_n21342.n123 2.199
R9087 a_1657_n21342.n123 a_1657_n21342.n122 2.199
R9088 a_1657_n21342.n59 a_1657_n21342.n48 2.199
R9089 a_1657_n21342.n67 a_1657_n21342.n59 2.199
R9090 a_1657_n21342.n139 a_1657_n21342.n67 2.199
R9091 a_1657_n21342.n139 a_1657_n21342.n43 2.199
R9092 a_1657_n21342.n43 a_1657_n21342.n38 2.199
R9093 a_1657_n21342.n38 a_1657_n21342.n12 2.199
R9094 a_1657_n21342.n12 a_1657_n21342.n7 2.199
R9095 a_1657_n21342.n120 a_1657_n21342.n119 2.199
R9096 a_1657_n21342.n121 a_1657_n21342.n120 2.199
R9097 a_1657_n21342.n124 a_1657_n21342.n121 2.199
R9098 a_1657_n21342.n96 a_1657_n21342.n95 1.121
R9099 a_1657_n21342.n117 a_1657_n21342.n116 1.121
R9100 a_1657_n21342.n78 a_1657_n21342.n77 1.121
R9101 a_1657_n21342.n114 a_1657_n21342.n113 1.121
R9102 a_1657_n21342.n72 a_1657_n21342.n71 1.121
R9103 a_1657_n21342.n75 a_1657_n21342.n74 1.121
R9104 a_1657_n21342.n111 a_1657_n21342.n110 1.121
R9105 a_1657_n21342.n25 a_1657_n21342.n24 1.121
R9106 a_1657_n21342.n28 a_1657_n21342.n27 1.121
R9107 a_1657_n21342.n31 a_1657_n21342.n30 1.121
R9108 a_1657_n21342.n84 a_1657_n21342.n83 1.121
R9109 a_1657_n21342.n87 a_1657_n21342.n86 1.121
R9110 a_1657_n21342.n90 a_1657_n21342.n89 1.121
R9111 a_1657_n21342.n52 a_1657_n21342.n51 1.121
R9112 a_1657_n21342.n45 a_1657_n21342.n44 1.121
R9113 a_1657_n21342.n126 a_1657_n21342.n125 1.121
R9114 a_1657_n21342.n129 a_1657_n21342.n128 1.121
R9115 a_1657_n21342.n132 a_1657_n21342.n131 1.121
R9116 a_1657_n21342.n135 a_1657_n21342.n134 1.121
R9117 a_1657_n21342.n138 a_1657_n21342.n137 1.121
R9118 a_1657_n21342.n141 a_1657_n21342.n140 1.121
R9119 a_1657_n21342.n40 a_1657_n21342.n39 1.121
R9120 a_1657_n21342.n42 a_1657_n21342.n41 1.121
R9121 a_1657_n21342.n69 a_1657_n21342.n68 1.121
R9122 a_1657_n21342.n81 a_1657_n21342.n80 1.121
R9123 a_1657_n21342.n14 a_1657_n21342.n13 1.121
R9124 a_1657_n21342.n37 a_1657_n21342.n36 1.121
R9125 a_1657_n21342.n34 a_1657_n21342.n33 1.121
R9126 a_1657_n21342.n50 a_1657_n21342.n49 1.121
R9127 a_1657_n21342.n58 a_1657_n21342.n57 1.121
R9128 a_1657_n21342.n55 a_1657_n21342.n54 1.121
R9129 a_1657_n21342.n93 a_1657_n21342.n92 1.121
R9130 a_1657_n21342.n99 a_1657_n21342.n98 1.121
R9131 a_1657_n21342.n9 a_1657_n21342.n8 1.121
R9132 a_1657_n21342.n11 a_1657_n21342.n10 1.121
R9133 a_1657_n21342.n61 a_1657_n21342.n60 1.121
R9134 a_1657_n21342.n66 a_1657_n21342.n65 1.121
R9135 a_1657_n21342.n63 a_1657_n21342.n62 1.121
R9136 a_1657_n21342.n108 a_1657_n21342.n107 1.121
R9137 a_1657_n21342.n105 a_1657_n21342.n104 1.121
R9138 a_1657_n21342.n102 a_1657_n21342.n101 1.121
R9139 a_1657_n21342.n47 a_1657_n21342.n46 1.121
R9140 a_1657_n21342.n1 a_1657_n21342.n0 1.121
R9141 a_1657_n21342.n6 a_1657_n21342.n5 1.121
R9142 a_1657_n21342.n3 a_1657_n21342.n2 1.121
R9143 a_1657_n21342.n22 a_1657_n21342.n21 1.121
R9144 a_1657_n21342.n19 a_1657_n21342.n18 1.121
R9145 a_1657_n21342.n16 a_1657_n21342.n15 1.121
R9146 a_1657_n21342.n97 a_1657_n21342.n96 0.552
R9147 a_1657_n21342.n118 a_1657_n21342.n117 0.552
R9148 a_1657_n21342.n79 a_1657_n21342.n78 0.552
R9149 a_1657_n21342.n43 a_1657_n21342.n42 0.552
R9150 a_1657_n21342.n70 a_1657_n21342.n69 0.552
R9151 a_1657_n21342.n82 a_1657_n21342.n81 0.552
R9152 a_1657_n21342.n115 a_1657_n21342.n114 0.552
R9153 a_1657_n21342.n73 a_1657_n21342.n72 0.552
R9154 a_1657_n21342.n76 a_1657_n21342.n75 0.552
R9155 a_1657_n21342.n38 a_1657_n21342.n37 0.552
R9156 a_1657_n21342.n35 a_1657_n21342.n34 0.552
R9157 a_1657_n21342.n59 a_1657_n21342.n58 0.552
R9158 a_1657_n21342.n56 a_1657_n21342.n55 0.552
R9159 a_1657_n21342.n94 a_1657_n21342.n93 0.552
R9160 a_1657_n21342.n100 a_1657_n21342.n99 0.552
R9161 a_1657_n21342.n112 a_1657_n21342.n111 0.552
R9162 a_1657_n21342.n26 a_1657_n21342.n25 0.552
R9163 a_1657_n21342.n29 a_1657_n21342.n28 0.552
R9164 a_1657_n21342.n32 a_1657_n21342.n31 0.552
R9165 a_1657_n21342.n12 a_1657_n21342.n11 0.552
R9166 a_1657_n21342.n67 a_1657_n21342.n66 0.552
R9167 a_1657_n21342.n64 a_1657_n21342.n63 0.552
R9168 a_1657_n21342.n109 a_1657_n21342.n108 0.552
R9169 a_1657_n21342.n106 a_1657_n21342.n105 0.552
R9170 a_1657_n21342.n103 a_1657_n21342.n102 0.552
R9171 a_1657_n21342.n85 a_1657_n21342.n84 0.552
R9172 a_1657_n21342.n88 a_1657_n21342.n87 0.552
R9173 a_1657_n21342.n91 a_1657_n21342.n90 0.552
R9174 a_1657_n21342.n53 a_1657_n21342.n52 0.552
R9175 a_1657_n21342.n48 a_1657_n21342.n45 0.552
R9176 a_1657_n21342.n7 a_1657_n21342.n6 0.552
R9177 a_1657_n21342.n4 a_1657_n21342.n3 0.552
R9178 a_1657_n21342.n23 a_1657_n21342.n22 0.552
R9179 a_1657_n21342.n20 a_1657_n21342.n19 0.552
R9180 a_1657_n21342.n17 a_1657_n21342.n16 0.552
R9181 a_1657_n21342.n127 a_1657_n21342.n126 0.552
R9182 a_1657_n21342.n130 a_1657_n21342.n129 0.552
R9183 a_1657_n21342.n133 a_1657_n21342.n132 0.552
R9184 a_1657_n21342.n136 a_1657_n21342.n135 0.552
R9185 a_1657_n21342.n139 a_1657_n21342.n138 0.552
R9186 a_1657_n21342.n43 a_1657_n21342.n40 0.278
R9187 a_1657_n21342.n80 a_1657_n21342.n79 0.278
R9188 a_1657_n21342.n74 a_1657_n21342.n73 0.278
R9189 a_1657_n21342.n38 a_1657_n21342.n14 0.278
R9190 a_1657_n21342.n36 a_1657_n21342.n35 0.278
R9191 a_1657_n21342.n59 a_1657_n21342.n50 0.278
R9192 a_1657_n21342.n57 a_1657_n21342.n56 0.278
R9193 a_1657_n21342.n98 a_1657_n21342.n97 0.278
R9194 a_1657_n21342.n27 a_1657_n21342.n26 0.278
R9195 a_1657_n21342.n30 a_1657_n21342.n29 0.278
R9196 a_1657_n21342.n12 a_1657_n21342.n9 0.278
R9197 a_1657_n21342.n67 a_1657_n21342.n61 0.278
R9198 a_1657_n21342.n65 a_1657_n21342.n64 0.278
R9199 a_1657_n21342.n107 a_1657_n21342.n106 0.278
R9200 a_1657_n21342.n104 a_1657_n21342.n103 0.278
R9201 a_1657_n21342.n86 a_1657_n21342.n85 0.278
R9202 a_1657_n21342.n89 a_1657_n21342.n88 0.278
R9203 a_1657_n21342.n48 a_1657_n21342.n47 0.278
R9204 a_1657_n21342.n7 a_1657_n21342.n1 0.278
R9205 a_1657_n21342.n5 a_1657_n21342.n4 0.278
R9206 a_1657_n21342.n21 a_1657_n21342.n20 0.278
R9207 a_1657_n21342.n18 a_1657_n21342.n17 0.278
R9208 a_1657_n21342.n125 a_1657_n21342.n124 0.278
R9209 a_1657_n21342.n128 a_1657_n21342.n127 0.278
R9210 a_1657_n21342.n131 a_1657_n21342.n130 0.278
R9211 a_1657_n21342.n134 a_1657_n21342.n133 0.278
R9212 a_1657_n21342.n137 a_1657_n21342.n136 0.278
R9213 a_1657_n21342.n140 a_1657_n21342.n139 0.278
R9214 casc_p.n361 casc_p.t34 48.207
R9215 casc_p.n364 casc_p.t31 48.207
R9216 casc_p.n367 casc_p.t4 48.207
R9217 casc_p.n370 casc_p.t61 48.207
R9218 casc_p.n330 casc_p.t37 48.207
R9219 casc_p.n333 casc_p.t7 48.207
R9220 casc_p.n284 casc_p.t10 48.207
R9221 casc_p.n287 casc_p.t40 48.207
R9222 casc_p.n238 casc_p.t46 48.207
R9223 casc_p.n241 casc_p.t13 48.207
R9224 casc_p.n192 casc_p.t22 48.207
R9225 casc_p.n195 casc_p.t49 48.207
R9226 casc_p.n146 casc_p.t52 48.207
R9227 casc_p.n149 casc_p.t19 48.207
R9228 casc_p.n88 casc_p.t28 48.207
R9229 casc_p.n91 casc_p.t16 48.207
R9230 casc_p.n94 casc_p.t58 48.207
R9231 casc_p.n97 casc_p.t43 48.207
R9232 casc_p.n100 casc_p.t25 48.207
R9233 casc_p.n103 casc_p.t55 48.207
R9234 casc_p.n2 casc_p.t222 48.207
R9235 casc_p.n1 casc_p.t319 48.207
R9236 casc_p.n334 casc_p.t230 24.628
R9237 casc_p.n299 casc_p.t202 24.628
R9238 casc_p.n288 casc_p.t358 24.628
R9239 casc_p.n253 casc_p.t353 24.628
R9240 casc_p.n242 casc_p.t177 24.628
R9241 casc_p.n207 casc_p.t173 24.628
R9242 casc_p.n196 casc_p.t320 24.628
R9243 casc_p.n161 casc_p.t309 24.628
R9244 casc_p.n150 casc_p.t139 24.628
R9245 casc_p.n115 casc_p.t151 24.628
R9246 casc_p.n104 casc_p.t298 24.628
R9247 casc_p.n61 casc_p.t292 24.628
R9248 casc_p.n50 casc_p.t118 24.628
R9249 casc_p.n3 casc_p.t283 24.628
R9250 casc_p.n39 casc_p.t195 24.628
R9251 casc_p.n373 casc_p.t380 24.628
R9252 casc_p.n298 casc_p.t148 23.97
R9253 casc_p.n252 casc_p.t291 23.97
R9254 casc_p.n206 casc_p.t112 23.97
R9255 casc_p.n160 casc_p.t259 23.97
R9256 casc_p.n114 casc_p.t100 23.97
R9257 casc_p.n60 casc_p.t252 23.97
R9258 casc_p.n49 casc_p.t385 23.97
R9259 casc_p.n383 casc_p.t182 23.97
R9260 casc_p.n372 casc_p.t376 23.967
R9261 casc_p.n371 casc_p.t204 23.967
R9262 casc_p.n358 casc_p.t395 23.967
R9263 casc_p.n357 casc_p.t226 23.967
R9264 casc_p.n356 casc_p.t88 23.967
R9265 casc_p.n355 casc_p.t389 23.967
R9266 casc_p.n354 casc_p.t248 23.967
R9267 casc_p.n353 casc_p.t82 23.967
R9268 casc_p.n352 casc_p.t134 23.967
R9269 casc_p.n351 casc_p.t101 23.967
R9270 casc_p.n350 casc_p.t293 23.967
R9271 casc_p.n349 casc_p.t260 23.967
R9272 casc_p.n348 casc_p.t130 23.967
R9273 casc_p.n347 casc_p.t279 23.967
R9274 casc_p.n346 casc_p.t163 23.967
R9275 casc_p.n345 casc_p.t117 23.967
R9276 casc_p.n344 casc_p.t323 23.967
R9277 casc_p.n343 casc_p.t149 23.967
R9278 casc_p.n342 casc_p.t352 23.967
R9279 casc_p.n341 casc_p.t306 23.967
R9280 casc_p.n340 casc_p.t379 23.967
R9281 casc_p.n339 casc_p.t349 23.967
R9282 casc_p.n338 casc_p.t218 23.967
R9283 casc_p.n337 casc_p.t370 23.967
R9284 casc_p.n336 casc_p.t238 23.967
R9285 casc_p.n335 casc_p.t208 23.967
R9286 casc_p.n334 casc_p.t74 23.967
R9287 casc_p.n327 casc_p.t372 23.967
R9288 casc_p.n326 casc_p.t339 23.967
R9289 casc_p.n325 casc_p.t210 23.967
R9290 casc_p.n324 casc_p.t175 23.967
R9291 casc_p.n323 casc_p.t369 23.967
R9292 casc_p.n322 casc_p.t200 23.967
R9293 casc_p.n321 casc_p.t393 23.967
R9294 casc_p.n320 casc_p.t362 23.967
R9295 casc_p.n319 casc_p.t229 23.967
R9296 casc_p.n318 casc_p.t386 23.967
R9297 casc_p.n317 casc_p.t107 23.967
R9298 casc_p.n316 casc_p.t85 23.967
R9299 casc_p.n315 casc_p.t265 23.967
R9300 casc_p.n314 casc_p.t246 23.967
R9301 casc_p.n313 casc_p.t106 23.967
R9302 casc_p.n312 casc_p.t257 23.967
R9303 casc_p.n311 casc_p.t129 23.967
R9304 casc_p.n310 casc_p.t97 23.967
R9305 casc_p.n309 casc_p.t288 23.967
R9306 casc_p.n308 casc_p.t113 23.967
R9307 casc_p.n307 casc_p.t315 23.967
R9308 casc_p.n306 casc_p.t269 23.967
R9309 casc_p.n305 casc_p.t357 23.967
R9310 casc_p.n304 casc_p.t310 23.967
R9311 casc_p.n303 casc_p.t189 23.967
R9312 casc_p.n302 casc_p.t343 23.967
R9313 casc_p.n301 casc_p.t213 23.967
R9314 casc_p.n300 casc_p.t179 23.967
R9315 casc_p.n299 casc_p.t373 23.967
R9316 casc_p.n297 casc_p.t231 23.967
R9317 casc_p.n296 casc_p.t365 23.967
R9318 casc_p.n295 casc_p.t211 23.967
R9319 casc_p.n294 casc_p.t342 23.967
R9320 casc_p.n293 casc_p.t374 23.967
R9321 casc_p.n292 casc_p.t180 23.967
R9322 casc_p.n291 casc_p.t214 23.967
R9323 casc_p.n290 casc_p.t345 23.967
R9324 casc_p.n289 casc_p.t191 23.967
R9325 casc_p.n288 casc_p.t312 23.967
R9326 casc_p.n281 casc_p.t196 23.967
R9327 casc_p.n280 casc_p.t158 23.967
R9328 casc_p.n279 casc_p.t359 23.967
R9329 casc_p.n278 casc_p.t317 23.967
R9330 casc_p.n277 casc_p.t194 23.967
R9331 casc_p.n276 casc_p.t347 23.967
R9332 casc_p.n275 casc_p.t216 23.967
R9333 casc_p.n274 casc_p.t184 23.967
R9334 casc_p.n273 casc_p.t377 23.967
R9335 casc_p.n272 casc_p.t205 23.967
R9336 casc_p.n271 casc_p.t256 23.967
R9337 casc_p.n270 casc_p.t233 23.967
R9338 casc_p.n269 casc_p.t96 23.967
R9339 casc_p.n268 casc_p.t70 23.967
R9340 casc_p.n267 casc_p.t255 23.967
R9341 casc_p.n266 casc_p.t89 23.967
R9342 casc_p.n265 casc_p.t268 23.967
R9343 casc_p.n264 casc_p.t249 23.967
R9344 casc_p.n263 casc_p.t110 23.967
R9345 casc_p.n262 casc_p.t261 23.967
R9346 casc_p.n261 casc_p.t135 23.967
R9347 casc_p.n260 casc_p.t102 23.967
R9348 casc_p.n259 casc_p.t176 23.967
R9349 casc_p.n258 casc_p.t131 23.967
R9350 casc_p.n257 casc_p.t335 23.967
R9351 casc_p.n256 casc_p.t164 23.967
R9352 casc_p.n255 casc_p.t361 23.967
R9353 casc_p.n254 casc_p.t324 23.967
R9354 casc_p.n253 casc_p.t197 23.967
R9355 casc_p.n251 casc_p.t383 23.967
R9356 casc_p.n250 casc_p.t188 23.967
R9357 casc_p.n249 casc_p.t360 23.967
R9358 casc_p.n248 casc_p.t162 23.967
R9359 casc_p.n247 casc_p.t199 23.967
R9360 casc_p.n246 casc_p.t326 23.967
R9361 casc_p.n245 casc_p.t363 23.967
R9362 casc_p.n244 casc_p.t166 23.967
R9363 casc_p.n243 casc_p.t337 23.967
R9364 casc_p.n242 casc_p.t133 23.967
R9365 casc_p.n235 casc_p.t341 23.967
R9366 casc_p.n234 casc_p.t296 23.967
R9367 casc_p.n233 casc_p.t178 23.967
R9368 casc_p.n232 casc_p.t137 23.967
R9369 casc_p.n231 casc_p.t340 23.967
R9370 casc_p.n230 casc_p.t169 23.967
R9371 casc_p.n229 casc_p.t364 23.967
R9372 casc_p.n228 casc_p.t329 23.967
R9373 casc_p.n227 casc_p.t201 23.967
R9374 casc_p.n226 casc_p.t355 23.967
R9375 casc_p.n225 casc_p.t87 23.967
R9376 casc_p.n224 casc_p.t387 23.967
R9377 casc_p.n223 casc_p.t247 23.967
R9378 casc_p.n222 casc_p.t220 23.967
R9379 casc_p.n221 casc_p.t86 23.967
R9380 casc_p.n220 casc_p.t241 23.967
R9381 casc_p.n219 casc_p.t98 23.967
R9382 casc_p.n218 casc_p.t77 23.967
R9383 casc_p.n217 casc_p.t258 23.967
R9384 casc_p.n216 casc_p.t92 23.967
R9385 casc_p.n215 casc_p.t272 23.967
R9386 casc_p.n214 casc_p.t254 23.967
R9387 casc_p.n213 casc_p.t316 23.967
R9388 casc_p.n212 casc_p.t270 23.967
R9389 casc_p.n211 casc_p.t153 23.967
R9390 casc_p.n210 casc_p.t300 23.967
R9391 casc_p.n209 casc_p.t183 23.967
R9392 casc_p.n208 casc_p.t142 23.967
R9393 casc_p.n207 casc_p.t344 23.967
R9394 casc_p.n205 casc_p.t203 23.967
R9395 casc_p.n204 casc_p.t334 23.967
R9396 casc_p.n203 casc_p.t181 23.967
R9397 casc_p.n202 casc_p.t299 23.967
R9398 casc_p.n201 casc_p.t346 23.967
R9399 casc_p.n200 casc_p.t143 23.967
R9400 casc_p.n199 casc_p.t185 23.967
R9401 casc_p.n198 casc_p.t301 23.967
R9402 casc_p.n197 casc_p.t156 23.967
R9403 casc_p.n196 casc_p.t271 23.967
R9404 casc_p.n189 casc_p.t160 23.967
R9405 casc_p.n188 casc_p.t114 23.967
R9406 casc_p.n187 casc_p.t321 23.967
R9407 casc_p.n186 casc_p.t273 23.967
R9408 casc_p.n185 casc_p.t159 23.967
R9409 casc_p.n184 casc_p.t303 23.967
R9410 casc_p.n183 casc_p.t186 23.967
R9411 casc_p.n182 casc_p.t144 23.967
R9412 casc_p.n181 casc_p.t348 23.967
R9413 casc_p.n180 casc_p.t174 23.967
R9414 casc_p.n179 casc_p.t235 23.967
R9415 casc_p.n178 casc_p.t206 23.967
R9416 casc_p.n177 casc_p.t71 23.967
R9417 casc_p.n176 casc_p.t366 23.967
R9418 casc_p.n175 casc_p.t234 23.967
R9419 casc_p.n174 casc_p.t390 23.967
R9420 casc_p.n173 casc_p.t250 23.967
R9421 casc_p.n172 casc_p.t227 23.967
R9422 casc_p.n171 casc_p.t90 23.967
R9423 casc_p.n170 casc_p.t244 23.967
R9424 casc_p.n169 casc_p.t105 23.967
R9425 casc_p.n168 casc_p.t83 23.967
R9426 casc_p.n167 casc_p.t136 23.967
R9427 casc_p.n166 casc_p.t103 23.967
R9428 casc_p.n165 casc_p.t294 23.967
R9429 casc_p.n164 casc_p.t121 23.967
R9430 casc_p.n163 casc_p.t328 23.967
R9431 casc_p.n162 casc_p.t280 23.967
R9432 casc_p.n161 casc_p.t165 23.967
R9433 casc_p.n159 casc_p.t354 23.967
R9434 casc_p.n158 casc_p.t150 23.967
R9435 casc_p.n157 casc_p.t327 23.967
R9436 casc_p.n156 casc_p.t120 23.967
R9437 casc_p.n155 casc_p.t167 23.967
R9438 casc_p.n154 casc_p.t281 23.967
R9439 casc_p.n153 casc_p.t331 23.967
R9440 casc_p.n152 casc_p.t123 23.967
R9441 casc_p.n151 casc_p.t295 23.967
R9442 casc_p.n150 casc_p.t104 23.967
R9443 casc_p.n143 casc_p.t325 23.967
R9444 casc_p.n142 casc_p.t278 23.967
R9445 casc_p.n141 casc_p.t161 23.967
R9446 casc_p.n140 casc_p.t115 23.967
R9447 casc_p.n139 casc_p.t322 23.967
R9448 casc_p.n138 casc_p.t147 23.967
R9449 casc_p.n137 casc_p.t350 23.967
R9450 casc_p.n136 casc_p.t305 23.967
R9451 casc_p.n135 casc_p.t187 23.967
R9452 casc_p.n134 casc_p.t338 23.967
R9453 casc_p.n133 casc_p.t75 23.967
R9454 casc_p.n132 casc_p.t367 23.967
R9455 casc_p.n131 casc_p.t236 23.967
R9456 casc_p.n130 casc_p.t207 23.967
R9457 casc_p.n129 casc_p.t72 23.967
R9458 casc_p.n128 casc_p.t228 23.967
R9459 casc_p.n127 casc_p.t91 23.967
R9460 casc_p.n126 casc_p.t391 23.967
R9461 casc_p.n125 casc_p.t251 23.967
R9462 casc_p.n124 casc_p.t84 23.967
R9463 casc_p.n123 casc_p.t264 23.967
R9464 casc_p.n122 casc_p.t245 23.967
R9465 casc_p.n121 casc_p.t297 23.967
R9466 casc_p.n120 casc_p.t262 23.967
R9467 casc_p.n119 casc_p.t138 23.967
R9468 casc_p.n118 casc_p.t284 23.967
R9469 casc_p.n117 casc_p.t170 23.967
R9470 casc_p.n116 casc_p.t122 23.967
R9471 casc_p.n115 casc_p.t330 23.967
R9472 casc_p.n113 casc_p.t190 23.967
R9473 casc_p.n112 casc_p.t311 23.967
R9474 casc_p.n111 casc_p.t168 23.967
R9475 casc_p.n110 casc_p.t282 23.967
R9476 casc_p.n109 casc_p.t332 23.967
R9477 casc_p.n108 casc_p.t124 23.967
R9478 casc_p.n107 casc_p.t171 23.967
R9479 casc_p.n106 casc_p.t289 23.967
R9480 casc_p.n105 casc_p.t140 23.967
R9481 casc_p.n104 casc_p.t263 23.967
R9482 casc_p.n85 casc_p.t141 23.967
R9483 casc_p.n84 casc_p.t290 23.967
R9484 casc_p.n83 casc_p.t172 23.967
R9485 casc_p.n82 casc_p.t126 23.967
R9486 casc_p.n81 casc_p.t333 23.967
R9487 casc_p.n80 casc_p.t157 23.967
R9488 casc_p.n79 casc_p.t225 23.967
R9489 casc_p.n78 casc_p.t192 23.967
R9490 casc_p.n77 casc_p.t388 23.967
R9491 casc_p.n76 casc_p.t356 23.967
R9492 casc_p.n75 casc_p.t224 23.967
R9493 casc_p.n74 casc_p.t375 23.967
R9494 casc_p.n73 casc_p.t243 23.967
R9495 casc_p.n72 casc_p.t212 23.967
R9496 casc_p.n71 casc_p.t81 23.967
R9497 casc_p.n70 casc_p.t232 23.967
R9498 casc_p.n69 casc_p.t95 23.967
R9499 casc_p.n68 casc_p.t394 23.967
R9500 casc_p.n67 casc_p.t116 23.967
R9501 casc_p.n66 casc_p.t93 23.967
R9502 casc_p.n65 casc_p.t274 23.967
R9503 casc_p.n64 casc_p.t109 23.967
R9504 casc_p.n63 casc_p.t304 23.967
R9505 casc_p.n62 casc_p.t266 23.967
R9506 casc_p.n61 casc_p.t145 23.967
R9507 casc_p.n59 casc_p.t336 23.967
R9508 casc_p.n58 casc_p.t132 23.967
R9509 casc_p.n57 casc_p.t302 23.967
R9510 casc_p.n56 casc_p.t108 23.967
R9511 casc_p.n55 casc_p.t146 23.967
R9512 casc_p.n54 casc_p.t267 23.967
R9513 casc_p.n53 casc_p.t307 23.967
R9514 casc_p.n52 casc_p.t111 23.967
R9515 casc_p.n51 casc_p.t276 23.967
R9516 casc_p.n50 casc_p.t94 23.967
R9517 casc_p.n25 casc_p.t128 23.967
R9518 casc_p.n24 casc_p.t314 23.967
R9519 casc_p.n23 casc_p.t242 23.967
R9520 casc_p.n22 casc_p.t125 23.967
R9521 casc_p.n21 casc_p.t198 23.967
R9522 casc_p.n20 casc_p.t382 23.967
R9523 casc_p.n19 casc_p.t287 23.967
R9524 casc_p.n18 casc_p.t154 23.967
R9525 casc_p.n17 casc_p.t80 23.967
R9526 casc_p.n16 casc_p.t285 23.967
R9527 casc_p.n15 casc_p.t223 23.967
R9528 casc_p.n14 casc_p.t78 23.967
R9529 casc_p.n13 casc_p.t318 23.967
R9530 casc_p.n12 casc_p.t221 23.967
R9531 casc_p.n11 casc_p.t127 23.967
R9532 casc_p.n10 casc_p.t313 23.967
R9533 casc_p.n9 casc_p.t384 23.967
R9534 casc_p.n8 casc_p.t240 23.967
R9535 casc_p.n7 casc_p.t155 23.967
R9536 casc_p.n6 casc_p.t381 23.967
R9537 casc_p.n5 casc_p.t286 23.967
R9538 casc_p.n4 casc_p.t152 23.967
R9539 casc_p.n3 casc_p.t79 23.967
R9540 casc_p.n48 casc_p.t119 23.967
R9541 casc_p.n47 casc_p.t215 23.967
R9542 casc_p.n46 casc_p.t308 23.967
R9543 casc_p.n45 casc_p.t73 23.967
R9544 casc_p.n44 casc_p.t217 23.967
R9545 casc_p.n43 casc_p.t275 23.967
R9546 casc_p.n42 casc_p.t99 23.967
R9547 casc_p.n41 casc_p.t193 23.967
R9548 casc_p.n40 casc_p.t277 23.967
R9549 casc_p.n39 casc_p.t378 23.967
R9550 casc_p.n382 casc_p.t253 23.967
R9551 casc_p.n381 casc_p.t392 23.967
R9552 casc_p.n380 casc_p.t237 23.967
R9553 casc_p.n379 casc_p.t368 23.967
R9554 casc_p.n378 casc_p.t76 23.967
R9555 casc_p.n377 casc_p.t209 23.967
R9556 casc_p.n376 casc_p.t239 23.967
R9557 casc_p.n375 casc_p.t371 23.967
R9558 casc_p.n374 casc_p.t219 23.967
R9559 casc_p.n373 casc_p.t351 23.967
R9560 casc_p.n34 casc_p.t67 14.202
R9561 casc_p.n31 casc_p.t1 14.202
R9562 casc_p.n286 casc_p.t42 13.873
R9563 casc_p.n286 casc_p.t41 13.871
R9564 casc_p.n329 casc_p.t38 13.858
R9565 casc_p.n329 casc_p.t39 13.858
R9566 casc_p.n283 casc_p.t11 13.858
R9567 casc_p.n283 casc_p.t12 13.858
R9568 casc_p.n237 casc_p.t47 13.858
R9569 casc_p.n237 casc_p.t48 13.858
R9570 casc_p.n191 casc_p.t23 13.858
R9571 casc_p.n191 casc_p.t24 13.858
R9572 casc_p.n145 casc_p.t53 13.858
R9573 casc_p.n145 casc_p.t54 13.858
R9574 casc_p.n87 casc_p.t29 13.858
R9575 casc_p.n87 casc_p.t30 13.858
R9576 casc_p.n93 casc_p.t59 13.858
R9577 casc_p.n93 casc_p.t60 13.858
R9578 casc_p.n99 casc_p.t26 13.858
R9579 casc_p.n99 casc_p.t27 13.858
R9580 casc_p.n360 casc_p.t35 13.858
R9581 casc_p.n360 casc_p.t36 13.858
R9582 casc_p.n366 casc_p.t5 13.858
R9583 casc_p.n366 casc_p.t6 13.858
R9584 casc_p.n369 casc_p.t63 13.853
R9585 casc_p.n332 casc_p.t9 13.853
R9586 casc_p.n240 casc_p.t15 13.853
R9587 casc_p.n194 casc_p.t51 13.853
R9588 casc_p.n148 casc_p.t21 13.853
R9589 casc_p.n90 casc_p.t18 13.853
R9590 casc_p.n96 casc_p.t45 13.853
R9591 casc_p.n102 casc_p.t57 13.853
R9592 casc_p.n363 casc_p.t33 13.853
R9593 casc_p.n332 casc_p.t8 13.852
R9594 casc_p.n240 casc_p.t14 13.852
R9595 casc_p.n194 casc_p.t50 13.852
R9596 casc_p.n148 casc_p.t20 13.852
R9597 casc_p.n90 casc_p.t17 13.852
R9598 casc_p.n96 casc_p.t44 13.852
R9599 casc_p.n102 casc_p.t56 13.852
R9600 casc_p.n363 casc_p.t32 13.852
R9601 casc_p.n369 casc_p.t62 13.852
R9602 casc_p.n33 casc_p.t3 13.849
R9603 casc_p.n32 casc_p.t65 13.849
R9604 casc_p.n0 casc_p.t66 12.05
R9605 casc_p.n0 casc_p.t2 12.05
R9606 casc_p.n30 casc_p.t64 12.05
R9607 casc_p.n30 casc_p.t0 12.05
R9608 casc_p.n37 casc_p.n35 9.3
R9609 casc_p.n37 casc_p.n36 9.3
R9610 casc_p.n38 casc_p.t68 8.529
R9611 casc_p.n38 casc_p.t69 8.525
R9612 casc_p.n392 casc_p.n38 5.493
R9613 casc_p.n391 casc_p.n390 2.199
R9614 casc_p.n390 casc_p.n389 2.199
R9615 casc_p.n389 casc_p.n388 2.199
R9616 casc_p.n388 casc_p.n387 2.199
R9617 casc_p.n387 casc_p.n386 2.199
R9618 casc_p.n386 casc_p.n385 2.199
R9619 casc_p.n385 casc_p.n384 2.199
R9620 casc_p.n33 casc_p.n32 1.175
R9621 casc_p.n393 casc_p.n392 1.074
R9622 casc_p.n300 casc_p.n299 1.002
R9623 casc_p.n302 casc_p.n301 1.002
R9624 casc_p.n304 casc_p.n303 1.002
R9625 casc_p.n306 casc_p.n305 1.002
R9626 casc_p.n308 casc_p.n307 1.002
R9627 casc_p.n310 casc_p.n309 1.002
R9628 casc_p.n312 casc_p.n311 1.002
R9629 casc_p.n314 casc_p.n313 1.002
R9630 casc_p.n316 casc_p.n315 1.002
R9631 casc_p.n318 casc_p.n317 1.002
R9632 casc_p.n320 casc_p.n319 1.002
R9633 casc_p.n322 casc_p.n321 1.002
R9634 casc_p.n324 casc_p.n323 1.002
R9635 casc_p.n326 casc_p.n325 1.002
R9636 casc_p.n297 casc_p.n296 1.002
R9637 casc_p.n295 casc_p.n294 1.002
R9638 casc_p.n293 casc_p.n292 1.002
R9639 casc_p.n291 casc_p.n290 1.002
R9640 casc_p.n289 casc_p.n288 1.002
R9641 casc_p.n254 casc_p.n253 1.002
R9642 casc_p.n256 casc_p.n255 1.002
R9643 casc_p.n258 casc_p.n257 1.002
R9644 casc_p.n260 casc_p.n259 1.002
R9645 casc_p.n262 casc_p.n261 1.002
R9646 casc_p.n264 casc_p.n263 1.002
R9647 casc_p.n266 casc_p.n265 1.002
R9648 casc_p.n268 casc_p.n267 1.002
R9649 casc_p.n270 casc_p.n269 1.002
R9650 casc_p.n272 casc_p.n271 1.002
R9651 casc_p.n274 casc_p.n273 1.002
R9652 casc_p.n276 casc_p.n275 1.002
R9653 casc_p.n278 casc_p.n277 1.002
R9654 casc_p.n280 casc_p.n279 1.002
R9655 casc_p.n251 casc_p.n250 1.002
R9656 casc_p.n249 casc_p.n248 1.002
R9657 casc_p.n247 casc_p.n246 1.002
R9658 casc_p.n245 casc_p.n244 1.002
R9659 casc_p.n243 casc_p.n242 1.002
R9660 casc_p.n208 casc_p.n207 1.002
R9661 casc_p.n210 casc_p.n209 1.002
R9662 casc_p.n212 casc_p.n211 1.002
R9663 casc_p.n214 casc_p.n213 1.002
R9664 casc_p.n216 casc_p.n215 1.002
R9665 casc_p.n218 casc_p.n217 1.002
R9666 casc_p.n220 casc_p.n219 1.002
R9667 casc_p.n222 casc_p.n221 1.002
R9668 casc_p.n224 casc_p.n223 1.002
R9669 casc_p.n226 casc_p.n225 1.002
R9670 casc_p.n228 casc_p.n227 1.002
R9671 casc_p.n230 casc_p.n229 1.002
R9672 casc_p.n232 casc_p.n231 1.002
R9673 casc_p.n234 casc_p.n233 1.002
R9674 casc_p.n205 casc_p.n204 1.002
R9675 casc_p.n203 casc_p.n202 1.002
R9676 casc_p.n201 casc_p.n200 1.002
R9677 casc_p.n199 casc_p.n198 1.002
R9678 casc_p.n197 casc_p.n196 1.002
R9679 casc_p.n162 casc_p.n161 1.002
R9680 casc_p.n164 casc_p.n163 1.002
R9681 casc_p.n166 casc_p.n165 1.002
R9682 casc_p.n168 casc_p.n167 1.002
R9683 casc_p.n170 casc_p.n169 1.002
R9684 casc_p.n172 casc_p.n171 1.002
R9685 casc_p.n174 casc_p.n173 1.002
R9686 casc_p.n176 casc_p.n175 1.002
R9687 casc_p.n178 casc_p.n177 1.002
R9688 casc_p.n180 casc_p.n179 1.002
R9689 casc_p.n182 casc_p.n181 1.002
R9690 casc_p.n184 casc_p.n183 1.002
R9691 casc_p.n186 casc_p.n185 1.002
R9692 casc_p.n188 casc_p.n187 1.002
R9693 casc_p.n159 casc_p.n158 1.002
R9694 casc_p.n157 casc_p.n156 1.002
R9695 casc_p.n155 casc_p.n154 1.002
R9696 casc_p.n153 casc_p.n152 1.002
R9697 casc_p.n151 casc_p.n150 1.002
R9698 casc_p.n116 casc_p.n115 1.002
R9699 casc_p.n118 casc_p.n117 1.002
R9700 casc_p.n120 casc_p.n119 1.002
R9701 casc_p.n122 casc_p.n121 1.002
R9702 casc_p.n124 casc_p.n123 1.002
R9703 casc_p.n126 casc_p.n125 1.002
R9704 casc_p.n128 casc_p.n127 1.002
R9705 casc_p.n130 casc_p.n129 1.002
R9706 casc_p.n132 casc_p.n131 1.002
R9707 casc_p.n134 casc_p.n133 1.002
R9708 casc_p.n136 casc_p.n135 1.002
R9709 casc_p.n138 casc_p.n137 1.002
R9710 casc_p.n140 casc_p.n139 1.002
R9711 casc_p.n142 casc_p.n141 1.002
R9712 casc_p.n113 casc_p.n112 1.002
R9713 casc_p.n111 casc_p.n110 1.002
R9714 casc_p.n109 casc_p.n108 1.002
R9715 casc_p.n107 casc_p.n106 1.002
R9716 casc_p.n105 casc_p.n104 1.002
R9717 casc_p.n62 casc_p.n61 1.002
R9718 casc_p.n64 casc_p.n63 1.002
R9719 casc_p.n66 casc_p.n65 1.002
R9720 casc_p.n68 casc_p.n67 1.002
R9721 casc_p.n70 casc_p.n69 1.002
R9722 casc_p.n72 casc_p.n71 1.002
R9723 casc_p.n74 casc_p.n73 1.002
R9724 casc_p.n76 casc_p.n75 1.002
R9725 casc_p.n78 casc_p.n77 1.002
R9726 casc_p.n80 casc_p.n79 1.002
R9727 casc_p.n82 casc_p.n81 1.002
R9728 casc_p.n84 casc_p.n83 1.002
R9729 casc_p.n59 casc_p.n58 1.002
R9730 casc_p.n57 casc_p.n56 1.002
R9731 casc_p.n55 casc_p.n54 1.002
R9732 casc_p.n53 casc_p.n52 1.002
R9733 casc_p.n51 casc_p.n50 1.002
R9734 casc_p.n4 casc_p.n3 1.002
R9735 casc_p.n6 casc_p.n5 1.002
R9736 casc_p.n8 casc_p.n7 1.002
R9737 casc_p.n10 casc_p.n9 1.002
R9738 casc_p.n12 casc_p.n11 1.002
R9739 casc_p.n14 casc_p.n13 1.002
R9740 casc_p.n16 casc_p.n15 1.002
R9741 casc_p.n18 casc_p.n17 1.002
R9742 casc_p.n20 casc_p.n19 1.002
R9743 casc_p.n22 casc_p.n21 1.002
R9744 casc_p.n24 casc_p.n23 1.002
R9745 casc_p.n48 casc_p.n47 1.002
R9746 casc_p.n46 casc_p.n45 1.002
R9747 casc_p.n44 casc_p.n43 1.002
R9748 casc_p.n42 casc_p.n41 1.002
R9749 casc_p.n40 casc_p.n39 1.002
R9750 casc_p.n382 casc_p.n381 1.002
R9751 casc_p.n380 casc_p.n379 1.002
R9752 casc_p.n378 casc_p.n377 1.002
R9753 casc_p.n376 casc_p.n375 1.002
R9754 casc_p.n374 casc_p.n373 1.002
R9755 casc_p.n335 casc_p.n334 1.002
R9756 casc_p.n337 casc_p.n336 1.002
R9757 casc_p.n339 casc_p.n338 1.002
R9758 casc_p.n341 casc_p.n340 1.002
R9759 casc_p.n343 casc_p.n342 1.002
R9760 casc_p.n345 casc_p.n344 1.002
R9761 casc_p.n347 casc_p.n346 1.002
R9762 casc_p.n349 casc_p.n348 1.002
R9763 casc_p.n351 casc_p.n350 1.002
R9764 casc_p.n353 casc_p.n352 1.002
R9765 casc_p.n355 casc_p.n354 1.002
R9766 casc_p.n357 casc_p.n356 1.002
R9767 casc_p.n392 casc_p.n391 0.84
R9768 casc_p.n392 casc_p.n0 0.779
R9769 casc_p.n0 casc_p.n29 0.752
R9770 casc_p.n2 casc_p.n394 0.75
R9771 casc_p.n1 casc_p.n27 0.75
R9772 casc_p.n328 casc_p.n327 0.728
R9773 casc_p.n282 casc_p.n281 0.728
R9774 casc_p.n236 casc_p.n235 0.728
R9775 casc_p.n190 casc_p.n189 0.728
R9776 casc_p.n144 casc_p.n143 0.728
R9777 casc_p.n86 casc_p.n85 0.728
R9778 casc_p.n26 casc_p.n25 0.728
R9779 casc_p.n359 casc_p.n358 0.728
R9780 casc_p.n371 casc_p.n370 0.728
R9781 casc_p.n301 casc_p.n300 0.66
R9782 casc_p.n303 casc_p.n302 0.66
R9783 casc_p.n305 casc_p.n304 0.66
R9784 casc_p.n307 casc_p.n306 0.66
R9785 casc_p.n309 casc_p.n308 0.66
R9786 casc_p.n311 casc_p.n310 0.66
R9787 casc_p.n313 casc_p.n312 0.66
R9788 casc_p.n315 casc_p.n314 0.66
R9789 casc_p.n317 casc_p.n316 0.66
R9790 casc_p.n319 casc_p.n318 0.66
R9791 casc_p.n321 casc_p.n320 0.66
R9792 casc_p.n323 casc_p.n322 0.66
R9793 casc_p.n325 casc_p.n324 0.66
R9794 casc_p.n327 casc_p.n326 0.66
R9795 casc_p.n296 casc_p.n295 0.66
R9796 casc_p.n294 casc_p.n293 0.66
R9797 casc_p.n292 casc_p.n291 0.66
R9798 casc_p.n290 casc_p.n289 0.66
R9799 casc_p.n255 casc_p.n254 0.66
R9800 casc_p.n257 casc_p.n256 0.66
R9801 casc_p.n259 casc_p.n258 0.66
R9802 casc_p.n261 casc_p.n260 0.66
R9803 casc_p.n263 casc_p.n262 0.66
R9804 casc_p.n265 casc_p.n264 0.66
R9805 casc_p.n267 casc_p.n266 0.66
R9806 casc_p.n269 casc_p.n268 0.66
R9807 casc_p.n271 casc_p.n270 0.66
R9808 casc_p.n273 casc_p.n272 0.66
R9809 casc_p.n275 casc_p.n274 0.66
R9810 casc_p.n277 casc_p.n276 0.66
R9811 casc_p.n279 casc_p.n278 0.66
R9812 casc_p.n281 casc_p.n280 0.66
R9813 casc_p.n250 casc_p.n249 0.66
R9814 casc_p.n248 casc_p.n247 0.66
R9815 casc_p.n246 casc_p.n245 0.66
R9816 casc_p.n244 casc_p.n243 0.66
R9817 casc_p.n209 casc_p.n208 0.66
R9818 casc_p.n211 casc_p.n210 0.66
R9819 casc_p.n213 casc_p.n212 0.66
R9820 casc_p.n215 casc_p.n214 0.66
R9821 casc_p.n217 casc_p.n216 0.66
R9822 casc_p.n219 casc_p.n218 0.66
R9823 casc_p.n221 casc_p.n220 0.66
R9824 casc_p.n223 casc_p.n222 0.66
R9825 casc_p.n225 casc_p.n224 0.66
R9826 casc_p.n227 casc_p.n226 0.66
R9827 casc_p.n229 casc_p.n228 0.66
R9828 casc_p.n231 casc_p.n230 0.66
R9829 casc_p.n233 casc_p.n232 0.66
R9830 casc_p.n235 casc_p.n234 0.66
R9831 casc_p.n204 casc_p.n203 0.66
R9832 casc_p.n202 casc_p.n201 0.66
R9833 casc_p.n200 casc_p.n199 0.66
R9834 casc_p.n198 casc_p.n197 0.66
R9835 casc_p.n163 casc_p.n162 0.66
R9836 casc_p.n165 casc_p.n164 0.66
R9837 casc_p.n167 casc_p.n166 0.66
R9838 casc_p.n169 casc_p.n168 0.66
R9839 casc_p.n171 casc_p.n170 0.66
R9840 casc_p.n173 casc_p.n172 0.66
R9841 casc_p.n175 casc_p.n174 0.66
R9842 casc_p.n177 casc_p.n176 0.66
R9843 casc_p.n179 casc_p.n178 0.66
R9844 casc_p.n181 casc_p.n180 0.66
R9845 casc_p.n183 casc_p.n182 0.66
R9846 casc_p.n185 casc_p.n184 0.66
R9847 casc_p.n187 casc_p.n186 0.66
R9848 casc_p.n189 casc_p.n188 0.66
R9849 casc_p.n158 casc_p.n157 0.66
R9850 casc_p.n156 casc_p.n155 0.66
R9851 casc_p.n154 casc_p.n153 0.66
R9852 casc_p.n152 casc_p.n151 0.66
R9853 casc_p.n117 casc_p.n116 0.66
R9854 casc_p.n119 casc_p.n118 0.66
R9855 casc_p.n121 casc_p.n120 0.66
R9856 casc_p.n123 casc_p.n122 0.66
R9857 casc_p.n125 casc_p.n124 0.66
R9858 casc_p.n127 casc_p.n126 0.66
R9859 casc_p.n129 casc_p.n128 0.66
R9860 casc_p.n131 casc_p.n130 0.66
R9861 casc_p.n133 casc_p.n132 0.66
R9862 casc_p.n135 casc_p.n134 0.66
R9863 casc_p.n137 casc_p.n136 0.66
R9864 casc_p.n139 casc_p.n138 0.66
R9865 casc_p.n141 casc_p.n140 0.66
R9866 casc_p.n143 casc_p.n142 0.66
R9867 casc_p.n112 casc_p.n111 0.66
R9868 casc_p.n110 casc_p.n109 0.66
R9869 casc_p.n108 casc_p.n107 0.66
R9870 casc_p.n106 casc_p.n105 0.66
R9871 casc_p.n63 casc_p.n62 0.66
R9872 casc_p.n65 casc_p.n64 0.66
R9873 casc_p.n67 casc_p.n66 0.66
R9874 casc_p.n69 casc_p.n68 0.66
R9875 casc_p.n71 casc_p.n70 0.66
R9876 casc_p.n73 casc_p.n72 0.66
R9877 casc_p.n75 casc_p.n74 0.66
R9878 casc_p.n77 casc_p.n76 0.66
R9879 casc_p.n79 casc_p.n78 0.66
R9880 casc_p.n81 casc_p.n80 0.66
R9881 casc_p.n83 casc_p.n82 0.66
R9882 casc_p.n85 casc_p.n84 0.66
R9883 casc_p.n58 casc_p.n57 0.66
R9884 casc_p.n56 casc_p.n55 0.66
R9885 casc_p.n54 casc_p.n53 0.66
R9886 casc_p.n52 casc_p.n51 0.66
R9887 casc_p.n5 casc_p.n4 0.66
R9888 casc_p.n7 casc_p.n6 0.66
R9889 casc_p.n9 casc_p.n8 0.66
R9890 casc_p.n11 casc_p.n10 0.66
R9891 casc_p.n13 casc_p.n12 0.66
R9892 casc_p.n15 casc_p.n14 0.66
R9893 casc_p.n17 casc_p.n16 0.66
R9894 casc_p.n19 casc_p.n18 0.66
R9895 casc_p.n21 casc_p.n20 0.66
R9896 casc_p.n23 casc_p.n22 0.66
R9897 casc_p.n25 casc_p.n24 0.66
R9898 casc_p.n47 casc_p.n46 0.66
R9899 casc_p.n45 casc_p.n44 0.66
R9900 casc_p.n43 casc_p.n42 0.66
R9901 casc_p.n41 casc_p.n40 0.66
R9902 casc_p.n381 casc_p.n380 0.66
R9903 casc_p.n379 casc_p.n378 0.66
R9904 casc_p.n377 casc_p.n376 0.66
R9905 casc_p.n375 casc_p.n374 0.66
R9906 casc_p.n336 casc_p.n335 0.66
R9907 casc_p.n338 casc_p.n337 0.66
R9908 casc_p.n340 casc_p.n339 0.66
R9909 casc_p.n342 casc_p.n341 0.66
R9910 casc_p.n344 casc_p.n343 0.66
R9911 casc_p.n346 casc_p.n345 0.66
R9912 casc_p.n348 casc_p.n347 0.66
R9913 casc_p.n350 casc_p.n349 0.66
R9914 casc_p.n352 casc_p.n351 0.66
R9915 casc_p.n354 casc_p.n353 0.66
R9916 casc_p.n356 casc_p.n355 0.66
R9917 casc_p.n358 casc_p.n357 0.66
R9918 casc_p.n372 casc_p.n371 0.66
R9919 casc_p.n298 casc_p.n297 0.655
R9920 casc_p.n252 casc_p.n251 0.655
R9921 casc_p.n206 casc_p.n205 0.655
R9922 casc_p.n160 casc_p.n159 0.655
R9923 casc_p.n114 casc_p.n113 0.655
R9924 casc_p.n60 casc_p.n59 0.655
R9925 casc_p.n49 casc_p.n48 0.655
R9926 casc_p.n383 casc_p.n382 0.655
R9927 casc_p.n384 casc_p.n372 0.599
R9928 casc_p.n92 casc_p.n91 0.454
R9929 casc_p.n98 casc_p.n97 0.454
R9930 casc_p.n365 casc_p.n364 0.454
R9931 casc_p casc_p.n26 0.438
R9932 casc_p.n385 casc_p.n298 0.369
R9933 casc_p.n386 casc_p.n252 0.369
R9934 casc_p.n387 casc_p.n206 0.369
R9935 casc_p.n388 casc_p.n160 0.369
R9936 casc_p.n389 casc_p.n114 0.369
R9937 casc_p.n390 casc_p.n60 0.369
R9938 casc_p.n391 casc_p.n49 0.369
R9939 casc_p.n384 casc_p.n383 0.369
R9940 casc_p.n32 casc_p.n31 0.353
R9941 casc_p.n34 casc_p.n33 0.353
R9942 casc_p.n385 casc_p.n333 0.325
R9943 casc_p.n386 casc_p.n287 0.325
R9944 casc_p.n387 casc_p.n241 0.325
R9945 casc_p.n388 casc_p.n195 0.325
R9946 casc_p.n389 casc_p.n149 0.325
R9947 casc_p.n390 casc_p.n103 0.325
R9948 casc_p.n286 casc_p.n285 0.292
R9949 casc_p.n31 casc_p.n30 0.29
R9950 casc_p.n330 casc_p.n329 0.282
R9951 casc_p.n284 casc_p.n283 0.282
R9952 casc_p.n238 casc_p.n237 0.282
R9953 casc_p.n192 casc_p.n191 0.282
R9954 casc_p.n146 casc_p.n145 0.282
R9955 casc_p.n88 casc_p.n87 0.282
R9956 casc_p.n94 casc_p.n93 0.282
R9957 casc_p.n100 casc_p.n99 0.282
R9958 casc_p.n361 casc_p.n360 0.282
R9959 casc_p.n367 casc_p.n366 0.282
R9960 casc_p.n0 casc_p.n37 0.281
R9961 casc_p.n333 casc_p.n332 0.278
R9962 casc_p.n241 casc_p.n240 0.278
R9963 casc_p.n195 casc_p.n194 0.278
R9964 casc_p.n149 casc_p.n148 0.278
R9965 casc_p.n91 casc_p.n90 0.278
R9966 casc_p.n97 casc_p.n96 0.278
R9967 casc_p.n103 casc_p.n102 0.278
R9968 casc_p.n364 casc_p.n363 0.278
R9969 casc_p.n370 casc_p.n369 0.278
R9970 casc_p.n332 casc_p.n331 0.271
R9971 casc_p.n240 casc_p.n239 0.271
R9972 casc_p.n194 casc_p.n193 0.271
R9973 casc_p.n148 casc_p.n147 0.271
R9974 casc_p.n90 casc_p.n89 0.271
R9975 casc_p.n96 casc_p.n95 0.271
R9976 casc_p.n102 casc_p.n101 0.271
R9977 casc_p.n363 casc_p.n362 0.271
R9978 casc_p.n369 casc_p.n368 0.271
R9979 casc_p.n329 casc_p.n328 0.267
R9980 casc_p.n283 casc_p.n282 0.267
R9981 casc_p.n237 casc_p.n236 0.267
R9982 casc_p.n191 casc_p.n190 0.267
R9983 casc_p.n145 casc_p.n144 0.267
R9984 casc_p.n87 casc_p.n86 0.267
R9985 casc_p.n93 casc_p.n92 0.267
R9986 casc_p.n99 casc_p.n98 0.267
R9987 casc_p.n360 casc_p.n359 0.267
R9988 casc_p.n366 casc_p.n365 0.267
R9989 casc_p.n287 casc_p.n286 0.257
R9990 casc_p casc_p.n395 0.155
R9991 casc_p.n331 casc_p.n330 0.112
R9992 casc_p.n285 casc_p.n284 0.112
R9993 casc_p.n239 casc_p.n238 0.112
R9994 casc_p.n193 casc_p.n192 0.112
R9995 casc_p.n147 casc_p.n146 0.112
R9996 casc_p.n89 casc_p.n88 0.112
R9997 casc_p.n95 casc_p.n94 0.112
R9998 casc_p.n101 casc_p.n100 0.112
R9999 casc_p.n362 casc_p.n361 0.112
R10000 casc_p.n368 casc_p.n367 0.112
R10001 casc_p.n2 casc_p.n393 0.046
R10002 casc_p.n393 casc_p.n1 0.045
R10003 casc_p.n395 casc_p.n2 0.019
R10004 casc_p.n1 casc_p.n28 0.019
R10005 casc_p.n37 casc_p.n34 0.015
R10006 a_2458_5328.n5 a_2458_5328.t68 13.849
R10007 a_2458_5328.n5 a_2458_5328.t102 13.849
R10008 a_2458_5328.n4 a_2458_5328.t30 13.849
R10009 a_2458_5328.n4 a_2458_5328.t177 13.849
R10010 a_2458_5328.n7 a_2458_5328.t57 13.849
R10011 a_2458_5328.n7 a_2458_5328.t117 13.849
R10012 a_2458_5328.n6 a_2458_5328.t53 13.849
R10013 a_2458_5328.n6 a_2458_5328.t124 13.849
R10014 a_2458_5328.n9 a_2458_5328.t80 13.849
R10015 a_2458_5328.n9 a_2458_5328.t132 13.849
R10016 a_2458_5328.n8 a_2458_5328.t86 13.849
R10017 a_2458_5328.n8 a_2458_5328.t166 13.849
R10018 a_2458_5328.n11 a_2458_5328.t24 13.849
R10019 a_2458_5328.n11 a_2458_5328.t112 13.849
R10020 a_2458_5328.n10 a_2458_5328.t54 13.849
R10021 a_2458_5328.n10 a_2458_5328.t122 13.849
R10022 a_2458_5328.n13 a_2458_5328.t73 13.849
R10023 a_2458_5328.n13 a_2458_5328.t127 13.849
R10024 a_2458_5328.n12 a_2458_5328.t89 13.849
R10025 a_2458_5328.n12 a_2458_5328.t138 13.849
R10026 a_2458_5328.n15 a_2458_5328.t37 13.849
R10027 a_2458_5328.n15 a_2458_5328.t147 13.849
R10028 a_2458_5328.n14 a_2458_5328.t23 13.849
R10029 a_2458_5328.n14 a_2458_5328.t113 13.849
R10030 a_2458_5328.n17 a_2458_5328.t38 13.849
R10031 a_2458_5328.n17 a_2458_5328.t106 13.849
R10032 a_2458_5328.n16 a_2458_5328.t36 13.849
R10033 a_2458_5328.n16 a_2458_5328.t128 13.849
R10034 a_2458_5328.n19 a_2458_5328.t58 13.849
R10035 a_2458_5328.n19 a_2458_5328.t100 13.849
R10036 a_2458_5328.n18 a_2458_5328.t67 13.849
R10037 a_2458_5328.n18 a_2458_5328.t108 13.849
R10038 a_2458_5328.n28 a_2458_5328.t76 13.849
R10039 a_2458_5328.n28 a_2458_5328.t136 13.849
R10040 a_2458_5328.n27 a_2458_5328.t26 13.849
R10041 a_2458_5328.n27 a_2458_5328.t111 13.849
R10042 a_2458_5328.n30 a_2458_5328.t72 13.849
R10043 a_2458_5328.n30 a_2458_5328.t130 13.849
R10044 a_2458_5328.n29 a_2458_5328.t87 13.849
R10045 a_2458_5328.n29 a_2458_5328.t165 13.849
R10046 a_2458_5328.n32 a_2458_5328.t35 13.849
R10047 a_2458_5328.n32 a_2458_5328.t149 13.849
R10048 a_2458_5328.n31 a_2458_5328.t21 13.849
R10049 a_2458_5328.n31 a_2458_5328.t116 13.849
R10050 a_2458_5328.n34 a_2458_5328.t75 13.849
R10051 a_2458_5328.n34 a_2458_5328.t110 13.849
R10052 a_2458_5328.n33 a_2458_5328.t78 13.849
R10053 a_2458_5328.n33 a_2458_5328.t134 13.849
R10054 a_2458_5328.n39 a_2458_5328.t92 13.849
R10055 a_2458_5328.n39 a_2458_5328.t143 13.849
R10056 a_2458_5328.n38 a_2458_5328.t3 13.849
R10057 a_2458_5328.n38 a_2458_5328.t163 13.849
R10058 a_2458_5328.n41 a_2458_5328.t183 13.849
R10059 a_2458_5328.n41 a_2458_5328.t148 13.849
R10060 a_2458_5328.n40 a_2458_5328.t196 13.849
R10061 a_2458_5328.n40 a_2458_5328.t115 13.849
R10062 a_2458_5328.n43 a_2458_5328.t193 13.849
R10063 a_2458_5328.n43 a_2458_5328.t107 13.849
R10064 a_2458_5328.n42 a_2458_5328.t180 13.849
R10065 a_2458_5328.n42 a_2458_5328.t129 13.849
R10066 a_2458_5328.n45 a_2458_5328.t2 13.849
R10067 a_2458_5328.n45 a_2458_5328.t145 13.849
R10068 a_2458_5328.n44 a_2458_5328.t182 13.849
R10069 a_2458_5328.n44 a_2458_5328.t150 13.849
R10070 a_2458_5328.n49 a_2458_5328.t46 13.849
R10071 a_2458_5328.n49 a_2458_5328.t103 13.849
R10072 a_2458_5328.n48 a_2458_5328.t181 13.849
R10073 a_2458_5328.n48 a_2458_5328.t109 13.849
R10074 a_2458_5328.n47 a_2458_5328.t4 13.849
R10075 a_2458_5328.n47 a_2458_5328.t161 13.849
R10076 a_2458_5328.n46 a_2458_5328.t45 13.849
R10077 a_2458_5328.n46 a_2458_5328.t104 13.849
R10078 a_2458_5328.n53 a_2458_5328.t95 13.849
R10079 a_2458_5328.n53 a_2458_5328.t141 13.849
R10080 a_2458_5328.n52 a_2458_5328.t184 13.849
R10081 a_2458_5328.n52 a_2458_5328.t146 13.849
R10082 a_2458_5328.n51 a_2458_5328.t49 13.849
R10083 a_2458_5328.n51 a_2458_5328.t172 13.849
R10084 a_2458_5328.n50 a_2458_5328.t94 13.849
R10085 a_2458_5328.n50 a_2458_5328.t142 13.849
R10086 a_2458_5328.n57 a_2458_5328.t48 13.849
R10087 a_2458_5328.n57 a_2458_5328.t162 13.849
R10088 a_2458_5328.n56 a_2458_5328.t93 13.849
R10089 a_2458_5328.n56 a_2458_5328.t105 13.849
R10090 a_2458_5328.n55 a_2458_5328.t50 13.849
R10091 a_2458_5328.n55 a_2458_5328.t123 13.849
R10092 a_2458_5328.n54 a_2458_5328.t47 13.849
R10093 a_2458_5328.n54 a_2458_5328.t164 13.849
R10094 a_2458_5328.n61 a_2458_5328.t70 13.849
R10095 a_2458_5328.n61 a_2458_5328.t152 13.849
R10096 a_2458_5328.n60 a_2458_5328.t12 13.849
R10097 a_2458_5328.n60 a_2458_5328.t98 13.849
R10098 a_2458_5328.n59 a_2458_5328.t71 13.849
R10099 a_2458_5328.n59 a_2458_5328.t119 13.849
R10100 a_2458_5328.n58 a_2458_5328.t5 13.849
R10101 a_2458_5328.n58 a_2458_5328.t153 13.849
R10102 a_2458_5328.n103 a_2458_5328.t60 13.849
R10103 a_2458_5328.n103 a_2458_5328.t160 13.849
R10104 a_2458_5328.n102 a_2458_5328.t90 13.849
R10105 a_2458_5328.n102 a_2458_5328.t137 13.849
R10106 a_2458_5328.n105 a_2458_5328.t28 13.849
R10107 a_2458_5328.n105 a_2458_5328.t140 13.849
R10108 a_2458_5328.n104 a_2458_5328.t69 13.849
R10109 a_2458_5328.n104 a_2458_5328.t101 13.849
R10110 a_2458_5328.n107 a_2458_5328.t61 13.849
R10111 a_2458_5328.n107 a_2458_5328.t159 13.849
R10112 a_2458_5328.n106 a_2458_5328.t29 13.849
R10113 a_2458_5328.n106 a_2458_5328.t139 13.849
R10114 a_2458_5328.n109 a_2458_5328.t32 13.849
R10115 a_2458_5328.n109 a_2458_5328.t175 13.849
R10116 a_2458_5328.n108 a_2458_5328.t59 13.849
R10117 a_2458_5328.n108 a_2458_5328.t99 13.849
R10118 a_2458_5328.n111 a_2458_5328.t64 13.849
R10119 a_2458_5328.n111 a_2458_5328.t156 13.849
R10120 a_2458_5328.n110 a_2458_5328.t33 13.849
R10121 a_2458_5328.n110 a_2458_5328.t174 13.849
R10122 a_2458_5328.n113 a_2458_5328.t83 13.849
R10123 a_2458_5328.n113 a_2458_5328.t170 13.849
R10124 a_2458_5328.n112 a_2458_5328.t65 13.849
R10125 a_2458_5328.n112 a_2458_5328.t155 13.849
R10126 a_2458_5328.n115 a_2458_5328.t88 13.849
R10127 a_2458_5328.n115 a_2458_5328.t121 13.849
R10128 a_2458_5328.n114 a_2458_5328.t55 13.849
R10129 a_2458_5328.n114 a_2458_5328.t169 13.849
R10130 a_2458_5328.n117 a_2458_5328.t22 13.849
R10131 a_2458_5328.n117 a_2458_5328.t114 13.849
R10132 a_2458_5328.n116 a_2458_5328.t77 13.849
R10133 a_2458_5328.n116 a_2458_5328.t135 13.849
R10134 a_2458_5328.n80 a_2458_5328.t81 13.849
R10135 a_2458_5328.n80 a_2458_5328.t131 13.849
R10136 a_2458_5328.n79 a_2458_5328.t39 13.849
R10137 a_2458_5328.n79 a_2458_5328.t144 13.849
R10138 a_2458_5328.n82 a_2458_5328.t62 13.849
R10139 a_2458_5328.n82 a_2458_5328.t158 13.849
R10140 a_2458_5328.n81 a_2458_5328.t31 13.849
R10141 a_2458_5328.n81 a_2458_5328.t176 13.849
R10142 a_2458_5328.n84 a_2458_5328.t82 13.849
R10143 a_2458_5328.n84 a_2458_5328.t171 13.849
R10144 a_2458_5328.n83 a_2458_5328.t63 13.849
R10145 a_2458_5328.n83 a_2458_5328.t157 13.849
R10146 a_2458_5328.n86 a_2458_5328.t66 13.849
R10147 a_2458_5328.n86 a_2458_5328.t154 13.849
R10148 a_2458_5328.n85 a_2458_5328.t34 13.849
R10149 a_2458_5328.n85 a_2458_5328.t173 13.849
R10150 a_2458_5328.n88 a_2458_5328.t84 13.849
R10151 a_2458_5328.n88 a_2458_5328.t168 13.849
R10152 a_2458_5328.n87 a_2458_5328.t52 13.849
R10153 a_2458_5328.n87 a_2458_5328.t125 13.849
R10154 a_2458_5328.n90 a_2458_5328.t56 13.849
R10155 a_2458_5328.n90 a_2458_5328.t120 13.849
R10156 a_2458_5328.n89 a_2458_5328.t85 13.849
R10157 a_2458_5328.n89 a_2458_5328.t167 13.849
R10158 a_2458_5328.n92 a_2458_5328.t25 13.849
R10159 a_2458_5328.n92 a_2458_5328.t133 13.849
R10160 a_2458_5328.n91 a_2458_5328.t79 13.849
R10161 a_2458_5328.n91 a_2458_5328.t118 13.849
R10162 a_2458_5328.n94 a_2458_5328.t74 13.849
R10163 a_2458_5328.n94 a_2458_5328.t126 13.849
R10164 a_2458_5328.n93 a_2458_5328.t27 13.849
R10165 a_2458_5328.n93 a_2458_5328.t151 13.849
R10166 a_2458_5328.n72 a_2458_5328.t198 10.905
R10167 a_2458_5328.n75 a_2458_5328.t44 8.979
R10168 a_2458_5328.n69 a_2458_5328.t96 8.265
R10169 a_2458_5328.n69 a_2458_5328.t91 8.265
R10170 a_2458_5328.n70 a_2458_5328.t199 8.265
R10171 a_2458_5328.n70 a_2458_5328.t97 8.265
R10172 a_2458_5328.n71 a_2458_5328.t186 8.265
R10173 a_2458_5328.n71 a_2458_5328.t43 8.265
R10174 a_2458_5328.n129 a_2458_5328.n128 7.826
R10175 a_2458_5328.n169 a_2458_5328.n168 7.774
R10176 a_2458_5328.n152 a_2458_5328.n151 7.773
R10177 a_2458_5328.n138 a_2458_5328.n137 7.773
R10178 a_2458_5328.n76 a_2458_5328.n75 7.361
R10179 a_2458_5328.n150 a_2458_5328.n149 4.514
R10180 a_2458_5328.n145 a_2458_5328.n144 4.514
R10181 a_2458_5328.n136 a_2458_5328.n135 4.514
R10182 a_2458_5328.n155 a_2458_5328.n3 4.513
R10183 a_2458_5328.n78 a_2458_5328.n26 3.568
R10184 a_2458_5328.n77 a_2458_5328.n37 3.568
R10185 a_2458_5328.n76 a_2458_5328.n68 3.568
R10186 a_2458_5328.n125 a_2458_5328.n124 3.568
R10187 a_2458_5328.n126 a_2458_5328.n101 3.568
R10188 a_2458_5328.n20 a_2458_5328.n19 2.739
R10189 a_2458_5328.n35 a_2458_5328.n34 2.739
R10190 a_2458_5328.n62 a_2458_5328.n61 2.739
R10191 a_2458_5328.n118 a_2458_5328.n117 2.739
R10192 a_2458_5328.n95 a_2458_5328.n94 2.739
R10193 a_2458_5328.n131 a_2458_5328.n127 2.648
R10194 a_2458_5328.n21 a_2458_5328.n20 2.199
R10195 a_2458_5328.n22 a_2458_5328.n21 2.199
R10196 a_2458_5328.n23 a_2458_5328.n22 2.199
R10197 a_2458_5328.n24 a_2458_5328.n23 2.199
R10198 a_2458_5328.n25 a_2458_5328.n24 2.199
R10199 a_2458_5328.n26 a_2458_5328.n25 2.199
R10200 a_2458_5328.n36 a_2458_5328.n35 2.199
R10201 a_2458_5328.n37 a_2458_5328.n36 2.199
R10202 a_2458_5328.n63 a_2458_5328.n62 2.199
R10203 a_2458_5328.n64 a_2458_5328.n63 2.199
R10204 a_2458_5328.n65 a_2458_5328.n64 2.199
R10205 a_2458_5328.n66 a_2458_5328.n65 2.199
R10206 a_2458_5328.n67 a_2458_5328.n66 2.199
R10207 a_2458_5328.n68 a_2458_5328.n67 2.199
R10208 a_2458_5328.n119 a_2458_5328.n118 2.199
R10209 a_2458_5328.n120 a_2458_5328.n119 2.199
R10210 a_2458_5328.n121 a_2458_5328.n120 2.199
R10211 a_2458_5328.n122 a_2458_5328.n121 2.199
R10212 a_2458_5328.n123 a_2458_5328.n122 2.199
R10213 a_2458_5328.n124 a_2458_5328.n123 2.199
R10214 a_2458_5328.n96 a_2458_5328.n95 2.199
R10215 a_2458_5328.n97 a_2458_5328.n96 2.199
R10216 a_2458_5328.n98 a_2458_5328.n97 2.199
R10217 a_2458_5328.n99 a_2458_5328.n98 2.199
R10218 a_2458_5328.n100 a_2458_5328.n99 2.199
R10219 a_2458_5328.n101 a_2458_5328.n100 2.199
R10220 a_2458_5328.n159 a_2458_5328.t179 2.153
R10221 a_2458_5328.n128 a_2458_5328.t17 2.153
R10222 a_2458_5328.n129 a_2458_5328.t6 2.153
R10223 a_2458_5328.n130 a_2458_5328.t16 2.153
R10224 a_2458_5328.t0 a_2458_5328.n169 2.142
R10225 a_2458_5328.n156 a_2458_5328.t18 2.142
R10226 a_2458_5328.n3 a_2458_5328.t15 2.142
R10227 a_2458_5328.n2 a_2458_5328.t192 2.142
R10228 a_2458_5328.n1 a_2458_5328.t40 2.142
R10229 a_2458_5328.n0 a_2458_5328.t189 2.142
R10230 a_2458_5328.n167 a_2458_5328.t190 2.142
R10231 a_2458_5328.n168 a_2458_5328.t185 2.142
R10232 a_2458_5328.n157 a_2458_5328.t8 2.142
R10233 a_2458_5328.n151 a_2458_5328.t13 2.142
R10234 a_2458_5328.n152 a_2458_5328.t178 2.142
R10235 a_2458_5328.n153 a_2458_5328.t10 2.142
R10236 a_2458_5328.n146 a_2458_5328.t51 2.142
R10237 a_2458_5328.n147 a_2458_5328.t1 2.142
R10238 a_2458_5328.n148 a_2458_5328.t41 2.142
R10239 a_2458_5328.n149 a_2458_5328.t11 2.142
R10240 a_2458_5328.n141 a_2458_5328.t20 2.142
R10241 a_2458_5328.n142 a_2458_5328.t188 2.142
R10242 a_2458_5328.n143 a_2458_5328.t7 2.142
R10243 a_2458_5328.n144 a_2458_5328.t194 2.142
R10244 a_2458_5328.n158 a_2458_5328.t9 2.142
R10245 a_2458_5328.n137 a_2458_5328.t42 2.142
R10246 a_2458_5328.n138 a_2458_5328.t195 2.142
R10247 a_2458_5328.n139 a_2458_5328.t197 2.142
R10248 a_2458_5328.n132 a_2458_5328.t14 2.142
R10249 a_2458_5328.n133 a_2458_5328.t191 2.142
R10250 a_2458_5328.n134 a_2458_5328.t187 2.142
R10251 a_2458_5328.n135 a_2458_5328.t19 2.142
R10252 a_2458_5328.n74 a_2458_5328.n69 1.827
R10253 a_2458_5328.n73 a_2458_5328.n70 1.827
R10254 a_2458_5328.n72 a_2458_5328.n71 1.827
R10255 a_2458_5328.n167 a_2458_5328.n166 1.808
R10256 a_2458_5328.n160 a_2458_5328.n159 1.646
R10257 a_2458_5328.n165 a_2458_5328.n157 1.62
R10258 a_2458_5328.n162 a_2458_5328.n158 1.62
R10259 a_2458_5328.n156 a_2458_5328.n155 1.496
R10260 a_2458_5328.n130 a_2458_5328.n129 1.414
R10261 a_2458_5328.n3 a_2458_5328.n2 1.361
R10262 a_2458_5328.n2 a_2458_5328.n1 1.361
R10263 a_2458_5328.n1 a_2458_5328.n0 1.361
R10264 a_2458_5328.n168 a_2458_5328.n167 1.361
R10265 a_2458_5328.n153 a_2458_5328.n152 1.361
R10266 a_2458_5328.n147 a_2458_5328.n146 1.361
R10267 a_2458_5328.n148 a_2458_5328.n147 1.361
R10268 a_2458_5328.n149 a_2458_5328.n148 1.361
R10269 a_2458_5328.n142 a_2458_5328.n141 1.361
R10270 a_2458_5328.n143 a_2458_5328.n142 1.361
R10271 a_2458_5328.n144 a_2458_5328.n143 1.361
R10272 a_2458_5328.n139 a_2458_5328.n138 1.361
R10273 a_2458_5328.n133 a_2458_5328.n132 1.361
R10274 a_2458_5328.n134 a_2458_5328.n133 1.361
R10275 a_2458_5328.n135 a_2458_5328.n134 1.361
R10276 a_2458_5328.n169 a_2458_5328.n156 1.361
R10277 a_2458_5328.n131 a_2458_5328.n130 1.335
R10278 a_2458_5328.n154 a_2458_5328.n153 1.308
R10279 a_2458_5328.n140 a_2458_5328.n139 1.308
R10280 a_2458_5328.n75 a_2458_5328.n74 0.908
R10281 a_2458_5328.n48 a_2458_5328.n47 0.868
R10282 a_2458_5328.n52 a_2458_5328.n51 0.868
R10283 a_2458_5328.n56 a_2458_5328.n55 0.868
R10284 a_2458_5328.n60 a_2458_5328.n59 0.868
R10285 a_2458_5328.n73 a_2458_5328.n72 0.812
R10286 a_2458_5328.n74 a_2458_5328.n73 0.796
R10287 a_2458_5328.n77 a_2458_5328.n76 0.752
R10288 a_2458_5328.n78 a_2458_5328.n77 0.752
R10289 a_2458_5328.n126 a_2458_5328.n125 0.752
R10290 a_2458_5328.n26 a_2458_5328.n5 0.54
R10291 a_2458_5328.n25 a_2458_5328.n7 0.54
R10292 a_2458_5328.n24 a_2458_5328.n9 0.54
R10293 a_2458_5328.n23 a_2458_5328.n11 0.54
R10294 a_2458_5328.n22 a_2458_5328.n13 0.54
R10295 a_2458_5328.n21 a_2458_5328.n15 0.54
R10296 a_2458_5328.n20 a_2458_5328.n17 0.54
R10297 a_2458_5328.n37 a_2458_5328.n28 0.54
R10298 a_2458_5328.n36 a_2458_5328.n30 0.54
R10299 a_2458_5328.n35 a_2458_5328.n32 0.54
R10300 a_2458_5328.n68 a_2458_5328.n39 0.54
R10301 a_2458_5328.n67 a_2458_5328.n41 0.54
R10302 a_2458_5328.n66 a_2458_5328.n43 0.54
R10303 a_2458_5328.n65 a_2458_5328.n45 0.54
R10304 a_2458_5328.n64 a_2458_5328.n49 0.54
R10305 a_2458_5328.n63 a_2458_5328.n53 0.54
R10306 a_2458_5328.n62 a_2458_5328.n57 0.54
R10307 a_2458_5328.n124 a_2458_5328.n103 0.54
R10308 a_2458_5328.n123 a_2458_5328.n105 0.54
R10309 a_2458_5328.n122 a_2458_5328.n107 0.54
R10310 a_2458_5328.n121 a_2458_5328.n109 0.54
R10311 a_2458_5328.n120 a_2458_5328.n111 0.54
R10312 a_2458_5328.n119 a_2458_5328.n113 0.54
R10313 a_2458_5328.n118 a_2458_5328.n115 0.54
R10314 a_2458_5328.n101 a_2458_5328.n80 0.54
R10315 a_2458_5328.n100 a_2458_5328.n82 0.54
R10316 a_2458_5328.n99 a_2458_5328.n84 0.54
R10317 a_2458_5328.n98 a_2458_5328.n86 0.54
R10318 a_2458_5328.n97 a_2458_5328.n88 0.54
R10319 a_2458_5328.n96 a_2458_5328.n90 0.54
R10320 a_2458_5328.n95 a_2458_5328.n92 0.54
R10321 a_2458_5328.n5 a_2458_5328.n4 0.464
R10322 a_2458_5328.n7 a_2458_5328.n6 0.464
R10323 a_2458_5328.n9 a_2458_5328.n8 0.464
R10324 a_2458_5328.n11 a_2458_5328.n10 0.464
R10325 a_2458_5328.n13 a_2458_5328.n12 0.464
R10326 a_2458_5328.n15 a_2458_5328.n14 0.464
R10327 a_2458_5328.n17 a_2458_5328.n16 0.464
R10328 a_2458_5328.n19 a_2458_5328.n18 0.464
R10329 a_2458_5328.n28 a_2458_5328.n27 0.464
R10330 a_2458_5328.n30 a_2458_5328.n29 0.464
R10331 a_2458_5328.n32 a_2458_5328.n31 0.464
R10332 a_2458_5328.n34 a_2458_5328.n33 0.464
R10333 a_2458_5328.n39 a_2458_5328.n38 0.464
R10334 a_2458_5328.n41 a_2458_5328.n40 0.464
R10335 a_2458_5328.n43 a_2458_5328.n42 0.464
R10336 a_2458_5328.n45 a_2458_5328.n44 0.464
R10337 a_2458_5328.n47 a_2458_5328.n46 0.464
R10338 a_2458_5328.n49 a_2458_5328.n48 0.464
R10339 a_2458_5328.n51 a_2458_5328.n50 0.464
R10340 a_2458_5328.n53 a_2458_5328.n52 0.464
R10341 a_2458_5328.n55 a_2458_5328.n54 0.464
R10342 a_2458_5328.n57 a_2458_5328.n56 0.464
R10343 a_2458_5328.n59 a_2458_5328.n58 0.464
R10344 a_2458_5328.n61 a_2458_5328.n60 0.464
R10345 a_2458_5328.n103 a_2458_5328.n102 0.464
R10346 a_2458_5328.n105 a_2458_5328.n104 0.464
R10347 a_2458_5328.n107 a_2458_5328.n106 0.464
R10348 a_2458_5328.n109 a_2458_5328.n108 0.464
R10349 a_2458_5328.n111 a_2458_5328.n110 0.464
R10350 a_2458_5328.n113 a_2458_5328.n112 0.464
R10351 a_2458_5328.n115 a_2458_5328.n114 0.464
R10352 a_2458_5328.n117 a_2458_5328.n116 0.464
R10353 a_2458_5328.n80 a_2458_5328.n79 0.464
R10354 a_2458_5328.n82 a_2458_5328.n81 0.464
R10355 a_2458_5328.n84 a_2458_5328.n83 0.464
R10356 a_2458_5328.n86 a_2458_5328.n85 0.464
R10357 a_2458_5328.n88 a_2458_5328.n87 0.464
R10358 a_2458_5328.n90 a_2458_5328.n89 0.464
R10359 a_2458_5328.n92 a_2458_5328.n91 0.464
R10360 a_2458_5328.n94 a_2458_5328.n93 0.464
R10361 a_2458_5328.n127 a_2458_5328.n126 0.411
R10362 a_2458_5328.n127 a_2458_5328.n78 0.34
R10363 a_2458_5328.n166 a_2458_5328.n165 0.188
R10364 a_2458_5328.n165 a_2458_5328.n164 0.188
R10365 a_2458_5328.n164 a_2458_5328.n163 0.188
R10366 a_2458_5328.n163 a_2458_5328.n162 0.188
R10367 a_2458_5328.n162 a_2458_5328.n161 0.188
R10368 a_2458_5328.n161 a_2458_5328.n160 0.188
R10369 a_2458_5328.n155 a_2458_5328.n154 0.188
R10370 a_2458_5328.n154 a_2458_5328.n150 0.188
R10371 a_2458_5328.n150 a_2458_5328.n145 0.188
R10372 a_2458_5328.n145 a_2458_5328.n140 0.188
R10373 a_2458_5328.n140 a_2458_5328.n136 0.188
R10374 a_2458_5328.n136 a_2458_5328.n131 0.188
R10375 Vom.n49 Vom.t124 57.533
R10376 Vom.n104 Vom.t49 14.623
R10377 Vom.n105 Vom.t28 14.623
R10378 Vom.n106 Vom.t64 14.623
R10379 Vom.n107 Vom.t26 14.623
R10380 Vom.n108 Vom.t60 14.623
R10381 Vom.n109 Vom.t15 14.623
R10382 Vom.n110 Vom.t55 14.623
R10383 Vom.n111 Vom.t47 14.623
R10384 Vom.n139 Vom.t50 14.598
R10385 Vom.n138 Vom.t8 14.598
R10386 Vom.n137 Vom.t52 14.598
R10387 Vom.n136 Vom.t10 14.598
R10388 Vom.n135 Vom.t63 14.598
R10389 Vom.n82 Vom.t69 14.598
R10390 Vom.n83 Vom.t62 14.598
R10391 Vom.n84 Vom.t17 14.598
R10392 Vom.n85 Vom.t59 14.598
R10393 Vom.n86 Vom.t11 14.598
R10394 Vom.n87 Vom.t53 14.598
R10395 Vom.n88 Vom.t4 14.598
R10396 Vom.n89 Vom.t76 14.598
R10397 Vom.n72 Vom.t77 14.598
R10398 Vom.n73 Vom.t51 14.598
R10399 Vom.n74 Vom.t2 14.598
R10400 Vom.n75 Vom.t46 14.598
R10401 Vom.n12 Vom.t23 14.598
R10402 Vom.n13 Vom.t1 14.598
R10403 Vom.n14 Vom.t41 14.598
R10404 Vom.n15 Vom.t75 14.598
R10405 Vom.n16 Vom.t31 14.598
R10406 Vom.n19 Vom.t67 14.598
R10407 Vom.n22 Vom.t24 14.598
R10408 Vom.n25 Vom.t13 14.598
R10409 Vom.n140 Vom.t40 14.598
R10410 Vom.n141 Vom.t35 14.598
R10411 Vom.n143 Vom.t79 14.598
R10412 Vom.n143 Vom.t72 13.849
R10413 Vom.n139 Vom.t39 13.849
R10414 Vom.n138 Vom.t78 13.849
R10415 Vom.n137 Vom.t44 13.849
R10416 Vom.n136 Vom.t3 13.849
R10417 Vom.n135 Vom.t29 13.849
R10418 Vom.n104 Vom.t20 13.849
R10419 Vom.n105 Vom.t65 13.849
R10420 Vom.n106 Vom.t19 13.849
R10421 Vom.n107 Vom.t61 13.849
R10422 Vom.n108 Vom.t16 13.849
R10423 Vom.n109 Vom.t56 13.849
R10424 Vom.n110 Vom.t7 13.849
R10425 Vom.n111 Vom.t0 13.849
R10426 Vom.n82 Vom.t43 13.849
R10427 Vom.n83 Vom.t18 13.849
R10428 Vom.n84 Vom.t57 13.849
R10429 Vom.n85 Vom.t14 13.849
R10430 Vom.n86 Vom.t54 13.849
R10431 Vom.n87 Vom.t6 13.849
R10432 Vom.n88 Vom.t45 13.849
R10433 Vom.n89 Vom.t38 13.849
R10434 Vom.n72 Vom.t48 13.849
R10435 Vom.n73 Vom.t42 13.849
R10436 Vom.n74 Vom.t74 13.849
R10437 Vom.n75 Vom.t37 13.849
R10438 Vom.n12 Vom.t68 13.849
R10439 Vom.n13 Vom.t73 13.849
R10440 Vom.n14 Vom.t34 13.849
R10441 Vom.n15 Vom.t70 13.849
R10442 Vom.n18 Vom.t30 13.849
R10443 Vom.n17 Vom.t36 13.849
R10444 Vom.n16 Vom.t21 13.849
R10445 Vom.n21 Vom.t66 13.849
R10446 Vom.n20 Vom.t71 13.849
R10447 Vom.n19 Vom.t58 13.849
R10448 Vom.n24 Vom.t22 13.849
R10449 Vom.n23 Vom.t32 13.849
R10450 Vom.n22 Vom.t9 13.849
R10451 Vom.n27 Vom.t12 13.849
R10452 Vom.n26 Vom.t25 13.849
R10453 Vom.n25 Vom.t5 13.849
R10454 Vom.n140 Vom.t33 13.849
R10455 Vom.n141 Vom.t27 13.849
R10456 Vom.n0 Vom.t132 12.05
R10457 Vom.n0 Vom.t143 12.05
R10458 Vom.n1 Vom.t133 12.05
R10459 Vom.n1 Vom.t125 12.05
R10460 Vom.n2 Vom.t128 12.05
R10461 Vom.n2 Vom.t120 12.05
R10462 Vom.n3 Vom.t129 12.05
R10463 Vom.n3 Vom.t141 12.05
R10464 Vom.n4 Vom.t123 12.05
R10465 Vom.n4 Vom.t137 12.05
R10466 Vom.n5 Vom.t139 12.05
R10467 Vom.n5 Vom.t127 12.05
R10468 Vom.n6 Vom.t138 12.05
R10469 Vom.n6 Vom.t121 12.05
R10470 Vom.n7 Vom.t122 12.05
R10471 Vom.n7 Vom.t135 12.05
R10472 Vom.n8 Vom.t136 12.05
R10473 Vom.n8 Vom.t131 12.05
R10474 Vom.n9 Vom.t140 12.05
R10475 Vom.n9 Vom.t134 12.05
R10476 Vom.n10 Vom.t126 12.05
R10477 Vom.n10 Vom.t142 12.05
R10478 Vom.n11 Vom.t144 12.05
R10479 Vom.n11 Vom.t130 12.05
R10480 Vom.n119 Vom.t90 8.857
R10481 Vom.n120 Vom.t118 8.857
R10482 Vom.n121 Vom.t91 8.857
R10483 Vom.n122 Vom.t112 8.857
R10484 Vom.n97 Vom.t110 8.857
R10485 Vom.n98 Vom.t81 8.857
R10486 Vom.n99 Vom.t111 8.857
R10487 Vom.n100 Vom.t101 8.857
R10488 Vom.n79 Vom.t116 8.857
R10489 Vom.n80 Vom.t87 8.857
R10490 Vom.n35 Vom.t105 8.857
R10491 Vom.n128 Vom.t107 8.857
R10492 Vom.n129 Vom.t80 8.857
R10493 Vom.n130 Vom.t108 8.857
R10494 Vom.n131 Vom.t85 8.857
R10495 Vom.n36 Vom.t109 8.8
R10496 Vom.n37 Vom.t86 8.8
R10497 Vom.n40 Vom.t117 8.8
R10498 Vom.n119 Vom.t96 8.266
R10499 Vom.n120 Vom.t119 8.266
R10500 Vom.n121 Vom.t98 8.266
R10501 Vom.n122 Vom.t102 8.266
R10502 Vom.n97 Vom.t82 8.266
R10503 Vom.n98 Vom.t113 8.266
R10504 Vom.n99 Vom.t83 8.266
R10505 Vom.n100 Vom.t89 8.266
R10506 Vom.n79 Vom.t84 8.266
R10507 Vom.n80 Vom.t115 8.266
R10508 Vom.n35 Vom.t92 8.266
R10509 Vom.n36 Vom.t104 8.266
R10510 Vom.n39 Vom.t93 8.266
R10511 Vom.n38 Vom.t106 8.266
R10512 Vom.n37 Vom.t114 8.266
R10513 Vom.n42 Vom.t100 8.266
R10514 Vom.n41 Vom.t95 8.266
R10515 Vom.n40 Vom.t97 8.266
R10516 Vom.n128 Vom.t99 8.266
R10517 Vom.n129 Vom.t94 8.266
R10518 Vom.n130 Vom.t103 8.266
R10519 Vom.n131 Vom.t88 8.266
R10520 Vom.n112 Vom.n111 2.632
R10521 Vom.n90 Vom.n89 2.609
R10522 Vom.n76 Vom.n75 2.609
R10523 Vom.n28 Vom.n27 2.609
R10524 Vom.n142 Vom.n141 2.609
R10525 Vom.n123 Vom.n122 2.597
R10526 Vom.n101 Vom.n100 2.597
R10527 Vom.n81 Vom.n80 2.597
R10528 Vom.n132 Vom.n131 2.597
R10529 Vom.n43 Vom.n42 2.559
R10530 Vom.n126 Vom.n118 2.506
R10531 Vom.n127 Vom.n96 2.506
R10532 Vom.n151 Vom.n78 2.506
R10533 Vom.n63 Vom.n34 2.506
R10534 Vom.n150 Vom.n149 2.506
R10535 Vom.n44 Vom.n43 2.22
R10536 Vom.n124 Vom.n123 2.219
R10537 Vom.n125 Vom.n124 2.219
R10538 Vom.n102 Vom.n101 2.219
R10539 Vom.n103 Vom.n102 2.219
R10540 Vom.n45 Vom.n44 2.219
R10541 Vom.n133 Vom.n132 2.219
R10542 Vom.n134 Vom.n133 2.219
R10543 Vom.n113 Vom.n112 2.199
R10544 Vom.n114 Vom.n113 2.199
R10545 Vom.n115 Vom.n114 2.199
R10546 Vom.n116 Vom.n115 2.199
R10547 Vom.n117 Vom.n116 2.199
R10548 Vom.n118 Vom.n117 2.199
R10549 Vom.n91 Vom.n90 2.199
R10550 Vom.n92 Vom.n91 2.199
R10551 Vom.n93 Vom.n92 2.199
R10552 Vom.n94 Vom.n93 2.199
R10553 Vom.n95 Vom.n94 2.199
R10554 Vom.n96 Vom.n95 2.199
R10555 Vom.n77 Vom.n76 2.199
R10556 Vom.n78 Vom.n77 2.199
R10557 Vom.n29 Vom.n28 2.199
R10558 Vom.n30 Vom.n29 2.199
R10559 Vom.n31 Vom.n30 2.199
R10560 Vom.n32 Vom.n31 2.199
R10561 Vom.n33 Vom.n32 2.199
R10562 Vom.n34 Vom.n33 2.199
R10563 Vom.n149 Vom.n148 2.199
R10564 Vom.n148 Vom.n147 2.199
R10565 Vom.n147 Vom.n146 2.199
R10566 Vom.n146 Vom.n145 2.199
R10567 Vom.n145 Vom.n144 2.199
R10568 Vom.n144 Vom.n142 2.199
R10569 Vom.n62 Vom.n6 2.042
R10570 Vom.n71 Vom.n10 2.042
R10571 Vom.n49 Vom.n0 2.042
R10572 Vom.n126 Vom.n125 1.528
R10573 Vom.n127 Vom.n103 1.528
R10574 Vom.n151 Vom.n81 1.528
R10575 Vom.n63 Vom.n45 1.528
R10576 Vom.n150 Vom.n134 1.528
R10577 Vom.n17 Vom.n16 1.159
R10578 Vom.n20 Vom.n19 1.159
R10579 Vom.n23 Vom.n22 1.159
R10580 Vom.n26 Vom.n25 1.159
R10581 Vom.n59 Vom.n9 1.151
R10582 Vom.n60 Vom.n8 1.151
R10583 Vom.n61 Vom.n7 1.151
R10584 Vom.n68 Vom.n3 1.151
R10585 Vom.n69 Vom.n4 1.151
R10586 Vom.n70 Vom.n5 1.151
R10587 Vom.n54 Vom.n1 1.151
R10588 Vom.n55 Vom.n2 1.151
R10589 Vom.n48 Vom.n11 1.151
R10590 Vom.n38 Vom.n37 0.859
R10591 Vom.n41 Vom.n40 0.859
R10592 Vom.n151 Vom.n150 0.752
R10593 Vom.n150 Vom.n127 0.752
R10594 Vom.n127 Vom.n126 0.752
R10595 Vom.n18 Vom.n17 0.749
R10596 Vom.n21 Vom.n20 0.749
R10597 Vom.n24 Vom.n23 0.749
R10598 Vom.n27 Vom.n26 0.749
R10599 Vom.n39 Vom.n38 0.534
R10600 Vom.n42 Vom.n41 0.534
R10601 Vom.n9 Vom.n58 0.455
R10602 Vom.n8 Vom.n59 0.455
R10603 Vom.n7 Vom.n60 0.455
R10604 Vom.n6 Vom.n61 0.455
R10605 Vom.n4 Vom.n68 0.455
R10606 Vom.n5 Vom.n69 0.455
R10607 Vom.n10 Vom.n70 0.455
R10608 Vom.n2 Vom.n54 0.455
R10609 Vom.n0 Vom.n48 0.455
R10610 Vom Vom.n71 0.437
R10611 Vom.n118 Vom.n104 0.433
R10612 Vom.n117 Vom.n105 0.433
R10613 Vom.n116 Vom.n106 0.433
R10614 Vom.n115 Vom.n107 0.433
R10615 Vom.n114 Vom.n108 0.433
R10616 Vom.n113 Vom.n109 0.433
R10617 Vom.n112 Vom.n110 0.433
R10618 Vom.n145 Vom.n139 0.41
R10619 Vom.n146 Vom.n138 0.41
R10620 Vom.n147 Vom.n137 0.41
R10621 Vom.n148 Vom.n136 0.41
R10622 Vom.n149 Vom.n135 0.41
R10623 Vom.n96 Vom.n82 0.41
R10624 Vom.n95 Vom.n83 0.41
R10625 Vom.n94 Vom.n84 0.41
R10626 Vom.n93 Vom.n85 0.41
R10627 Vom.n92 Vom.n86 0.41
R10628 Vom.n91 Vom.n87 0.41
R10629 Vom.n90 Vom.n88 0.41
R10630 Vom.n78 Vom.n72 0.41
R10631 Vom.n77 Vom.n73 0.41
R10632 Vom.n76 Vom.n74 0.41
R10633 Vom.n34 Vom.n12 0.41
R10634 Vom.n33 Vom.n13 0.41
R10635 Vom.n32 Vom.n14 0.41
R10636 Vom.n31 Vom.n15 0.41
R10637 Vom.n30 Vom.n18 0.41
R10638 Vom.n29 Vom.n21 0.41
R10639 Vom.n28 Vom.n24 0.41
R10640 Vom.n142 Vom.n140 0.41
R10641 Vom.n144 Vom.n143 0.41
R10642 Vom.n125 Vom.n119 0.378
R10643 Vom.n124 Vom.n120 0.378
R10644 Vom.n123 Vom.n121 0.378
R10645 Vom.n103 Vom.n97 0.378
R10646 Vom.n102 Vom.n98 0.378
R10647 Vom.n101 Vom.n99 0.378
R10648 Vom.n81 Vom.n79 0.378
R10649 Vom.n45 Vom.n35 0.378
R10650 Vom.n134 Vom.n128 0.378
R10651 Vom.n133 Vom.n129 0.378
R10652 Vom.n132 Vom.n130 0.378
R10653 Vom.n60 Vom.n55 0.376
R10654 Vom.n62 Vom.n49 0.376
R10655 Vom.n44 Vom.n36 0.338
R10656 Vom.n43 Vom.n39 0.338
R10657 Vom.n11 Vom.n47 0.246
R10658 Vom.n10 Vom.n64 0.246
R10659 Vom.n9 Vom.n57 0.246
R10660 Vom.n8 Vom.n56 0.246
R10661 Vom.n7 Vom.n51 0.246
R10662 Vom.n6 Vom.n50 0.246
R10663 Vom.n5 Vom.n65 0.246
R10664 Vom.n4 Vom.n66 0.246
R10665 Vom.n3 Vom.n67 0.246
R10666 Vom.n2 Vom.n52 0.246
R10667 Vom.n1 Vom.n53 0.246
R10668 Vom.n0 Vom.n46 0.246
R10669 Vom.n71 Vom.n63 0.211
R10670 Vom.n63 Vom.n62 0.164
R10671 Vom Vom.n151 0.102
R10672 a_12760_n20342.n19 a_12760_n20342.t4 17.971
R10673 a_12760_n20342.t0 a_12760_n20342.n19 14.431
R10674 a_12760_n20342.n20 a_12760_n20342.t1 14.13
R10675 a_12760_n20342.n19 a_12760_n20342.t3 13.849
R10676 a_12760_n20342.n20 a_12760_n20342.t2 13.849
R10677 a_12760_n20342.n78 a_12760_n20342.t107 12.05
R10678 a_12760_n20342.n78 a_12760_n20342.t92 12.05
R10679 a_12760_n20342.n77 a_12760_n20342.t42 12.05
R10680 a_12760_n20342.n77 a_12760_n20342.t32 12.05
R10681 a_12760_n20342.n79 a_12760_n20342.t24 12.05
R10682 a_12760_n20342.n79 a_12760_n20342.t11 12.05
R10683 a_12760_n20342.n82 a_12760_n20342.t83 12.05
R10684 a_12760_n20342.n82 a_12760_n20342.t69 12.05
R10685 a_12760_n20342.n49 a_12760_n20342.t28 12.05
R10686 a_12760_n20342.n49 a_12760_n20342.t86 12.05
R10687 a_12760_n20342.n50 a_12760_n20342.t94 12.05
R10688 a_12760_n20342.n50 a_12760_n20342.t29 12.05
R10689 a_12760_n20342.n52 a_12760_n20342.t103 12.05
R10690 a_12760_n20342.n52 a_12760_n20342.t38 12.05
R10691 a_12760_n20342.n54 a_12760_n20342.t48 12.05
R10692 a_12760_n20342.n54 a_12760_n20342.t110 12.05
R10693 a_12760_n20342.n58 a_12760_n20342.t85 12.05
R10694 a_12760_n20342.n58 a_12760_n20342.t71 12.05
R10695 a_12760_n20342.n57 a_12760_n20342.t17 12.05
R10696 a_12760_n20342.n57 a_12760_n20342.t6 12.05
R10697 a_12760_n20342.n56 a_12760_n20342.t7 12.05
R10698 a_12760_n20342.n56 a_12760_n20342.t124 12.05
R10699 a_12760_n20342.n55 a_12760_n20342.t65 12.05
R10700 a_12760_n20342.n55 a_12760_n20342.t54 12.05
R10701 a_12760_n20342.n26 a_12760_n20342.t125 12.05
R10702 a_12760_n20342.n26 a_12760_n20342.t111 12.05
R10703 a_12760_n20342.n23 a_12760_n20342.t62 12.05
R10704 a_12760_n20342.n23 a_12760_n20342.t47 12.05
R10705 a_12760_n20342.n24 a_12760_n20342.t121 12.05
R10706 a_12760_n20342.n24 a_12760_n20342.t101 12.05
R10707 a_12760_n20342.n47 a_12760_n20342.t21 12.05
R10708 a_12760_n20342.n47 a_12760_n20342.t105 12.05
R10709 a_12760_n20342.n46 a_12760_n20342.t77 12.05
R10710 a_12760_n20342.n46 a_12760_n20342.t15 12.05
R10711 a_12760_n20342.n43 a_12760_n20342.t23 12.05
R10712 a_12760_n20342.n43 a_12760_n20342.t79 12.05
R10713 a_12760_n20342.n21 a_12760_n20342.t90 12.05
R10714 a_12760_n20342.n21 a_12760_n20342.t78 12.05
R10715 a_12760_n20342.n75 a_12760_n20342.t35 12.05
R10716 a_12760_n20342.n75 a_12760_n20342.t25 12.05
R10717 a_12760_n20342.n76 a_12760_n20342.t102 12.05
R10718 a_12760_n20342.n76 a_12760_n20342.t89 12.05
R10719 a_12760_n20342.n51 a_12760_n20342.t118 12.05
R10720 a_12760_n20342.n51 a_12760_n20342.t100 12.05
R10721 a_12760_n20342.n73 a_12760_n20342.t53 12.05
R10722 a_12760_n20342.n73 a_12760_n20342.t113 12.05
R10723 a_12760_n20342.n70 a_12760_n20342.t40 12.05
R10724 a_12760_n20342.n70 a_12760_n20342.t97 12.05
R10725 a_12760_n20342.n68 a_12760_n20342.t96 12.05
R10726 a_12760_n20342.n68 a_12760_n20342.t33 12.05
R10727 a_12760_n20342.n42 a_12760_n20342.t30 12.05
R10728 a_12760_n20342.n42 a_12760_n20342.t88 12.05
R10729 a_12760_n20342.n35 a_12760_n20342.t91 12.05
R10730 a_12760_n20342.n35 a_12760_n20342.t27 12.05
R10731 a_12760_n20342.n36 a_12760_n20342.t109 12.05
R10732 a_12760_n20342.n36 a_12760_n20342.t93 12.05
R10733 a_12760_n20342.n40 a_12760_n20342.t95 12.05
R10734 a_12760_n20342.n40 a_12760_n20342.t41 12.05
R10735 a_12760_n20342.n33 a_12760_n20342.t52 12.05
R10736 a_12760_n20342.n33 a_12760_n20342.t37 12.05
R10737 a_12760_n20342.n34 a_12760_n20342.t116 12.05
R10738 a_12760_n20342.n34 a_12760_n20342.t98 12.05
R10739 a_12760_n20342.n67 a_12760_n20342.t59 12.05
R10740 a_12760_n20342.n67 a_12760_n20342.t43 12.05
R10741 a_12760_n20342.n69 a_12760_n20342.t128 12.05
R10742 a_12760_n20342.n69 a_12760_n20342.t114 12.05
R10743 a_12760_n20342.n63 a_12760_n20342.t64 12.05
R10744 a_12760_n20342.n63 a_12760_n20342.t49 12.05
R10745 a_12760_n20342.n59 a_12760_n20342.t58 12.05
R10746 a_12760_n20342.n59 a_12760_n20342.t119 12.05
R10747 a_12760_n20342.n30 a_12760_n20342.t115 12.05
R10748 a_12760_n20342.n30 a_12760_n20342.t46 12.05
R10749 a_12760_n20342.n27 a_12760_n20342.t51 12.05
R10750 a_12760_n20342.n27 a_12760_n20342.t112 12.05
R10751 a_12760_n20342.n28 a_12760_n20342.t108 12.05
R10752 a_12760_n20342.n28 a_12760_n20342.t39 12.05
R10753 a_12760_n20342.n29 a_12760_n20342.t56 12.05
R10754 a_12760_n20342.n29 a_12760_n20342.t13 12.05
R10755 a_12760_n20342.n60 a_12760_n20342.t127 12.05
R10756 a_12760_n20342.n60 a_12760_n20342.t61 12.05
R10757 a_12760_n20342.n61 a_12760_n20342.t8 12.05
R10758 a_12760_n20342.n61 a_12760_n20342.t67 12.05
R10759 a_12760_n20342.n65 a_12760_n20342.t75 12.05
R10760 a_12760_n20342.n65 a_12760_n20342.t12 12.05
R10761 a_12760_n20342.n62 a_12760_n20342.t122 12.05
R10762 a_12760_n20342.n62 a_12760_n20342.t104 12.05
R10763 a_12760_n20342.n32 a_12760_n20342.t50 12.05
R10764 a_12760_n20342.n32 a_12760_n20342.t36 12.05
R10765 a_12760_n20342.n31 a_12760_n20342.t117 12.05
R10766 a_12760_n20342.n31 a_12760_n20342.t99 12.05
R10767 a_12760_n20342.n37 a_12760_n20342.t44 12.05
R10768 a_12760_n20342.n37 a_12760_n20342.t34 12.05
R10769 a_12760_n20342.n39 a_12760_n20342.t14 12.05
R10770 a_12760_n20342.n39 a_12760_n20342.t80 12.05
R10771 a_12760_n20342.n64 a_12760_n20342.t68 12.05
R10772 a_12760_n20342.n64 a_12760_n20342.t63 12.05
R10773 a_12760_n20342.n66 a_12760_n20342.t16 12.05
R10774 a_12760_n20342.n66 a_12760_n20342.t5 12.05
R10775 a_12760_n20342.n71 a_12760_n20342.t9 12.05
R10776 a_12760_n20342.n71 a_12760_n20342.t126 12.05
R10777 a_12760_n20342.n72 a_12760_n20342.t76 12.05
R10778 a_12760_n20342.n72 a_12760_n20342.t66 12.05
R10779 a_12760_n20342.n44 a_12760_n20342.t87 12.05
R10780 a_12760_n20342.n44 a_12760_n20342.t73 12.05
R10781 a_12760_n20342.n45 a_12760_n20342.t74 12.05
R10782 a_12760_n20342.n45 a_12760_n20342.t20 12.05
R10783 a_12760_n20342.n22 a_12760_n20342.t31 12.05
R10784 a_12760_n20342.n22 a_12760_n20342.t19 12.05
R10785 a_12760_n20342.n38 a_12760_n20342.t26 12.05
R10786 a_12760_n20342.n38 a_12760_n20342.t81 12.05
R10787 a_12760_n20342.n41 a_12760_n20342.t120 12.05
R10788 a_12760_n20342.n41 a_12760_n20342.t72 12.05
R10789 a_12760_n20342.n74 a_12760_n20342.t123 12.05
R10790 a_12760_n20342.n74 a_12760_n20342.t57 12.05
R10791 a_12760_n20342.n53 a_12760_n20342.t60 12.05
R10792 a_12760_n20342.n53 a_12760_n20342.t45 12.05
R10793 a_12760_n20342.n81 a_12760_n20342.t84 12.05
R10794 a_12760_n20342.n81 a_12760_n20342.t70 12.05
R10795 a_12760_n20342.n80 a_12760_n20342.t22 12.05
R10796 a_12760_n20342.n80 a_12760_n20342.t10 12.05
R10797 a_12760_n20342.n48 a_12760_n20342.t82 12.05
R10798 a_12760_n20342.n48 a_12760_n20342.t18 12.05
R10799 a_12760_n20342.n25 a_12760_n20342.t106 12.05
R10800 a_12760_n20342.n25 a_12760_n20342.t55 12.05
R10801 a_12760_n20342.n19 a_12760_n20342.n89 9.462
R10802 a_12760_n20342.n78 a_12760_n20342.n87 9.3
R10803 a_12760_n20342.n78 a_12760_n20342.n88 9.3
R10804 a_12760_n20342.n77 a_12760_n20342.n84 9.3
R10805 a_12760_n20342.n77 a_12760_n20342.n85 9.3
R10806 a_12760_n20342.n79 a_12760_n20342.n91 9.3
R10807 a_12760_n20342.n79 a_12760_n20342.n92 9.3
R10808 a_12760_n20342.n82 a_12760_n20342.n190 9.3
R10809 a_12760_n20342.n82 a_12760_n20342.n191 9.3
R10810 a_12760_n20342.n49 a_12760_n20342.n193 9.3
R10811 a_12760_n20342.n49 a_12760_n20342.n194 9.3
R10812 a_12760_n20342.n50 a_12760_n20342.n196 9.3
R10813 a_12760_n20342.n50 a_12760_n20342.n197 9.3
R10814 a_12760_n20342.n52 a_12760_n20342.n202 9.3
R10815 a_12760_n20342.n52 a_12760_n20342.n203 9.3
R10816 a_12760_n20342.n54 a_12760_n20342.n209 9.3
R10817 a_12760_n20342.n54 a_12760_n20342.n210 9.3
R10818 a_12760_n20342.n58 a_12760_n20342.n222 9.3
R10819 a_12760_n20342.n58 a_12760_n20342.n223 9.3
R10820 a_12760_n20342.n57 a_12760_n20342.n219 9.3
R10821 a_12760_n20342.n57 a_12760_n20342.n220 9.3
R10822 a_12760_n20342.n56 a_12760_n20342.n216 9.3
R10823 a_12760_n20342.n56 a_12760_n20342.n217 9.3
R10824 a_12760_n20342.n55 a_12760_n20342.n213 9.3
R10825 a_12760_n20342.n55 a_12760_n20342.n214 9.3
R10826 a_12760_n20342.n26 a_12760_n20342.n117 9.3
R10827 a_12760_n20342.n26 a_12760_n20342.n118 9.3
R10828 a_12760_n20342.n23 a_12760_n20342.n106 9.3
R10829 a_12760_n20342.n23 a_12760_n20342.n107 9.3
R10830 a_12760_n20342.n24 a_12760_n20342.n109 9.3
R10831 a_12760_n20342.n24 a_12760_n20342.n110 9.3
R10832 a_12760_n20342.n47 a_12760_n20342.n183 9.3
R10833 a_12760_n20342.n47 a_12760_n20342.n184 9.3
R10834 a_12760_n20342.n46 a_12760_n20342.n180 9.3
R10835 a_12760_n20342.n46 a_12760_n20342.n181 9.3
R10836 a_12760_n20342.n43 a_12760_n20342.n170 9.3
R10837 a_12760_n20342.n43 a_12760_n20342.n171 9.3
R10838 a_12760_n20342.n21 a_12760_n20342.n100 9.3
R10839 a_12760_n20342.n21 a_12760_n20342.n101 9.3
R10840 a_12760_n20342.n75 a_12760_n20342.n286 9.3
R10841 a_12760_n20342.n75 a_12760_n20342.n287 9.3
R10842 a_12760_n20342.n76 a_12760_n20342.n289 9.3
R10843 a_12760_n20342.n76 a_12760_n20342.n290 9.3
R10844 a_12760_n20342.n51 a_12760_n20342.n199 9.3
R10845 a_12760_n20342.n51 a_12760_n20342.n200 9.3
R10846 a_12760_n20342.n73 a_12760_n20342.n278 9.3
R10847 a_12760_n20342.n73 a_12760_n20342.n279 9.3
R10848 a_12760_n20342.n70 a_12760_n20342.n267 9.3
R10849 a_12760_n20342.n70 a_12760_n20342.n268 9.3
R10850 a_12760_n20342.n68 a_12760_n20342.n261 9.3
R10851 a_12760_n20342.n68 a_12760_n20342.n262 9.3
R10852 a_12760_n20342.n42 a_12760_n20342.n167 9.3
R10853 a_12760_n20342.n42 a_12760_n20342.n168 9.3
R10854 a_12760_n20342.n35 a_12760_n20342.n146 9.3
R10855 a_12760_n20342.n35 a_12760_n20342.n147 9.3
R10856 a_12760_n20342.n36 a_12760_n20342.n149 9.3
R10857 a_12760_n20342.n36 a_12760_n20342.n150 9.3
R10858 a_12760_n20342.n40 a_12760_n20342.n161 9.3
R10859 a_12760_n20342.n40 a_12760_n20342.n162 9.3
R10860 a_12760_n20342.n33 a_12760_n20342.n140 9.3
R10861 a_12760_n20342.n33 a_12760_n20342.n141 9.3
R10862 a_12760_n20342.n34 a_12760_n20342.n143 9.3
R10863 a_12760_n20342.n34 a_12760_n20342.n144 9.3
R10864 a_12760_n20342.n67 a_12760_n20342.n258 9.3
R10865 a_12760_n20342.n67 a_12760_n20342.n259 9.3
R10866 a_12760_n20342.n69 a_12760_n20342.n264 9.3
R10867 a_12760_n20342.n69 a_12760_n20342.n265 9.3
R10868 a_12760_n20342.n63 a_12760_n20342.n242 9.3
R10869 a_12760_n20342.n63 a_12760_n20342.n243 9.3
R10870 a_12760_n20342.n59 a_12760_n20342.n228 9.3
R10871 a_12760_n20342.n59 a_12760_n20342.n229 9.3
R10872 a_12760_n20342.n30 a_12760_n20342.n131 9.3
R10873 a_12760_n20342.n30 a_12760_n20342.n132 9.3
R10874 a_12760_n20342.n27 a_12760_n20342.n120 9.3
R10875 a_12760_n20342.n27 a_12760_n20342.n121 9.3
R10876 a_12760_n20342.n28 a_12760_n20342.n123 9.3
R10877 a_12760_n20342.n28 a_12760_n20342.n124 9.3
R10878 a_12760_n20342.n29 a_12760_n20342.n126 9.3
R10879 a_12760_n20342.n29 a_12760_n20342.n127 9.3
R10880 a_12760_n20342.n60 a_12760_n20342.n231 9.3
R10881 a_12760_n20342.n60 a_12760_n20342.n232 9.3
R10882 a_12760_n20342.n61 a_12760_n20342.n234 9.3
R10883 a_12760_n20342.n61 a_12760_n20342.n235 9.3
R10884 a_12760_n20342.n65 a_12760_n20342.n248 9.3
R10885 a_12760_n20342.n65 a_12760_n20342.n249 9.3
R10886 a_12760_n20342.n62 a_12760_n20342.n239 9.3
R10887 a_12760_n20342.n62 a_12760_n20342.n240 9.3
R10888 a_12760_n20342.n32 a_12760_n20342.n137 9.3
R10889 a_12760_n20342.n32 a_12760_n20342.n138 9.3
R10890 a_12760_n20342.n31 a_12760_n20342.n134 9.3
R10891 a_12760_n20342.n31 a_12760_n20342.n135 9.3
R10892 a_12760_n20342.n37 a_12760_n20342.n152 9.3
R10893 a_12760_n20342.n37 a_12760_n20342.n153 9.3
R10894 a_12760_n20342.n39 a_12760_n20342.n158 9.3
R10895 a_12760_n20342.n39 a_12760_n20342.n159 9.3
R10896 a_12760_n20342.n64 a_12760_n20342.n245 9.3
R10897 a_12760_n20342.n64 a_12760_n20342.n246 9.3
R10898 a_12760_n20342.n66 a_12760_n20342.n252 9.3
R10899 a_12760_n20342.n66 a_12760_n20342.n253 9.3
R10900 a_12760_n20342.n71 a_12760_n20342.n270 9.3
R10901 a_12760_n20342.n71 a_12760_n20342.n271 9.3
R10902 a_12760_n20342.n72 a_12760_n20342.n273 9.3
R10903 a_12760_n20342.n72 a_12760_n20342.n274 9.3
R10904 a_12760_n20342.n44 a_12760_n20342.n173 9.3
R10905 a_12760_n20342.n44 a_12760_n20342.n174 9.3
R10906 a_12760_n20342.n45 a_12760_n20342.n176 9.3
R10907 a_12760_n20342.n45 a_12760_n20342.n177 9.3
R10908 a_12760_n20342.n22 a_12760_n20342.n103 9.3
R10909 a_12760_n20342.n22 a_12760_n20342.n104 9.3
R10910 a_12760_n20342.n38 a_12760_n20342.n155 9.3
R10911 a_12760_n20342.n38 a_12760_n20342.n156 9.3
R10912 a_12760_n20342.n41 a_12760_n20342.n164 9.3
R10913 a_12760_n20342.n41 a_12760_n20342.n165 9.3
R10914 a_12760_n20342.n74 a_12760_n20342.n281 9.3
R10915 a_12760_n20342.n74 a_12760_n20342.n282 9.3
R10916 a_12760_n20342.n53 a_12760_n20342.n205 9.3
R10917 a_12760_n20342.n53 a_12760_n20342.n206 9.3
R10918 a_12760_n20342.n81 a_12760_n20342.n97 9.3
R10919 a_12760_n20342.n81 a_12760_n20342.n98 9.3
R10920 a_12760_n20342.n80 a_12760_n20342.n94 9.3
R10921 a_12760_n20342.n80 a_12760_n20342.n95 9.3
R10922 a_12760_n20342.n48 a_12760_n20342.n187 9.3
R10923 a_12760_n20342.n48 a_12760_n20342.n188 9.3
R10924 a_12760_n20342.n25 a_12760_n20342.n112 9.3
R10925 a_12760_n20342.n25 a_12760_n20342.n113 9.3
R10926 a_12760_n20342.n89 a_12760_n20342.n78 1.423
R10927 a_12760_n20342.n15 a_12760_n20342.n14 1.251
R10928 a_12760_n20342.n28 a_12760_n20342.n128 1.228
R10929 a_12760_n20342.n27 a_12760_n20342.n129 1.228
R10930 a_12760_n20342.n9 a_12760_n20342.n30 1.228
R10931 a_12760_n20342.n14 a_12760_n20342.n59 1.228
R10932 a_12760_n20342.n6 a_12760_n20342.n65 1.228
R10933 a_12760_n20342.n236 a_12760_n20342.n61 1.228
R10934 a_12760_n20342.n237 a_12760_n20342.n60 1.228
R10935 a_12760_n20342.n9 a_12760_n20342.n32 1.228
R10936 a_12760_n20342.n15 a_12760_n20342.n62 1.228
R10937 a_12760_n20342.n256 a_12760_n20342.n63 1.228
R10938 a_12760_n20342.n6 a_12760_n20342.n66 1.228
R10939 a_12760_n20342.n255 a_12760_n20342.n64 1.228
R10940 a_12760_n20342.n276 a_12760_n20342.n72 1.228
R10941 a_12760_n20342.n1 a_12760_n20342.n71 1.228
R10942 a_12760_n20342.n0 a_12760_n20342.n69 1.228
R10943 a_12760_n20342.n15 a_12760_n20342.n67 1.228
R10944 a_12760_n20342.n10 a_12760_n20342.n34 1.228
R10945 a_12760_n20342.n44 a_12760_n20342.n178 1.228
R10946 a_12760_n20342.n38 a_12760_n20342.n13 1.228
R10947 a_12760_n20342.n35 a_12760_n20342.n4 1.228
R10948 a_12760_n20342.n10 a_12760_n20342.n42 1.228
R10949 a_12760_n20342.n16 a_12760_n20342.n68 1.228
R10950 a_12760_n20342.n0 a_12760_n20342.n70 1.228
R10951 a_12760_n20342.n1 a_12760_n20342.n73 1.228
R10952 a_12760_n20342.n284 a_12760_n20342.n74 1.228
R10953 a_12760_n20342.n7 a_12760_n20342.n53 1.228
R10954 a_12760_n20342.n2 a_12760_n20342.n51 1.228
R10955 a_12760_n20342.n291 a_12760_n20342.n76 1.228
R10956 a_12760_n20342.n16 a_12760_n20342.n75 1.228
R10957 a_12760_n20342.n11 a_12760_n20342.n21 1.228
R10958 a_12760_n20342.n11 a_12760_n20342.n48 1.228
R10959 a_12760_n20342.n43 a_12760_n20342.n5 1.228
R10960 a_12760_n20342.n46 a_12760_n20342.n185 1.228
R10961 a_12760_n20342.n24 a_12760_n20342.n114 1.228
R10962 a_12760_n20342.n23 a_12760_n20342.n115 1.228
R10963 a_12760_n20342.n8 a_12760_n20342.n26 1.228
R10964 a_12760_n20342.n14 a_12760_n20342.n55 1.228
R10965 a_12760_n20342.n226 a_12760_n20342.n56 1.228
R10966 a_12760_n20342.n225 a_12760_n20342.n57 1.228
R10967 a_12760_n20342.n224 a_12760_n20342.n58 1.228
R10968 a_12760_n20342.n7 a_12760_n20342.n54 1.228
R10969 a_12760_n20342.n2 a_12760_n20342.n52 1.228
R10970 a_12760_n20342.n211 a_12760_n20342.n50 1.228
R10971 a_12760_n20342.n17 a_12760_n20342.n49 1.228
R10972 a_12760_n20342.n18 a_12760_n20342.n80 1.212
R10973 a_12760_n20342.n18 a_12760_n20342.n82 1.212
R10974 a_12760_n20342.n89 a_12760_n20342.n77 1.183
R10975 a_12760_n20342.n52 a_12760_n20342.n7 1.18
R10976 a_12760_n20342.n64 a_12760_n20342.n6 1.18
R10977 a_12760_n20342.n5 a_12760_n20342.n46 1.18
R10978 a_12760_n20342.n50 a_12760_n20342.n2 1.18
R10979 a_12760_n20342.n70 a_12760_n20342.n1 1.18
R10980 a_12760_n20342.n68 a_12760_n20342.n0 1.18
R10981 a_12760_n20342.n19 a_12760_n20342.n20 1.177
R10982 a_12760_n20342.n76 a_12760_n20342.n288 1.037
R10983 a_12760_n20342.n69 a_12760_n20342.n263 1.037
R10984 a_12760_n20342.n67 a_12760_n20342.n257 1.037
R10985 a_12760_n20342.n61 a_12760_n20342.n233 1.037
R10986 a_12760_n20342.n58 a_12760_n20342.n221 1.037
R10987 a_12760_n20342.n54 a_12760_n20342.n208 1.037
R10988 a_12760_n20342.n51 a_12760_n20342.n198 1.037
R10989 a_12760_n20342.n48 a_12760_n20342.n186 1.037
R10990 a_12760_n20342.n42 a_12760_n20342.n166 1.037
R10991 a_12760_n20342.n34 a_12760_n20342.n142 1.037
R10992 a_12760_n20342.n32 a_12760_n20342.n136 1.037
R10993 a_12760_n20342.n30 a_12760_n20342.n130 1.037
R10994 a_12760_n20342.n26 a_12760_n20342.n116 1.037
R10995 a_12760_n20342.n21 a_12760_n20342.n99 1.037
R10996 a_12760_n20342.n82 a_12760_n20342.n189 1.033
R10997 a_12760_n20342.n80 a_12760_n20342.n93 1.033
R10998 a_12760_n20342.n78 a_12760_n20342.n86 1.033
R10999 a_12760_n20342.n77 a_12760_n20342.n83 1.033
R11000 a_12760_n20342.n20 a_12760_n20342.n79 0.965
R11001 a_12760_n20342.n82 a_12760_n20342.n17 0.838
R11002 a_12760_n20342.n16 a_12760_n20342.n15 0.834
R11003 a_12760_n20342.n13 a_12760_n20342.n12 0.834
R11004 a_12760_n20342.n11 a_12760_n20342.n10 0.834
R11005 a_12760_n20342.n10 a_12760_n20342.n9 0.834
R11006 a_12760_n20342.n9 a_12760_n20342.n8 0.834
R11007 a_12760_n20342.n4 a_12760_n20342.n3 0.834
R11008 a_12760_n20342.n17 a_12760_n20342.n16 0.831
R11009 a_12760_n20342.n18 a_12760_n20342.n11 0.79
R11010 a_12760_n20342.n75 a_12760_n20342.n291 0.763
R11011 a_12760_n20342.n74 a_12760_n20342.n283 0.763
R11012 a_12760_n20342.n73 a_12760_n20342.n284 0.763
R11013 a_12760_n20342.n72 a_12760_n20342.n275 0.763
R11014 a_12760_n20342.n71 a_12760_n20342.n276 0.763
R11015 a_12760_n20342.n66 a_12760_n20342.n254 0.763
R11016 a_12760_n20342.n65 a_12760_n20342.n250 0.763
R11017 a_12760_n20342.n63 a_12760_n20342.n255 0.763
R11018 a_12760_n20342.n62 a_12760_n20342.n256 0.763
R11019 a_12760_n20342.n60 a_12760_n20342.n236 0.763
R11020 a_12760_n20342.n59 a_12760_n20342.n237 0.763
R11021 a_12760_n20342.n57 a_12760_n20342.n224 0.763
R11022 a_12760_n20342.n56 a_12760_n20342.n225 0.763
R11023 a_12760_n20342.n55 a_12760_n20342.n226 0.763
R11024 a_12760_n20342.n53 a_12760_n20342.n207 0.763
R11025 a_12760_n20342.n49 a_12760_n20342.n211 0.763
R11026 a_12760_n20342.n185 a_12760_n20342.n47 0.763
R11027 a_12760_n20342.n178 a_12760_n20342.n45 0.763
R11028 a_12760_n20342.n5 a_12760_n20342.n44 0.763
R11029 a_12760_n20342.n11 a_12760_n20342.n43 0.763
R11030 a_12760_n20342.n13 a_12760_n20342.n41 0.763
R11031 a_12760_n20342.n13 a_12760_n20342.n40 0.763
R11032 a_12760_n20342.n12 a_12760_n20342.n39 0.763
R11033 a_12760_n20342.n4 a_12760_n20342.n38 0.763
R11034 a_12760_n20342.n3 a_12760_n20342.n37 0.763
R11035 a_12760_n20342.n4 a_12760_n20342.n36 0.763
R11036 a_12760_n20342.n10 a_12760_n20342.n35 0.763
R11037 a_12760_n20342.n10 a_12760_n20342.n33 0.763
R11038 a_12760_n20342.n9 a_12760_n20342.n31 0.763
R11039 a_12760_n20342.n128 a_12760_n20342.n29 0.763
R11040 a_12760_n20342.n129 a_12760_n20342.n28 0.763
R11041 a_12760_n20342.n9 a_12760_n20342.n27 0.763
R11042 a_12760_n20342.n114 a_12760_n20342.n25 0.763
R11043 a_12760_n20342.n115 a_12760_n20342.n24 0.763
R11044 a_12760_n20342.n8 a_12760_n20342.n23 0.763
R11045 a_12760_n20342.n11 a_12760_n20342.n22 0.763
R11046 a_12760_n20342.n79 a_12760_n20342.n90 0.752
R11047 a_12760_n20342.n49 a_12760_n20342.n192 0.752
R11048 a_12760_n20342.n50 a_12760_n20342.n195 0.752
R11049 a_12760_n20342.n52 a_12760_n20342.n201 0.752
R11050 a_12760_n20342.n57 a_12760_n20342.n218 0.752
R11051 a_12760_n20342.n56 a_12760_n20342.n215 0.752
R11052 a_12760_n20342.n55 a_12760_n20342.n212 0.752
R11053 a_12760_n20342.n23 a_12760_n20342.n105 0.752
R11054 a_12760_n20342.n24 a_12760_n20342.n108 0.752
R11055 a_12760_n20342.n47 a_12760_n20342.n182 0.752
R11056 a_12760_n20342.n46 a_12760_n20342.n179 0.752
R11057 a_12760_n20342.n43 a_12760_n20342.n169 0.752
R11058 a_12760_n20342.n75 a_12760_n20342.n285 0.752
R11059 a_12760_n20342.n73 a_12760_n20342.n277 0.752
R11060 a_12760_n20342.n70 a_12760_n20342.n266 0.752
R11061 a_12760_n20342.n68 a_12760_n20342.n260 0.752
R11062 a_12760_n20342.n35 a_12760_n20342.n145 0.752
R11063 a_12760_n20342.n36 a_12760_n20342.n148 0.752
R11064 a_12760_n20342.n40 a_12760_n20342.n160 0.752
R11065 a_12760_n20342.n33 a_12760_n20342.n139 0.752
R11066 a_12760_n20342.n63 a_12760_n20342.n241 0.752
R11067 a_12760_n20342.n59 a_12760_n20342.n227 0.752
R11068 a_12760_n20342.n27 a_12760_n20342.n119 0.752
R11069 a_12760_n20342.n28 a_12760_n20342.n122 0.752
R11070 a_12760_n20342.n29 a_12760_n20342.n125 0.752
R11071 a_12760_n20342.n60 a_12760_n20342.n230 0.752
R11072 a_12760_n20342.n65 a_12760_n20342.n247 0.752
R11073 a_12760_n20342.n62 a_12760_n20342.n238 0.752
R11074 a_12760_n20342.n31 a_12760_n20342.n133 0.752
R11075 a_12760_n20342.n37 a_12760_n20342.n151 0.752
R11076 a_12760_n20342.n39 a_12760_n20342.n157 0.752
R11077 a_12760_n20342.n64 a_12760_n20342.n244 0.752
R11078 a_12760_n20342.n66 a_12760_n20342.n251 0.752
R11079 a_12760_n20342.n71 a_12760_n20342.n269 0.752
R11080 a_12760_n20342.n72 a_12760_n20342.n272 0.752
R11081 a_12760_n20342.n44 a_12760_n20342.n172 0.752
R11082 a_12760_n20342.n45 a_12760_n20342.n175 0.752
R11083 a_12760_n20342.n22 a_12760_n20342.n102 0.752
R11084 a_12760_n20342.n38 a_12760_n20342.n154 0.752
R11085 a_12760_n20342.n41 a_12760_n20342.n163 0.752
R11086 a_12760_n20342.n74 a_12760_n20342.n280 0.752
R11087 a_12760_n20342.n53 a_12760_n20342.n204 0.752
R11088 a_12760_n20342.n81 a_12760_n20342.n96 0.752
R11089 a_12760_n20342.n25 a_12760_n20342.n111 0.752
R11090 a_12760_n20342.n18 a_12760_n20342.n81 0.743
R11091 a_12760_n20342.n79 a_12760_n20342.n18 0.743
R11092 a_2370_n29452.n4 a_2370_n29452.t8 145.713
R11093 a_2370_n29452.n3 a_2370_n29452.t11 145.462
R11094 a_2370_n29452.n4 a_2370_n29452.t10 140.804
R11095 a_2370_n29452.n3 a_2370_n29452.t9 140.553
R11096 a_2370_n29452.n5 a_2370_n29452.n4 9.199
R11097 a_2370_n29452.n6 a_2370_n29452.n5 8.276
R11098 a_2370_n29452.n8 a_2370_n29452.n7 5.784
R11099 a_2370_n29452.n5 a_2370_n29452.n3 4.589
R11100 a_2370_n29452.n0 a_2370_n29452.t4 4.132
R11101 a_2370_n29452.n0 a_2370_n29452.t3 4.132
R11102 a_2370_n29452.n1 a_2370_n29452.t2 4.132
R11103 a_2370_n29452.n1 a_2370_n29452.t1 4.132
R11104 a_2370_n29452.n2 a_2370_n29452.t7 4.132
R11105 a_2370_n29452.n2 a_2370_n29452.t6 4.132
R11106 a_2370_n29452.t0 a_2370_n29452.n9 4.132
R11107 a_2370_n29452.n9 a_2370_n29452.t5 4.132
R11108 a_2370_n29452.n9 a_2370_n29452.n8 2.723
R11109 a_2370_n29452.n8 a_2370_n29452.n0 2.126
R11110 a_2370_n29452.n7 a_2370_n29452.n1 2.126
R11111 a_2370_n29452.n6 a_2370_n29452.n2 2.126
R11112 a_2370_n29452.n7 a_2370_n29452.n6 0.597
R11113 Vfold_bot_m Vfold_bot_m.n6 12.649
R11114 Vfold_bot_m.n3 Vfold_bot_m.t109 9.688
R11115 Vfold_bot_m.n6 Vfold_bot_m.t54 9.038
R11116 Vfold_bot_m.n103 Vfold_bot_m.t27 8.266
R11117 Vfold_bot_m.n98 Vfold_bot_m.t83 8.266
R11118 Vfold_bot_m.n98 Vfold_bot_m.t112 8.266
R11119 Vfold_bot_m.n97 Vfold_bot_m.t103 8.266
R11120 Vfold_bot_m.n97 Vfold_bot_m.t14 8.266
R11121 Vfold_bot_m.n100 Vfold_bot_m.t11 8.266
R11122 Vfold_bot_m.n100 Vfold_bot_m.t87 8.266
R11123 Vfold_bot_m.n99 Vfold_bot_m.t73 8.266
R11124 Vfold_bot_m.n99 Vfold_bot_m.t36 8.266
R11125 Vfold_bot_m.n96 Vfold_bot_m.t81 8.266
R11126 Vfold_bot_m.n96 Vfold_bot_m.t33 8.266
R11127 Vfold_bot_m.n95 Vfold_bot_m.t102 8.266
R11128 Vfold_bot_m.n95 Vfold_bot_m.t113 8.266
R11129 Vfold_bot_m.n70 Vfold_bot_m.t94 8.266
R11130 Vfold_bot_m.n70 Vfold_bot_m.t55 8.266
R11131 Vfold_bot_m.n69 Vfold_bot_m.t71 8.266
R11132 Vfold_bot_m.n69 Vfold_bot_m.t28 8.266
R11133 Vfold_bot_m.n72 Vfold_bot_m.t74 8.266
R11134 Vfold_bot_m.n72 Vfold_bot_m.t39 8.266
R11135 Vfold_bot_m.n71 Vfold_bot_m.t93 8.266
R11136 Vfold_bot_m.n71 Vfold_bot_m.t15 8.266
R11137 Vfold_bot_m.n74 Vfold_bot_m.t95 8.266
R11138 Vfold_bot_m.n74 Vfold_bot_m.t56 8.266
R11139 Vfold_bot_m.n73 Vfold_bot_m.t72 8.266
R11140 Vfold_bot_m.n73 Vfold_bot_m.t40 8.266
R11141 Vfold_bot_m.n76 Vfold_bot_m.t101 8.266
R11142 Vfold_bot_m.n76 Vfold_bot_m.t4 8.266
R11143 Vfold_bot_m.n75 Vfold_bot_m.t86 8.266
R11144 Vfold_bot_m.n75 Vfold_bot_m.t29 8.266
R11145 Vfold_bot_m.n28 Vfold_bot_m.t84 8.266
R11146 Vfold_bot_m.n28 Vfold_bot_m.t13 8.266
R11147 Vfold_bot_m.n27 Vfold_bot_m.t68 8.266
R11148 Vfold_bot_m.n27 Vfold_bot_m.t25 8.266
R11149 Vfold_bot_m.n30 Vfold_bot_m.t67 8.266
R11150 Vfold_bot_m.n30 Vfold_bot_m.t26 8.266
R11151 Vfold_bot_m.n29 Vfold_bot_m.t92 8.266
R11152 Vfold_bot_m.n29 Vfold_bot_m.t59 8.266
R11153 Vfold_bot_m.n32 Vfold_bot_m.t88 8.266
R11154 Vfold_bot_m.n32 Vfold_bot_m.t3 8.266
R11155 Vfold_bot_m.n31 Vfold_bot_m.t69 8.266
R11156 Vfold_bot_m.n31 Vfold_bot_m.t57 8.266
R11157 Vfold_bot_m.n34 Vfold_bot_m.t100 8.266
R11158 Vfold_bot_m.n34 Vfold_bot_m.t35 8.266
R11159 Vfold_bot_m.n33 Vfold_bot_m.t97 8.266
R11160 Vfold_bot_m.n33 Vfold_bot_m.t58 8.266
R11161 Vfold_bot_m.n23 Vfold_bot_m.t96 8.266
R11162 Vfold_bot_m.n23 Vfold_bot_m.t12 8.266
R11163 Vfold_bot_m.n22 Vfold_bot_m.t77 8.266
R11164 Vfold_bot_m.n22 Vfold_bot_m.t37 8.266
R11165 Vfold_bot_m.n25 Vfold_bot_m.t76 8.266
R11166 Vfold_bot_m.n25 Vfold_bot_m.t38 8.266
R11167 Vfold_bot_m.n24 Vfold_bot_m.t99 8.266
R11168 Vfold_bot_m.n24 Vfold_bot_m.t114 8.266
R11169 Vfold_bot_m.n8 Vfold_bot_m.t65 8.266
R11170 Vfold_bot_m.n8 Vfold_bot_m.t42 8.266
R11171 Vfold_bot_m.n7 Vfold_bot_m.t90 8.266
R11172 Vfold_bot_m.n7 Vfold_bot_m.t51 8.266
R11173 Vfold_bot_m.n10 Vfold_bot_m.t89 8.266
R11174 Vfold_bot_m.n10 Vfold_bot_m.t50 8.266
R11175 Vfold_bot_m.n9 Vfold_bot_m.t70 8.266
R11176 Vfold_bot_m.n9 Vfold_bot_m.t44 8.266
R11177 Vfold_bot_m.n14 Vfold_bot_m.t66 8.266
R11178 Vfold_bot_m.n14 Vfold_bot_m.t43 8.266
R11179 Vfold_bot_m.n13 Vfold_bot_m.t91 8.266
R11180 Vfold_bot_m.n13 Vfold_bot_m.t47 8.266
R11181 Vfold_bot_m.n12 Vfold_bot_m.t75 8.266
R11182 Vfold_bot_m.n12 Vfold_bot_m.t48 8.266
R11183 Vfold_bot_m.n11 Vfold_bot_m.t98 8.266
R11184 Vfold_bot_m.n11 Vfold_bot_m.t52 8.266
R11185 Vfold_bot_m.n18 Vfold_bot_m.t85 8.266
R11186 Vfold_bot_m.n18 Vfold_bot_m.t41 8.266
R11187 Vfold_bot_m.n17 Vfold_bot_m.t80 8.266
R11188 Vfold_bot_m.n17 Vfold_bot_m.t45 8.266
R11189 Vfold_bot_m.n16 Vfold_bot_m.t82 8.266
R11190 Vfold_bot_m.n16 Vfold_bot_m.t46 8.266
R11191 Vfold_bot_m.n15 Vfold_bot_m.t78 8.266
R11192 Vfold_bot_m.n15 Vfold_bot_m.t49 8.266
R11193 Vfold_bot_m.n102 Vfold_bot_m.t79 8.266
R11194 Vfold_bot_m.n102 Vfold_bot_m.t34 8.266
R11195 Vfold_bot_m.n103 Vfold_bot_m.t104 8.266
R11196 Vfold_bot_m.n106 Vfold_bot_m.n94 8.129
R11197 Vfold_bot_m.n2 Vfold_bot_m.t60 6.923
R11198 Vfold_bot_m.n2 Vfold_bot_m.t64 6.923
R11199 Vfold_bot_m.n1 Vfold_bot_m.t53 6.923
R11200 Vfold_bot_m.n1 Vfold_bot_m.t63 6.923
R11201 Vfold_bot_m.n0 Vfold_bot_m.t119 6.923
R11202 Vfold_bot_m.n0 Vfold_bot_m.t108 6.923
R11203 Vfold_bot_m.n67 Vfold_bot_m.n43 4.849
R11204 Vfold_bot_m.n108 Vfold_bot_m.n68 4.848
R11205 Vfold_bot_m.n62 Vfold_bot_m.n61 4.827
R11206 Vfold_bot_m.n64 Vfold_bot_m.n53 4.826
R11207 Vfold_bot_m.n65 Vfold_bot_m.n49 4.826
R11208 Vfold_bot_m.n45 Vfold_bot_m.t16 3.557
R11209 Vfold_bot_m.n44 Vfold_bot_m.t118 3.557
R11210 Vfold_bot_m.n88 Vfold_bot_m.t116 3.557
R11211 Vfold_bot_m.n89 Vfold_bot_m.t17 3.557
R11212 Vfold_bot_m.n43 Vfold_bot_m.t22 3.557
R11213 Vfold_bot_m.n42 Vfold_bot_m.t61 3.557
R11214 Vfold_bot_m.n41 Vfold_bot_m.t111 3.557
R11215 Vfold_bot_m.n40 Vfold_bot_m.t32 3.557
R11216 Vfold_bot_m.n39 Vfold_bot_m.t115 3.557
R11217 Vfold_bot_m.n38 Vfold_bot_m.t2 3.557
R11218 Vfold_bot_m.n92 Vfold_bot_m.t110 3.557
R11219 Vfold_bot_m.n93 Vfold_bot_m.t105 3.557
R11220 Vfold_bot_m.n58 Vfold_bot_m.t23 3.536
R11221 Vfold_bot_m.n59 Vfold_bot_m.t8 3.536
R11222 Vfold_bot_m.n60 Vfold_bot_m.t24 3.536
R11223 Vfold_bot_m.n61 Vfold_bot_m.t21 3.536
R11224 Vfold_bot_m.n57 Vfold_bot_m.t6 3.536
R11225 Vfold_bot_m.n56 Vfold_bot_m.t20 3.536
R11226 Vfold_bot_m.n80 Vfold_bot_m.t0 3.536
R11227 Vfold_bot_m.n81 Vfold_bot_m.t117 3.536
R11228 Vfold_bot_m.n55 Vfold_bot_m.t19 3.536
R11229 Vfold_bot_m.n54 Vfold_bot_m.t62 3.536
R11230 Vfold_bot_m.n83 Vfold_bot_m.t31 3.536
R11231 Vfold_bot_m.n84 Vfold_bot_m.t18 3.536
R11232 Vfold_bot_m.n53 Vfold_bot_m.t5 3.536
R11233 Vfold_bot_m.n52 Vfold_bot_m.t107 3.536
R11234 Vfold_bot_m.n51 Vfold_bot_m.t9 3.536
R11235 Vfold_bot_m.n50 Vfold_bot_m.t106 3.536
R11236 Vfold_bot_m.n49 Vfold_bot_m.t10 3.536
R11237 Vfold_bot_m.n48 Vfold_bot_m.t1 3.536
R11238 Vfold_bot_m.n47 Vfold_bot_m.t30 3.536
R11239 Vfold_bot_m.n46 Vfold_bot_m.t7 3.536
R11240 Vfold_bot_m.n19 Vfold_bot_m.n18 2.67
R11241 Vfold_bot_m.n101 Vfold_bot_m.n100 2.668
R11242 Vfold_bot_m.n77 Vfold_bot_m.n76 2.668
R11243 Vfold_bot_m.n35 Vfold_bot_m.n34 2.668
R11244 Vfold_bot_m.n26 Vfold_bot_m.n25 2.668
R11245 Vfold_bot_m.n20 Vfold_bot_m.n19 2.22
R11246 Vfold_bot_m.n104 Vfold_bot_m.n101 2.219
R11247 Vfold_bot_m.n78 Vfold_bot_m.n77 2.219
R11248 Vfold_bot_m.n79 Vfold_bot_m.n78 2.219
R11249 Vfold_bot_m.n36 Vfold_bot_m.n35 2.219
R11250 Vfold_bot_m.n37 Vfold_bot_m.n36 2.219
R11251 Vfold_bot_m.n21 Vfold_bot_m.n20 2.219
R11252 Vfold_bot_m.n105 Vfold_bot_m.n104 2.219
R11253 Vfold_bot_m.n3 Vfold_bot_m.n2 2.115
R11254 Vfold_bot_m.n4 Vfold_bot_m.n1 2.115
R11255 Vfold_bot_m.n5 Vfold_bot_m.n0 2.115
R11256 Vfold_bot_m.n62 Vfold_bot_m.n57 1.808
R11257 Vfold_bot_m.n66 Vfold_bot_m.n45 1.643
R11258 Vfold_bot_m.n68 Vfold_bot_m.n39 1.643
R11259 Vfold_bot_m.n63 Vfold_bot_m.n55 1.62
R11260 Vfold_bot_m.n82 Vfold_bot_m.n81 1.496
R11261 Vfold_bot_m.n45 Vfold_bot_m.n44 1.414
R11262 Vfold_bot_m.n89 Vfold_bot_m.n88 1.414
R11263 Vfold_bot_m.n43 Vfold_bot_m.n42 1.414
R11264 Vfold_bot_m.n42 Vfold_bot_m.n41 1.414
R11265 Vfold_bot_m.n41 Vfold_bot_m.n40 1.414
R11266 Vfold_bot_m.n39 Vfold_bot_m.n38 1.414
R11267 Vfold_bot_m.n93 Vfold_bot_m.n92 1.414
R11268 Vfold_bot_m.n59 Vfold_bot_m.n58 1.361
R11269 Vfold_bot_m.n60 Vfold_bot_m.n59 1.361
R11270 Vfold_bot_m.n61 Vfold_bot_m.n60 1.361
R11271 Vfold_bot_m.n57 Vfold_bot_m.n56 1.361
R11272 Vfold_bot_m.n81 Vfold_bot_m.n80 1.361
R11273 Vfold_bot_m.n55 Vfold_bot_m.n54 1.361
R11274 Vfold_bot_m.n84 Vfold_bot_m.n83 1.361
R11275 Vfold_bot_m.n53 Vfold_bot_m.n52 1.361
R11276 Vfold_bot_m.n52 Vfold_bot_m.n51 1.361
R11277 Vfold_bot_m.n51 Vfold_bot_m.n50 1.361
R11278 Vfold_bot_m.n49 Vfold_bot_m.n48 1.361
R11279 Vfold_bot_m.n48 Vfold_bot_m.n47 1.361
R11280 Vfold_bot_m.n47 Vfold_bot_m.n46 1.361
R11281 Vfold_bot_m.n90 Vfold_bot_m.n89 1.338
R11282 Vfold_bot_m.n94 Vfold_bot_m.n93 1.338
R11283 Vfold_bot_m Vfold_bot_m.n111 1.317
R11284 Vfold_bot_m.n85 Vfold_bot_m.n84 1.308
R11285 Vfold_bot_m.n107 Vfold_bot_m.n79 1.116
R11286 Vfold_bot_m.n109 Vfold_bot_m.n37 1.116
R11287 Vfold_bot_m.n110 Vfold_bot_m.n26 1.116
R11288 Vfold_bot_m.n111 Vfold_bot_m.n21 1.116
R11289 Vfold_bot_m.n106 Vfold_bot_m.n105 1.116
R11290 Vfold_bot_m.n111 Vfold_bot_m.n110 0.752
R11291 Vfold_bot_m.n110 Vfold_bot_m.n109 0.752
R11292 Vfold_bot_m.n107 Vfold_bot_m.n106 0.752
R11293 Vfold_bot_m.n13 Vfold_bot_m.n12 0.687
R11294 Vfold_bot_m.n17 Vfold_bot_m.n16 0.687
R11295 Vfold_bot_m.n5 Vfold_bot_m.n4 0.65
R11296 Vfold_bot_m.n6 Vfold_bot_m.n5 0.65
R11297 Vfold_bot_m.n4 Vfold_bot_m.n3 0.637
R11298 Vfold_bot_m.n108 Vfold_bot_m.n107 0.592
R11299 Vfold_bot_m.n101 Vfold_bot_m.n98 0.449
R11300 Vfold_bot_m.n105 Vfold_bot_m.n96 0.449
R11301 Vfold_bot_m.n79 Vfold_bot_m.n70 0.449
R11302 Vfold_bot_m.n78 Vfold_bot_m.n72 0.449
R11303 Vfold_bot_m.n77 Vfold_bot_m.n74 0.449
R11304 Vfold_bot_m.n37 Vfold_bot_m.n28 0.449
R11305 Vfold_bot_m.n36 Vfold_bot_m.n30 0.449
R11306 Vfold_bot_m.n35 Vfold_bot_m.n32 0.449
R11307 Vfold_bot_m.n26 Vfold_bot_m.n23 0.449
R11308 Vfold_bot_m.n21 Vfold_bot_m.n8 0.449
R11309 Vfold_bot_m.n20 Vfold_bot_m.n10 0.449
R11310 Vfold_bot_m.n19 Vfold_bot_m.n14 0.449
R11311 Vfold_bot_m.n104 Vfold_bot_m.n103 0.449
R11312 Vfold_bot_m.n98 Vfold_bot_m.n97 0.365
R11313 Vfold_bot_m.n100 Vfold_bot_m.n99 0.365
R11314 Vfold_bot_m.n96 Vfold_bot_m.n95 0.365
R11315 Vfold_bot_m.n70 Vfold_bot_m.n69 0.365
R11316 Vfold_bot_m.n72 Vfold_bot_m.n71 0.365
R11317 Vfold_bot_m.n74 Vfold_bot_m.n73 0.365
R11318 Vfold_bot_m.n76 Vfold_bot_m.n75 0.365
R11319 Vfold_bot_m.n28 Vfold_bot_m.n27 0.365
R11320 Vfold_bot_m.n30 Vfold_bot_m.n29 0.365
R11321 Vfold_bot_m.n32 Vfold_bot_m.n31 0.365
R11322 Vfold_bot_m.n34 Vfold_bot_m.n33 0.365
R11323 Vfold_bot_m.n23 Vfold_bot_m.n22 0.365
R11324 Vfold_bot_m.n25 Vfold_bot_m.n24 0.365
R11325 Vfold_bot_m.n8 Vfold_bot_m.n7 0.365
R11326 Vfold_bot_m.n10 Vfold_bot_m.n9 0.365
R11327 Vfold_bot_m.n12 Vfold_bot_m.n11 0.365
R11328 Vfold_bot_m.n14 Vfold_bot_m.n13 0.365
R11329 Vfold_bot_m.n16 Vfold_bot_m.n15 0.365
R11330 Vfold_bot_m.n18 Vfold_bot_m.n17 0.365
R11331 Vfold_bot_m.n103 Vfold_bot_m.n102 0.365
R11332 Vfold_bot_m.n68 Vfold_bot_m.n67 0.188
R11333 Vfold_bot_m.n67 Vfold_bot_m.n66 0.188
R11334 Vfold_bot_m.n66 Vfold_bot_m.n65 0.188
R11335 Vfold_bot_m.n65 Vfold_bot_m.n64 0.188
R11336 Vfold_bot_m.n64 Vfold_bot_m.n63 0.188
R11337 Vfold_bot_m.n63 Vfold_bot_m.n62 0.188
R11338 Vfold_bot_m.n94 Vfold_bot_m.n91 0.188
R11339 Vfold_bot_m.n91 Vfold_bot_m.n90 0.188
R11340 Vfold_bot_m.n90 Vfold_bot_m.n87 0.188
R11341 Vfold_bot_m.n87 Vfold_bot_m.n86 0.188
R11342 Vfold_bot_m.n86 Vfold_bot_m.n85 0.188
R11343 Vfold_bot_m.n85 Vfold_bot_m.n82 0.188
R11344 Vfold_bot_m.n109 Vfold_bot_m.n108 0.159
R11345 a_2467_n29152.n3 a_2467_n29152.t7 14.598
R11346 a_2467_n29152.n8 a_2467_n29152.t14 14.598
R11347 a_2467_n29152.n7 a_2467_n29152.t9 13.849
R11348 a_2467_n29152.n6 a_2467_n29152.t15 13.849
R11349 a_2467_n29152.n5 a_2467_n29152.t6 13.849
R11350 a_2467_n29152.n4 a_2467_n29152.t10 13.849
R11351 a_2467_n29152.n3 a_2467_n29152.t12 13.849
R11352 a_2467_n29152.n12 a_2467_n29152.t16 13.849
R11353 a_2467_n29152.n11 a_2467_n29152.t11 13.849
R11354 a_2467_n29152.n10 a_2467_n29152.t13 13.849
R11355 a_2467_n29152.n9 a_2467_n29152.t17 13.849
R11356 a_2467_n29152.n8 a_2467_n29152.t8 13.849
R11357 a_2467_n29152.n14 a_2467_n29152.n13 10.655
R11358 a_2467_n29152.t5 a_2467_n29152.n17 8.564
R11359 a_2467_n29152.n0 a_2467_n29152.t2 8.535
R11360 a_2467_n29152.n17 a_2467_n29152.t0 8.376
R11361 a_2467_n29152.n16 a_2467_n29152.t19 8.376
R11362 a_2467_n29152.n15 a_2467_n29152.t3 8.376
R11363 a_2467_n29152.n0 a_2467_n29152.t18 8.347
R11364 a_2467_n29152.n1 a_2467_n29152.t1 8.347
R11365 a_2467_n29152.n2 a_2467_n29152.t4 8.347
R11366 a_2467_n29152.n15 a_2467_n29152.n14 5.589
R11367 a_2467_n29152.n13 a_2467_n29152.n12 2.584
R11368 a_2467_n29152.n4 a_2467_n29152.n3 1.159
R11369 a_2467_n29152.n6 a_2467_n29152.n5 1.159
R11370 a_2467_n29152.n9 a_2467_n29152.n8 1.159
R11371 a_2467_n29152.n11 a_2467_n29152.n10 1.159
R11372 a_2467_n29152.n5 a_2467_n29152.n4 0.749
R11373 a_2467_n29152.n7 a_2467_n29152.n6 0.749
R11374 a_2467_n29152.n10 a_2467_n29152.n9 0.749
R11375 a_2467_n29152.n12 a_2467_n29152.n11 0.749
R11376 a_2467_n29152.n14 a_2467_n29152.n2 0.683
R11377 a_2467_n29152.n13 a_2467_n29152.n7 0.385
R11378 a_2467_n29152.n2 a_2467_n29152.n1 0.188
R11379 a_2467_n29152.n1 a_2467_n29152.n0 0.188
R11380 a_2467_n29152.n16 a_2467_n29152.n15 0.188
R11381 a_2467_n29152.n17 a_2467_n29152.n16 0.188
R11382 a_2458_6128.n170 a_2458_6128.t116 13.849
R11383 a_2458_6128.n169 a_2458_6128.t55 13.849
R11384 a_2458_6128.n169 a_2458_6128.t98 13.849
R11385 a_2458_6128.n6 a_2458_6128.t9 13.849
R11386 a_2458_6128.n6 a_2458_6128.t157 13.849
R11387 a_2458_6128.n5 a_2458_6128.t60 13.849
R11388 a_2458_6128.n5 a_2458_6128.t112 13.849
R11389 a_2458_6128.n8 a_2458_6128.t1 13.849
R11390 a_2458_6128.n8 a_2458_6128.t128 13.849
R11391 a_2458_6128.n7 a_2458_6128.t86 13.849
R11392 a_2458_6128.n7 a_2458_6128.t151 13.849
R11393 a_2458_6128.n10 a_2458_6128.t41 13.849
R11394 a_2458_6128.n10 a_2458_6128.t136 13.849
R11395 a_2458_6128.n9 a_2458_6128.t35 13.849
R11396 a_2458_6128.n9 a_2458_6128.t115 13.849
R11397 a_2458_6128.n12 a_2458_6128.t180 13.849
R11398 a_2458_6128.n12 a_2458_6128.t152 13.849
R11399 a_2458_6128.n11 a_2458_6128.t186 13.849
R11400 a_2458_6128.n11 a_2458_6128.t118 13.849
R11401 a_2458_6128.n14 a_2458_6128.t185 13.849
R11402 a_2458_6128.n14 a_2458_6128.t102 13.849
R11403 a_2458_6128.n13 a_2458_6128.t178 13.849
R11404 a_2458_6128.n13 a_2458_6128.t160 13.849
R11405 a_2458_6128.n16 a_2458_6128.t179 13.849
R11406 a_2458_6128.n16 a_2458_6128.t156 13.849
R11407 a_2458_6128.n15 a_2458_6128.t184 13.849
R11408 a_2458_6128.n15 a_2458_6128.t133 13.849
R11409 a_2458_6128.n18 a_2458_6128.t194 13.849
R11410 a_2458_6128.n18 a_2458_6128.t134 13.849
R11411 a_2458_6128.n17 a_2458_6128.t77 13.849
R11412 a_2458_6128.n17 a_2458_6128.t166 13.849
R11413 a_2458_6128.n20 a_2458_6128.t3 13.849
R11414 a_2458_6128.n20 a_2458_6128.t124 13.849
R11415 a_2458_6128.n19 a_2458_6128.t76 13.849
R11416 a_2458_6128.n19 a_2458_6128.t140 13.849
R11417 a_2458_6128.n22 a_2458_6128.t40 13.849
R11418 a_2458_6128.n22 a_2458_6128.t135 13.849
R11419 a_2458_6128.n21 a_2458_6128.t56 13.849
R11420 a_2458_6128.n21 a_2458_6128.t110 13.849
R11421 a_2458_6128.n24 a_2458_6128.t17 13.849
R11422 a_2458_6128.n24 a_2458_6128.t139 13.849
R11423 a_2458_6128.n23 a_2458_6128.t48 13.849
R11424 a_2458_6128.n23 a_2458_6128.t149 13.849
R11425 a_2458_6128.n26 a_2458_6128.t43 13.849
R11426 a_2458_6128.n26 a_2458_6128.t159 13.849
R11427 a_2458_6128.n25 a_2458_6128.t15 13.849
R11428 a_2458_6128.n25 a_2458_6128.t137 13.849
R11429 a_2458_6128.n28 a_2458_6128.t13 13.849
R11430 a_2458_6128.n28 a_2458_6128.t164 13.849
R11431 a_2458_6128.n27 a_2458_6128.t44 13.849
R11432 a_2458_6128.n27 a_2458_6128.t144 13.849
R11433 a_2458_6128.n30 a_2458_6128.t39 13.849
R11434 a_2458_6128.n30 a_2458_6128.t106 13.849
R11435 a_2458_6128.n29 a_2458_6128.t10 13.849
R11436 a_2458_6128.n29 a_2458_6128.t161 13.849
R11437 a_2458_6128.n32 a_2458_6128.t7 13.849
R11438 a_2458_6128.n32 a_2458_6128.t155 13.849
R11439 a_2458_6128.n31 a_2458_6128.t36 13.849
R11440 a_2458_6128.n31 a_2458_6128.t103 13.849
R11441 a_2458_6128.n34 a_2458_6128.t59 13.849
R11442 a_2458_6128.n34 a_2458_6128.t130 13.849
R11443 a_2458_6128.n33 a_2458_6128.t33 13.849
R11444 a_2458_6128.n33 a_2458_6128.t153 13.849
R11445 a_2458_6128.n36 a_2458_6128.t29 13.849
R11446 a_2458_6128.n36 a_2458_6128.t97 13.849
R11447 a_2458_6128.n35 a_2458_6128.t57 13.849
R11448 a_2458_6128.n35 a_2458_6128.t111 13.849
R11449 a_2458_6128.n141 a_2458_6128.t193 13.849
R11450 a_2458_6128.n141 a_2458_6128.t147 13.849
R11451 a_2458_6128.n140 a_2458_6128.t177 13.849
R11452 a_2458_6128.n140 a_2458_6128.t162 13.849
R11453 a_2458_6128.n143 a_2458_6128.t2 13.849
R11454 a_2458_6128.n143 a_2458_6128.t126 13.849
R11455 a_2458_6128.n142 a_2458_6128.t187 13.849
R11456 a_2458_6128.n142 a_2458_6128.t117 13.849
R11457 a_2458_6128.n145 a_2458_6128.t66 13.849
R11458 a_2458_6128.n145 a_2458_6128.t108 13.849
R11459 a_2458_6128.n144 a_2458_6128.t87 13.849
R11460 a_2458_6128.n144 a_2458_6128.t113 13.849
R11461 a_2458_6128.n147 a_2458_6128.t92 13.849
R11462 a_2458_6128.n147 a_2458_6128.t95 13.849
R11463 a_2458_6128.n146 a_2458_6128.t0 13.849
R11464 a_2458_6128.n146 a_2458_6128.t131 13.849
R11465 a_2458_6128.n99 a_2458_6128.t30 13.849
R11466 a_2458_6128.n99 a_2458_6128.t99 13.849
R11467 a_2458_6128.n98 a_2458_6128.t53 13.849
R11468 a_2458_6128.n98 a_2458_6128.t125 13.849
R11469 a_2458_6128.n101 a_2458_6128.t25 13.849
R11470 a_2458_6128.n101 a_2458_6128.t170 13.849
R11471 a_2458_6128.n100 a_2458_6128.t31 13.849
R11472 a_2458_6128.n100 a_2458_6128.t100 13.849
R11473 a_2458_6128.n103 a_2458_6128.t51 13.849
R11474 a_2458_6128.n103 a_2458_6128.t121 13.849
R11475 a_2458_6128.n102 a_2458_6128.t54 13.849
R11476 a_2458_6128.n102 a_2458_6128.t107 13.849
R11477 a_2458_6128.n105 a_2458_6128.t23 13.849
R11478 a_2458_6128.n105 a_2458_6128.t168 13.849
R11479 a_2458_6128.n104 a_2458_6128.t27 13.849
R11480 a_2458_6128.n104 a_2458_6128.t173 13.849
R11481 a_2458_6128.n107 a_2458_6128.t50 13.849
R11482 a_2458_6128.n107 a_2458_6128.t119 13.849
R11483 a_2458_6128.n106 a_2458_6128.t52 13.849
R11484 a_2458_6128.n106 a_2458_6128.t122 13.849
R11485 a_2458_6128.n109 a_2458_6128.t18 13.849
R11486 a_2458_6128.n109 a_2458_6128.t141 13.849
R11487 a_2458_6128.n108 a_2458_6128.t24 13.849
R11488 a_2458_6128.n108 a_2458_6128.t169 13.849
R11489 a_2458_6128.n111 a_2458_6128.t11 13.849
R11490 a_2458_6128.n111 a_2458_6128.t94 13.849
R11491 a_2458_6128.n110 a_2458_6128.t19 13.849
R11492 a_2458_6128.n110 a_2458_6128.t120 13.849
R11493 a_2458_6128.n113 a_2458_6128.t37 13.849
R11494 a_2458_6128.n113 a_2458_6128.t104 13.849
R11495 a_2458_6128.n112 a_2458_6128.t45 13.849
R11496 a_2458_6128.n112 a_2458_6128.t145 13.849
R11497 a_2458_6128.n76 a_2458_6128.t21 13.849
R11498 a_2458_6128.n76 a_2458_6128.t143 13.849
R11499 a_2458_6128.n75 a_2458_6128.t47 13.849
R11500 a_2458_6128.n75 a_2458_6128.t148 13.849
R11501 a_2458_6128.n78 a_2458_6128.t16 13.849
R11502 a_2458_6128.n78 a_2458_6128.t138 13.849
R11503 a_2458_6128.n77 a_2458_6128.t22 13.849
R11504 a_2458_6128.n77 a_2458_6128.t167 13.849
R11505 a_2458_6128.n80 a_2458_6128.t42 13.849
R11506 a_2458_6128.n80 a_2458_6128.t158 13.849
R11507 a_2458_6128.n79 a_2458_6128.t49 13.849
R11508 a_2458_6128.n79 a_2458_6128.t150 13.849
R11509 a_2458_6128.n82 a_2458_6128.t12 13.849
R11510 a_2458_6128.n82 a_2458_6128.t163 13.849
R11511 a_2458_6128.n81 a_2458_6128.t20 13.849
R11512 a_2458_6128.n81 a_2458_6128.t142 13.849
R11513 a_2458_6128.n84 a_2458_6128.t38 13.849
R11514 a_2458_6128.n84 a_2458_6128.t105 13.849
R11515 a_2458_6128.n83 a_2458_6128.t46 13.849
R11516 a_2458_6128.n83 a_2458_6128.t146 13.849
R11517 a_2458_6128.n86 a_2458_6128.t6 13.849
R11518 a_2458_6128.n86 a_2458_6128.t154 13.849
R11519 a_2458_6128.n85 a_2458_6128.t14 13.849
R11520 a_2458_6128.n85 a_2458_6128.t165 13.849
R11521 a_2458_6128.n88 a_2458_6128.t58 13.849
R11522 a_2458_6128.n88 a_2458_6128.t129 13.849
R11523 a_2458_6128.n87 a_2458_6128.t8 13.849
R11524 a_2458_6128.n87 a_2458_6128.t132 13.849
R11525 a_2458_6128.n90 a_2458_6128.t28 13.849
R11526 a_2458_6128.n90 a_2458_6128.t96 13.849
R11527 a_2458_6128.n89 a_2458_6128.t34 13.849
R11528 a_2458_6128.n89 a_2458_6128.t114 13.849
R11529 a_2458_6128.n1 a_2458_6128.t32 13.849
R11530 a_2458_6128.n1 a_2458_6128.t101 13.849
R11531 a_2458_6128.n0 a_2458_6128.t26 13.849
R11532 a_2458_6128.n0 a_2458_6128.t171 13.849
R11533 a_2458_6128.n3 a_2458_6128.t4 13.849
R11534 a_2458_6128.n3 a_2458_6128.t123 13.849
R11535 a_2458_6128.n2 a_2458_6128.t191 13.849
R11536 a_2458_6128.n2 a_2458_6128.t172 13.849
R11537 a_2458_6128.n167 a_2458_6128.t190 13.849
R11538 a_2458_6128.n167 a_2458_6128.t109 13.849
R11539 a_2458_6128.n166 a_2458_6128.t81 13.849
R11540 a_2458_6128.n166 a_2458_6128.t127 13.849
R11541 a_2458_6128.t61 a_2458_6128.n170 13.849
R11542 a_2458_6128.n154 a_2458_6128.t196 10.855
R11543 a_2458_6128.n158 a_2458_6128.n157 8.834
R11544 a_2458_6128.n157 a_2458_6128.t91 8.266
R11545 a_2458_6128.n153 a_2458_6128.t64 8.265
R11546 a_2458_6128.n153 a_2458_6128.t65 8.265
R11547 a_2458_6128.n152 a_2458_6128.t197 8.265
R11548 a_2458_6128.n152 a_2458_6128.t198 8.265
R11549 a_2458_6128.n151 a_2458_6128.t195 8.265
R11550 a_2458_6128.n151 a_2458_6128.t189 8.265
R11551 a_2458_6128.n136 a_2458_6128.n135 6.78
R11552 a_2458_6128.n64 a_2458_6128.n63 5.009
R11553 a_2458_6128.n74 a_2458_6128.n73 4.822
R11554 a_2458_6128.n68 a_2458_6128.n49 4.821
R11555 a_2458_6128.n65 a_2458_6128.n57 4.821
R11556 a_2458_6128.n138 a_2458_6128.n74 3.31
R11557 a_2458_6128.n37 a_2458_6128.n36 2.739
R11558 a_2458_6128.n148 a_2458_6128.n147 2.739
R11559 a_2458_6128.n114 a_2458_6128.n113 2.739
R11560 a_2458_6128.n91 a_2458_6128.n90 2.739
R11561 a_2458_6128.n38 a_2458_6128.n37 2.199
R11562 a_2458_6128.n39 a_2458_6128.n38 2.199
R11563 a_2458_6128.n40 a_2458_6128.n39 2.199
R11564 a_2458_6128.n41 a_2458_6128.n40 2.199
R11565 a_2458_6128.n42 a_2458_6128.n41 2.199
R11566 a_2458_6128.n43 a_2458_6128.n42 2.199
R11567 a_2458_6128.n149 a_2458_6128.n148 2.199
R11568 a_2458_6128.n150 a_2458_6128.n149 2.199
R11569 a_2458_6128.n115 a_2458_6128.n114 2.199
R11570 a_2458_6128.n116 a_2458_6128.n115 2.199
R11571 a_2458_6128.n117 a_2458_6128.n116 2.199
R11572 a_2458_6128.n118 a_2458_6128.n117 2.199
R11573 a_2458_6128.n119 a_2458_6128.n118 2.199
R11574 a_2458_6128.n120 a_2458_6128.n119 2.199
R11575 a_2458_6128.n92 a_2458_6128.n91 2.199
R11576 a_2458_6128.n93 a_2458_6128.n92 2.199
R11577 a_2458_6128.n94 a_2458_6128.n93 2.199
R11578 a_2458_6128.n95 a_2458_6128.n94 2.199
R11579 a_2458_6128.n96 a_2458_6128.n95 2.199
R11580 a_2458_6128.n97 a_2458_6128.n96 2.199
R11581 a_2458_6128.n161 a_2458_6128.n160 2.199
R11582 a_2458_6128.n162 a_2458_6128.n161 2.199
R11583 a_2458_6128.n163 a_2458_6128.n162 2.199
R11584 a_2458_6128.n164 a_2458_6128.n163 2.199
R11585 a_2458_6128.n165 a_2458_6128.n164 2.199
R11586 a_2458_6128.n168 a_2458_6128.n165 2.199
R11587 a_2458_6128.n168 a_2458_6128.n4 2.199
R11588 a_2458_6128.n70 a_2458_6128.t188 2.067
R11589 a_2458_6128.n71 a_2458_6128.t199 2.067
R11590 a_2458_6128.n72 a_2458_6128.t63 2.067
R11591 a_2458_6128.n73 a_2458_6128.t67 2.067
R11592 a_2458_6128.n63 a_2458_6128.t79 2.067
R11593 a_2458_6128.n62 a_2458_6128.t175 2.067
R11594 a_2458_6128.n61 a_2458_6128.t80 2.067
R11595 a_2458_6128.n60 a_2458_6128.t89 2.067
R11596 a_2458_6128.n45 a_2458_6128.t174 2.067
R11597 a_2458_6128.n44 a_2458_6128.t83 2.067
R11598 a_2458_6128.n132 a_2458_6128.t74 2.067
R11599 a_2458_6128.n133 a_2458_6128.t72 2.067
R11600 a_2458_6128.n49 a_2458_6128.t75 2.067
R11601 a_2458_6128.n48 a_2458_6128.t5 2.067
R11602 a_2458_6128.n47 a_2458_6128.t62 2.067
R11603 a_2458_6128.n46 a_2458_6128.t78 2.067
R11604 a_2458_6128.n51 a_2458_6128.t182 2.067
R11605 a_2458_6128.n50 a_2458_6128.t68 2.067
R11606 a_2458_6128.n128 a_2458_6128.t176 2.067
R11607 a_2458_6128.n129 a_2458_6128.t192 2.067
R11608 a_2458_6128.n53 a_2458_6128.t181 2.067
R11609 a_2458_6128.n52 a_2458_6128.t93 2.067
R11610 a_2458_6128.n125 a_2458_6128.t69 2.067
R11611 a_2458_6128.n126 a_2458_6128.t183 2.067
R11612 a_2458_6128.n57 a_2458_6128.t82 2.067
R11613 a_2458_6128.n56 a_2458_6128.t85 2.067
R11614 a_2458_6128.n55 a_2458_6128.t88 2.067
R11615 a_2458_6128.n54 a_2458_6128.t70 2.067
R11616 a_2458_6128.n59 a_2458_6128.t73 2.067
R11617 a_2458_6128.n58 a_2458_6128.t71 2.067
R11618 a_2458_6128.n121 a_2458_6128.t84 2.067
R11619 a_2458_6128.n122 a_2458_6128.t90 2.067
R11620 a_2458_6128.n154 a_2458_6128.n153 1.777
R11621 a_2458_6128.n155 a_2458_6128.n152 1.777
R11622 a_2458_6128.n156 a_2458_6128.n151 1.777
R11623 a_2458_6128.n69 a_2458_6128.n45 1.615
R11624 a_2458_6128.n67 a_2458_6128.n51 1.615
R11625 a_2458_6128.n66 a_2458_6128.n53 1.615
R11626 a_2458_6128.n64 a_2458_6128.n59 1.615
R11627 a_2458_6128.n61 a_2458_6128.n60 1.352
R11628 a_2458_6128.n62 a_2458_6128.n61 1.352
R11629 a_2458_6128.n63 a_2458_6128.n62 1.352
R11630 a_2458_6128.n133 a_2458_6128.n132 1.352
R11631 a_2458_6128.n45 a_2458_6128.n44 1.352
R11632 a_2458_6128.n47 a_2458_6128.n46 1.352
R11633 a_2458_6128.n48 a_2458_6128.n47 1.352
R11634 a_2458_6128.n49 a_2458_6128.n48 1.352
R11635 a_2458_6128.n129 a_2458_6128.n128 1.352
R11636 a_2458_6128.n51 a_2458_6128.n50 1.352
R11637 a_2458_6128.n126 a_2458_6128.n125 1.352
R11638 a_2458_6128.n53 a_2458_6128.n52 1.352
R11639 a_2458_6128.n55 a_2458_6128.n54 1.352
R11640 a_2458_6128.n56 a_2458_6128.n55 1.352
R11641 a_2458_6128.n57 a_2458_6128.n56 1.352
R11642 a_2458_6128.n122 a_2458_6128.n121 1.352
R11643 a_2458_6128.n59 a_2458_6128.n58 1.352
R11644 a_2458_6128.n73 a_2458_6128.n72 1.352
R11645 a_2458_6128.n72 a_2458_6128.n71 1.352
R11646 a_2458_6128.n71 a_2458_6128.n70 1.352
R11647 a_2458_6128.n134 a_2458_6128.n133 1.303
R11648 a_2458_6128.n130 a_2458_6128.n129 1.303
R11649 a_2458_6128.n127 a_2458_6128.n126 1.303
R11650 a_2458_6128.n123 a_2458_6128.n122 1.303
R11651 a_2458_6128.n139 a_2458_6128.n43 1.068
R11652 a_2458_6128.n158 a_2458_6128.n150 1.068
R11653 a_2458_6128.n136 a_2458_6128.n120 1.068
R11654 a_2458_6128.n137 a_2458_6128.n97 1.068
R11655 a_2458_6128.n160 a_2458_6128.n159 1.068
R11656 a_2458_6128.n157 a_2458_6128.n156 1.053
R11657 a_2458_6128.n155 a_2458_6128.n154 0.812
R11658 a_2458_6128.n156 a_2458_6128.n155 0.796
R11659 a_2458_6128.n159 a_2458_6128.n158 0.752
R11660 a_2458_6128.n159 a_2458_6128.n139 0.752
R11661 a_2458_6128.n137 a_2458_6128.n136 0.752
R11662 a_2458_6128.n165 a_2458_6128.n8 0.54
R11663 a_2458_6128.n164 a_2458_6128.n12 0.54
R11664 a_2458_6128.n163 a_2458_6128.n14 0.54
R11665 a_2458_6128.n162 a_2458_6128.n16 0.54
R11666 a_2458_6128.n161 a_2458_6128.n18 0.54
R11667 a_2458_6128.n160 a_2458_6128.n20 0.54
R11668 a_2458_6128.n43 a_2458_6128.n22 0.54
R11669 a_2458_6128.n42 a_2458_6128.n24 0.54
R11670 a_2458_6128.n41 a_2458_6128.n26 0.54
R11671 a_2458_6128.n40 a_2458_6128.n28 0.54
R11672 a_2458_6128.n39 a_2458_6128.n30 0.54
R11673 a_2458_6128.n38 a_2458_6128.n32 0.54
R11674 a_2458_6128.n37 a_2458_6128.n34 0.54
R11675 a_2458_6128.n150 a_2458_6128.n141 0.54
R11676 a_2458_6128.n149 a_2458_6128.n143 0.54
R11677 a_2458_6128.n148 a_2458_6128.n145 0.54
R11678 a_2458_6128.n120 a_2458_6128.n99 0.54
R11679 a_2458_6128.n119 a_2458_6128.n101 0.54
R11680 a_2458_6128.n118 a_2458_6128.n103 0.54
R11681 a_2458_6128.n117 a_2458_6128.n105 0.54
R11682 a_2458_6128.n116 a_2458_6128.n107 0.54
R11683 a_2458_6128.n115 a_2458_6128.n109 0.54
R11684 a_2458_6128.n114 a_2458_6128.n111 0.54
R11685 a_2458_6128.n97 a_2458_6128.n76 0.54
R11686 a_2458_6128.n96 a_2458_6128.n78 0.54
R11687 a_2458_6128.n95 a_2458_6128.n80 0.54
R11688 a_2458_6128.n94 a_2458_6128.n82 0.54
R11689 a_2458_6128.n93 a_2458_6128.n84 0.54
R11690 a_2458_6128.n92 a_2458_6128.n86 0.54
R11691 a_2458_6128.n91 a_2458_6128.n88 0.54
R11692 a_2458_6128.n4 a_2458_6128.n3 0.54
R11693 a_2458_6128.n168 a_2458_6128.n167 0.54
R11694 a_2458_6128.n170 a_2458_6128.n169 0.464
R11695 a_2458_6128.n6 a_2458_6128.n5 0.464
R11696 a_2458_6128.n8 a_2458_6128.n7 0.464
R11697 a_2458_6128.n10 a_2458_6128.n9 0.464
R11698 a_2458_6128.n12 a_2458_6128.n11 0.464
R11699 a_2458_6128.n14 a_2458_6128.n13 0.464
R11700 a_2458_6128.n16 a_2458_6128.n15 0.464
R11701 a_2458_6128.n18 a_2458_6128.n17 0.464
R11702 a_2458_6128.n20 a_2458_6128.n19 0.464
R11703 a_2458_6128.n22 a_2458_6128.n21 0.464
R11704 a_2458_6128.n24 a_2458_6128.n23 0.464
R11705 a_2458_6128.n26 a_2458_6128.n25 0.464
R11706 a_2458_6128.n28 a_2458_6128.n27 0.464
R11707 a_2458_6128.n30 a_2458_6128.n29 0.464
R11708 a_2458_6128.n32 a_2458_6128.n31 0.464
R11709 a_2458_6128.n34 a_2458_6128.n33 0.464
R11710 a_2458_6128.n36 a_2458_6128.n35 0.464
R11711 a_2458_6128.n141 a_2458_6128.n140 0.464
R11712 a_2458_6128.n143 a_2458_6128.n142 0.464
R11713 a_2458_6128.n145 a_2458_6128.n144 0.464
R11714 a_2458_6128.n147 a_2458_6128.n146 0.464
R11715 a_2458_6128.n99 a_2458_6128.n98 0.464
R11716 a_2458_6128.n101 a_2458_6128.n100 0.464
R11717 a_2458_6128.n103 a_2458_6128.n102 0.464
R11718 a_2458_6128.n105 a_2458_6128.n104 0.464
R11719 a_2458_6128.n107 a_2458_6128.n106 0.464
R11720 a_2458_6128.n109 a_2458_6128.n108 0.464
R11721 a_2458_6128.n111 a_2458_6128.n110 0.464
R11722 a_2458_6128.n113 a_2458_6128.n112 0.464
R11723 a_2458_6128.n76 a_2458_6128.n75 0.464
R11724 a_2458_6128.n78 a_2458_6128.n77 0.464
R11725 a_2458_6128.n80 a_2458_6128.n79 0.464
R11726 a_2458_6128.n82 a_2458_6128.n81 0.464
R11727 a_2458_6128.n84 a_2458_6128.n83 0.464
R11728 a_2458_6128.n86 a_2458_6128.n85 0.464
R11729 a_2458_6128.n88 a_2458_6128.n87 0.464
R11730 a_2458_6128.n90 a_2458_6128.n89 0.464
R11731 a_2458_6128.n1 a_2458_6128.n0 0.464
R11732 a_2458_6128.n3 a_2458_6128.n2 0.464
R11733 a_2458_6128.n167 a_2458_6128.n166 0.464
R11734 a_2458_6128.n138 a_2458_6128.n137 0.401
R11735 a_2458_6128.n139 a_2458_6128.n138 0.35
R11736 a_2458_6128.n165 a_2458_6128.n6 0.277
R11737 a_2458_6128.n164 a_2458_6128.n10 0.277
R11738 a_2458_6128.n4 a_2458_6128.n1 0.277
R11739 a_2458_6128.n170 a_2458_6128.n168 0.277
R11740 a_2458_6128.n65 a_2458_6128.n64 0.188
R11741 a_2458_6128.n66 a_2458_6128.n65 0.188
R11742 a_2458_6128.n67 a_2458_6128.n66 0.188
R11743 a_2458_6128.n68 a_2458_6128.n67 0.188
R11744 a_2458_6128.n69 a_2458_6128.n68 0.188
R11745 a_2458_6128.n74 a_2458_6128.n69 0.188
R11746 a_2458_6128.n124 a_2458_6128.n123 0.188
R11747 a_2458_6128.n127 a_2458_6128.n124 0.188
R11748 a_2458_6128.n130 a_2458_6128.n127 0.188
R11749 a_2458_6128.n131 a_2458_6128.n130 0.188
R11750 a_2458_6128.n134 a_2458_6128.n131 0.188
R11751 a_2458_6128.n135 a_2458_6128.n134 0.188
R11752 Vop.n40 Vop.t120 57.198
R11753 Vop.n64 Vop.t14 14.623
R11754 Vop.n65 Vop.t55 14.623
R11755 Vop.n66 Vop.t15 14.623
R11756 Vop.n67 Vop.t49 14.623
R11757 Vop.n68 Vop.t11 14.623
R11758 Vop.n69 Vop.t45 14.623
R11759 Vop.n70 Vop.t9 14.623
R11760 Vop.n71 Vop.t2 14.623
R11761 Vop.n96 Vop.t6 14.598
R11762 Vop.n95 Vop.t18 14.598
R11763 Vop.n33 Vop.t31 14.598
R11764 Vop.n34 Vop.t66 14.598
R11765 Vop.n35 Vop.t21 14.598
R11766 Vop.n36 Vop.t62 14.598
R11767 Vop.n42 Vop.t5 14.598
R11768 Vop.n43 Vop.t43 14.598
R11769 Vop.n44 Vop.t7 14.598
R11770 Vop.n45 Vop.t41 14.598
R11771 Vop.n46 Vop.t3 14.598
R11772 Vop.n47 Vop.t34 14.598
R11773 Vop.n48 Vop.t73 14.598
R11774 Vop.n49 Vop.t63 14.598
R11775 Vop.n0 Vop.t39 14.598
R11776 Vop.n1 Vop.t35 14.598
R11777 Vop.n2 Vop.t74 14.598
R11778 Vop.n3 Vop.t29 14.598
R11779 Vop.n4 Vop.t64 14.598
R11780 Vop.n5 Vop.t67 14.598
R11781 Vop.n6 Vop.t20 14.598
R11782 Vop.n7 Vop.t22 14.598
R11783 Vop.n8 Vop.t53 14.598
R11784 Vop.n9 Vop.t58 14.598
R11785 Vop.n10 Vop.t47 14.598
R11786 Vop.n11 Vop.t48 14.598
R11787 Vop.n97 Vop.t1 14.598
R11788 Vop.n98 Vop.t30 14.598
R11789 Vop.n99 Vop.t69 14.598
R11790 Vop.n100 Vop.t24 14.598
R11791 Vop.n101 Vop.t19 14.598
R11792 Vop.n106 Vop.t36 14.598
R11793 Vop.n96 Vop.t38 13.849
R11794 Vop.n95 Vop.t76 13.849
R11795 Vop.n33 Vop.t4 13.849
R11796 Vop.n34 Vop.t57 13.849
R11797 Vop.n35 Vop.t16 13.849
R11798 Vop.n36 Vop.t50 13.849
R11799 Vop.n64 Vop.t54 13.849
R11800 Vop.n65 Vop.t46 13.849
R11801 Vop.n66 Vop.t10 13.849
R11802 Vop.n67 Vop.t44 13.849
R11803 Vop.n68 Vop.t8 13.849
R11804 Vop.n69 Vop.t40 13.849
R11805 Vop.n70 Vop.t0 13.849
R11806 Vop.n71 Vop.t70 13.849
R11807 Vop.n42 Vop.t42 13.849
R11808 Vop.n43 Vop.t37 13.849
R11809 Vop.n44 Vop.t78 13.849
R11810 Vop.n45 Vop.t32 13.849
R11811 Vop.n46 Vop.t71 13.849
R11812 Vop.n47 Vop.t25 13.849
R11813 Vop.n48 Vop.t60 13.849
R11814 Vop.n49 Vop.t51 13.849
R11815 Vop.n0 Vop.t13 13.849
R11816 Vop.n1 Vop.t75 13.849
R11817 Vop.n2 Vop.t27 13.849
R11818 Vop.n3 Vop.t68 13.849
R11819 Vop.n4 Vop.t77 13.849
R11820 Vop.n5 Vop.t23 13.849
R11821 Vop.n6 Vop.t28 13.849
R11822 Vop.n7 Vop.t59 13.849
R11823 Vop.n8 Vop.t65 13.849
R11824 Vop.n9 Vop.t17 13.849
R11825 Vop.n10 Vop.t56 13.849
R11826 Vop.n11 Vop.t12 13.849
R11827 Vop.n97 Vop.t33 13.849
R11828 Vop.n98 Vop.t72 13.849
R11829 Vop.n99 Vop.t26 13.849
R11830 Vop.n100 Vop.t61 13.849
R11831 Vop.n101 Vop.t52 13.849
R11832 Vop.n106 Vop.t79 13.849
R11833 Vop.n30 Vop.t97 8.857
R11834 Vop.n31 Vop.t111 8.857
R11835 Vop.n79 Vop.t88 8.857
R11836 Vop.n80 Vop.t92 8.857
R11837 Vop.n81 Vop.t81 8.857
R11838 Vop.n82 Vop.t86 8.857
R11839 Vop.n57 Vop.t113 8.857
R11840 Vop.n58 Vop.t108 8.857
R11841 Vop.n59 Vop.t114 8.857
R11842 Vop.n60 Vop.t119 8.857
R11843 Vop.n20 Vop.t106 8.857
R11844 Vop.n21 Vop.t115 8.857
R11845 Vop.n22 Vop.t85 8.857
R11846 Vop.n24 Vop.t102 8.857
R11847 Vop.n25 Vop.t94 8.857
R11848 Vop.n88 Vop.t82 8.857
R11849 Vop.n89 Vop.t101 8.857
R11850 Vop.n90 Vop.t83 8.857
R11851 Vop.n91 Vop.t98 8.857
R11852 Vop.n23 Vop.t107 8.8
R11853 Vop.n30 Vop.t105 8.266
R11854 Vop.n31 Vop.t96 8.266
R11855 Vop.n79 Vop.t80 8.266
R11856 Vop.n80 Vop.t87 8.266
R11857 Vop.n81 Vop.t91 8.266
R11858 Vop.n82 Vop.t90 8.266
R11859 Vop.n57 Vop.t99 8.266
R11860 Vop.n58 Vop.t112 8.266
R11861 Vop.n59 Vop.t100 8.266
R11862 Vop.n60 Vop.t89 8.266
R11863 Vop.n20 Vop.t116 8.266
R11864 Vop.n21 Vop.t109 8.266
R11865 Vop.n22 Vop.t110 8.266
R11866 Vop.n23 Vop.t118 8.266
R11867 Vop.n24 Vop.t93 8.266
R11868 Vop.n25 Vop.t117 8.266
R11869 Vop.n88 Vop.t103 8.266
R11870 Vop.n89 Vop.t84 8.266
R11871 Vop.n90 Vop.t104 8.266
R11872 Vop.n91 Vop.t95 8.266
R11873 Vop.n72 Vop.n71 2.632
R11874 Vop.n37 Vop.n36 2.609
R11875 Vop.n50 Vop.n49 2.609
R11876 Vop.n102 Vop.n101 2.609
R11877 Vop.n32 Vop.n31 2.597
R11878 Vop.n83 Vop.n82 2.597
R11879 Vop.n61 Vop.n60 2.597
R11880 Vop.n92 Vop.n91 2.597
R11881 Vop.n41 Vop.n29 2.529
R11882 Vop.n40 Vop.n32 2.528
R11883 Vop.n86 Vop.n85 2.528
R11884 Vop.n87 Vop.n63 2.528
R11885 Vop.n110 Vop.n94 2.528
R11886 Vop.n29 Vop.n28 2.221
R11887 Vop.n28 Vop.n27 2.22
R11888 Vop.n84 Vop.n83 2.219
R11889 Vop.n85 Vop.n84 2.219
R11890 Vop.n62 Vop.n61 2.219
R11891 Vop.n63 Vop.n62 2.219
R11892 Vop.n27 Vop.n26 2.219
R11893 Vop.n93 Vop.n92 2.219
R11894 Vop.n94 Vop.n93 2.219
R11895 Vop.n38 Vop.n37 2.199
R11896 Vop.n39 Vop.n38 2.199
R11897 Vop.n73 Vop.n72 2.199
R11898 Vop.n74 Vop.n73 2.199
R11899 Vop.n75 Vop.n74 2.199
R11900 Vop.n76 Vop.n75 2.199
R11901 Vop.n77 Vop.n76 2.199
R11902 Vop.n78 Vop.n77 2.199
R11903 Vop.n51 Vop.n50 2.199
R11904 Vop.n52 Vop.n51 2.199
R11905 Vop.n53 Vop.n52 2.199
R11906 Vop.n54 Vop.n53 2.199
R11907 Vop.n55 Vop.n54 2.199
R11908 Vop.n56 Vop.n55 2.199
R11909 Vop.n13 Vop.n12 2.199
R11910 Vop.n14 Vop.n13 2.199
R11911 Vop.n15 Vop.n14 2.199
R11912 Vop.n16 Vop.n15 2.199
R11913 Vop.n17 Vop.n16 2.199
R11914 Vop.n18 Vop.n17 2.199
R11915 Vop.n19 Vop.n18 2.199
R11916 Vop.n109 Vop.n108 2.199
R11917 Vop.n108 Vop.n107 2.199
R11918 Vop.n103 Vop.n102 2.199
R11919 Vop.n104 Vop.n103 2.199
R11920 Vop.n105 Vop.n104 2.199
R11921 Vop.n107 Vop.n105 2.199
R11922 Vop.n40 Vop.n39 1.506
R11923 Vop.n86 Vop.n78 1.506
R11924 Vop.n87 Vop.n56 1.506
R11925 Vop.n41 Vop.n19 1.506
R11926 Vop.n110 Vop.n109 1.506
R11927 Vop.n110 Vop.n87 0.752
R11928 Vop.n87 Vop.n86 0.752
R11929 Vop.n41 Vop.n40 0.72
R11930 Vop.n15 Vop.n4 0.697
R11931 Vop.n14 Vop.n6 0.697
R11932 Vop.n13 Vop.n8 0.697
R11933 Vop.n12 Vop.n10 0.697
R11934 Vop.n26 Vop.n24 0.591
R11935 Vop.n27 Vop.n22 0.581
R11936 Vop Vop.n110 0.487
R11937 Vop.n78 Vop.n64 0.433
R11938 Vop.n77 Vop.n65 0.433
R11939 Vop.n76 Vop.n66 0.433
R11940 Vop.n75 Vop.n67 0.433
R11941 Vop.n74 Vop.n68 0.433
R11942 Vop.n73 Vop.n69 0.433
R11943 Vop.n72 Vop.n70 0.433
R11944 Vop.n108 Vop.n96 0.41
R11945 Vop.n109 Vop.n95 0.41
R11946 Vop.n39 Vop.n33 0.41
R11947 Vop.n38 Vop.n34 0.41
R11948 Vop.n37 Vop.n35 0.41
R11949 Vop.n56 Vop.n42 0.41
R11950 Vop.n55 Vop.n43 0.41
R11951 Vop.n54 Vop.n44 0.41
R11952 Vop.n53 Vop.n45 0.41
R11953 Vop.n52 Vop.n46 0.41
R11954 Vop.n51 Vop.n47 0.41
R11955 Vop.n50 Vop.n48 0.41
R11956 Vop.n19 Vop.n0 0.41
R11957 Vop.n18 Vop.n1 0.41
R11958 Vop.n17 Vop.n2 0.41
R11959 Vop.n16 Vop.n3 0.41
R11960 Vop.n15 Vop.n5 0.41
R11961 Vop.n14 Vop.n7 0.41
R11962 Vop.n13 Vop.n9 0.41
R11963 Vop.n12 Vop.n11 0.41
R11964 Vop.n105 Vop.n97 0.41
R11965 Vop.n104 Vop.n98 0.41
R11966 Vop.n103 Vop.n99 0.41
R11967 Vop.n102 Vop.n100 0.41
R11968 Vop.n107 Vop.n106 0.41
R11969 Vop.n32 Vop.n30 0.378
R11970 Vop.n85 Vop.n79 0.378
R11971 Vop.n84 Vop.n80 0.378
R11972 Vop.n83 Vop.n81 0.378
R11973 Vop.n63 Vop.n57 0.378
R11974 Vop.n62 Vop.n58 0.378
R11975 Vop.n61 Vop.n59 0.378
R11976 Vop.n29 Vop.n20 0.378
R11977 Vop.n28 Vop.n21 0.378
R11978 Vop.n26 Vop.n25 0.378
R11979 Vop.n94 Vop.n88 0.378
R11980 Vop.n93 Vop.n89 0.378
R11981 Vop.n92 Vop.n90 0.378
R11982 Vop.n27 Vop.n23 0.338
R11983 Vop Vop.n41 0.264
R11984 Vxp.n45 Vxp.t116 14.528
R11985 Vxp.n42 Vxp.t75 14.528
R11986 Vxp.n39 Vxp.t128 14.528
R11987 Vxp.n36 Vxp.t85 14.528
R11988 Vxp.n33 Vxp.t132 14.528
R11989 Vxp.n30 Vxp.t87 14.528
R11990 Vxp.n48 Vxp.t105 14.528
R11991 Vxp.n27 Vxp.t42 14.528
R11992 Vxp.n54 Vxp.t68 13.849
R11993 Vxp.n28 Vxp.t93 13.849
R11994 Vxp.n145 Vxp.t99 13.849
R11995 Vxp.n164 Vxp.t45 13.849
R11996 Vxp.n163 Vxp.t79 13.849
R11997 Vxp.n197 Vxp.t100 13.849
R11998 Vxp.n196 Vxp.t133 13.849
R11999 Vxp.n80 Vxp.t81 13.849
R12000 Vxp.n78 Vxp.t135 13.849
R12001 Vxp.n74 Vxp.t48 13.849
R12002 Vxp.n52 Vxp.t130 13.849
R12003 Vxp.n82 Vxp.t117 13.849
R12004 Vxp.n83 Vxp.t83 13.849
R12005 Vxp.n199 Vxp.t69 13.849
R12006 Vxp.n200 Vxp.t129 13.849
R12007 Vxp.n166 Vxp.t80 13.849
R12008 Vxp.n161 Vxp.t54 13.849
R12009 Vxp.n158 Vxp.t44 13.849
R12010 Vxp.n162 Vxp.t91 13.849
R12011 Vxp.n208 Vxp.t47 13.849
R12012 Vxp.n186 Vxp.t56 13.849
R12013 Vxp.n181 Vxp.t101 13.849
R12014 Vxp.n182 Vxp.t66 13.849
R12015 Vxp.n156 Vxp.t52 13.849
R12016 Vxp.n187 Vxp.t94 13.849
R12017 Vxp.n98 Vxp.t107 13.849
R12018 Vxp.n97 Vxp.t46 13.849
R12019 Vxp.n71 Vxp.t57 13.849
R12020 Vxp.n70 Vxp.t95 13.849
R12021 Vxp.n46 Vxp.t49 13.849
R12022 Vxp.n45 Vxp.t90 13.849
R12023 Vxp.n188 Vxp.t112 13.849
R12024 Vxp.n178 Vxp.t58 13.849
R12025 Vxp.n179 Vxp.t121 13.849
R12026 Vxp.n154 Vxp.t108 13.849
R12027 Vxp.n189 Vxp.t50 13.849
R12028 Vxp.n95 Vxp.t64 13.849
R12029 Vxp.n94 Vxp.t98 13.849
R12030 Vxp.n68 Vxp.t113 13.849
R12031 Vxp.n67 Vxp.t51 13.849
R12032 Vxp.n43 Vxp.t103 13.849
R12033 Vxp.n42 Vxp.t43 13.849
R12034 Vxp.n190 Vxp.t71 13.849
R12035 Vxp.n175 Vxp.t114 13.849
R12036 Vxp.n176 Vxp.t82 13.849
R12037 Vxp.n152 Vxp.t65 13.849
R12038 Vxp.n191 Vxp.t104 13.849
R12039 Vxp.n92 Vxp.t118 13.849
R12040 Vxp.n91 Vxp.t55 13.849
R12041 Vxp.n65 Vxp.t72 13.849
R12042 Vxp.n64 Vxp.t106 13.849
R12043 Vxp.n40 Vxp.t60 13.849
R12044 Vxp.n39 Vxp.t97 13.849
R12045 Vxp.n192 Vxp.t124 13.849
R12046 Vxp.n172 Vxp.t74 13.849
R12047 Vxp.n173 Vxp.t131 13.849
R12048 Vxp.n150 Vxp.t120 13.849
R12049 Vxp.n193 Vxp.t62 13.849
R12050 Vxp.n89 Vxp.t78 13.849
R12051 Vxp.n88 Vxp.t111 13.849
R12052 Vxp.n62 Vxp.t125 13.849
R12053 Vxp.n61 Vxp.t63 13.849
R12054 Vxp.n37 Vxp.t115 13.849
R12055 Vxp.n36 Vxp.t53 13.849
R12056 Vxp.n194 Vxp.t76 13.849
R12057 Vxp.n169 Vxp.t119 13.849
R12058 Vxp.n170 Vxp.t84 13.849
R12059 Vxp.n148 Vxp.t73 13.849
R12060 Vxp.n195 Vxp.t109 13.849
R12061 Vxp.n86 Vxp.t123 13.849
R12062 Vxp.n85 Vxp.t61 13.849
R12063 Vxp.n59 Vxp.t77 13.849
R12064 Vxp.n58 Vxp.t110 13.849
R12065 Vxp.n34 Vxp.t67 13.849
R12066 Vxp.n33 Vxp.t102 13.849
R12067 Vxp.n207 Vxp.t88 13.849
R12068 Vxp.n77 Vxp.t96 13.849
R12069 Vxp.n167 Vxp.t134 13.849
R12070 Vxp.n146 Vxp.t127 13.849
R12071 Vxp.n53 Vxp.t70 13.849
R12072 Vxp.n31 Vxp.t122 13.849
R12073 Vxp.n30 Vxp.t59 13.849
R12074 Vxp.n73 Vxp.t89 13.849
R12075 Vxp.n49 Vxp.t41 13.849
R12076 Vxp.n48 Vxp.t86 13.849
R12077 Vxp.n79 Vxp.t92 13.849
R12078 Vxp.n27 Vxp.t126 13.849
R12079 Vxp.n55 Vxp.t136 13.849
R12080 Vxp.n106 Vxp.t140 3.473
R12081 Vxp.n105 Vxp.t29 3.473
R12082 Vxp.n104 Vxp.t23 3.473
R12083 Vxp.n103 Vxp.t12 3.473
R12084 Vxp.n102 Vxp.t24 3.473
R12085 Vxp.n17 Vxp.t21 3.473
R12086 Vxp.n18 Vxp.t37 3.473
R12087 Vxp.n19 Vxp.t5 3.473
R12088 Vxp.n16 Vxp.t7 3.473
R12089 Vxp.n15 Vxp.t20 3.473
R12090 Vxp.n14 Vxp.t34 3.473
R12091 Vxp.n107 Vxp.t15 3.473
R12092 Vxp.n108 Vxp.t27 3.473
R12093 Vxp.n109 Vxp.t14 3.473
R12094 Vxp.n110 Vxp.t0 3.473
R12095 Vxp.n111 Vxp.t148 3.473
R12096 Vxp.n13 Vxp.t138 3.473
R12097 Vxp.n12 Vxp.t139 3.473
R12098 Vxp.n113 Vxp.t150 3.473
R12099 Vxp.n114 Vxp.t30 3.473
R12100 Vxp.n115 Vxp.t11 3.473
R12101 Vxp.n116 Vxp.t32 3.473
R12102 Vxp.n11 Vxp.t40 3.473
R12103 Vxp.n10 Vxp.t6 3.473
R12104 Vxp.n118 Vxp.t143 3.473
R12105 Vxp.n119 Vxp.t17 3.473
R12106 Vxp.n120 Vxp.t142 3.473
R12107 Vxp.n121 Vxp.t151 3.473
R12108 Vxp.n9 Vxp.t16 3.473
R12109 Vxp.n8 Vxp.t18 3.473
R12110 Vxp.n123 Vxp.t1 3.473
R12111 Vxp.n124 Vxp.t31 3.473
R12112 Vxp.n125 Vxp.t8 3.473
R12113 Vxp.n126 Vxp.t26 3.473
R12114 Vxp.n7 Vxp.t149 3.473
R12115 Vxp.n6 Vxp.t13 3.473
R12116 Vxp.n128 Vxp.t4 3.473
R12117 Vxp.n129 Vxp.t35 3.473
R12118 Vxp.n130 Vxp.t3 3.473
R12119 Vxp.n131 Vxp.t147 3.473
R12120 Vxp.n5 Vxp.t36 3.473
R12121 Vxp.n4 Vxp.t25 3.473
R12122 Vxp.n3 Vxp.t22 3.473
R12123 Vxp.n133 Vxp.t137 3.473
R12124 Vxp.n134 Vxp.t145 3.473
R12125 Vxp.n135 Vxp.t33 3.473
R12126 Vxp.n136 Vxp.t19 3.473
R12127 Vxp.n137 Vxp.t10 3.473
R12128 Vxp.n2 Vxp.t146 3.473
R12129 Vxp.n1 Vxp.t2 3.473
R12130 Vxp.n0 Vxp.t28 3.473
R12131 Vxp.n139 Vxp.t39 3.473
R12132 Vxp.n140 Vxp.t9 3.473
R12133 Vxp.n141 Vxp.t38 3.473
R12134 Vxp.n142 Vxp.t144 3.473
R12135 Vxp.n143 Vxp.t141 3.473
R12136 Vxp.n160 Vxp.n159 3.311
R12137 Vxp.n210 Vxp.n209 3.206
R12138 Vxp.n185 Vxp.n184 3.206
R12139 Vxp.n76 Vxp.n75 3.206
R12140 Vxp.n101 Vxp.n100 3.206
R12141 Vxp.n51 Vxp.n50 3.206
R12142 Vxp.n51 Vxp.n26 2.969
R12143 Vxp.n147 Vxp.n145 2.849
R12144 Vxp.n117 Vxp.n116 2.66
R12145 Vxp.n21 Vxp.n13 2.66
R12146 Vxp.n122 Vxp.n121 2.66
R12147 Vxp.n22 Vxp.n11 2.66
R12148 Vxp.n127 Vxp.n126 2.66
R12149 Vxp.n23 Vxp.n9 2.66
R12150 Vxp.n132 Vxp.n131 2.66
R12151 Vxp.n24 Vxp.n7 2.66
R12152 Vxp.n168 Vxp.n165 2.199
R12153 Vxp.n201 Vxp.n198 2.199
R12154 Vxp.n202 Vxp.n201 2.199
R12155 Vxp.n203 Vxp.n202 2.199
R12156 Vxp.n204 Vxp.n203 2.199
R12157 Vxp.n205 Vxp.n204 2.199
R12158 Vxp.n206 Vxp.n205 2.199
R12159 Vxp.n209 Vxp.n206 2.199
R12160 Vxp.n184 Vxp.n183 2.199
R12161 Vxp.n183 Vxp.n180 2.199
R12162 Vxp.n180 Vxp.n177 2.199
R12163 Vxp.n177 Vxp.n174 2.199
R12164 Vxp.n174 Vxp.n171 2.199
R12165 Vxp.n171 Vxp.n168 2.199
R12166 Vxp.n57 Vxp.n56 2.199
R12167 Vxp.n60 Vxp.n57 2.199
R12168 Vxp.n63 Vxp.n60 2.199
R12169 Vxp.n66 Vxp.n63 2.199
R12170 Vxp.n69 Vxp.n66 2.199
R12171 Vxp.n72 Vxp.n69 2.199
R12172 Vxp.n75 Vxp.n72 2.199
R12173 Vxp.n100 Vxp.n99 2.199
R12174 Vxp.n99 Vxp.n96 2.199
R12175 Vxp.n96 Vxp.n93 2.199
R12176 Vxp.n93 Vxp.n90 2.199
R12177 Vxp.n90 Vxp.n87 2.199
R12178 Vxp.n87 Vxp.n84 2.199
R12179 Vxp.n84 Vxp.n81 2.199
R12180 Vxp.n149 Vxp.n147 2.199
R12181 Vxp.n151 Vxp.n149 2.199
R12182 Vxp.n153 Vxp.n151 2.199
R12183 Vxp.n155 Vxp.n153 2.199
R12184 Vxp.n157 Vxp.n155 2.199
R12185 Vxp.n159 Vxp.n157 2.199
R12186 Vxp.n50 Vxp.n47 2.199
R12187 Vxp.n47 Vxp.n44 2.199
R12188 Vxp.n44 Vxp.n41 2.199
R12189 Vxp.n41 Vxp.n38 2.199
R12190 Vxp.n38 Vxp.n35 2.199
R12191 Vxp.n35 Vxp.n32 2.199
R12192 Vxp.n32 Vxp.n29 2.199
R12193 Vxp.n111 Vxp.n110 1.246
R12194 Vxp.n110 Vxp.n109 1.246
R12195 Vxp.n109 Vxp.n108 1.246
R12196 Vxp.n108 Vxp.n107 1.246
R12197 Vxp.n15 Vxp.n14 1.246
R12198 Vxp.n16 Vxp.n15 1.246
R12199 Vxp.n116 Vxp.n115 1.246
R12200 Vxp.n115 Vxp.n114 1.246
R12201 Vxp.n114 Vxp.n113 1.246
R12202 Vxp.n13 Vxp.n12 1.246
R12203 Vxp.n121 Vxp.n120 1.246
R12204 Vxp.n120 Vxp.n119 1.246
R12205 Vxp.n119 Vxp.n118 1.246
R12206 Vxp.n11 Vxp.n10 1.246
R12207 Vxp.n126 Vxp.n125 1.246
R12208 Vxp.n125 Vxp.n124 1.246
R12209 Vxp.n124 Vxp.n123 1.246
R12210 Vxp.n9 Vxp.n8 1.246
R12211 Vxp.n131 Vxp.n130 1.246
R12212 Vxp.n130 Vxp.n129 1.246
R12213 Vxp.n129 Vxp.n128 1.246
R12214 Vxp.n7 Vxp.n6 1.246
R12215 Vxp.n137 Vxp.n136 1.246
R12216 Vxp.n136 Vxp.n135 1.246
R12217 Vxp.n135 Vxp.n134 1.246
R12218 Vxp.n134 Vxp.n133 1.246
R12219 Vxp.n4 Vxp.n3 1.246
R12220 Vxp.n5 Vxp.n4 1.246
R12221 Vxp.n143 Vxp.n142 1.246
R12222 Vxp.n142 Vxp.n141 1.246
R12223 Vxp.n141 Vxp.n140 1.246
R12224 Vxp.n140 Vxp.n139 1.246
R12225 Vxp.n1 Vxp.n0 1.246
R12226 Vxp.n2 Vxp.n1 1.246
R12227 Vxp.n19 Vxp.n18 1.246
R12228 Vxp.n18 Vxp.n17 1.246
R12229 Vxp.n103 Vxp.n102 1.246
R12230 Vxp.n104 Vxp.n103 1.246
R12231 Vxp.n105 Vxp.n104 1.246
R12232 Vxp.n106 Vxp.n105 1.246
R12233 Vxp.n20 Vxp.n16 1.124
R12234 Vxp.n112 Vxp.n111 1.124
R12235 Vxp.n138 Vxp.n137 0.936
R12236 Vxp.n25 Vxp.n5 0.936
R12237 Vxp.n144 Vxp.n143 0.936
R12238 Vxp.n26 Vxp.n2 0.936
R12239 Vxp.n20 Vxp.n19 0.936
R12240 Vxp.n112 Vxp.n106 0.936
R12241 Vxp.n159 Vxp.n158 0.65
R12242 Vxp.n157 Vxp.n156 0.65
R12243 Vxp.n183 Vxp.n181 0.65
R12244 Vxp.n47 Vxp.n45 0.65
R12245 Vxp.n72 Vxp.n70 0.65
R12246 Vxp.n99 Vxp.n97 0.65
R12247 Vxp.n206 Vxp.n187 0.65
R12248 Vxp.n155 Vxp.n154 0.65
R12249 Vxp.n180 Vxp.n178 0.65
R12250 Vxp.n44 Vxp.n42 0.65
R12251 Vxp.n69 Vxp.n67 0.65
R12252 Vxp.n96 Vxp.n94 0.65
R12253 Vxp.n205 Vxp.n189 0.65
R12254 Vxp.n153 Vxp.n152 0.65
R12255 Vxp.n177 Vxp.n175 0.65
R12256 Vxp.n41 Vxp.n39 0.65
R12257 Vxp.n66 Vxp.n64 0.65
R12258 Vxp.n93 Vxp.n91 0.65
R12259 Vxp.n204 Vxp.n191 0.65
R12260 Vxp.n151 Vxp.n150 0.65
R12261 Vxp.n174 Vxp.n172 0.65
R12262 Vxp.n38 Vxp.n36 0.65
R12263 Vxp.n63 Vxp.n61 0.65
R12264 Vxp.n90 Vxp.n88 0.65
R12265 Vxp.n203 Vxp.n193 0.65
R12266 Vxp.n149 Vxp.n148 0.65
R12267 Vxp.n171 Vxp.n169 0.65
R12268 Vxp.n35 Vxp.n33 0.65
R12269 Vxp.n60 Vxp.n58 0.65
R12270 Vxp.n87 Vxp.n85 0.65
R12271 Vxp.n202 Vxp.n195 0.65
R12272 Vxp.n209 Vxp.n207 0.65
R12273 Vxp.n184 Vxp.n162 0.65
R12274 Vxp.n147 Vxp.n146 0.65
R12275 Vxp.n168 Vxp.n166 0.65
R12276 Vxp.n201 Vxp.n199 0.65
R12277 Vxp.n84 Vxp.n82 0.65
R12278 Vxp.n32 Vxp.n30 0.65
R12279 Vxp.n57 Vxp.n53 0.65
R12280 Vxp.n50 Vxp.n48 0.65
R12281 Vxp.n75 Vxp.n73 0.65
R12282 Vxp.n100 Vxp.n78 0.65
R12283 Vxp.n81 Vxp.n79 0.65
R12284 Vxp.n198 Vxp.n196 0.65
R12285 Vxp.n165 Vxp.n163 0.65
R12286 Vxp.n29 Vxp.n27 0.65
R12287 Vxp.n56 Vxp.n54 0.65
R12288 Vxp.n160 Vxp.n144 0.401
R12289 Vxp.n184 Vxp.n161 0.387
R12290 Vxp.n183 Vxp.n182 0.387
R12291 Vxp.n206 Vxp.n186 0.387
R12292 Vxp.n47 Vxp.n46 0.387
R12293 Vxp.n72 Vxp.n71 0.387
R12294 Vxp.n99 Vxp.n98 0.387
R12295 Vxp.n180 Vxp.n179 0.387
R12296 Vxp.n205 Vxp.n188 0.387
R12297 Vxp.n44 Vxp.n43 0.387
R12298 Vxp.n69 Vxp.n68 0.387
R12299 Vxp.n96 Vxp.n95 0.387
R12300 Vxp.n177 Vxp.n176 0.387
R12301 Vxp.n204 Vxp.n190 0.387
R12302 Vxp.n41 Vxp.n40 0.387
R12303 Vxp.n66 Vxp.n65 0.387
R12304 Vxp.n93 Vxp.n92 0.387
R12305 Vxp.n174 Vxp.n173 0.387
R12306 Vxp.n203 Vxp.n192 0.387
R12307 Vxp.n38 Vxp.n37 0.387
R12308 Vxp.n63 Vxp.n62 0.387
R12309 Vxp.n90 Vxp.n89 0.387
R12310 Vxp.n171 Vxp.n170 0.387
R12311 Vxp.n202 Vxp.n194 0.387
R12312 Vxp.n35 Vxp.n34 0.387
R12313 Vxp.n60 Vxp.n59 0.387
R12314 Vxp.n87 Vxp.n86 0.387
R12315 Vxp.n100 Vxp.n77 0.387
R12316 Vxp.n209 Vxp.n208 0.387
R12317 Vxp.n168 Vxp.n167 0.387
R12318 Vxp.n201 Vxp.n200 0.387
R12319 Vxp.n84 Vxp.n83 0.387
R12320 Vxp.n57 Vxp.n52 0.387
R12321 Vxp.n32 Vxp.n31 0.387
R12322 Vxp.n50 Vxp.n49 0.387
R12323 Vxp.n75 Vxp.n74 0.387
R12324 Vxp.n81 Vxp.n80 0.387
R12325 Vxp.n198 Vxp.n197 0.387
R12326 Vxp.n165 Vxp.n164 0.387
R12327 Vxp.n29 Vxp.n28 0.387
R12328 Vxp.n56 Vxp.n55 0.387
R12329 Vxp.n76 Vxp.n51 0.376
R12330 Vxp.n101 Vxp.n76 0.376
R12331 Vxp.n210 Vxp.n185 0.376
R12332 Vxp.n185 Vxp.n160 0.27
R12333 Vxp Vxp.n101 0.196
R12334 Vxp.n26 Vxp.n25 0.188
R12335 Vxp.n25 Vxp.n24 0.188
R12336 Vxp.n24 Vxp.n23 0.188
R12337 Vxp.n23 Vxp.n22 0.188
R12338 Vxp.n22 Vxp.n21 0.188
R12339 Vxp.n21 Vxp.n20 0.188
R12340 Vxp.n144 Vxp.n138 0.188
R12341 Vxp.n138 Vxp.n132 0.188
R12342 Vxp.n132 Vxp.n127 0.188
R12343 Vxp.n127 Vxp.n122 0.188
R12344 Vxp.n122 Vxp.n117 0.188
R12345 Vxp.n117 Vxp.n112 0.188
R12346 Vxp Vxp.n210 0.179
R12347 level_shifter_up_8.x_hv.n1 level_shifter_up_8.x_hv.t7 224.138
R12348 level_shifter_up_8.x_hv.n2 level_shifter_up_8.x_hv.t9 224.127
R12349 level_shifter_up_8.x_hv.n0 level_shifter_up_8.x_hv.t4 224.127
R12350 level_shifter_up_8.x_hv.n0 level_shifter_up_8.x_hv.t3 224.124
R12351 level_shifter_up_8.x_hv.n1 level_shifter_up_8.x_hv.t6 223.679
R12352 level_shifter_up_8.x_hv.n2 level_shifter_up_8.x_hv.t1 223.679
R12353 level_shifter_up_8.x_hv.n0 level_shifter_up_8.x_hv.t2 223.679
R12354 level_shifter_up_8.x_hv.n0 level_shifter_up_8.x_hv.t5 223.679
R12355 level_shifter_up_8.x_hv.n3 level_shifter_up_8.x_hv.t8 65.158
R12356 level_shifter_up_8.x_hv.n3 level_shifter_up_8.x_hv.t0 13.87
R12357 level_shifter_up_8.x_hv.n3 level_shifter_up_8.x_hv.n2 8.169
R12358 level_shifter_up_8.x_hv.n2 level_shifter_up_8.x_hv.n0 4.523
R12359 level_shifter_up_8.x_hv level_shifter_up_8.x_hv.n3 0.584
R12360 level_shifter_up_8.x_hv.n2 level_shifter_up_8.x_hv.n1 0.343
R12361 a_33657_n21342.n3 a_33657_n21342.t7 13.849
R12362 a_33657_n21342.n2 a_33657_n21342.t0 13.849
R12363 a_33657_n21342.n2 a_33657_n21342.t4 13.849
R12364 a_33657_n21342.n1 a_33657_n21342.t5 13.849
R12365 a_33657_n21342.n1 a_33657_n21342.t6 13.849
R12366 a_33657_n21342.n0 a_33657_n21342.t1 13.849
R12367 a_33657_n21342.n0 a_33657_n21342.t3 13.849
R12368 a_33657_n21342.t2 a_33657_n21342.n3 13.849
R12369 a_33657_n21342.n3 a_33657_n21342.n2 0.868
R12370 a_33657_n21342.n2 a_33657_n21342.n1 0.464
R12371 a_33657_n21342.n3 a_33657_n21342.n0 0.464
R12372 a_23013_n25097.n0 a_23013_n25097.t13 14.598
R12373 a_23013_n25097.n5 a_23013_n25097.t10 14.598
R12374 a_23013_n25097.n4 a_23013_n25097.t19 13.849
R12375 a_23013_n25097.n3 a_23013_n25097.t17 13.849
R12376 a_23013_n25097.n2 a_23013_n25097.t12 13.849
R12377 a_23013_n25097.n1 a_23013_n25097.t14 13.849
R12378 a_23013_n25097.n0 a_23013_n25097.t15 13.849
R12379 a_23013_n25097.n9 a_23013_n25097.t11 13.849
R12380 a_23013_n25097.n8 a_23013_n25097.t18 13.849
R12381 a_23013_n25097.n7 a_23013_n25097.t9 13.849
R12382 a_23013_n25097.n6 a_23013_n25097.t16 13.849
R12383 a_23013_n25097.n5 a_23013_n25097.t8 13.849
R12384 a_23013_n25097.n15 a_23013_n25097.t7 7.181
R12385 a_23013_n25097.t22 a_23013_n25097.n10 7.039
R12386 a_23013_n25097.n19 a_23013_n25097.t21 6.584
R12387 a_23013_n25097.n17 a_23013_n25097.t1 6.584
R12388 a_23013_n25097.n16 a_23013_n25097.t6 6.584
R12389 a_23013_n25097.n20 a_23013_n25097.n19 5.451
R12390 a_23013_n25097.t22 a_23013_n25097.n21 4.454
R12391 a_23013_n25097.n11 a_23013_n25097.t2 4.132
R12392 a_23013_n25097.n11 a_23013_n25097.t24 4.132
R12393 a_23013_n25097.n12 a_23013_n25097.t23 4.132
R12394 a_23013_n25097.n12 a_23013_n25097.t3 4.132
R12395 a_23013_n25097.n13 a_23013_n25097.t0 4.132
R12396 a_23013_n25097.n13 a_23013_n25097.t20 4.132
R12397 a_23013_n25097.n14 a_23013_n25097.t5 4.132
R12398 a_23013_n25097.n14 a_23013_n25097.t4 4.132
R12399 a_23013_n25097.n10 a_23013_n25097.n9 2.909
R12400 a_23013_n25097.n21 a_23013_n25097.n11 2.452
R12401 a_23013_n25097.n20 a_23013_n25097.n12 2.452
R12402 a_23013_n25097.n18 a_23013_n25097.n13 2.452
R12403 a_23013_n25097.n15 a_23013_n25097.n14 2.452
R12404 a_23013_n25097.n1 a_23013_n25097.n0 1.159
R12405 a_23013_n25097.n3 a_23013_n25097.n2 1.159
R12406 a_23013_n25097.n6 a_23013_n25097.n5 1.159
R12407 a_23013_n25097.n8 a_23013_n25097.n7 1.159
R12408 a_23013_n25097.n17 a_23013_n25097.n16 0.795
R12409 a_23013_n25097.n2 a_23013_n25097.n1 0.749
R12410 a_23013_n25097.n4 a_23013_n25097.n3 0.749
R12411 a_23013_n25097.n7 a_23013_n25097.n6 0.749
R12412 a_23013_n25097.n9 a_23013_n25097.n8 0.749
R12413 a_23013_n25097.n10 a_23013_n25097.n4 0.71
R12414 a_23013_n25097.n16 a_23013_n25097.n15 0.597
R12415 a_23013_n25097.n18 a_23013_n25097.n17 0.597
R12416 a_23013_n25097.n19 a_23013_n25097.n18 0.597
R12417 a_23013_n25097.n21 a_23013_n25097.n20 0.597
R12418 bias_p.n215 bias_p.n214 15.3
R12419 bias_p.n216 bias_p.t2 13.849
R12420 bias_p.n36 bias_p.t44 12.05
R12421 bias_p.n36 bias_p.t37 12.05
R12422 bias_p.n29 bias_p.t88 12.05
R12423 bias_p.n29 bias_p.t84 12.05
R12424 bias_p.n28 bias_p.t86 12.05
R12425 bias_p.n28 bias_p.t71 12.05
R12426 bias_p.n27 bias_p.t32 12.05
R12427 bias_p.n27 bias_p.t15 12.05
R12428 bias_p.n26 bias_p.t73 12.05
R12429 bias_p.n26 bias_p.t59 12.05
R12430 bias_p.n25 bias_p.t27 12.05
R12431 bias_p.n25 bias_p.t12 12.05
R12432 bias_p.n24 bias_p.t64 12.05
R12433 bias_p.n24 bias_p.t56 12.05
R12434 bias_p.n114 bias_p.t50 12.05
R12435 bias_p.n114 bias_p.t20 12.05
R12436 bias_p.n6 bias_p.t77 12.05
R12437 bias_p.n6 bias_p.t25 12.05
R12438 bias_p.n5 bias_p.t36 12.05
R12439 bias_p.n5 bias_p.t79 12.05
R12440 bias_p.n10 bias_p.t54 12.05
R12441 bias_p.n10 bias_p.t98 12.05
R12442 bias_p.n11 bias_p.t102 12.05
R12443 bias_p.n11 bias_p.t55 12.05
R12444 bias_p.n12 bias_p.t63 12.05
R12445 bias_p.n12 bias_p.t11 12.05
R12446 bias_p.n13 bias_p.t75 12.05
R12447 bias_p.n13 bias_p.t23 12.05
R12448 bias_p.n14 bias_p.t34 12.05
R12449 bias_p.n14 bias_p.t78 12.05
R12450 bias_p.n22 bias_p.t38 12.05
R12451 bias_p.n22 bias_p.t29 12.05
R12452 bias_p.n34 bias_p.t40 12.05
R12453 bias_p.n34 bias_p.t87 12.05
R12454 bias_p.n35 bias_p.t91 12.05
R12455 bias_p.n35 bias_p.t41 12.05
R12456 bias_p.n32 bias_p.t47 12.05
R12457 bias_p.n32 bias_p.t39 12.05
R12458 bias_p.n33 bias_p.t96 12.05
R12459 bias_p.n33 bias_p.t90 12.05
R12460 bias_p.n30 bias_p.t93 12.05
R12461 bias_p.n30 bias_p.t43 12.05
R12462 bias_p.n31 bias_p.t49 12.05
R12463 bias_p.n31 bias_p.t94 12.05
R12464 bias_p.n21 bias_p.t85 12.05
R12465 bias_p.n21 bias_p.t69 12.05
R12466 bias_p.n20 bias_p.t72 12.05
R12467 bias_p.n20 bias_p.t58 12.05
R12468 bias_p.n19 bias_p.t16 12.05
R12469 bias_p.n19 bias_p.t101 12.05
R12470 bias_p.n18 bias_p.t60 12.05
R12471 bias_p.n18 bias_p.t52 12.05
R12472 bias_p.n17 bias_p.t13 12.05
R12473 bias_p.n17 bias_p.t99 12.05
R12474 bias_p.n1 bias_p.t28 12.05
R12475 bias_p.n1 bias_p.t14 12.05
R12476 bias_p.n116 bias_p.t22 12.05
R12477 bias_p.n116 bias_p.t80 12.05
R12478 bias_p.n2 bias_p.t83 12.05
R12479 bias_p.n2 bias_p.t67 12.05
R12480 bias_p.n99 bias_p.t35 12.05
R12481 bias_p.n99 bias_p.t19 12.05
R12482 bias_p.n3 bias_p.t17 12.05
R12483 bias_p.n3 bias_p.t62 12.05
R12484 bias_p.n118 bias_p.t81 12.05
R12485 bias_p.n118 bias_p.t45 12.05
R12486 bias_p.n4 bias_p.t74 12.05
R12487 bias_p.n4 bias_p.t21 12.05
R12488 bias_p.n101 bias_p.t26 12.05
R12489 bias_p.n101 bias_p.t66 12.05
R12490 bias_p.n8 bias_p.t51 12.05
R12491 bias_p.n8 bias_p.t95 12.05
R12492 bias_p.n7 bias_p.t33 12.05
R12493 bias_p.n7 bias_p.t92 12.05
R12494 bias_p.n9 bias_p.t100 12.05
R12495 bias_p.n9 bias_p.t53 12.05
R12496 bias_p.n16 bias_p.t57 12.05
R12497 bias_p.n16 bias_p.t48 12.05
R12498 bias_p.n15 bias_p.t68 12.05
R12499 bias_p.n15 bias_p.t31 12.05
R12500 bias_p.n38 bias_p.t70 12.05
R12501 bias_p.n38 bias_p.t18 12.05
R12502 bias_p.n39 bias_p.t24 12.05
R12503 bias_p.n39 bias_p.t65 12.05
R12504 bias_p.n37 bias_p.t42 12.05
R12505 bias_p.n37 bias_p.t89 12.05
R12506 bias_p.n97 bias_p.t82 12.05
R12507 bias_p.n97 bias_p.t30 12.05
R12508 bias_p.n23 bias_p.t46 12.05
R12509 bias_p.n23 bias_p.t97 12.05
R12510 bias_p.n215 bias_p.n44 9.619
R12511 bias_p.n53 bias_p.n51 9.3
R12512 bias_p.n53 bias_p.n52 9.3
R12513 bias_p.n84 bias_p.n82 9.3
R12514 bias_p.n84 bias_p.n83 9.3
R12515 bias_p.n88 bias_p.n86 9.3
R12516 bias_p.n88 bias_p.n87 9.3
R12517 bias_p.n92 bias_p.n90 9.3
R12518 bias_p.n92 bias_p.n91 9.3
R12519 bias_p.n96 bias_p.n94 9.3
R12520 bias_p.n96 bias_p.n95 9.3
R12521 bias_p.n106 bias_p.n104 9.3
R12522 bias_p.n106 bias_p.n105 9.3
R12523 bias_p.n113 bias_p.n111 9.3
R12524 bias_p.n113 bias_p.n112 9.3
R12525 bias_p.n192 bias_p.n190 9.3
R12526 bias_p.n192 bias_p.n191 9.3
R12527 bias_p.n188 bias_p.n186 9.3
R12528 bias_p.n188 bias_p.n187 9.3
R12529 bias_p.n184 bias_p.n182 9.3
R12530 bias_p.n184 bias_p.n183 9.3
R12531 bias_p.n180 bias_p.n178 9.3
R12532 bias_p.n180 bias_p.n179 9.3
R12533 bias_p.n176 bias_p.n174 9.3
R12534 bias_p.n176 bias_p.n175 9.3
R12535 bias_p.n134 bias_p.n132 9.3
R12536 bias_p.n134 bias_p.n133 9.3
R12537 bias_p.n61 bias_p.n59 9.3
R12538 bias_p.n61 bias_p.n60 9.3
R12539 bias_p.n57 bias_p.n55 9.3
R12540 bias_p.n57 bias_p.n56 9.3
R12541 bias_p.n69 bias_p.n67 9.3
R12542 bias_p.n69 bias_p.n68 9.3
R12543 bias_p.n65 bias_p.n63 9.3
R12544 bias_p.n65 bias_p.n64 9.3
R12545 bias_p.n77 bias_p.n75 9.3
R12546 bias_p.n77 bias_p.n76 9.3
R12547 bias_p.n73 bias_p.n71 9.3
R12548 bias_p.n73 bias_p.n72 9.3
R12549 bias_p.n138 bias_p.n136 9.3
R12550 bias_p.n138 bias_p.n137 9.3
R12551 bias_p.n142 bias_p.n140 9.3
R12552 bias_p.n142 bias_p.n141 9.3
R12553 bias_p.n146 bias_p.n144 9.3
R12554 bias_p.n146 bias_p.n145 9.3
R12555 bias_p.n150 bias_p.n148 9.3
R12556 bias_p.n150 bias_p.n149 9.3
R12557 bias_p.n154 bias_p.n152 9.3
R12558 bias_p.n154 bias_p.n153 9.3
R12559 bias_p.n200 bias_p.n198 9.3
R12560 bias_p.n200 bias_p.n199 9.3
R12561 bias_p.n204 bias_p.n202 9.3
R12562 bias_p.n204 bias_p.n203 9.3
R12563 bias_p.n196 bias_p.n194 9.3
R12564 bias_p.n196 bias_p.n195 9.3
R12565 bias_p.n158 bias_p.n156 9.3
R12566 bias_p.n158 bias_p.n157 9.3
R12567 bias_p.n162 bias_p.n160 9.3
R12568 bias_p.n162 bias_p.n161 9.3
R12569 bias_p.n43 bias_p.n41 9.3
R12570 bias_p.n43 bias_p.n42 9.3
R12571 bias_p.n48 bias_p.n46 9.3
R12572 bias_p.n48 bias_p.n47 9.3
R12573 bias_p.n123 bias_p.n121 9.3
R12574 bias_p.n123 bias_p.n122 9.3
R12575 bias_p.n44 bias_p.t10 8.857
R12576 bias_p.n44 bias_p.t9 8.266
R12577 bias_p.n172 bias_p.t8 7.482
R12578 bias_p.n170 bias_p.t5 7.48
R12579 bias_p.n49 bias_p.t6 6.923
R12580 bias_p.n49 bias_p.t7 6.923
R12581 bias_p.n214 bias_p.n213 5.786
R12582 bias_p.n39 bias_p.n38 1.738
R12583 bias_p.t1 bias_p.n39 1.73
R12584 bias_p.n80 bias_p.n35 1.228
R12585 bias_p.n79 bias_p.n33 1.228
R12586 bias_p.n78 bias_p.n31 1.228
R12587 bias_p.n8 bias_p.n205 1.228
R12588 bias_p.n9 bias_p.n206 1.228
R12589 bias_p.n16 bias_p.n163 1.228
R12590 bias_p.n17 bias_p.n164 1.228
R12591 bias_p.n18 bias_p.n165 1.228
R12592 bias_p.n19 bias_p.n166 1.228
R12593 bias_p.n20 bias_p.n167 1.228
R12594 bias_p.n21 bias_p.n168 1.228
R12595 bias_p.n22 bias_p.n169 1.228
R12596 bias_p.n14 bias_p.n211 1.228
R12597 bias_p.n13 bias_p.n210 1.228
R12598 bias_p.n12 bias_p.n209 1.228
R12599 bias_p.n11 bias_p.n208 1.228
R12600 bias_p.n10 bias_p.n207 1.228
R12601 bias_p.n24 bias_p.n124 1.228
R12602 bias_p.n25 bias_p.n125 1.228
R12603 bias_p.n26 bias_p.n126 1.228
R12604 bias_p.n27 bias_p.n127 1.228
R12605 bias_p.n28 bias_p.n128 1.228
R12606 bias_p.n29 bias_p.n129 1.228
R12607 bias_p.n36 bias_p.n130 1.228
R12608 bias_p.n100 bias_p.n99 1.22
R12609 bias_p.n102 bias_p.n101 1.22
R12610 bias_p.n98 bias_p.n97 1.22
R12611 bias_p.n214 bias_p.n37 1.085
R12612 bias_p.n36 bias_p.n50 0.752
R12613 bias_p.n29 bias_p.n81 0.752
R12614 bias_p.n28 bias_p.n85 0.752
R12615 bias_p.n27 bias_p.n89 0.752
R12616 bias_p.n26 bias_p.n93 0.752
R12617 bias_p.n25 bias_p.n103 0.752
R12618 bias_p.n24 bias_p.n110 0.752
R12619 bias_p.n10 bias_p.n189 0.752
R12620 bias_p.n11 bias_p.n185 0.752
R12621 bias_p.n12 bias_p.n181 0.752
R12622 bias_p.n13 bias_p.n177 0.752
R12623 bias_p.n14 bias_p.n173 0.752
R12624 bias_p.n22 bias_p.n131 0.752
R12625 bias_p.n34 bias_p.n58 0.752
R12626 bias_p.n35 bias_p.n54 0.752
R12627 bias_p.n32 bias_p.n66 0.752
R12628 bias_p.n33 bias_p.n62 0.752
R12629 bias_p.n30 bias_p.n74 0.752
R12630 bias_p.n31 bias_p.n70 0.752
R12631 bias_p.n21 bias_p.n135 0.752
R12632 bias_p.n20 bias_p.n139 0.752
R12633 bias_p.n19 bias_p.n143 0.752
R12634 bias_p.n18 bias_p.n147 0.752
R12635 bias_p.n17 bias_p.n151 0.752
R12636 bias_p.n8 bias_p.n197 0.752
R12637 bias_p.n7 bias_p.n201 0.752
R12638 bias_p.n9 bias_p.n193 0.752
R12639 bias_p.n16 bias_p.n155 0.752
R12640 bias_p.n15 bias_p.n159 0.752
R12641 bias_p.n38 bias_p.n40 0.752
R12642 bias_p.n37 bias_p.n45 0.752
R12643 bias_p.n23 bias_p.n120 0.752
R12644 bias_p.n0 bias_p.n36 0.704
R12645 bias_p.n107 bias_p.n6 0.633
R12646 bias_p.n98 bias_p.n5 0.633
R12647 bias_p.n102 bias_p.n4 0.633
R12648 bias_p.n109 bias_p.n3 0.633
R12649 bias_p.n100 bias_p.n2 0.633
R12650 bias_p.n108 bias_p.n1 0.633
R12651 bias_p.n171 bias_p.n49 0.591
R12652 bias_p.n115 bias_p.n114 0.589
R12653 bias_p.n117 bias_p.n116 0.589
R12654 bias_p.n119 bias_p.n118 0.589
R12655 bias_p.n213 bias_p.n212 0.512
R12656 bias_p.n80 bias_p.n34 0.478
R12657 bias_p.n79 bias_p.n32 0.478
R12658 bias_p.n78 bias_p.n30 0.478
R12659 bias_p.n205 bias_p.n7 0.478
R12660 bias_p.n206 bias_p.n8 0.478
R12661 bias_p.n207 bias_p.n9 0.478
R12662 bias_p.n163 bias_p.n15 0.478
R12663 bias_p.n164 bias_p.n16 0.478
R12664 bias_p.n165 bias_p.n17 0.478
R12665 bias_p.n166 bias_p.n18 0.478
R12666 bias_p.n167 bias_p.n19 0.478
R12667 bias_p.n168 bias_p.n20 0.478
R12668 bias_p.n169 bias_p.n21 0.478
R12669 bias_p.n0 bias_p.n22 0.478
R12670 bias_p.n212 bias_p.n14 0.478
R12671 bias_p.n211 bias_p.n13 0.478
R12672 bias_p.n210 bias_p.n12 0.478
R12673 bias_p.n209 bias_p.n11 0.478
R12674 bias_p.n208 bias_p.n10 0.478
R12675 bias_p.n124 bias_p.n23 0.478
R12676 bias_p.n125 bias_p.n24 0.478
R12677 bias_p.n126 bias_p.n25 0.478
R12678 bias_p.n127 bias_p.n26 0.478
R12679 bias_p.n128 bias_p.n27 0.478
R12680 bias_p.n129 bias_p.n28 0.478
R12681 bias_p.n130 bias_p.n29 0.478
R12682 bias_p.n170 bias_p.n0 0.47
R12683 bias_p.n79 bias_p.n78 0.417
R12684 bias_p.n80 bias_p.n79 0.417
R12685 bias_p.n130 bias_p.n80 0.417
R12686 bias_p.n108 bias_p.n107 0.417
R12687 bias_p.n109 bias_p.n108 0.417
R12688 bias_p.n125 bias_p.n109 0.417
R12689 bias_p.n100 bias_p.n98 0.417
R12690 bias_p.n102 bias_p.n100 0.417
R12691 bias_p.n126 bias_p.n102 0.417
R12692 bias_p.n117 bias_p.n115 0.417
R12693 bias_p.n119 bias_p.n117 0.417
R12694 bias_p.n124 bias_p.n119 0.417
R12695 bias_p.n216 bias_p.n215 0.361
R12696 bias_p bias_p.n216 0.314
R12697 bias_p.n37 bias_p.n48 0.285
R12698 bias_p.n36 bias_p.n53 0.285
R12699 bias_p.n35 bias_p.n57 0.285
R12700 bias_p.n34 bias_p.n61 0.285
R12701 bias_p.n33 bias_p.n65 0.285
R12702 bias_p.n32 bias_p.n69 0.285
R12703 bias_p.n31 bias_p.n73 0.285
R12704 bias_p.n30 bias_p.n77 0.285
R12705 bias_p.n29 bias_p.n84 0.285
R12706 bias_p.n28 bias_p.n88 0.285
R12707 bias_p.n27 bias_p.n92 0.285
R12708 bias_p.n26 bias_p.n96 0.285
R12709 bias_p.n25 bias_p.n106 0.285
R12710 bias_p.n24 bias_p.n113 0.285
R12711 bias_p.n23 bias_p.n123 0.285
R12712 bias_p.n22 bias_p.n134 0.285
R12713 bias_p.n21 bias_p.n138 0.285
R12714 bias_p.n20 bias_p.n142 0.285
R12715 bias_p.n19 bias_p.n146 0.285
R12716 bias_p.n18 bias_p.n150 0.285
R12717 bias_p.n17 bias_p.n154 0.285
R12718 bias_p.n16 bias_p.n158 0.285
R12719 bias_p.n15 bias_p.n162 0.285
R12720 bias_p.n14 bias_p.n176 0.285
R12721 bias_p.n13 bias_p.n180 0.285
R12722 bias_p.n12 bias_p.n184 0.285
R12723 bias_p.n11 bias_p.n188 0.285
R12724 bias_p.n10 bias_p.n192 0.285
R12725 bias_p.n9 bias_p.n196 0.285
R12726 bias_p.n8 bias_p.n200 0.285
R12727 bias_p.n7 bias_p.n204 0.285
R12728 bias_p.n38 bias_p.n43 0.281
R12729 bias_p bias_p.t1 0.274
R12730 bias_p.n213 bias_p.n172 0.166
R12731 bias_p.n171 bias_p.n170 0.145
R12732 bias_p.n172 bias_p.n171 0.145
R12733 a_2467_n30310.n98 a_2467_n30310.n97 11.662
R12734 a_2467_n30310.n94 a_2467_n30310.t117 9.546
R12735 a_2467_n30310.n97 a_2467_n30310.t60 8.896
R12736 a_2467_n30310.n112 a_2467_n30310.t50 8.266
R12737 a_2467_n30310.n102 a_2467_n30310.t80 8.266
R12738 a_2467_n30310.n102 a_2467_n30310.t19 8.266
R12739 a_2467_n30310.n101 a_2467_n30310.t99 8.266
R12740 a_2467_n30310.n101 a_2467_n30310.t36 8.266
R12741 a_2467_n30310.n104 a_2467_n30310.t88 8.266
R12742 a_2467_n30310.n104 a_2467_n30310.t57 8.266
R12743 a_2467_n30310.n103 a_2467_n30310.t106 8.266
R12744 a_2467_n30310.n103 a_2467_n30310.t51 8.266
R12745 a_2467_n30310.n106 a_2467_n30310.t72 8.266
R12746 a_2467_n30310.n106 a_2467_n30310.t114 8.266
R12747 a_2467_n30310.n105 a_2467_n30310.t76 8.266
R12748 a_2467_n30310.n105 a_2467_n30310.t43 8.266
R12749 a_2467_n30310.n108 a_2467_n30310.t87 8.266
R12750 a_2467_n30310.n108 a_2467_n30310.t54 8.266
R12751 a_2467_n30310.n107 a_2467_n30310.t73 8.266
R12752 a_2467_n30310.n107 a_2467_n30310.t49 8.266
R12753 a_2467_n30310.n2 a_2467_n30310.t86 8.266
R12754 a_2467_n30310.n2 a_2467_n30310.t56 8.266
R12755 a_2467_n30310.n1 a_2467_n30310.t105 8.266
R12756 a_2467_n30310.n1 a_2467_n30310.t48 8.266
R12757 a_2467_n30310.n57 a_2467_n30310.t69 8.266
R12758 a_2467_n30310.n57 a_2467_n30310.t28 8.266
R12759 a_2467_n30310.n56 a_2467_n30310.t92 8.266
R12760 a_2467_n30310.n56 a_2467_n30310.t62 8.266
R12761 a_2467_n30310.n59 a_2467_n30310.t91 8.266
R12762 a_2467_n30310.n59 a_2467_n30310.t63 8.266
R12763 a_2467_n30310.n58 a_2467_n30310.t71 8.266
R12764 a_2467_n30310.n58 a_2467_n30310.t31 8.266
R12765 a_2467_n30310.n61 a_2467_n30310.t70 8.266
R12766 a_2467_n30310.n61 a_2467_n30310.t20 8.266
R12767 a_2467_n30310.n60 a_2467_n30310.t95 8.266
R12768 a_2467_n30310.n60 a_2467_n30310.t22 8.266
R12769 a_2467_n30310.n63 a_2467_n30310.t35 8.266
R12770 a_2467_n30310.n63 a_2467_n30310.t94 8.266
R12771 a_2467_n30310.n62 a_2467_n30310.t90 8.266
R12772 a_2467_n30310.n62 a_2467_n30310.t5 8.266
R12773 a_2467_n30310.n46 a_2467_n30310.t103 8.266
R12774 a_2467_n30310.n46 a_2467_n30310.t13 8.266
R12775 a_2467_n30310.n45 a_2467_n30310.t83 8.266
R12776 a_2467_n30310.n45 a_2467_n30310.t112 8.266
R12777 a_2467_n30310.n48 a_2467_n30310.t82 8.266
R12778 a_2467_n30310.n48 a_2467_n30310.t113 8.266
R12779 a_2467_n30310.n47 a_2467_n30310.t107 8.266
R12780 a_2467_n30310.n47 a_2467_n30310.t109 8.266
R12781 a_2467_n30310.n50 a_2467_n30310.t104 8.266
R12782 a_2467_n30310.n50 a_2467_n30310.t115 8.266
R12783 a_2467_n30310.n49 a_2467_n30310.t84 8.266
R12784 a_2467_n30310.n49 a_2467_n30310.t4 8.266
R12785 a_2467_n30310.n52 a_2467_n30310.t93 8.266
R12786 a_2467_n30310.n52 a_2467_n30310.t40 8.266
R12787 a_2467_n30310.n51 a_2467_n30310.t89 8.266
R12788 a_2467_n30310.n51 a_2467_n30310.t34 8.266
R12789 a_2467_n30310.n4 a_2467_n30310.t77 8.266
R12790 a_2467_n30310.n4 a_2467_n30310.t41 8.266
R12791 a_2467_n30310.n3 a_2467_n30310.t96 8.266
R12792 a_2467_n30310.n3 a_2467_n30310.t23 8.266
R12793 a_2467_n30310.n6 a_2467_n30310.t98 8.266
R12794 a_2467_n30310.n6 a_2467_n30310.t61 8.266
R12795 a_2467_n30310.n5 a_2467_n30310.t75 8.266
R12796 a_2467_n30310.n5 a_2467_n30310.t42 8.266
R12797 a_2467_n30310.n8 a_2467_n30310.t78 8.266
R12798 a_2467_n30310.n8 a_2467_n30310.t14 8.266
R12799 a_2467_n30310.n7 a_2467_n30310.t97 8.266
R12800 a_2467_n30310.n7 a_2467_n30310.t37 8.266
R12801 a_2467_n30310.n10 a_2467_n30310.t74 8.266
R12802 a_2467_n30310.n10 a_2467_n30310.t24 8.266
R12803 a_2467_n30310.n9 a_2467_n30310.t102 8.266
R12804 a_2467_n30310.n9 a_2467_n30310.t30 8.266
R12805 a_2467_n30310.n87 a_2467_n30310.t79 8.266
R12806 a_2467_n30310.n87 a_2467_n30310.t52 8.266
R12807 a_2467_n30310.n86 a_2467_n30310.t101 8.266
R12808 a_2467_n30310.n86 a_2467_n30310.t47 8.266
R12809 a_2467_n30310.n89 a_2467_n30310.t100 8.266
R12810 a_2467_n30310.n89 a_2467_n30310.t46 8.266
R12811 a_2467_n30310.n88 a_2467_n30310.t81 8.266
R12812 a_2467_n30310.n88 a_2467_n30310.t53 8.266
R12813 a_2467_n30310.n0 a_2467_n30310.t85 8.266
R12814 a_2467_n30310.n0 a_2467_n30310.t55 8.266
R12815 a_2467_n30310.t108 a_2467_n30310.n112 8.266
R12816 a_2467_n30310.n82 a_2467_n30310.n81 8.096
R12817 a_2467_n30310.n91 a_2467_n30310.t111 6.923
R12818 a_2467_n30310.n91 a_2467_n30310.t116 6.923
R12819 a_2467_n30310.n92 a_2467_n30310.t59 6.923
R12820 a_2467_n30310.n92 a_2467_n30310.t15 6.923
R12821 a_2467_n30310.n93 a_2467_n30310.t3 6.923
R12822 a_2467_n30310.n93 a_2467_n30310.t16 6.923
R12823 a_2467_n30310.n24 a_2467_n30310.n21 4.696
R12824 a_2467_n30310.n44 a_2467_n30310.n17 4.508
R12825 a_2467_n30310.n40 a_2467_n30310.n39 4.508
R12826 a_2467_n30310.n29 a_2467_n30310.n28 4.508
R12827 a_2467_n30310.n84 a_2467_n30310.n44 4.307
R12828 a_2467_n30310.n100 a_2467_n30310.n99 3.617
R12829 a_2467_n30310.n82 a_2467_n30310.n66 3.616
R12830 a_2467_n30310.n83 a_2467_n30310.n55 3.616
R12831 a_2467_n30310.n85 a_2467_n30310.n13 3.616
R12832 a_2467_n30310.n98 a_2467_n30310.n90 3.616
R12833 a_2467_n30310.n17 a_2467_n30310.t29 3.463
R12834 a_2467_n30310.n16 a_2467_n30310.t64 3.463
R12835 a_2467_n30310.n15 a_2467_n30310.t6 3.463
R12836 a_2467_n30310.n14 a_2467_n30310.t58 3.463
R12837 a_2467_n30310.n18 a_2467_n30310.t10 3.463
R12838 a_2467_n30310.n19 a_2467_n30310.t27 3.463
R12839 a_2467_n30310.n20 a_2467_n30310.t11 3.463
R12840 a_2467_n30310.n21 a_2467_n30310.t38 3.463
R12841 a_2467_n30310.n68 a_2467_n30310.t7 3.463
R12842 a_2467_n30310.n67 a_2467_n30310.t21 3.463
R12843 a_2467_n30310.n41 a_2467_n30310.t25 3.463
R12844 a_2467_n30310.n42 a_2467_n30310.t44 3.463
R12845 a_2467_n30310.n36 a_2467_n30310.t0 3.463
R12846 a_2467_n30310.n37 a_2467_n30310.t39 3.463
R12847 a_2467_n30310.n38 a_2467_n30310.t1 3.463
R12848 a_2467_n30310.n39 a_2467_n30310.t9 3.463
R12849 a_2467_n30310.n70 a_2467_n30310.t110 3.463
R12850 a_2467_n30310.n69 a_2467_n30310.t26 3.463
R12851 a_2467_n30310.n33 a_2467_n30310.t12 3.463
R12852 a_2467_n30310.n34 a_2467_n30310.t18 3.463
R12853 a_2467_n30310.n72 a_2467_n30310.t17 3.463
R12854 a_2467_n30310.n71 a_2467_n30310.t119 3.463
R12855 a_2467_n30310.n30 a_2467_n30310.t65 3.463
R12856 a_2467_n30310.n31 a_2467_n30310.t68 3.463
R12857 a_2467_n30310.n25 a_2467_n30310.t8 3.463
R12858 a_2467_n30310.n26 a_2467_n30310.t33 3.463
R12859 a_2467_n30310.n27 a_2467_n30310.t118 3.463
R12860 a_2467_n30310.n28 a_2467_n30310.t66 3.463
R12861 a_2467_n30310.n74 a_2467_n30310.t67 3.463
R12862 a_2467_n30310.n73 a_2467_n30310.t32 3.463
R12863 a_2467_n30310.n22 a_2467_n30310.t45 3.463
R12864 a_2467_n30310.n23 a_2467_n30310.t2 3.463
R12865 a_2467_n30310.n64 a_2467_n30310.n63 2.668
R12866 a_2467_n30310.n53 a_2467_n30310.n52 2.668
R12867 a_2467_n30310.n11 a_2467_n30310.n10 2.668
R12868 a_2467_n30310.n90 a_2467_n30310.n89 2.668
R12869 a_2467_n30310.n111 a_2467_n30310.n100 2.221
R12870 a_2467_n30310.n111 a_2467_n30310.n110 2.22
R12871 a_2467_n30310.n110 a_2467_n30310.n109 2.219
R12872 a_2467_n30310.n65 a_2467_n30310.n64 2.219
R12873 a_2467_n30310.n66 a_2467_n30310.n65 2.219
R12874 a_2467_n30310.n54 a_2467_n30310.n53 2.219
R12875 a_2467_n30310.n55 a_2467_n30310.n54 2.219
R12876 a_2467_n30310.n12 a_2467_n30310.n11 2.219
R12877 a_2467_n30310.n13 a_2467_n30310.n12 2.219
R12878 a_2467_n30310.n96 a_2467_n30310.n91 1.973
R12879 a_2467_n30310.n95 a_2467_n30310.n92 1.973
R12880 a_2467_n30310.n94 a_2467_n30310.n93 1.973
R12881 a_2467_n30310.n80 a_2467_n30310.n68 1.617
R12882 a_2467_n30310.n78 a_2467_n30310.n70 1.617
R12883 a_2467_n30310.n77 a_2467_n30310.n72 1.617
R12884 a_2467_n30310.n75 a_2467_n30310.n74 1.617
R12885 a_2467_n30310.n19 a_2467_n30310.n18 1.352
R12886 a_2467_n30310.n20 a_2467_n30310.n19 1.352
R12887 a_2467_n30310.n21 a_2467_n30310.n20 1.352
R12888 a_2467_n30310.n42 a_2467_n30310.n41 1.352
R12889 a_2467_n30310.n68 a_2467_n30310.n67 1.352
R12890 a_2467_n30310.n39 a_2467_n30310.n38 1.352
R12891 a_2467_n30310.n38 a_2467_n30310.n37 1.352
R12892 a_2467_n30310.n37 a_2467_n30310.n36 1.352
R12893 a_2467_n30310.n34 a_2467_n30310.n33 1.352
R12894 a_2467_n30310.n70 a_2467_n30310.n69 1.352
R12895 a_2467_n30310.n31 a_2467_n30310.n30 1.352
R12896 a_2467_n30310.n72 a_2467_n30310.n71 1.352
R12897 a_2467_n30310.n28 a_2467_n30310.n27 1.352
R12898 a_2467_n30310.n27 a_2467_n30310.n26 1.352
R12899 a_2467_n30310.n26 a_2467_n30310.n25 1.352
R12900 a_2467_n30310.n23 a_2467_n30310.n22 1.352
R12901 a_2467_n30310.n74 a_2467_n30310.n73 1.352
R12902 a_2467_n30310.n17 a_2467_n30310.n16 1.352
R12903 a_2467_n30310.n16 a_2467_n30310.n15 1.352
R12904 a_2467_n30310.n15 a_2467_n30310.n14 1.352
R12905 a_2467_n30310.n43 a_2467_n30310.n42 1.302
R12906 a_2467_n30310.n35 a_2467_n30310.n34 1.302
R12907 a_2467_n30310.n32 a_2467_n30310.n31 1.302
R12908 a_2467_n30310.n24 a_2467_n30310.n23 1.302
R12909 a_2467_n30310.n99 a_2467_n30310.n98 0.752
R12910 a_2467_n30310.n99 a_2467_n30310.n85 0.752
R12911 a_2467_n30310.n83 a_2467_n30310.n82 0.749
R12912 a_2467_n30310.n85 a_2467_n30310.n84 0.714
R12913 a_2467_n30310.n96 a_2467_n30310.n95 0.65
R12914 a_2467_n30310.n97 a_2467_n30310.n96 0.65
R12915 a_2467_n30310.n95 a_2467_n30310.n94 0.637
R12916 a_2467_n30310.n110 a_2467_n30310.n104 0.449
R12917 a_2467_n30310.n109 a_2467_n30310.n108 0.449
R12918 a_2467_n30310.n100 a_2467_n30310.n2 0.449
R12919 a_2467_n30310.n66 a_2467_n30310.n57 0.449
R12920 a_2467_n30310.n65 a_2467_n30310.n59 0.449
R12921 a_2467_n30310.n64 a_2467_n30310.n61 0.449
R12922 a_2467_n30310.n55 a_2467_n30310.n46 0.449
R12923 a_2467_n30310.n54 a_2467_n30310.n48 0.449
R12924 a_2467_n30310.n53 a_2467_n30310.n50 0.449
R12925 a_2467_n30310.n13 a_2467_n30310.n4 0.449
R12926 a_2467_n30310.n12 a_2467_n30310.n6 0.449
R12927 a_2467_n30310.n11 a_2467_n30310.n8 0.449
R12928 a_2467_n30310.n90 a_2467_n30310.n87 0.449
R12929 a_2467_n30310.n112 a_2467_n30310.n111 0.449
R12930 a_2467_n30310.n102 a_2467_n30310.n101 0.365
R12931 a_2467_n30310.n104 a_2467_n30310.n103 0.365
R12932 a_2467_n30310.n106 a_2467_n30310.n105 0.365
R12933 a_2467_n30310.n108 a_2467_n30310.n107 0.365
R12934 a_2467_n30310.n2 a_2467_n30310.n1 0.365
R12935 a_2467_n30310.n57 a_2467_n30310.n56 0.365
R12936 a_2467_n30310.n59 a_2467_n30310.n58 0.365
R12937 a_2467_n30310.n61 a_2467_n30310.n60 0.365
R12938 a_2467_n30310.n63 a_2467_n30310.n62 0.365
R12939 a_2467_n30310.n46 a_2467_n30310.n45 0.365
R12940 a_2467_n30310.n48 a_2467_n30310.n47 0.365
R12941 a_2467_n30310.n50 a_2467_n30310.n49 0.365
R12942 a_2467_n30310.n52 a_2467_n30310.n51 0.365
R12943 a_2467_n30310.n4 a_2467_n30310.n3 0.365
R12944 a_2467_n30310.n6 a_2467_n30310.n5 0.365
R12945 a_2467_n30310.n8 a_2467_n30310.n7 0.365
R12946 a_2467_n30310.n10 a_2467_n30310.n9 0.365
R12947 a_2467_n30310.n87 a_2467_n30310.n86 0.365
R12948 a_2467_n30310.n89 a_2467_n30310.n88 0.365
R12949 a_2467_n30310.n112 a_2467_n30310.n0 0.365
R12950 a_2467_n30310.n110 a_2467_n30310.n102 0.237
R12951 a_2467_n30310.n109 a_2467_n30310.n106 0.237
R12952 a_2467_n30310.n81 a_2467_n30310.n80 0.188
R12953 a_2467_n30310.n80 a_2467_n30310.n79 0.188
R12954 a_2467_n30310.n79 a_2467_n30310.n78 0.188
R12955 a_2467_n30310.n78 a_2467_n30310.n77 0.188
R12956 a_2467_n30310.n77 a_2467_n30310.n76 0.188
R12957 a_2467_n30310.n76 a_2467_n30310.n75 0.188
R12958 a_2467_n30310.n44 a_2467_n30310.n43 0.188
R12959 a_2467_n30310.n43 a_2467_n30310.n40 0.188
R12960 a_2467_n30310.n40 a_2467_n30310.n35 0.188
R12961 a_2467_n30310.n35 a_2467_n30310.n32 0.188
R12962 a_2467_n30310.n32 a_2467_n30310.n29 0.188
R12963 a_2467_n30310.n29 a_2467_n30310.n24 0.188
R12964 a_2467_n30310.n84 a_2467_n30310.n83 0.034
R12965 level_shifter_up_0.xb_hv.n1 level_shifter_up_0.xb_hv.t2 132.104
R12966 level_shifter_up_0.xb_hv.n2 level_shifter_up_0.xb_hv.t4 132.103
R12967 level_shifter_up_0.xb_hv.n0 level_shifter_up_0.xb_hv.t14 132.101
R12968 level_shifter_up_0.xb_hv.n0 level_shifter_up_0.xb_hv.t12 129.855
R12969 level_shifter_up_0.xb_hv.n1 level_shifter_up_0.xb_hv.t6 129.816
R12970 level_shifter_up_0.xb_hv.n8 level_shifter_up_0.xb_hv.t9 127.45
R12971 level_shifter_up_0.xb_hv.n9 level_shifter_up_0.xb_hv.t15 127.45
R12972 level_shifter_up_0.xb_hv.n7 level_shifter_up_0.xb_hv.t16 127.45
R12973 level_shifter_up_0.xb_hv.n1 level_shifter_up_0.xb_hv.t17 66.731
R12974 level_shifter_up_0.xb_hv.n18 level_shifter_up_0.xb_hv.t3 66.726
R12975 level_shifter_up_0.xb_hv.n0 level_shifter_up_0.xb_hv.t18 66.085
R12976 level_shifter_up_0.xb_hv.n3 level_shifter_up_0.xb_hv.t8 66.069
R12977 level_shifter_up_0.xb_hv.n2 level_shifter_up_0.xb_hv.t10 66.068
R12978 level_shifter_up_0.xb_hv.n1 level_shifter_up_0.xb_hv.t13 66.065
R12979 level_shifter_up_0.xb_hv.n18 level_shifter_up_0.xb_hv.t7 66.057
R12980 level_shifter_up_0.xb_hv.n2 level_shifter_up_0.xb_hv.t11 66.009
R12981 level_shifter_up_0.xb_hv.n10 level_shifter_up_0.xb_hv.t5 65.149
R12982 level_shifter_up_0.xb_hv level_shifter_up_0.xb_hv.t1 17.195
R12983 hyst1b_hv level_shifter_up_0.xb_hv.n18 13.918
R12984 level_shifter_up_0.xb_hv.n10 level_shifter_up_0.xb_hv.t0 13.866
R12985 level_shifter_up_0.xb_hv.n3 level_shifter_up_0.xb_hv.n7 4.654
R12986 level_shifter_up_0.xb_hv.n0 level_shifter_up_0.xb_hv.n9 4.653
R12987 level_shifter_up_0.xb_hv.n2 level_shifter_up_0.xb_hv.n8 4.651
R12988 level_shifter_up_0.xb_hv.n3 level_shifter_up_0.xb_hv.n16 4.5
R12989 level_shifter_up_0.xb_hv.n0 level_shifter_up_0.xb_hv.n15 4.5
R12990 level_shifter_up_0.xb_hv.n0 level_shifter_up_0.xb_hv.n14 4.5
R12991 level_shifter_up_0.xb_hv.n2 level_shifter_up_0.xb_hv.n13 4.5
R12992 level_shifter_up_0.xb_hv.n2 level_shifter_up_0.xb_hv.n17 4.5
R12993 level_shifter_up_0.xb_hv.n1 level_shifter_up_0.xb_hv.n12 4.5
R12994 hyst1b_hv level_shifter_up_0.xb_hv.n11 2.126
R12995 level_shifter_up_0.xb_hv.n11 level_shifter_up_0.xb_hv.n10 0.46
R12996 level_shifter_up_0.xb_hv.n0 level_shifter_up_0.xb_hv.n5 0.436
R12997 level_shifter_up_0.xb_hv.n2 level_shifter_up_0.xb_hv.n6 0.41
R12998 level_shifter_up_0.xb_hv.n18 level_shifter_up_0.xb_hv.n1 0.39
R12999 level_shifter_up_0.xb_hv.n11 level_shifter_up_0.xb_hv 0.321
R13000 level_shifter_up_0.xb_hv.n0 level_shifter_up_0.xb_hv.n3 0.279
R13001 level_shifter_up_0.xb_hv.n1 level_shifter_up_0.xb_hv.n2 0.259
R13002 level_shifter_up_0.xb_hv.n2 level_shifter_up_0.xb_hv.n0 0.256
R13003 level_shifter_up_0.xb_hv.n0 level_shifter_up_0.xb_hv.n4 0.249
R13004 a_32057_n15000.n4 a_32057_n15000.t9 14.718
R13005 a_32057_n15000.n7 a_32057_n15000.t16 14.718
R13006 a_32057_n15000.n8 a_32057_n15000.t1 14.718
R13007 a_32057_n15000.n11 a_32057_n15000.t8 14.718
R13008 a_32057_n15000.n12 a_32057_n15000.t4 14.718
R13009 a_32057_n15000.n15 a_32057_n15000.t10 14.718
R13010 a_32057_n15000.n6 a_32057_n15000.t3 13.849
R13011 a_32057_n15000.n5 a_32057_n15000.t15 13.849
R13012 a_32057_n15000.n4 a_32057_n15000.t12 13.849
R13013 a_32057_n15000.n7 a_32057_n15000.t7 13.849
R13014 a_32057_n15000.n10 a_32057_n15000.t2 13.849
R13015 a_32057_n15000.n9 a_32057_n15000.t6 13.849
R13016 a_32057_n15000.n8 a_32057_n15000.t11 13.849
R13017 a_32057_n15000.n11 a_32057_n15000.t14 13.849
R13018 a_32057_n15000.n14 a_32057_n15000.t5 13.849
R13019 a_32057_n15000.n13 a_32057_n15000.t17 13.849
R13020 a_32057_n15000.n12 a_32057_n15000.t13 13.849
R13021 a_32057_n15000.n15 a_32057_n15000.t0 13.849
R13022 a_32057_n15000.n1 a_32057_n15000.t23 13.847
R13023 a_32057_n15000.n1 a_32057_n15000.t33 13.847
R13024 a_32057_n15000.n2 a_32057_n15000.t27 13.847
R13025 a_32057_n15000.n2 a_32057_n15000.t25 13.847
R13026 a_32057_n15000.n3 a_32057_n15000.t26 13.847
R13027 a_32057_n15000.n3 a_32057_n15000.t31 13.847
R13028 a_32057_n15000.n19 a_32057_n15000.t21 13.847
R13029 a_32057_n15000.n19 a_32057_n15000.t18 13.847
R13030 a_32057_n15000.n20 a_32057_n15000.t24 13.847
R13031 a_32057_n15000.n20 a_32057_n15000.t22 13.847
R13032 a_32057_n15000.n21 a_32057_n15000.t20 13.847
R13033 a_32057_n15000.n21 a_32057_n15000.t28 13.847
R13034 a_32057_n15000.n0 a_32057_n15000.t30 13.847
R13035 a_32057_n15000.n0 a_32057_n15000.t19 13.847
R13036 a_32057_n15000.t32 a_32057_n15000.n29 13.847
R13037 a_32057_n15000.n29 a_32057_n15000.t29 13.847
R13038 a_32057_n15000.n24 a_32057_n15000.n18 12.108
R13039 a_32057_n15000.n17 a_32057_n15000.n16 2.199
R13040 a_32057_n15000.n18 a_32057_n15000.n17 2.199
R13041 a_32057_n15000.n29 a_32057_n15000.n28 1.598
R13042 a_32057_n15000.n22 a_32057_n15000.n21 1.582
R13043 a_32057_n15000.n5 a_32057_n15000.n4 1.325
R13044 a_32057_n15000.n9 a_32057_n15000.n8 1.325
R13045 a_32057_n15000.n13 a_32057_n15000.n12 1.325
R13046 a_32057_n15000.n27 a_32057_n15000.n1 1.098
R13047 a_32057_n15000.n26 a_32057_n15000.n2 1.098
R13048 a_32057_n15000.n25 a_32057_n15000.n3 1.098
R13049 a_32057_n15000.n23 a_32057_n15000.n19 1.098
R13050 a_32057_n15000.n22 a_32057_n15000.n20 1.098
R13051 a_32057_n15000.n28 a_32057_n15000.n0 1.098
R13052 a_32057_n15000.n6 a_32057_n15000.n5 0.869
R13053 a_32057_n15000.n10 a_32057_n15000.n9 0.869
R13054 a_32057_n15000.n14 a_32057_n15000.n13 0.869
R13055 a_32057_n15000.n18 a_32057_n15000.n6 0.759
R13056 a_32057_n15000.n17 a_32057_n15000.n10 0.759
R13057 a_32057_n15000.n16 a_32057_n15000.n14 0.759
R13058 a_32057_n15000.n23 a_32057_n15000.n22 0.5
R13059 a_32057_n15000.n26 a_32057_n15000.n25 0.5
R13060 a_32057_n15000.n27 a_32057_n15000.n26 0.5
R13061 a_32057_n15000.n18 a_32057_n15000.n7 0.495
R13062 a_32057_n15000.n17 a_32057_n15000.n11 0.495
R13063 a_32057_n15000.n16 a_32057_n15000.n15 0.495
R13064 a_32057_n15000.n28 a_32057_n15000.n27 0.489
R13065 a_32057_n15000.n24 a_32057_n15000.n23 0.445
R13066 a_32057_n15000.n25 a_32057_n15000.n24 0.039
R13067 a_2458_6570.n8 a_2458_6570.n7 8.96
R13068 a_2458_6570.n3 a_2458_6570.t10 8.857
R13069 a_2458_6570.n7 a_2458_6570.t11 8.266
R13070 a_2458_6570.n6 a_2458_6570.t8 8.266
R13071 a_2458_6570.n5 a_2458_6570.t9 8.266
R13072 a_2458_6570.n4 a_2458_6570.t6 8.266
R13073 a_2458_6570.n3 a_2458_6570.t7 8.266
R13074 a_2458_6570.n0 a_2458_6570.t2 7.196
R13075 a_2458_6570.t0 a_2458_6570.n11 7.188
R13076 a_2458_6570.n0 a_2458_6570.t3 7.008
R13077 a_2458_6570.n1 a_2458_6570.t4 7.008
R13078 a_2458_6570.n2 a_2458_6570.t13 7.008
R13079 a_2458_6570.n9 a_2458_6570.t1 7
R13080 a_2458_6570.n10 a_2458_6570.t12 7
R13081 a_2458_6570.n11 a_2458_6570.t5 7
R13082 a_2458_6570.n9 a_2458_6570.n8 5.589
R13083 a_2458_6570.n4 a_2458_6570.n3 0.97
R13084 a_2458_6570.n6 a_2458_6570.n5 0.97
R13085 a_2458_6570.n8 a_2458_6570.n2 0.683
R13086 a_2458_6570.n5 a_2458_6570.n4 0.591
R13087 a_2458_6570.n7 a_2458_6570.n6 0.591
R13088 a_2458_6570.n1 a_2458_6570.n0 0.188
R13089 a_2458_6570.n2 a_2458_6570.n1 0.188
R13090 a_2458_6570.n11 a_2458_6570.n10 0.188
R13091 a_2458_6570.n10 a_2458_6570.n9 0.188
R13092 a_32059_n897.n5 a_32059_n897.t2 8.266
R13093 a_32059_n897.n4 a_32059_n897.t7 8.266
R13094 a_32059_n897.n4 a_32059_n897.t3 8.266
R13095 a_32059_n897.n3 a_32059_n897.t6 8.266
R13096 a_32059_n897.n3 a_32059_n897.t4 8.266
R13097 a_32059_n897.n2 a_32059_n897.t9 8.266
R13098 a_32059_n897.n2 a_32059_n897.t5 8.266
R13099 a_32059_n897.n1 a_32059_n897.t8 8.266
R13100 a_32059_n897.n1 a_32059_n897.t1 8.266
R13101 a_32059_n897.n0 a_32059_n897.t0 8.266
R13102 a_32059_n897.n0 a_32059_n897.t11 8.266
R13103 a_32059_n897.t10 a_32059_n897.n5 8.266
R13104 a_32059_n897.n2 a_32059_n897.n1 0.687
R13105 a_32059_n897.n4 a_32059_n897.n3 0.687
R13106 a_32059_n897.n1 a_32059_n897.n0 0.365
R13107 a_32059_n897.n3 a_32059_n897.n2 0.365
R13108 a_32059_n897.n5 a_32059_n897.n4 0.365
R13109 Vinp.n110 Vinp.t4 150.133
R13110 Vinp.n55 Vinp.t20 149.252
R13111 Vinp.n64 Vinp.t33 140.488
R13112 Vinp.n7 Vinp.t32 140.028
R13113 Vinp.n62 Vinp.t28 139.094
R13114 Vinp.n68 Vinp.t22 139.094
R13115 Vinp.n65 Vinp.t42 139.094
R13116 Vinp.n74 Vinp.t54 139.094
R13117 Vinp.n76 Vinp.t27 139.094
R13118 Vinp.n78 Vinp.t10 139.094
R13119 Vinp.n84 Vinp.t6 139.094
R13120 Vinp.n82 Vinp.t31 139.094
R13121 Vinp.n90 Vinp.t15 139.094
R13122 Vinp.n92 Vinp.t53 139.094
R13123 Vinp.n94 Vinp.t35 139.094
R13124 Vinp.n110 Vinp.t40 139.094
R13125 Vinp.n96 Vinp.t18 139.094
R13126 Vinp.n105 Vinp.t39 139.094
R13127 Vinp.n98 Vinp.t30 139.094
R13128 Vinp.n99 Vinp.t5 139.094
R13129 Vinp.n106 Vinp.t16 139.094
R13130 Vinp.n104 Vinp.t26 139.094
R13131 Vinp.n108 Vinp.t1 139.094
R13132 Vinp.n101 Vinp.t48 139.094
R13133 Vinp.n88 Vinp.t11 139.094
R13134 Vinp.n80 Vinp.t21 139.094
R13135 Vinp.n86 Vinp.t49 139.094
R13136 Vinp.n72 Vinp.t47 139.094
R13137 Vinp.n70 Vinp.t7 139.094
R13138 Vinp.n58 Vinp.t56 139.094
R13139 Vinp.n49 Vinp.t43 138.461
R13140 Vinp.n15 Vinp.t45 138.461
R13141 Vinp.n1 Vinp.t51 138.461
R13142 Vinp.n11 Vinp.t19 138.29
R13143 Vinp.n8 Vinp.t41 138.29
R13144 Vinp.n16 Vinp.t55 138.29
R13145 Vinp.n18 Vinp.t29 138.29
R13146 Vinp.n20 Vinp.t38 138.29
R13147 Vinp.n27 Vinp.t9 138.29
R13148 Vinp.n25 Vinp.t34 138.29
R13149 Vinp.n23 Vinp.t23 138.29
R13150 Vinp.n32 Vinp.t13 138.29
R13151 Vinp.n34 Vinp.t24 138.29
R13152 Vinp.n36 Vinp.t2 138.29
R13153 Vinp.n38 Vinp.t8 138.29
R13154 Vinp.n44 Vinp.t17 138.29
R13155 Vinp.n43 Vinp.t46 138.29
R13156 Vinp.n41 Vinp.t37 138.29
R13157 Vinp.n50 Vinp.t50 138.29
R13158 Vinp.n51 Vinp.t36 138.29
R13159 Vinp.n52 Vinp.t3 138.29
R13160 Vinp.n55 Vinp.t12 138.29
R13161 Vinp.n46 Vinp.t25 138.29
R13162 Vinp.n29 Vinp.t14 138.29
R13163 Vinp.n13 Vinp.t0 138.29
R13164 Vinp.n4 Vinp.t44 138.29
R13165 Vinp.n32 Vinp.t52 132.598
R13166 Vinp Vinp.n111 16.797
R13167 Vinp Vinp.n56 12.157
R13168 Vinp.n51 Vinp.n50 4.698
R13169 Vinp.n3 Vinp.n2 4.698
R13170 Vinp.n106 Vinp.n105 4.698
R13171 Vinp.n60 Vinp.n59 4.698
R13172 Vinp.n95 Vinp.n94 3.877
R13173 Vinp.n87 Vinp.n86 3.877
R13174 Vinp.n79 Vinp.n78 3.877
R13175 Vinp.n63 Vinp.n57 3.497
R13176 Vinp.n31 Vinp.n30 3.252
R13177 Vinp.n40 Vinp.n39 3.252
R13178 Vinp.n22 Vinp.n21 3.252
R13179 Vinp.n52 Vinp.n51 3.132
R13180 Vinp.n2 Vinp.n1 3.132
R13181 Vinp.n105 Vinp.n104 3.132
R13182 Vinp.n61 Vinp.n60 3.132
R13183 Vinp.n50 Vinp.n49 2.96
R13184 Vinp.n38 Vinp.n37 2.96
R13185 Vinp.n34 Vinp.n33 2.96
R13186 Vinp.n25 Vinp.n24 2.96
R13187 Vinp.n29 Vinp.n28 2.96
R13188 Vinp.n20 Vinp.n19 2.96
R13189 Vinp.n16 Vinp.n15 2.96
R13190 Vinp.n4 Vinp.n3 2.96
R13191 Vinp.n107 Vinp.n106 2.96
R13192 Vinp.n93 Vinp.n92 2.96
R13193 Vinp.n89 Vinp.n88 2.96
R13194 Vinp.n81 Vinp.n80 2.96
R13195 Vinp.n85 Vinp.n84 2.96
R13196 Vinp.n77 Vinp.n76 2.96
R13197 Vinp.n73 Vinp.n72 2.96
R13198 Vinp.n59 Vinp.n58 2.96
R13199 Vinp.n6 Vinp.n0 2.742
R13200 Vinp.n103 Vinp.n102 2.483
R13201 Vinp.n111 Vinp.n110 2.353
R13202 Vinp.n109 Vinp.n108 2.311
R13203 Vinp.n71 Vinp.n70 2.311
R13204 Vinp.n63 Vinp.n62 2.311
R13205 Vinp.n14 Vinp.n13 1.858
R13206 Vinp.n56 Vinp.n55 1.858
R13207 Vinp.n47 Vinp.n46 1.738
R13208 Vinp.n42 Vinp.n41 1.738
R13209 Vinp.n45 Vinp.n44 1.738
R13210 Vinp.n9 Vinp.n8 1.738
R13211 Vinp.n12 Vinp.n11 1.738
R13212 Vinp.n101 Vinp.n100 1.738
R13213 Vinp.n98 Vinp.n97 1.738
R13214 Vinp.n65 Vinp.n64 1.738
R13215 Vinp.n68 Vinp.n67 1.738
R13216 Vinp.n70 Vinp.n69 1.738
R13217 Vinp.n48 Vinp.n47 1.686
R13218 Vinp.n54 Vinp.n53 1.686
R13219 Vinp.n6 Vinp.n5 1.686
R13220 Vinp.n44 Vinp.n43 1.566
R13221 Vinp.n10 Vinp.n9 1.566
R13222 Vinp.n99 Vinp.n98 1.566
R13223 Vinp.n67 Vinp.n66 1.566
R13224 Vinp.n43 Vinp.n42 1.394
R13225 Vinp.n46 Vinp.n45 1.394
R13226 Vinp.n36 Vinp.n35 1.394
R13227 Vinp.n27 Vinp.n26 1.394
R13228 Vinp.n18 Vinp.n17 1.394
R13229 Vinp.n8 Vinp.n7 1.394
R13230 Vinp.n11 Vinp.n10 1.394
R13231 Vinp.n13 Vinp.n12 1.394
R13232 Vinp.n100 Vinp.n99 1.394
R13233 Vinp.n97 Vinp.n96 1.394
R13234 Vinp.n102 Vinp.n101 1.394
R13235 Vinp.n91 Vinp.n90 1.394
R13236 Vinp.n83 Vinp.n82 1.394
R13237 Vinp.n75 Vinp.n74 1.394
R13238 Vinp.n66 Vinp.n65 1.394
R13239 Vinp.n69 Vinp.n68 1.394
R13240 Vinp.n14 Vinp.n6 1.014
R13241 Vinp.n22 Vinp.n14 1.014
R13242 Vinp.n31 Vinp.n22 1.014
R13243 Vinp.n40 Vinp.n31 1.014
R13244 Vinp.n48 Vinp.n40 1.014
R13245 Vinp.n54 Vinp.n48 1.014
R13246 Vinp.n56 Vinp.n54 1.014
R13247 Vinp.n71 Vinp.n63 1.014
R13248 Vinp.n79 Vinp.n71 1.014
R13249 Vinp.n87 Vinp.n79 1.014
R13250 Vinp.n95 Vinp.n87 1.014
R13251 Vinp.n103 Vinp.n95 1.014
R13252 Vinp.n109 Vinp.n103 1.014
R13253 Vinp.n111 Vinp.n109 1.014
R13254 Vinp.n53 Vinp.n52 0.171
R13255 Vinp.n39 Vinp.n38 0.171
R13256 Vinp.n37 Vinp.n36 0.171
R13257 Vinp.n35 Vinp.n34 0.171
R13258 Vinp.n33 Vinp.n32 0.171
R13259 Vinp.n24 Vinp.n23 0.171
R13260 Vinp.n26 Vinp.n25 0.171
R13261 Vinp.n28 Vinp.n27 0.171
R13262 Vinp.n30 Vinp.n29 0.171
R13263 Vinp.n21 Vinp.n20 0.171
R13264 Vinp.n19 Vinp.n18 0.171
R13265 Vinp.n17 Vinp.n16 0.171
R13266 Vinp.n5 Vinp.n4 0.171
R13267 Vinp.n108 Vinp.n107 0.171
R13268 Vinp.n94 Vinp.n93 0.171
R13269 Vinp.n92 Vinp.n91 0.171
R13270 Vinp.n90 Vinp.n89 0.171
R13271 Vinp.n82 Vinp.n81 0.171
R13272 Vinp.n84 Vinp.n83 0.171
R13273 Vinp.n86 Vinp.n85 0.171
R13274 Vinp.n78 Vinp.n77 0.171
R13275 Vinp.n76 Vinp.n75 0.171
R13276 Vinp.n74 Vinp.n73 0.171
R13277 Vinp.n62 Vinp.n61 0.171
R13278 bias_var_n.n9 bias_var_n.n45 21.009
R13279 bias_var_n.n43 bias_var_n.t3 14.676
R13280 bias_var_n.n44 bias_var_n.t5 13.849
R13281 bias_var_n.n45 bias_var_n.t4 13.849
R13282 bias_var_n.n43 bias_var_n.t2 13.849
R13283 bias_var_n.n42 bias_var_n.t59 12.058
R13284 bias_var_n.n9 bias_var_n.t25 12.05
R13285 bias_var_n.n9 bias_var_n.t56 12.05
R13286 bias_var_n.n10 bias_var_n.t52 12.05
R13287 bias_var_n.n10 bias_var_n.t26 12.05
R13288 bias_var_n.n11 bias_var_n.t54 12.05
R13289 bias_var_n.n11 bias_var_n.t24 12.05
R13290 bias_var_n.n12 bias_var_n.t51 12.05
R13291 bias_var_n.n12 bias_var_n.t15 12.05
R13292 bias_var_n.n13 bias_var_n.t33 12.05
R13293 bias_var_n.n13 bias_var_n.t20 12.05
R13294 bias_var_n.n14 bias_var_n.t23 12.05
R13295 bias_var_n.n14 bias_var_n.t9 12.05
R13296 bias_var_n.n15 bias_var_n.t7 12.05
R13297 bias_var_n.n15 bias_var_n.t46 12.05
R13298 bias_var_n.n16 bias_var_n.t58 12.05
R13299 bias_var_n.n16 bias_var_n.t29 12.05
R13300 bias_var_n.n17 bias_var_n.t41 12.05
R13301 bias_var_n.n17 bias_var_n.t28 12.05
R13302 bias_var_n.n18 bias_var_n.t32 12.05
R13303 bias_var_n.n18 bias_var_n.t18 12.05
R13304 bias_var_n.n19 bias_var_n.t30 12.05
R13305 bias_var_n.n19 bias_var_n.t53 12.05
R13306 bias_var_n.n20 bias_var_n.t22 12.05
R13307 bias_var_n.n20 bias_var_n.t49 12.05
R13308 bias_var_n.n21 bias_var_n.t50 12.05
R13309 bias_var_n.n21 bias_var_n.t14 12.05
R13310 bias_var_n.n22 bias_var_n.t17 12.05
R13311 bias_var_n.n22 bias_var_n.t62 12.05
R13312 bias_var_n.n23 bias_var_n.t27 12.05
R13313 bias_var_n.n23 bias_var_n.t13 12.05
R13314 bias_var_n.n24 bias_var_n.t42 12.05
R13315 bias_var_n.n24 bias_var_n.t11 12.05
R13316 bias_var_n.n25 bias_var_n.t12 12.05
R13317 bias_var_n.n25 bias_var_n.t45 12.05
R13318 bias_var_n.n26 bias_var_n.t60 12.05
R13319 bias_var_n.n26 bias_var_n.t38 12.05
R13320 bias_var_n.n27 bias_var_n.t63 12.05
R13321 bias_var_n.n27 bias_var_n.t43 12.05
R13322 bias_var_n.n28 bias_var_n.t61 12.05
R13323 bias_var_n.n28 bias_var_n.t36 12.05
R13324 bias_var_n.n29 bias_var_n.t37 12.05
R13325 bias_var_n.n29 bias_var_n.t57 12.05
R13326 bias_var_n.n30 bias_var_n.t35 12.05
R13327 bias_var_n.n30 bias_var_n.t21 12.05
R13328 bias_var_n.n31 bias_var_n.t44 12.05
R13329 bias_var_n.n31 bias_var_n.t31 12.05
R13330 bias_var_n.n32 bias_var_n.t39 12.05
R13331 bias_var_n.n32 bias_var_n.t10 12.05
R13332 bias_var_n.n33 bias_var_n.t8 12.05
R13333 bias_var_n.n33 bias_var_n.t40 12.05
R13334 bias_var_n.n34 bias_var_n.t19 12.05
R13335 bias_var_n.n34 bias_var_n.t48 12.05
R13336 bias_var_n.n35 bias_var_n.t16 12.05
R13337 bias_var_n.n35 bias_var_n.t47 12.05
R13338 bias_var_n.n42 bias_var_n.t34 12.05
R13339 bias_var_n.n13 bias_var_n.n36 1.715
R13340 bias_var_n.n44 bias_var_n.n43 1.283
R13341 bias_var_n.n7 bias_var_n.n17 1.142
R13342 bias_var_n.n4 bias_var_n.n18 1.142
R13343 bias_var_n.n6 bias_var_n.n23 1.142
R13344 bias_var_n.n3 bias_var_n.n22 1.142
R13345 bias_var_n.n40 bias_var_n.n25 1.142
R13346 bias_var_n.n3 bias_var_n.n26 1.142
R13347 bias_var_n.n37 bias_var_n.n31 1.142
R13348 bias_var_n.n2 bias_var_n.n30 1.142
R13349 bias_var_n.n29 bias_var_n.n38 1.142
R13350 bias_var_n.n7 bias_var_n.n34 1.142
R13351 bias_var_n.n4 bias_var_n.n33 1.142
R13352 bias_var_n.n32 bias_var_n.n1 1.142
R13353 bias_var_n.n8 bias_var_n.n13 1.142
R13354 bias_var_n.n5 bias_var_n.n14 1.142
R13355 bias_var_n.n35 bias_var_n.n41 1.142
R13356 bias_var_n.n8 bias_var_n.n42 1.142
R13357 bias_var_n.n5 bias_var_n.n11 1.142
R13358 bias_var_n.n10 bias_var_n.n46 1.142
R13359 bias_var_n.n11 bias_var_n.n8 0.881
R13360 bias_var_n.n0 bias_var_n.n20 0.881
R13361 bias_var_n.n7 bias_var_n.n6 0.834
R13362 bias_var_n.n5 bias_var_n.n4 0.834
R13363 bias_var_n.n4 bias_var_n.n3 0.834
R13364 bias_var_n.n3 bias_var_n.n2 0.834
R13365 bias_var_n.n1 bias_var_n.n0 0.834
R13366 bias_var_n.n45 bias_var_n.n44 0.827
R13367 bias_var_n bias_var_n.n5 0.473
R13368 bias_var_n.n4 bias_var_n.n19 0.464
R13369 bias_var_n.n1 bias_var_n.n16 0.464
R13370 bias_var_n.n3 bias_var_n.n21 0.464
R13371 bias_var_n.n25 bias_var_n.n39 0.464
R13372 bias_var_n.n26 bias_var_n.n40 0.464
R13373 bias_var_n.n3 bias_var_n.n27 0.464
R13374 bias_var_n.n0 bias_var_n.n24 0.464
R13375 bias_var_n.n30 bias_var_n.n37 0.464
R13376 bias_var_n.n2 bias_var_n.n29 0.464
R13377 bias_var_n.n38 bias_var_n.n28 0.464
R13378 bias_var_n.n33 bias_var_n.n7 0.464
R13379 bias_var_n.n4 bias_var_n.n32 0.464
R13380 bias_var_n.n1 bias_var_n.n15 0.464
R13381 bias_var_n.n5 bias_var_n.n35 0.464
R13382 bias_var_n.n41 bias_var_n.n12 0.464
R13383 bias_var_n.n5 bias_var_n.n10 0.464
R13384 bias_var_n.n46 bias_var_n.n9 0.464
R13385 a_32057_n8742.n5 a_32057_n8742.t1 13.849
R13386 a_32057_n8742.n4 a_32057_n8742.t0 13.849
R13387 a_32057_n8742.n4 a_32057_n8742.t11 13.849
R13388 a_32057_n8742.n3 a_32057_n8742.t8 13.849
R13389 a_32057_n8742.n3 a_32057_n8742.t5 13.849
R13390 a_32057_n8742.n2 a_32057_n8742.t4 13.849
R13391 a_32057_n8742.n2 a_32057_n8742.t9 13.849
R13392 a_32057_n8742.n1 a_32057_n8742.t3 13.849
R13393 a_32057_n8742.n1 a_32057_n8742.t10 13.849
R13394 a_32057_n8742.n0 a_32057_n8742.t2 13.849
R13395 a_32057_n8742.n0 a_32057_n8742.t7 13.849
R13396 a_32057_n8742.t6 a_32057_n8742.n5 13.849
R13397 a_32057_n8742.n5 a_32057_n8742.n4 0.868
R13398 a_32057_n8742.n2 a_32057_n8742.n1 0.868
R13399 a_32057_n8742.n4 a_32057_n8742.n3 0.464
R13400 a_32057_n8742.n1 a_32057_n8742.n0 0.464
R13401 a_32057_n8742.n5 a_32057_n8742.n2 0.464
R13402 a_32057_n13616.n27 a_32057_n13616.n21 16.083
R13403 a_32057_n13616.n9 a_32057_n13616.t29 14.598
R13404 a_32057_n13616.n4 a_32057_n13616.t25 14.598
R13405 a_32057_n13616.n22 a_32057_n13616.t19 14.598
R13406 a_32057_n13616.n37 a_32057_n13616.t13 14.598
R13407 a_32057_n13616.n35 a_32057_n13616.t15 13.849
R13408 a_32057_n13616.n34 a_32057_n13616.t12 13.849
R13409 a_32057_n13616.n33 a_32057_n13616.t11 13.849
R13410 a_32057_n13616.n32 a_32057_n13616.t14 13.849
R13411 a_32057_n13616.n23 a_32057_n13616.t24 13.849
R13412 a_32057_n13616.n24 a_32057_n13616.t27 13.849
R13413 a_32057_n13616.n25 a_32057_n13616.t18 13.849
R13414 a_32057_n13616.n26 a_32057_n13616.t21 13.849
R13415 a_32057_n13616.n8 a_32057_n13616.t26 13.849
R13416 a_32057_n13616.n7 a_32057_n13616.t9 13.849
R13417 a_32057_n13616.n6 a_32057_n13616.t20 13.849
R13418 a_32057_n13616.n5 a_32057_n13616.t31 13.849
R13419 a_32057_n13616.n9 a_32057_n13616.t17 13.849
R13420 a_32057_n13616.n3 a_32057_n13616.t8 13.849
R13421 a_32057_n13616.n2 a_32057_n13616.t23 13.849
R13422 a_32057_n13616.n1 a_32057_n13616.t28 13.849
R13423 a_32057_n13616.n0 a_32057_n13616.t22 13.849
R13424 a_32057_n13616.n4 a_32057_n13616.t30 13.849
R13425 a_32057_n13616.n22 a_32057_n13616.t10 13.849
R13426 a_32057_n13616.t16 a_32057_n13616.n37 13.849
R13427 a_32057_n13616.n17 a_32057_n13616.t38 6.923
R13428 a_32057_n13616.n17 a_32057_n13616.t6 6.923
R13429 a_32057_n13616.n16 a_32057_n13616.t34 6.923
R13430 a_32057_n13616.n16 a_32057_n13616.t4 6.923
R13431 a_32057_n13616.n15 a_32057_n13616.t1 6.923
R13432 a_32057_n13616.n15 a_32057_n13616.t36 6.923
R13433 a_32057_n13616.n14 a_32057_n13616.t32 6.923
R13434 a_32057_n13616.n14 a_32057_n13616.t37 6.923
R13435 a_32057_n13616.n13 a_32057_n13616.t2 6.923
R13436 a_32057_n13616.n13 a_32057_n13616.t5 6.923
R13437 a_32057_n13616.n12 a_32057_n13616.t33 6.923
R13438 a_32057_n13616.n12 a_32057_n13616.t3 6.923
R13439 a_32057_n13616.n11 a_32057_n13616.t39 6.923
R13440 a_32057_n13616.n11 a_32057_n13616.t0 6.923
R13441 a_32057_n13616.n10 a_32057_n13616.t35 6.923
R13442 a_32057_n13616.n10 a_32057_n13616.t7 6.923
R13443 a_32057_n13616.n32 a_32057_n13616.n31 2.609
R13444 a_32057_n13616.n36 a_32057_n13616.n29 2.199
R13445 a_32057_n13616.n29 a_32057_n13616.n28 2.199
R13446 a_32057_n13616.n28 a_32057_n13616.n27 2.199
R13447 a_32057_n13616.n31 a_32057_n13616.n30 2.199
R13448 a_32057_n13616.n18 a_32057_n13616.n16 1.848
R13449 a_32057_n13616.n19 a_32057_n13616.n14 1.848
R13450 a_32057_n13616.n20 a_32057_n13616.n12 1.848
R13451 a_32057_n13616.n21 a_32057_n13616.n10 1.848
R13452 a_32057_n13616.n18 a_32057_n13616.n17 1.823
R13453 a_32057_n13616.n19 a_32057_n13616.n15 1.823
R13454 a_32057_n13616.n20 a_32057_n13616.n13 1.823
R13455 a_32057_n13616.n21 a_32057_n13616.n11 1.823
R13456 a_32057_n13616.n7 a_32057_n13616.n6 1.159
R13457 a_32057_n13616.n2 a_32057_n13616.n1 1.159
R13458 a_32057_n13616.n25 a_32057_n13616.n24 1.159
R13459 a_32057_n13616.n34 a_32057_n13616.n33 1.159
R13460 a_32057_n13616.n6 a_32057_n13616.n5 0.749
R13461 a_32057_n13616.n8 a_32057_n13616.n7 0.749
R13462 a_32057_n13616.n1 a_32057_n13616.n0 0.749
R13463 a_32057_n13616.n3 a_32057_n13616.n2 0.749
R13464 a_32057_n13616.n26 a_32057_n13616.n25 0.749
R13465 a_32057_n13616.n24 a_32057_n13616.n23 0.749
R13466 a_32057_n13616.n33 a_32057_n13616.n32 0.749
R13467 a_32057_n13616.n35 a_32057_n13616.n34 0.749
R13468 a_32057_n13616.n28 a_32057_n13616.n9 0.685
R13469 a_32057_n13616.n29 a_32057_n13616.n4 0.685
R13470 a_32057_n13616.n27 a_32057_n13616.n22 0.685
R13471 a_32057_n13616.n37 a_32057_n13616.n36 0.685
R13472 a_32057_n13616.n28 a_32057_n13616.n8 0.422
R13473 a_32057_n13616.n29 a_32057_n13616.n3 0.422
R13474 a_32057_n13616.n27 a_32057_n13616.n26 0.422
R13475 a_32057_n13616.n36 a_32057_n13616.n35 0.422
R13476 a_32057_n13616.n21 a_32057_n13616.n20 0.361
R13477 a_32057_n13616.n19 a_32057_n13616.n18 0.361
R13478 a_32057_n13616.n20 a_32057_n13616.n19 0.354
R13479 a_11160_n9542.n4 a_11160_n9542.t6 48.207
R13480 a_11160_n9542.n2 a_11160_n9542.t0 48.207
R13481 a_11160_n9542.n2 a_11160_n9542.t10 48.207
R13482 a_11160_n9542.n3 a_11160_n9542.t4 48.207
R13483 a_11160_n9542.n0 a_11160_n9542.t8 24.204
R13484 a_11160_n9542.n6 a_11160_n9542.t2 24.204
R13485 a_11160_n9542.n0 a_11160_n9542.t12 14.666
R13486 a_11160_n9542.n0 a_11160_n9542.t9 14.124
R13487 a_11160_n9542.n6 a_11160_n9542.t3 14.124
R13488 a_11160_n9542.n0 a_11160_n9542.t7 13.849
R13489 a_11160_n9542.n2 a_11160_n9542.t11 13.849
R13490 a_11160_n9542.n5 a_11160_n9542.t5 13.849
R13491 a_11160_n9542.t1 a_11160_n9542.n10 13.849
R13492 a_11160_n9542.n1 a_11160_n9542.t13 12.05
R13493 a_11160_n9542.n1 a_11160_n9542.t14 12.05
R13494 a_11160_n9542.n1 a_11160_n9542.n8 9.3
R13495 a_11160_n9542.n1 a_11160_n9542.n9 9.3
R13496 a_11160_n9542.n0 a_11160_n9542.n1 1.257
R13497 a_11160_n9542.n10 a_11160_n9542.n0 1.159
R13498 a_11160_n9542.n2 a_11160_n9542.n5 1.159
R13499 a_11160_n9542.n1 a_11160_n9542.n7 1.033
R13500 a_11160_n9542.n2 a_11160_n9542.n4 0.777
R13501 a_11160_n9542.n2 a_11160_n9542.n3 0.777
R13502 a_11160_n9542.n10 a_11160_n9542.n2 0.608
R13503 a_11160_n9542.n3 a_11160_n9542.n6 0.48
R13504 a_11257_n8742.t5 a_11257_n8742.n10 15.074
R13505 a_11257_n8742.n4 a_11257_n8742.t10 14.964
R13506 a_11257_n8742.n10 a_11257_n8742.t2 13.849
R13507 a_11257_n8742.n9 a_11257_n8742.t1 13.849
R13508 a_11257_n8742.n8 a_11257_n8742.t4 13.849
R13509 a_11257_n8742.n0 a_11257_n8742.t3 13.849
R13510 a_11257_n8742.n2 a_11257_n8742.t6 13.849
R13511 a_11257_n8742.n1 a_11257_n8742.t7 13.849
R13512 a_11257_n8742.n3 a_11257_n8742.t0 13.849
R13513 a_11257_n8742.n6 a_11257_n8742.t9 13.849
R13514 a_11257_n8742.n5 a_11257_n8742.t11 13.849
R13515 a_11257_n8742.n4 a_11257_n8742.t8 13.849
R13516 a_11257_n8742.n10 a_11257_n8742.n9 1.909
R13517 a_11257_n8742.n5 a_11257_n8742.n4 1.701
R13518 a_11257_n8742.n7 a_11257_n8742.n6 1.366
R13519 a_11257_n8742.n0 a_11257_n8742.n3 1.225
R13520 a_11257_n8742.n9 a_11257_n8742.n8 1.225
R13521 a_11257_n8742.n6 a_11257_n8742.n5 1.115
R13522 a_11257_n8742.n2 a_11257_n8742.n1 0.948
R13523 a_11257_n8742.n7 a_11257_n8742.n0 0.743
R13524 a_11257_n8742.n8 a_11257_n8742.n7 0.735
R13525 a_11257_n8742.n0 a_11257_n8742.n2 0.355
R13526 level_shifter_up_8.xb_hv.n0 level_shifter_up_8.xb_hv.t8 224.141
R13527 level_shifter_up_8.xb_hv.n1 level_shifter_up_8.xb_hv.t9 224.139
R13528 level_shifter_up_8.xb_hv.n1 level_shifter_up_8.xb_hv.t1 224.139
R13529 level_shifter_up_8.xb_hv.n0 level_shifter_up_8.xb_hv.t4 224.138
R13530 level_shifter_up_8.xb_hv.n0 level_shifter_up_8.xb_hv.t6 223.679
R13531 level_shifter_up_8.xb_hv.n0 level_shifter_up_8.xb_hv.t5 223.679
R13532 level_shifter_up_8.xb_hv.n1 level_shifter_up_8.xb_hv.t3 223.679
R13533 level_shifter_up_8.xb_hv.n1 level_shifter_up_8.xb_hv.t2 223.679
R13534 level_shifter_up_8.xb_hv.n2 level_shifter_up_8.xb_hv.t7 65.02
R13535 level_shifter_up_8.xb_hv.n2 level_shifter_up_8.xb_hv.t0 13.86
R13536 level_shifter_up_8.xb_hv.n2 level_shifter_up_8.xb_hv.n3 10.169
R13537 level_shifter_up_8.xb_hv.n3 level_shifter_up_8.xb_hv.n1 4.6
R13538 level_shifter_up_8.xb_hv level_shifter_up_8.xb_hv.n2 0.733
R13539 level_shifter_up_8.xb_hv.n3 level_shifter_up_8.xb_hv.n0 0.554
R13540 a_2370_6628.n2 a_2370_6628.t9 144.451
R13541 a_2370_6628.n1 a_2370_6628.t11 143.858
R13542 a_2370_6628.n2 a_2370_6628.t10 139.542
R13543 a_2370_6628.n1 a_2370_6628.t8 138.949
R13544 a_2370_6628.n3 a_2370_6628.n2 9.011
R13545 a_2370_6628.n5 a_2370_6628.t7 6.923
R13546 a_2370_6628.n5 a_2370_6628.t6 6.923
R13547 a_2370_6628.n6 a_2370_6628.t5 6.923
R13548 a_2370_6628.n6 a_2370_6628.t4 6.923
R13549 a_2370_6628.n0 a_2370_6628.t3 6.923
R13550 a_2370_6628.n0 a_2370_6628.t2 6.923
R13551 a_2370_6628.n9 a_2370_6628.t1 6.923
R13552 a_2370_6628.t0 a_2370_6628.n9 6.923
R13553 a_2370_6628.n8 a_2370_6628.n7 5.784
R13554 a_2370_6628.n3 a_2370_6628.n1 4.777
R13555 a_2370_6628.n4 a_2370_6628.n3 4.213
R13556 a_2370_6628.n7 a_2370_6628.n6 2.696
R13557 a_2370_6628.n7 a_2370_6628.n5 2.099
R13558 a_2370_6628.n4 a_2370_6628.n0 2.099
R13559 a_2370_6628.n9 a_2370_6628.n8 2.099
R13560 a_2370_6628.n8 a_2370_6628.n4 0.597
R13561 a_23032_4566.n15 a_23032_4566.t4 9.348
R13562 a_23032_4566.n13 a_23032_4566.t7 9.348
R13563 a_23032_4566.n12 a_23032_4566.t17 9.348
R13564 a_23032_4566.n10 a_23032_4566.t16 9.348
R13565 a_23032_4566.n0 a_23032_4566.t10 8.857
R13566 a_23032_4566.n4 a_23032_4566.t13 8.266
R13567 a_23032_4566.n3 a_23032_4566.t11 8.266
R13568 a_23032_4566.n2 a_23032_4566.t14 8.266
R13569 a_23032_4566.n1 a_23032_4566.t12 8.266
R13570 a_23032_4566.n0 a_23032_4566.t9 8.266
R13571 a_23032_4566.n5 a_23032_4566.t6 6.923
R13572 a_23032_4566.n5 a_23032_4566.t5 6.923
R13573 a_23032_4566.n6 a_23032_4566.t15 6.923
R13574 a_23032_4566.n6 a_23032_4566.t18 6.923
R13575 a_23032_4566.n7 a_23032_4566.t8 6.923
R13576 a_23032_4566.n7 a_23032_4566.t0 6.923
R13577 a_23032_4566.n8 a_23032_4566.t2 6.923
R13578 a_23032_4566.n8 a_23032_4566.t1 6.923
R13579 a_23032_4566.t3 a_23032_4566.n4 6.309
R13580 a_23032_4566.n10 a_23032_4566.n9 5.451
R13581 a_23032_4566.n9 a_23032_4566.n8 3.022
R13582 a_23032_4566.n14 a_23032_4566.n5 2.425
R13583 a_23032_4566.n11 a_23032_4566.n6 2.425
R13584 a_23032_4566.n9 a_23032_4566.n7 2.425
R13585 a_23032_4566.t3 a_23032_4566.n15 2.322
R13586 a_23032_4566.n1 a_23032_4566.n0 0.97
R13587 a_23032_4566.n3 a_23032_4566.n2 0.97
R13588 a_23032_4566.n13 a_23032_4566.n12 0.795
R13589 a_23032_4566.n11 a_23032_4566.n10 0.597
R13590 a_23032_4566.n12 a_23032_4566.n11 0.597
R13591 a_23032_4566.n14 a_23032_4566.n13 0.597
R13592 a_23032_4566.n15 a_23032_4566.n14 0.597
R13593 a_23032_4566.n2 a_23032_4566.n1 0.591
R13594 a_23032_4566.n4 a_23032_4566.n3 0.591
R13595 level_shifter_up_5.xb_hv.n4 level_shifter_up_5.xb_hv.t3 66.232
R13596 level_shifter_up_5.xb_hv.n4 level_shifter_up_5.xb_hv.t2 66.111
R13597 level_shifter_up_5.xb_hv.n3 level_shifter_up_5.xb_hv.t4 65.149
R13598 level_shifter_up_5.xb_hv.n3 level_shifter_up_5.xb_hv.t0 13.866
R13599 hyst0b_hv level_shifter_up_5.xb_hv.n5 13.337
R13600 level_shifter_up_5.xb_hv.t8 level_shifter_up_5.xb_hv.n1 66.322
R13601 level_shifter_up_5.xb_hv.t1 hyst0b_hv 3.603
R13602 level_shifter_up_5.xb_hv level_shifter_up_5.xb_hv.n3 0.942
R13603 level_shifter_up_5.xb_hv.n2 level_shifter_up_5.xb_hv.n4 0.011
R13604 level_shifter_up_5.xb_hv.t5 level_shifter_up_5.xb_hv.n2 66.052
R13605 level_shifter_up_5.xb_hv.n0 level_shifter_up_5.xb_hv.n1 0.011
R13606 level_shifter_up_5.xb_hv.n1 level_shifter_up_5.xb_hv.t7 66.022
R13607 level_shifter_up_5.xb_hv.n5 level_shifter_up_5.xb_hv.n2 0.235
R13608 level_shifter_up_5.xb_hv.n5 level_shifter_up_5.xb_hv.n0 0.243
R13609 level_shifter_up_5.xb_hv level_shifter_up_5.xb_hv.t1 0.053
R13610 level_shifter_up_5.xb_hv.n0 level_shifter_up_5.xb_hv.t6 66.093
R13611 a_32057_n9600.n8 a_32057_n9600.n5 17.686
R13612 a_32057_n9600.n7 a_32057_n9600.t6 15.789
R13613 a_32057_n9600.t10 a_32057_n9600.n9 15.773
R13614 a_32057_n9600.n1 a_32057_n9600.t0 14.718
R13615 a_32057_n9600.n2 a_32057_n9600.t5 14.718
R13616 a_32057_n9600.n1 a_32057_n9600.t3 13.849
R13617 a_32057_n9600.n4 a_32057_n9600.t4 13.849
R13618 a_32057_n9600.n3 a_32057_n9600.t1 13.849
R13619 a_32057_n9600.n2 a_32057_n9600.t2 13.849
R13620 a_32057_n9600.n6 a_32057_n9600.t8 13.847
R13621 a_32057_n9600.n6 a_32057_n9600.t7 13.847
R13622 a_32057_n9600.n0 a_32057_n9600.t11 13.847
R13623 a_32057_n9600.n0 a_32057_n9600.t9 13.847
R13624 a_32057_n9600.n3 a_32057_n9600.n2 1.325
R13625 a_32057_n9600.n7 a_32057_n9600.n6 1.106
R13626 a_32057_n9600.n9 a_32057_n9600.n0 1.106
R13627 a_32057_n9600.n4 a_32057_n9600.n3 0.869
R13628 a_32057_n9600.n5 a_32057_n9600.n1 0.759
R13629 a_32057_n9600.n5 a_32057_n9600.n4 0.495
R13630 a_32057_n9600.n9 a_32057_n9600.n8 0.257
R13631 a_32057_n9600.n8 a_32057_n9600.n7 0.242
R13632 trim[5].n0 trim[5].t3 38.514
R13633 trim[5].n1 trim[5].t0 37.895
R13634 trim[5].n0 trim[5].t2 37.185
R13635 trim[5] trim[5].t1 3.676
R13636 trim[5].n2 trim[5] 1.353
R13637 trim[5].n2 trim[5].n1 0.568
R13638 trim[5].n1 trim[5].n0 0.432
R13639 trim[5] trim[5].n2 0.019
R13640 bias_n.n80 bias_n.t88 12.772
R13641 bias_n.n40 bias_n.t6 12.052
R13642 bias_n.n0 bias_n.t25 12.05
R13643 bias_n.n0 bias_n.t68 12.05
R13644 bias_n.n1 bias_n.t55 12.05
R13645 bias_n.n1 bias_n.t29 12.05
R13646 bias_n.n2 bias_n.t51 12.05
R13647 bias_n.n2 bias_n.t15 12.05
R13648 bias_n.n3 bias_n.t79 12.05
R13649 bias_n.n3 bias_n.t37 12.05
R13650 bias_n.n4 bias_n.t58 12.05
R13651 bias_n.n4 bias_n.t40 12.05
R13652 bias_n.n5 bias_n.t35 12.05
R13653 bias_n.n5 bias_n.t81 12.05
R13654 bias_n.n6 bias_n.t21 12.05
R13655 bias_n.n6 bias_n.t66 12.05
R13656 bias_n.n7 bias_n.t20 12.05
R13657 bias_n.n7 bias_n.t71 12.05
R13658 bias_n.n8 bias_n.t23 12.05
R13659 bias_n.n8 bias_n.t65 12.05
R13660 bias_n.n9 bias_n.t73 12.05
R13661 bias_n.n9 bias_n.t34 12.05
R13662 bias_n.n10 bias_n.t56 12.05
R13663 bias_n.n10 bias_n.t19 12.05
R13664 bias_n.n11 bias_n.t52 12.05
R13665 bias_n.n11 bias_n.t26 12.05
R13666 bias_n.n12 bias_n.t50 12.05
R13667 bias_n.n12 bias_n.t12 12.05
R13668 bias_n.n13 bias_n.t13 12.05
R13669 bias_n.n13 bias_n.t48 12.05
R13670 bias_n.n14 bias_n.t18 12.05
R13671 bias_n.n14 bias_n.t83 12.05
R13672 bias_n.n15 bias_n.t32 12.05
R13673 bias_n.n15 bias_n.t11 12.05
R13674 bias_n.n16 bias_n.t84 12.05
R13675 bias_n.n16 bias_n.t41 12.05
R13676 bias_n.n17 bias_n.t10 12.05
R13677 bias_n.n17 bias_n.t77 12.05
R13678 bias_n.n18 bias_n.t82 12.05
R13679 bias_n.n18 bias_n.t63 12.05
R13680 bias_n.n19 bias_n.t42 12.05
R13681 bias_n.n19 bias_n.t75 12.05
R13682 bias_n.n20 bias_n.t30 12.05
R13683 bias_n.n20 bias_n.t72 12.05
R13684 bias_n.n21 bias_n.t61 12.05
R13685 bias_n.n21 bias_n.t33 12.05
R13686 bias_n.n22 bias_n.t60 12.05
R13687 bias_n.n22 bias_n.t22 12.05
R13688 bias_n.n23 bias_n.t76 12.05
R13689 bias_n.n23 bias_n.t36 12.05
R13690 bias_n.n24 bias_n.t86 12.05
R13691 bias_n.n24 bias_n.t43 12.05
R13692 bias_n.n25 bias_n.t44 12.05
R13693 bias_n.n25 bias_n.t78 12.05
R13694 bias_n.n26 bias_n.t38 12.05
R13695 bias_n.n26 bias_n.t69 12.05
R13696 bias_n.n27 bias_n.t80 12.05
R13697 bias_n.n27 bias_n.t57 12.05
R13698 bias_n.n28 bias_n.t9 12.05
R13699 bias_n.n28 bias_n.t74 12.05
R13700 bias_n.n29 bias_n.t27 12.05
R13701 bias_n.n29 bias_n.t8 12.05
R13702 bias_n.n30 bias_n.t16 12.05
R13703 bias_n.n30 bias_n.t49 12.05
R13704 bias_n.n40 bias_n.t4 12.05
R13705 bias_n.n31 bias_n.t59 12.05
R13706 bias_n.n31 bias_n.t46 12.05
R13707 bias_n.n32 bias_n.t31 12.05
R13708 bias_n.n32 bias_n.t62 12.05
R13709 bias_n.n33 bias_n.t45 12.05
R13710 bias_n.n33 bias_n.t87 12.05
R13711 bias_n.n34 bias_n.t85 12.05
R13712 bias_n.n34 bias_n.t64 12.05
R13713 bias_n.n35 bias_n.t24 12.05
R13714 bias_n.n35 bias_n.t53 12.05
R13715 bias_n.n36 bias_n.t54 12.05
R13716 bias_n.n36 bias_n.t17 12.05
R13717 bias_n.n37 bias_n.t67 12.05
R13718 bias_n.n37 bias_n.t39 12.05
R13719 bias_n.n38 bias_n.t28 12.05
R13720 bias_n.n38 bias_n.t70 12.05
R13721 bias_n.n39 bias_n.t47 12.05
R13722 bias_n.n39 bias_n.t14 12.05
R13723 bias_n.n87 bias_n.t0 8.479
R13724 bias_n.n83 bias_n.n82 7.648
R13725 bias_n.n83 bias_n.t7 4.516
R13726 bias_n.n85 bias_n.t1 4.513
R13727 bias_n.n66 bias_n.t3 4.132
R13728 bias_n.n66 bias_n.t2 4.132
R13729 bias_n.n82 bias_n.n81 3.442
R13730 bias_n.n86 bias_n.n85 2.34
R13731 bias_n.n46 bias_n.n9 1.142
R13732 bias_n.n11 bias_n.n96 1.142
R13733 bias_n.n49 bias_n.n15 1.142
R13734 bias_n.n13 bias_n.n100 1.142
R13735 bias_n.n52 bias_n.n17 1.142
R13736 bias_n.n19 bias_n.n104 1.142
R13737 bias_n.n55 bias_n.n23 1.142
R13738 bias_n.n58 bias_n.n5 1.142
R13739 bias_n.n7 bias_n.n112 1.142
R13740 bias_n.n43 bias_n.n28 1.142
R13741 bias_n.n26 bias_n.n92 1.142
R13742 bias_n.n30 bias_n.n118 1.142
R13743 bias_n.n1 bias_n.n123 1.142
R13744 bias_n.n40 bias_n.n89 1.129
R13745 bias_n.n69 bias_n.n32 1.117
R13746 bias_n.n78 bias_n.n35 1.107
R13747 bias_n.n77 bias_n.n37 1.107
R13748 bias_n.n80 bias_n.n39 1.107
R13749 bias_n.n72 bias_n.n34 1.037
R13750 bias_n.n120 bias_n.n25 0.881
R13751 bias_n.n87 bias_n.n86 0.83
R13752 bias_n.n78 bias_n.n77 0.617
R13753 bias_n.n88 bias_n.n87 0.616
R13754 bias_n bias_n.n124 0.517
R13755 bias_n.n69 bias_n.n31 0.5
R13756 bias_n.n72 bias_n.n33 0.5
R13757 bias_n.n78 bias_n.n36 0.5
R13758 bias_n.n77 bias_n.n38 0.5
R13759 bias_n.n40 bias_n.n88 0.467
R13760 bias_n.n46 bias_n.n10 0.464
R13761 bias_n.n97 bias_n.n11 0.464
R13762 bias_n.n96 bias_n.n8 0.464
R13763 bias_n.n49 bias_n.n14 0.464
R13764 bias_n.n101 bias_n.n13 0.464
R13765 bias_n.n100 bias_n.n12 0.464
R13766 bias_n.n52 bias_n.n18 0.464
R13767 bias_n.n105 bias_n.n19 0.464
R13768 bias_n.n104 bias_n.n16 0.464
R13769 bias_n.n55 bias_n.n22 0.464
R13770 bias_n.n107 bias_n.n21 0.464
R13771 bias_n.n111 bias_n.n20 0.464
R13772 bias_n.n58 bias_n.n6 0.464
R13773 bias_n.n113 bias_n.n7 0.464
R13774 bias_n.n112 bias_n.n4 0.464
R13775 bias_n.n116 bias_n.n24 0.464
R13776 bias_n.n43 bias_n.n27 0.464
R13777 bias_n.n93 bias_n.n26 0.464
R13778 bias_n.n92 bias_n.n3 0.464
R13779 bias_n.n60 bias_n.n29 0.464
R13780 bias_n.n120 bias_n.n30 0.464
R13781 bias_n.n118 bias_n.n2 0.464
R13782 bias_n.n124 bias_n.n1 0.464
R13783 bias_n.n123 bias_n.n0 0.464
R13784 bias_n.n86 bias_n.n65 0.417
R13785 bias_n.n65 bias_n.n64 0.417
R13786 bias_n.n64 bias_n.n63 0.417
R13787 bias_n.n63 bias_n.n62 0.417
R13788 bias_n.n62 bias_n.n61 0.417
R13789 bias_n.n118 bias_n.n116 0.417
R13790 bias_n.n112 bias_n.n111 0.417
R13791 bias_n.n88 bias_n.n60 0.417
R13792 bias_n.n88 bias_n.n58 0.417
R13793 bias_n.n58 bias_n.n55 0.417
R13794 bias_n.n55 bias_n.n52 0.417
R13795 bias_n.n52 bias_n.n49 0.417
R13796 bias_n.n49 bias_n.n46 0.417
R13797 bias_n.n46 bias_n.n43 0.417
R13798 bias_n.n124 bias_n.n120 0.417
R13799 bias_n.n124 bias_n.n113 0.417
R13800 bias_n.n113 bias_n.n107 0.417
R13801 bias_n.n107 bias_n.n105 0.417
R13802 bias_n.n105 bias_n.n101 0.417
R13803 bias_n.n101 bias_n.n97 0.417
R13804 bias_n.n97 bias_n.n93 0.417
R13805 bias_n.n84 bias_n.n66 0.417
R13806 bias_n.n82 bias_n.n72 0.349
R13807 bias_n.n81 bias_n.n80 0.349
R13808 bias_n.n82 bias_n.n69 0.259
R13809 bias_n.n81 bias_n.n78 0.259
R13810 bias_n.n39 bias_n.n79 0.246
R13811 bias_n.n38 bias_n.n76 0.246
R13812 bias_n.n37 bias_n.n75 0.246
R13813 bias_n.n36 bias_n.n74 0.246
R13814 bias_n.n35 bias_n.n73 0.246
R13815 bias_n.n34 bias_n.n71 0.246
R13816 bias_n.n33 bias_n.n70 0.246
R13817 bias_n.n32 bias_n.n68 0.246
R13818 bias_n.n31 bias_n.n67 0.246
R13819 bias_n.n30 bias_n.n114 0.246
R13820 bias_n.n29 bias_n.n59 0.246
R13821 bias_n.n28 bias_n.n42 0.246
R13822 bias_n.n27 bias_n.n41 0.246
R13823 bias_n.n26 bias_n.n90 0.246
R13824 bias_n.n25 bias_n.n119 0.246
R13825 bias_n.n24 bias_n.n115 0.246
R13826 bias_n.n23 bias_n.n53 0.246
R13827 bias_n.n22 bias_n.n54 0.246
R13828 bias_n.n21 bias_n.n106 0.246
R13829 bias_n.n20 bias_n.n110 0.246
R13830 bias_n.n19 bias_n.n102 0.246
R13831 bias_n.n18 bias_n.n51 0.246
R13832 bias_n.n17 bias_n.n50 0.246
R13833 bias_n.n16 bias_n.n103 0.246
R13834 bias_n.n15 bias_n.n47 0.246
R13835 bias_n.n14 bias_n.n48 0.246
R13836 bias_n.n13 bias_n.n98 0.246
R13837 bias_n.n12 bias_n.n99 0.246
R13838 bias_n.n11 bias_n.n94 0.246
R13839 bias_n.n10 bias_n.n45 0.246
R13840 bias_n.n9 bias_n.n44 0.246
R13841 bias_n.n8 bias_n.n95 0.246
R13842 bias_n.n7 bias_n.n108 0.246
R13843 bias_n.n6 bias_n.n57 0.246
R13844 bias_n.n5 bias_n.n56 0.246
R13845 bias_n.n4 bias_n.n109 0.246
R13846 bias_n.n3 bias_n.n91 0.246
R13847 bias_n.n2 bias_n.n117 0.246
R13848 bias_n.n1 bias_n.n121 0.246
R13849 bias_n.n0 bias_n.n122 0.246
R13850 bias_n.t5 bias_n.n40 0.167
R13851 bias_n.n84 bias_n.n83 0.141
R13852 bias_n.n85 bias_n.n84 0.141
R13853 bias_n bias_n.t5 0.122
R13854 trim[3].n0 trim[3].t0 38.514
R13855 trim[3].n1 trim[3].t2 37.895
R13856 trim[3].n0 trim[3].t3 37.185
R13857 trim[3] trim[3].t1 3.65
R13858 trim[3].n2 trim[3] 1.34
R13859 trim[3].n2 trim[3].n1 0.6
R13860 trim[3].n1 trim[3].n0 0.432
R13861 trim[3] trim[3].n2 0.013
R13862 a_32057_n14142.n18 a_32057_n14142.t6 13.849
R13863 a_32057_n14142.n17 a_32057_n14142.t12 13.849
R13864 a_32057_n14142.n17 a_32057_n14142.t22 13.849
R13865 a_32057_n14142.n9 a_32057_n14142.t4 13.849
R13866 a_32057_n14142.n9 a_32057_n14142.t32 13.849
R13867 a_32057_n14142.n8 a_32057_n14142.t14 13.849
R13868 a_32057_n14142.n8 a_32057_n14142.t24 13.849
R13869 a_32057_n14142.n7 a_32057_n14142.t0 13.849
R13870 a_32057_n14142.n7 a_32057_n14142.t28 13.849
R13871 a_32057_n14142.n6 a_32057_n14142.t5 13.849
R13872 a_32057_n14142.n6 a_32057_n14142.t33 13.849
R13873 a_32057_n14142.n5 a_32057_n14142.t8 13.849
R13874 a_32057_n14142.n5 a_32057_n14142.t18 13.849
R13875 a_32057_n14142.n4 a_32057_n14142.t2 13.849
R13876 a_32057_n14142.n4 a_32057_n14142.t30 13.849
R13877 a_32057_n14142.n15 a_32057_n14142.t26 13.849
R13878 a_32057_n14142.n15 a_32057_n14142.t16 13.849
R13879 a_32057_n14142.n14 a_32057_n14142.t7 13.849
R13880 a_32057_n14142.n14 a_32057_n14142.t35 13.849
R13881 a_32057_n14142.n13 a_32057_n14142.t11 13.849
R13882 a_32057_n14142.n13 a_32057_n14142.t21 13.849
R13883 a_32057_n14142.n12 a_32057_n14142.t17 13.849
R13884 a_32057_n14142.n12 a_32057_n14142.t27 13.849
R13885 a_32057_n14142.n11 a_32057_n14142.t3 13.849
R13886 a_32057_n14142.n11 a_32057_n14142.t31 13.849
R13887 a_32057_n14142.n10 a_32057_n14142.t13 13.849
R13888 a_32057_n14142.n10 a_32057_n14142.t23 13.849
R13889 a_32057_n14142.n3 a_32057_n14142.t9 13.849
R13890 a_32057_n14142.n3 a_32057_n14142.t19 13.849
R13891 a_32057_n14142.n2 a_32057_n14142.t15 13.849
R13892 a_32057_n14142.n2 a_32057_n14142.t25 13.849
R13893 a_32057_n14142.n1 a_32057_n14142.t1 13.849
R13894 a_32057_n14142.n1 a_32057_n14142.t29 13.849
R13895 a_32057_n14142.n0 a_32057_n14142.t10 13.849
R13896 a_32057_n14142.n0 a_32057_n14142.t20 13.849
R13897 a_32057_n14142.t34 a_32057_n14142.n18 13.849
R13898 a_32057_n14142.n16 a_32057_n14142.n15 2.739
R13899 a_32057_n14142.n17 a_32057_n14142.n16 2.739
R13900 a_32057_n14142.n6 a_32057_n14142.n5 0.868
R13901 a_32057_n14142.n8 a_32057_n14142.n7 0.868
R13902 a_32057_n14142.n12 a_32057_n14142.n11 0.868
R13903 a_32057_n14142.n14 a_32057_n14142.n13 0.868
R13904 a_32057_n14142.n2 a_32057_n14142.n1 0.868
R13905 a_32057_n14142.n18 a_32057_n14142.n3 0.868
R13906 a_32057_n14142.n16 a_32057_n14142.n9 0.54
R13907 a_32057_n14142.n5 a_32057_n14142.n4 0.464
R13908 a_32057_n14142.n7 a_32057_n14142.n6 0.464
R13909 a_32057_n14142.n9 a_32057_n14142.n8 0.464
R13910 a_32057_n14142.n11 a_32057_n14142.n10 0.464
R13911 a_32057_n14142.n13 a_32057_n14142.n12 0.464
R13912 a_32057_n14142.n15 a_32057_n14142.n14 0.464
R13913 a_32057_n14142.n18 a_32057_n14142.n17 0.464
R13914 a_32057_n14142.n1 a_32057_n14142.n0 0.464
R13915 a_32057_n14142.n3 a_32057_n14142.n2 0.464
R13916 level_shifter_up_3.x_hv.n1 level_shifter_up_3.x_hv.t2 193.288
R13917 level_shifter_up_3.x_hv.n0 level_shifter_up_3.x_hv.t8 193.288
R13918 level_shifter_up_3.x_hv.n1 level_shifter_up_3.x_hv.t5 193.285
R13919 level_shifter_up_3.x_hv.n0 level_shifter_up_3.x_hv.t9 193.285
R13920 level_shifter_up_3.x_hv.n1 level_shifter_up_3.x_hv.t6 192.83
R13921 level_shifter_up_3.x_hv.n1 level_shifter_up_3.x_hv.t4 192.83
R13922 level_shifter_up_3.x_hv.n0 level_shifter_up_3.x_hv.t10 192.83
R13923 level_shifter_up_3.x_hv.n0 level_shifter_up_3.x_hv.t7 192.83
R13924 level_shifter_up_3.x_hv.n2 level_shifter_up_3.x_hv.t3 65.176
R13925 level_shifter_up_3.x_hv level_shifter_up_3.x_hv.t0 17.281
R13926 level_shifter_up_3.x_hv.n2 level_shifter_up_3.x_hv.t1 13.85
R13927 level_shifter_up_3.x_hv.n3 level_shifter_up_3.x_hv.n0 4.853
R13928 trim5_hv level_shifter_up_3.x_hv.n3 2.678
R13929 level_shifter_up_3.x_hv trim5_hv 1.714
R13930 level_shifter_up_3.x_hv level_shifter_up_3.x_hv.n2 0.763
R13931 level_shifter_up_3.x_hv.n3 level_shifter_up_3.x_hv.n1 0.636
R13932 a_2370_n28652.n3 a_2370_n28652.t8 142.545
R13933 a_2370_n28652.n4 a_2370_n28652.t9 141.963
R13934 a_2370_n28652.n3 a_2370_n28652.t10 140.969
R13935 a_2370_n28652.n4 a_2370_n28652.t11 140.387
R13936 a_2370_n28652.n5 a_2370_n28652.n4 11.699
R13937 a_2370_n28652.n6 a_2370_n28652.n5 11.25
R13938 a_2370_n28652.n5 a_2370_n28652.n3 7.089
R13939 a_2370_n28652.n1 a_2370_n28652.t5 4.132
R13940 a_2370_n28652.n1 a_2370_n28652.t7 4.132
R13941 a_2370_n28652.n2 a_2370_n28652.t4 4.132
R13942 a_2370_n28652.n2 a_2370_n28652.t6 4.132
R13943 a_2370_n28652.n0 a_2370_n28652.t0 4.132
R13944 a_2370_n28652.n0 a_2370_n28652.t1 4.132
R13945 a_2370_n28652.t3 a_2370_n28652.n9 4.132
R13946 a_2370_n28652.n9 a_2370_n28652.t2 4.132
R13947 a_2370_n28652.n8 a_2370_n28652.n0 2.397
R13948 a_2370_n28652.n7 a_2370_n28652.n1 1.8
R13949 a_2370_n28652.n6 a_2370_n28652.n2 1.8
R13950 a_2370_n28652.n9 a_2370_n28652.n8 1.8
R13951 a_2370_n28652.n8 a_2370_n28652.n7 1.44
R13952 a_2370_n28652.n7 a_2370_n28652.n6 0.607
R13953 Vinm.n110 Vinm.t37 147.437
R13954 Vinm.n55 Vinm.t56 145.662
R13955 Vinm.n96 Vinm.t47 140.946
R13956 Vinm.n41 Vinm.t7 139.57
R13957 Vinm.n62 Vinm.t53 139.552
R13958 Vinm.n82 Vinm.t1 139.552
R13959 Vinm.n84 Vinm.t39 139.552
R13960 Vinm.n92 Vinm.t32 139.552
R13961 Vinm.n90 Vinm.t44 139.552
R13962 Vinm.n97 Vinm.t0 139.552
R13963 Vinm.n100 Vinm.t38 139.552
R13964 Vinm.n106 Vinm.t40 139.552
R13965 Vinm.n105 Vinm.t13 139.552
R13966 Vinm.n110 Vinm.t8 139.552
R13967 Vinm.n104 Vinm.t5 139.552
R13968 Vinm.n108 Vinm.t30 139.552
R13969 Vinm.n102 Vinm.t25 139.552
R13970 Vinm.n88 Vinm.t36 139.552
R13971 Vinm.n94 Vinm.t14 139.552
R13972 Vinm.n86 Vinm.t26 139.552
R13973 Vinm.n80 Vinm.t49 139.552
R13974 Vinm.n64 Vinm.t12 139.552
R13975 Vinm.n74 Vinm.t24 139.552
R13976 Vinm.n66 Vinm.t20 139.552
R13977 Vinm.n67 Vinm.t50 139.552
R13978 Vinm.n76 Vinm.t6 139.552
R13979 Vinm.n72 Vinm.t16 139.552
R13980 Vinm.n78 Vinm.t43 139.552
R13981 Vinm.n69 Vinm.t34 139.552
R13982 Vinm.n58 Vinm.t33 139.552
R13983 Vinm.n49 Vinm.t22 138.003
R13984 Vinm.n33 Vinm.t41 138.003
R13985 Vinm.n1 Vinm.t27 138.003
R13986 Vinm.n4 Vinm.t21 137.832
R13987 Vinm.n10 Vinm.t48 137.832
R13988 Vinm.n9 Vinm.t19 137.832
R13989 Vinm.n7 Vinm.t10 137.832
R13990 Vinm.n24 Vinm.t52 137.832
R13991 Vinm.n36 Vinm.t35 137.832
R13992 Vinm.n34 Vinm.t51 137.832
R13993 Vinm.n42 Vinm.t15 137.832
R13994 Vinm.n45 Vinm.t54 137.832
R13995 Vinm.n51 Vinm.t3 137.832
R13996 Vinm.n50 Vinm.t29 137.832
R13997 Vinm.n55 Vinm.t46 137.832
R13998 Vinm.n52 Vinm.t11 137.832
R13999 Vinm.n47 Vinm.t45 137.832
R14000 Vinm.n38 Vinm.t31 137.832
R14001 Vinm.n21 Vinm.t17 137.832
R14002 Vinm.n28 Vinm.t42 137.832
R14003 Vinm.n19 Vinm.t9 137.832
R14004 Vinm.n26 Vinm.t2 137.832
R14005 Vinm.n17 Vinm.t23 137.832
R14006 Vinm.n30 Vinm.t28 137.832
R14007 Vinm.n15 Vinm.t18 137.832
R14008 Vinm.n12 Vinm.t55 137.832
R14009 Vinm.n24 Vinm.t4 130.574
R14010 Vinm Vinm.n111 16.792
R14011 Vinm Vinm.n56 12.654
R14012 Vinm.n6 Vinm.n0 4.944
R14013 Vinm.n36 Vinm.n35 4.526
R14014 Vinm.n19 Vinm.n18 4.526
R14015 Vinm.n28 Vinm.n27 4.526
R14016 Vinm.n91 Vinm.n90 4.526
R14017 Vinm.n83 Vinm.n82 4.526
R14018 Vinm.n75 Vinm.n74 4.526
R14019 Vinm.n63 Vinm.n57 4.438
R14020 Vinm.n56 Vinm.n55 4.049
R14021 Vinm.n54 Vinm.n53 3.877
R14022 Vinm.n6 Vinm.n5 3.877
R14023 Vinm.n111 Vinm.n110 3.305
R14024 Vinm.n109 Vinm.n108 3.252
R14025 Vinm.n63 Vinm.n62 3.252
R14026 Vinm.n52 Vinm.n51 3.132
R14027 Vinm.n2 Vinm.n1 3.132
R14028 Vinm.n105 Vinm.n104 3.132
R14029 Vinm.n61 Vinm.n60 3.132
R14030 Vinm.n50 Vinm.n49 2.96
R14031 Vinm.n34 Vinm.n33 2.96
R14032 Vinm.n38 Vinm.n37 2.96
R14033 Vinm.n17 Vinm.n16 2.96
R14034 Vinm.n21 Vinm.n20 2.96
R14035 Vinm.n30 Vinm.n29 2.96
R14036 Vinm.n26 Vinm.n25 2.96
R14037 Vinm.n4 Vinm.n3 2.96
R14038 Vinm.n107 Vinm.n106 2.96
R14039 Vinm.n89 Vinm.n88 2.96
R14040 Vinm.n93 Vinm.n92 2.96
R14041 Vinm.n85 Vinm.n84 2.96
R14042 Vinm.n81 Vinm.n80 2.96
R14043 Vinm.n73 Vinm.n72 2.96
R14044 Vinm.n77 Vinm.n76 2.96
R14045 Vinm.n59 Vinm.n58 2.96
R14046 Vinm.n48 Vinm.n47 2.483
R14047 Vinm.n40 Vinm.n39 2.311
R14048 Vinm.n14 Vinm.n13 2.311
R14049 Vinm.n23 Vinm.n22 2.311
R14050 Vinm.n32 Vinm.n31 2.311
R14051 Vinm.n71 Vinm.n70 1.858
R14052 Vinm.n46 Vinm.n45 1.738
R14053 Vinm.n43 Vinm.n42 1.738
R14054 Vinm.n13 Vinm.n12 1.738
R14055 Vinm.n8 Vinm.n7 1.738
R14056 Vinm.n11 Vinm.n10 1.738
R14057 Vinm.n102 Vinm.n101 1.738
R14058 Vinm.n100 Vinm.n99 1.738
R14059 Vinm.n97 Vinm.n96 1.738
R14060 Vinm.n69 Vinm.n68 1.738
R14061 Vinm.n66 Vinm.n65 1.738
R14062 Vinm.n103 Vinm.n102 1.686
R14063 Vinm.n95 Vinm.n94 1.686
R14064 Vinm.n87 Vinm.n86 1.686
R14065 Vinm.n79 Vinm.n78 1.686
R14066 Vinm.n51 Vinm.n50 1.566
R14067 Vinm.n44 Vinm.n43 1.566
R14068 Vinm.n10 Vinm.n9 1.566
R14069 Vinm.n3 Vinm.n2 1.566
R14070 Vinm.n106 Vinm.n105 1.566
R14071 Vinm.n99 Vinm.n98 1.566
R14072 Vinm.n67 Vinm.n66 1.566
R14073 Vinm.n60 Vinm.n59 1.566
R14074 Vinm.n47 Vinm.n46 1.394
R14075 Vinm.n45 Vinm.n44 1.394
R14076 Vinm.n42 Vinm.n41 1.394
R14077 Vinm.n9 Vinm.n8 1.394
R14078 Vinm.n12 Vinm.n11 1.394
R14079 Vinm.n101 Vinm.n100 1.394
R14080 Vinm.n98 Vinm.n97 1.394
R14081 Vinm.n68 Vinm.n67 1.394
R14082 Vinm.n65 Vinm.n64 1.394
R14083 Vinm.n70 Vinm.n69 1.394
R14084 Vinm.n14 Vinm.n6 1.014
R14085 Vinm.n23 Vinm.n14 1.014
R14086 Vinm.n32 Vinm.n23 1.014
R14087 Vinm.n40 Vinm.n32 1.014
R14088 Vinm.n48 Vinm.n40 1.014
R14089 Vinm.n54 Vinm.n48 1.014
R14090 Vinm.n56 Vinm.n54 1.014
R14091 Vinm.n71 Vinm.n63 1.014
R14092 Vinm.n79 Vinm.n71 1.014
R14093 Vinm.n87 Vinm.n79 1.014
R14094 Vinm.n95 Vinm.n87 1.014
R14095 Vinm.n103 Vinm.n95 1.014
R14096 Vinm.n109 Vinm.n103 1.014
R14097 Vinm.n111 Vinm.n109 1.014
R14098 Vinm.n53 Vinm.n52 0.171
R14099 Vinm.n35 Vinm.n34 0.171
R14100 Vinm.n37 Vinm.n36 0.171
R14101 Vinm.n39 Vinm.n38 0.171
R14102 Vinm.n18 Vinm.n17 0.171
R14103 Vinm.n20 Vinm.n19 0.171
R14104 Vinm.n22 Vinm.n21 0.171
R14105 Vinm.n31 Vinm.n30 0.171
R14106 Vinm.n29 Vinm.n28 0.171
R14107 Vinm.n27 Vinm.n26 0.171
R14108 Vinm.n25 Vinm.n24 0.171
R14109 Vinm.n16 Vinm.n15 0.171
R14110 Vinm.n5 Vinm.n4 0.171
R14111 Vinm.n108 Vinm.n107 0.171
R14112 Vinm.n90 Vinm.n89 0.171
R14113 Vinm.n92 Vinm.n91 0.171
R14114 Vinm.n94 Vinm.n93 0.171
R14115 Vinm.n86 Vinm.n85 0.171
R14116 Vinm.n84 Vinm.n83 0.171
R14117 Vinm.n82 Vinm.n81 0.171
R14118 Vinm.n74 Vinm.n73 0.171
R14119 Vinm.n76 Vinm.n75 0.171
R14120 Vinm.n78 Vinm.n77 0.171
R14121 Vinm.n62 Vinm.n61 0.171
R14122 level_shifter_up_4.xb_hv.n2 level_shifter_up_4.xb_hv.t3 219.677
R14123 level_shifter_up_4.xb_hv.n4 level_shifter_up_4.xb_hv.t2 219.328
R14124 level_shifter_up_4.xb_hv.n3 level_shifter_up_4.xb_hv.t9 219.328
R14125 level_shifter_up_4.xb_hv.n2 level_shifter_up_4.xb_hv.t5 219.328
R14126 level_shifter_up_4.xb_hv.t1 level_shifter_up_4.xb_hv.t7 65.004
R14127 level_shifter_up_4.xb_hv.n0 level_shifter_up_4.xb_hv.t10 62.556
R14128 level_shifter_up_4.xb_hv.n0 level_shifter_up_4.xb_hv.t6 61.993
R14129 level_shifter_up_4.xb_hv.n0 level_shifter_up_4.xb_hv.t4 61.993
R14130 level_shifter_up_4.xb_hv.n1 level_shifter_up_4.xb_hv.t8 61.946
R14131 enb_hv level_shifter_up_4.xb_hv.n5 25.827
R14132 level_shifter_up_4.xb_hv level_shifter_up_4.xb_hv.t0 17.195
R14133 level_shifter_up_4.xb_hv.n5 level_shifter_up_4.xb_hv.n1 8.684
R14134 level_shifter_up_4.xb_hv.n5 level_shifter_up_4.xb_hv.n4 7.034
R14135 level_shifter_up_4.xb_hv.t1 level_shifter_up_4.xb_hv 0.751
R14136 enb_hv level_shifter_up_4.xb_hv.t1 0.61
R14137 level_shifter_up_4.xb_hv.n1 level_shifter_up_4.xb_hv.n0 0.573
R14138 level_shifter_up_4.xb_hv.n3 level_shifter_up_4.xb_hv.n2 0.349
R14139 level_shifter_up_4.xb_hv.n4 level_shifter_up_4.xb_hv.n3 0.349
R14140 a_35086_7130.n41 a_35086_7130.t5 409.759
R14141 a_35086_7130.n38 a_35086_7130.t14 233.89
R14142 a_35086_7130.n1 a_35086_7130.t19 96.409
R14143 a_35086_7130.n2 a_35086_7130.t9 96.409
R14144 a_35086_7130.n0 a_35086_7130.t10 96.409
R14145 a_35086_7130.n12 a_35086_7130.t12 48.52
R14146 a_35086_7130.n13 a_35086_7130.t3 48.519
R14147 a_35086_7130.n15 a_35086_7130.t13 48.518
R14148 a_35086_7130.n16 a_35086_7130.t7 48.518
R14149 a_35086_7130.n14 a_35086_7130.t4 48.518
R14150 a_35086_7130.n6 a_35086_7130.t16 48.2
R14151 a_35086_7130.n8 a_35086_7130.t2 48.2
R14152 a_35086_7130.n10 a_35086_7130.t11 48.2
R14153 a_35086_7130.n7 a_35086_7130.t18 48.2
R14154 a_35086_7130.n11 a_35086_7130.t15 48.2
R14155 a_35086_7130.n3 a_35086_7130.t8 48.2
R14156 a_35086_7130.n4 a_35086_7130.t6 48.2
R14157 a_35086_7130.n5 a_35086_7130.t17 48.2
R14158 a_35086_7130.n37 a_35086_7130.t1 17.404
R14159 a_35086_7130.n36 a_35086_7130.n15 14.294
R14160 a_35086_7130.t0 a_35086_7130.n41 14.284
R14161 a_35086_7130.n6 a_35086_7130.n25 9.3
R14162 a_35086_7130.n8 a_35086_7130.n31 9.3
R14163 a_35086_7130.n10 a_35086_7130.n28 9.3
R14164 a_35086_7130.n7 a_35086_7130.n29 9.3
R14165 a_35086_7130.n11 a_35086_7130.n17 9.3
R14166 a_35086_7130.n3 a_35086_7130.n19 9.3
R14167 a_35086_7130.n4 a_35086_7130.n21 9.3
R14168 a_35086_7130.n5 a_35086_7130.n23 9.3
R14169 a_35086_7130.n41 a_35086_7130.n40 4.554
R14170 a_35086_7130.n11 a_35086_7130.n18 4.5
R14171 a_35086_7130.n3 a_35086_7130.n20 4.142
R14172 a_35086_7130.n4 a_35086_7130.n22 3.389
R14173 a_35086_7130.n40 a_35086_7130.n36 2.68
R14174 a_35086_7130.n5 a_35086_7130.n24 2.636
R14175 a_35086_7130.n6 a_35086_7130.n26 1.883
R14176 a_35086_7130.n8 a_35086_7130.n32 1.13
R14177 a_35086_7130.n0 a_35086_7130.n33 0.967
R14178 a_35086_7130.n1 a_35086_7130.n34 0.943
R14179 a_35086_7130.n2 a_35086_7130.n35 0.92
R14180 a_35086_7130.n39 a_35086_7130.n38 0.625
R14181 a_35086_7130.n39 a_35086_7130.n37 0.576
R14182 a_35086_7130.n10 a_35086_7130.n27 0.377
R14183 a_35086_7130.n7 a_35086_7130.n30 0.377
R14184 a_35086_7130.n4 a_35086_7130.n3 0.374
R14185 a_35086_7130.n40 a_35086_7130.n39 0.363
R14186 a_35086_7130.n7 a_35086_7130.n10 0.344
R14187 a_35086_7130.n3 a_35086_7130.n11 0.344
R14188 a_35086_7130.n9 a_35086_7130.n7 0.335
R14189 a_35086_7130.n5 a_35086_7130.n4 0.335
R14190 a_35086_7130.n6 a_35086_7130.n5 0.295
R14191 a_35086_7130.n16 a_35086_7130.n14 0.295
R14192 a_35086_7130.n2 a_35086_7130.n13 0.295
R14193 a_35086_7130.n1 a_35086_7130.n12 0.295
R14194 a_35086_7130.n12 a_35086_7130.n0 0.264
R14195 a_35086_7130.n13 a_35086_7130.n1 0.264
R14196 a_35086_7130.n14 a_35086_7130.n2 0.264
R14197 a_35086_7130.n15 a_35086_7130.n16 0.263
R14198 a_35086_7130.n36 a_35086_7130.n9 0.245
R14199 a_35086_7130.n9 a_35086_7130.n6 0.082
R14200 a_35086_7130.n9 a_35086_7130.n8 0.079
R14201 a_32059_n4755.n18 a_32059_n4755.n17 9.705
R14202 a_32059_n4755.n8 a_32059_n4755.t6 8.857
R14203 a_32059_n4755.n12 a_32059_n4755.t15 8.857
R14204 a_32059_n4755.n11 a_32059_n4755.t13 8.266
R14205 a_32059_n4755.n10 a_32059_n4755.t12 8.266
R14206 a_32059_n4755.n9 a_32059_n4755.t5 8.266
R14207 a_32059_n4755.n8 a_32059_n4755.t14 8.266
R14208 a_32059_n4755.n16 a_32059_n4755.t8 8.266
R14209 a_32059_n4755.n15 a_32059_n4755.t10 8.266
R14210 a_32059_n4755.n14 a_32059_n4755.t9 8.266
R14211 a_32059_n4755.n13 a_32059_n4755.t7 8.266
R14212 a_32059_n4755.n12 a_32059_n4755.t11 8.266
R14213 a_32059_n4755.n0 a_32059_n4755.t2 8.265
R14214 a_32059_n4755.n0 a_32059_n4755.t26 8.265
R14215 a_32059_n4755.n7 a_32059_n4755.t22 8.265
R14216 a_32059_n4755.n7 a_32059_n4755.t20 8.265
R14217 a_32059_n4755.n6 a_32059_n4755.t0 8.265
R14218 a_32059_n4755.n6 a_32059_n4755.t25 8.265
R14219 a_32059_n4755.n5 a_32059_n4755.t18 8.265
R14220 a_32059_n4755.n5 a_32059_n4755.t23 8.265
R14221 a_32059_n4755.n4 a_32059_n4755.t4 8.265
R14222 a_32059_n4755.n4 a_32059_n4755.t16 8.265
R14223 a_32059_n4755.n2 a_32059_n4755.t21 8.265
R14224 a_32059_n4755.n2 a_32059_n4755.t17 8.265
R14225 a_32059_n4755.n1 a_32059_n4755.t1 8.265
R14226 a_32059_n4755.n1 a_32059_n4755.t3 8.265
R14227 a_32059_n4755.t24 a_32059_n4755.n21 8.265
R14228 a_32059_n4755.n21 a_32059_n4755.t19 8.265
R14229 a_32059_n4755.n17 a_32059_n4755.n16 2.581
R14230 a_32059_n4755.n17 a_32059_n4755.n11 1.505
R14231 a_32059_n4755.n18 a_32059_n4755.n7 1.185
R14232 a_32059_n4755.n19 a_32059_n4755.n5 1.185
R14233 a_32059_n4755.n3 a_32059_n4755.n2 1.185
R14234 a_32059_n4755.n21 a_32059_n4755.n20 1.185
R14235 a_32059_n4755.n20 a_32059_n4755.n0 1.177
R14236 a_32059_n4755.n18 a_32059_n4755.n6 1.177
R14237 a_32059_n4755.n19 a_32059_n4755.n4 1.177
R14238 a_32059_n4755.n3 a_32059_n4755.n1 1.177
R14239 a_32059_n4755.n9 a_32059_n4755.n8 0.97
R14240 a_32059_n4755.n11 a_32059_n4755.n10 0.97
R14241 a_32059_n4755.n13 a_32059_n4755.n12 0.97
R14242 a_32059_n4755.n15 a_32059_n4755.n14 0.97
R14243 a_32059_n4755.n20 a_32059_n4755.n3 0.812
R14244 a_32059_n4755.n19 a_32059_n4755.n18 0.812
R14245 a_32059_n4755.n20 a_32059_n4755.n19 0.796
R14246 a_32059_n4755.n10 a_32059_n4755.n9 0.591
R14247 a_32059_n4755.n14 a_32059_n4755.n13 0.591
R14248 a_32059_n4755.n16 a_32059_n4755.n15 0.591
R14249 res_p_bot.n9 res_p_bot.t14 14.598
R14250 res_p_bot.n9 res_p_bot.t15 13.849
R14251 res_p_bot.n10 res_p_bot.n9 9.912
R14252 res_p_bot.n7 res_p_bot.t7 8.356
R14253 res_p_bot.n7 res_p_bot.t8 8.268
R14254 res_p_bot.n5 res_p_bot.t9 6.91
R14255 res_p_bot.n4 res_p_bot.t3 6.91
R14256 res_p_bot.n2 res_p_bot.t2 6.91
R14257 res_p_bot.n12 res_p_bot.t5 6.91
R14258 res_p_bot.n14 res_p_bot.t16 6.91
R14259 res_p_bot.n8 res_p_bot.t13 6.871
R14260 res_p_bot.n15 res_p_bot.n14 5.169
R14261 res_p_bot.n0 res_p_bot.t12 4.132
R14262 res_p_bot.n0 res_p_bot.t0 4.132
R14263 res_p_bot.n1 res_p_bot.t4 4.132
R14264 res_p_bot.n1 res_p_bot.t1 4.132
R14265 res_p_bot.n11 res_p_bot.t11 4.132
R14266 res_p_bot.n11 res_p_bot.t10 4.132
R14267 res_p_bot.n5 res_p_bot.n4 2.961
R14268 res_p_bot.n6 res_p_bot.n0 2.778
R14269 res_p_bot.n3 res_p_bot.n1 2.778
R14270 res_p_bot.n13 res_p_bot.n11 2.778
R14271 res_p_bot res_p_bot.n10 2.303
R14272 res_p_bot.n8 res_p_bot.n7 1.791
R14273 res_p_bot res_p_bot.n15 1.468
R14274 res_p_bot.n13 res_p_bot.n12 0.607
R14275 res_p_bot.n3 res_p_bot.n2 0.597
R14276 res_p_bot.n4 res_p_bot.n3 0.597
R14277 res_p_bot.n6 res_p_bot.n5 0.597
R14278 res_p_bot.n14 res_p_bot.n13 0.586
R14279 res_p_bot.n10 res_p_bot.n8 0.548
R14280 res_p_bot.n8 res_p_bot.n6 0.48
R14281 res_p_bot.n15 res_p_bot.t6 0.329
R14282 Vop_stg2.n1 Vop_stg2.t3 49.549
R14283 Vop_stg2.n2 Vop_stg2.t0 48.422
R14284 Vop_stg2.n0 Vop_stg2.t2 36.428
R14285 Vop_stg2.n1 Vop_stg2.t4 7.121
R14286 Vop_stg2.n0 Vop_stg2.t1 4.157
R14287 Vop_stg2.n2 Vop_stg2.n1 0.741
R14288 Vop_stg2 Vop_stg2.n0 0.442
R14289 Vop_stg2.n0 Vop_stg2.n2 0.264
R14290 a_31098_4670.n3 a_31098_4670.t8 409.142
R14291 a_31098_4670.n3 a_31098_4670.t7 234.473
R14292 a_31098_4670.n7 a_31098_4670.t2 13.057
R14293 a_31098_4670.n7 a_31098_4670.t4 9.275
R14294 a_31098_4670.n6 a_31098_4670.t3 9.275
R14295 a_31098_4670.n0 a_31098_4670.t1 8.413
R14296 a_31098_4670.n9 a_31098_4670.t5 8.265
R14297 a_31098_4670.t6 a_31098_4670.n9 8.265
R14298 a_31098_4670.n2 a_31098_4670.t0 7.141
R14299 a_31098_4670.n9 a_31098_4670.n8 1.01
R14300 a_31098_4670.n0 a_31098_4670.n2 0.802
R14301 a_31098_4670.n8 a_31098_4670.n6 0.363
R14302 a_31098_4670.n8 a_31098_4670.n7 0.363
R14303 a_31098_4670.n5 a_31098_4670.n1 0.305
R14304 a_31098_4670.n4 a_31098_4670.n3 0.25
R14305 a_31098_4670.n6 a_31098_4670.n5 0.21
R14306 a_31098_4670.n1 a_31098_4670.n4 0.156
R14307 a_31098_4670.n1 a_31098_4670.n0 0.081
R14308 Vom_stg2.n0 Vom_stg2.t4 49.543
R14309 Vom_stg2.n1 Vom_stg2.t0 48.423
R14310 Vom_stg2 Vom_stg2.t2 37.023
R14311 Vom_stg2.n0 Vom_stg2.t3 7.134
R14312 Vom_stg2 Vom_stg2.t1 4.132
R14313 Vom_stg2.n1 Vom_stg2.n0 0.747
R14314 Vom_stg2 Vom_stg2.n1 0.641
R14315 a_29757_7018.n0 a_29757_7018.t3 13.847
R14316 a_29757_7018.n0 a_29757_7018.t4 13.847
R14317 a_29757_7018.n1 a_29757_7018.t5 13.847
R14318 a_29757_7018.n1 a_29757_7018.t2 13.847
R14319 a_29757_7018.n2 a_29757_7018.t1 7.746
R14320 a_29757_7018.t0 a_29757_7018.n2 7.389
R14321 a_29757_7018.n0 a_29757_7018.n1 0.894
R14322 a_29757_7018.n2 a_29757_7018.n0 0.886
R14323 a_32059_n4497.n8 a_32059_n4497.t14 8.266
R14324 a_32059_n4497.n7 a_32059_n4497.t2 8.266
R14325 a_32059_n4497.n7 a_32059_n4497.t9 8.266
R14326 a_32059_n4497.n1 a_32059_n4497.t6 8.266
R14327 a_32059_n4497.n1 a_32059_n4497.t13 8.266
R14328 a_32059_n4497.n0 a_32059_n4497.t10 8.266
R14329 a_32059_n4497.n0 a_32059_n4497.t3 8.266
R14330 a_32059_n4497.n5 a_32059_n4497.t4 8.266
R14331 a_32059_n4497.n5 a_32059_n4497.t11 8.266
R14332 a_32059_n4497.n4 a_32059_n4497.t0 8.266
R14333 a_32059_n4497.n4 a_32059_n4497.t15 8.266
R14334 a_32059_n4497.n3 a_32059_n4497.t1 8.266
R14335 a_32059_n4497.n3 a_32059_n4497.t8 8.266
R14336 a_32059_n4497.n2 a_32059_n4497.t5 8.266
R14337 a_32059_n4497.n2 a_32059_n4497.t12 8.266
R14338 a_32059_n4497.t7 a_32059_n4497.n8 8.266
R14339 a_32059_n4497.n6 a_32059_n4497.n1 1.835
R14340 a_32059_n4497.n4 a_32059_n4497.n3 0.687
R14341 a_32059_n4497.n6 a_32059_n4497.n5 0.458
R14342 a_32059_n4497.n1 a_32059_n4497.n0 0.365
R14343 a_32059_n4497.n3 a_32059_n4497.n2 0.365
R14344 a_32059_n4497.n5 a_32059_n4497.n4 0.365
R14345 a_32059_n4497.n8 a_32059_n4497.n7 0.365
R14346 a_32059_n4497.n7 a_32059_n4497.n6 0.228
R14347 level_shifter_up_1.xb_hv.n0 level_shifter_up_1.xb_hv.t1 193.288
R14348 level_shifter_up_1.xb_hv.n0 level_shifter_up_1.xb_hv.t2 193.285
R14349 level_shifter_up_1.xb_hv.n0 level_shifter_up_1.xb_hv.t3 192.83
R14350 level_shifter_up_1.xb_hv.n0 level_shifter_up_1.xb_hv.t4 192.83
R14351 level_shifter_up_1.xb_hv.n2 level_shifter_up_1.xb_hv.t7 65.97
R14352 level_shifter_up_1.xb_hv.n2 level_shifter_up_1.xb_hv.t6 65.939
R14353 level_shifter_up_1.xb_hv.n1 level_shifter_up_1.xb_hv.t5 65.015
R14354 level_shifter_up_1.xb_hv.n1 level_shifter_up_1.xb_hv.t0 13.863
R14355 level_shifter_up_1.xb_hv.n3 level_shifter_up_1.xb_hv.n2 10.618
R14356 trim3b_hv level_shifter_up_1.xb_hv.n3 9.854
R14357 level_shifter_up_1.xb_hv.n1 trim3b_hv 4.783
R14358 level_shifter_up_1.xb_hv.n3 level_shifter_up_1.xb_hv.n0 1.261
R14359 level_shifter_up_1.xb_hv level_shifter_up_1.xb_hv.n1 0.724
R14360 a_27936_n27260.n1 a_27936_n27260.t2 6.203
R14361 a_27936_n27260.t3 a_27936_n27260.n5 5.606
R14362 a_27936_n27260.n2 a_27936_n27260.t4 4.132
R14363 a_27936_n27260.n2 a_27936_n27260.t5 4.132
R14364 a_27936_n27260.n3 a_27936_n27260.t7 4.132
R14365 a_27936_n27260.n3 a_27936_n27260.t6 4.132
R14366 a_27936_n27260.n0 a_27936_n27260.t0 4.132
R14367 a_27936_n27260.n0 a_27936_n27260.t1 4.132
R14368 a_27936_n27260.n4 a_27936_n27260.n3 2.071
R14369 a_27936_n27260.n4 a_27936_n27260.n2 1.474
R14370 a_27936_n27260.n1 a_27936_n27260.n0 1.474
R14371 a_27936_n27260.n5 a_27936_n27260.n4 1.117
R14372 a_27936_n27260.n5 a_27936_n27260.n1 0.607
R14373 a_12857_n14142.n1 a_12857_n14142.t2 13.851
R14374 a_12857_n14142.n3 a_12857_n14142.t0 13.851
R14375 a_12857_n14142.n2 a_12857_n14142.t1 13.849
R14376 a_12857_n14142.n2 a_12857_n14142.t7 13.849
R14377 a_12857_n14142.n1 a_12857_n14142.t4 13.849
R14378 a_12857_n14142.n0 a_12857_n14142.t3 13.849
R14379 a_12857_n14142.n0 a_12857_n14142.t5 13.849
R14380 a_12857_n14142.t6 a_12857_n14142.n3 13.849
R14381 a_12857_n14142.n1 a_12857_n14142.n0 1.121
R14382 a_12857_n14142.n3 a_12857_n14142.n2 1.121
R14383 a_12857_n14142.n2 a_12857_n14142.n1 0.762
R14384 a_25696_11382.n13 a_25696_11382.t11 21.212
R14385 a_25696_11382.n3 a_25696_11382.t7 14.402
R14386 a_25696_11382.n12 a_25696_11382.t9 9.675
R14387 a_25696_11382.n10 a_25696_11382.t0 9.674
R14388 a_25696_11382.n9 a_25696_11382.t12 9.674
R14389 a_25696_11382.n7 a_25696_11382.t13 9.674
R14390 a_25696_11382.n6 a_25696_11382.t5 9.674
R14391 a_25696_11382.n4 a_25696_11382.t4 9.674
R14392 a_25696_11382.n3 a_25696_11382.t8 7.599
R14393 a_25696_11382.n0 a_25696_11382.t10 6.923
R14394 a_25696_11382.n0 a_25696_11382.t2 6.923
R14395 a_25696_11382.n1 a_25696_11382.t15 6.923
R14396 a_25696_11382.n1 a_25696_11382.t14 6.923
R14397 a_25696_11382.n2 a_25696_11382.t6 6.923
R14398 a_25696_11382.n2 a_25696_11382.t3 6.923
R14399 a_25696_11382.n4 a_25696_11382.n3 6.218
R14400 a_25696_11382.n10 a_25696_11382.n9 2.961
R14401 a_25696_11382.n11 a_25696_11382.n0 2.751
R14402 a_25696_11382.n8 a_25696_11382.n1 2.751
R14403 a_25696_11382.n5 a_25696_11382.n2 2.751
R14404 a_25696_11382.n7 a_25696_11382.n6 0.784
R14405 a_25696_11382.n12 a_25696_11382.n11 0.619
R14406 a_25696_11382.n6 a_25696_11382.n5 0.607
R14407 a_25696_11382.n8 a_25696_11382.n7 0.597
R14408 a_25696_11382.n9 a_25696_11382.n8 0.597
R14409 a_25696_11382.n11 a_25696_11382.n10 0.597
R14410 a_25696_11382.n5 a_25696_11382.n4 0.586
R14411 a_25696_11382.n13 a_25696_11382.n12 0.443
R14412 a_25696_11382.t1 a_25696_11382.n13 0.361
R14413 a_11257_n14142.n0 a_11257_n14142.t0 15.112
R14414 a_11257_n14142.n0 a_11257_n14142.t3 14.777
R14415 a_11257_n14142.t2 a_11257_n14142.n0 14.403
R14416 a_11257_n14142.n0 a_11257_n14142.t1 13.85
R14417 a_9060_4530.n2 a_9060_4530.n0 19.412
R14418 a_9060_4530.n3 a_9060_4530.t6 14.842
R14419 a_9060_4530.n3 a_9060_4530.t7 14.842
R14420 a_9060_4530.n4 a_9060_4530.t2 13.851
R14421 a_9060_4530.n6 a_9060_4530.t0 13.851
R14422 a_9060_4530.n5 a_9060_4530.t3 13.849
R14423 a_9060_4530.n5 a_9060_4530.t9 13.849
R14424 a_9060_4530.n4 a_9060_4530.t8 13.849
R14425 a_9060_4530.n1 a_9060_4530.t11 13.849
R14426 a_9060_4530.n1 a_9060_4530.t1 13.849
R14427 a_9060_4530.t10 a_9060_4530.n6 13.849
R14428 a_9060_4530.n0 a_9060_4530.t4 4.428
R14429 a_9060_4530.n0 a_9060_4530.t5 2.066
R14430 a_9060_4530.n5 a_9060_4530.n4 1.121
R14431 a_9060_4530.n4 a_9060_4530.n3 1.062
R14432 a_9060_4530.n6 a_9060_4530.n2 0.905
R14433 a_9060_4530.n6 a_9060_4530.n5 0.762
R14434 a_9060_4530.n2 a_9060_4530.n1 0.183
R14435 a_9060_4172.n1 a_9060_4172.n0 10.477
R14436 a_9060_4172.n0 a_9060_4172.t3 8.857
R14437 a_9060_4172.n0 a_9060_4172.t2 8.266
R14438 a_9060_4172.n1 a_9060_4172.t1 3.187
R14439 a_9060_4172.t0 a_9060_4172.n1 3.187
R14440 level_shifter_up_5.x_hv.n0 level_shifter_up_5.x_hv.t5 65.176
R14441 level_shifter_up_5.x_hv.n1 level_shifter_up_5.x_hv.t4 64.991
R14442 level_shifter_up_5.x_hv.n2 level_shifter_up_5.x_hv.t3 63.577
R14443 level_shifter_up_5.x_hv.n1 level_shifter_up_5.x_hv.t2 63.013
R14444 hyst0_hv level_shifter_up_5.x_hv.n2 25.856
R14445 level_shifter_up_5.x_hv.n3 level_shifter_up_5.x_hv.t1 16.717
R14446 level_shifter_up_5.x_hv.n0 level_shifter_up_5.x_hv.t0 13.85
R14447 level_shifter_up_5.x_hv.n3 hyst0_hv 3.861
R14448 level_shifter_up_5.x_hv level_shifter_up_5.x_hv.n0 0.958
R14449 level_shifter_up_5.x_hv.n2 level_shifter_up_5.x_hv.n1 0.687
R14450 level_shifter_up_5.x_hv level_shifter_up_5.x_hv.n3 0.321
R14451 a_33659_n1551.n2 a_33659_n1551.t3 9.445
R14452 a_33659_n1551.n0 a_33659_n1551.t0 9.194
R14453 a_33659_n1551.n1 a_33659_n1551.t2 8.963
R14454 a_33659_n1551.n0 a_33659_n1551.t1 8.266
R14455 a_33659_n1551.n3 a_33659_n1551.t5 8.265
R14456 a_33659_n1551.t4 a_33659_n1551.n3 8.265
R14457 a_33659_n1551.n2 a_33659_n1551.n1 5.21
R14458 a_33659_n1551.n3 a_33659_n1551.n2 1.168
R14459 a_33659_n1551.n1 a_33659_n1551.n0 0.876
R14460 a_34666_7130.n40 a_34666_7130.t13 409.759
R14461 a_34666_7130.n37 a_34666_7130.t4 233.89
R14462 a_34666_7130.n7 a_34666_7130.t15 96.409
R14463 a_34666_7130.n8 a_34666_7130.t6 96.409
R14464 a_34666_7130.n6 a_34666_7130.t7 96.409
R14465 a_34666_7130.n11 a_34666_7130.t9 48.52
R14466 a_34666_7130.n12 a_34666_7130.t18 48.519
R14467 a_34666_7130.n14 a_34666_7130.t11 48.518
R14468 a_34666_7130.n15 a_34666_7130.t3 48.518
R14469 a_34666_7130.n13 a_34666_7130.t19 48.518
R14470 a_34666_7130.n2 a_34666_7130.t17 48.2
R14471 a_34666_7130.n1 a_34666_7130.t8 48.2
R14472 a_34666_7130.n9 a_34666_7130.t14 48.2
R14473 a_34666_7130.n0 a_34666_7130.t5 48.2
R14474 a_34666_7130.n10 a_34666_7130.t16 48.2
R14475 a_34666_7130.n5 a_34666_7130.t12 48.2
R14476 a_34666_7130.n4 a_34666_7130.t10 48.2
R14477 a_34666_7130.n3 a_34666_7130.t2 48.2
R14478 a_34666_7130.n36 a_34666_7130.t0 17.404
R14479 a_34666_7130.n35 a_34666_7130.n14 14.966
R14480 a_34666_7130.t1 a_34666_7130.n40 14.284
R14481 a_34666_7130.n2 a_34666_7130.n24 9.3
R14482 a_34666_7130.n1 a_34666_7130.n30 9.3
R14483 a_34666_7130.n9 a_34666_7130.n27 9.3
R14484 a_34666_7130.n0 a_34666_7130.n28 9.3
R14485 a_34666_7130.n10 a_34666_7130.n16 9.3
R14486 a_34666_7130.n5 a_34666_7130.n18 9.3
R14487 a_34666_7130.n4 a_34666_7130.n20 9.3
R14488 a_34666_7130.n3 a_34666_7130.n22 9.3
R14489 a_34666_7130.n10 a_34666_7130.n17 4.5
R14490 a_34666_7130.n5 a_34666_7130.n19 4.142
R14491 a_34666_7130.n40 a_34666_7130.n39 4.138
R14492 a_34666_7130.n4 a_34666_7130.n21 3.389
R14493 a_34666_7130.n39 a_34666_7130.n35 2.836
R14494 a_34666_7130.n3 a_34666_7130.n23 2.636
R14495 a_34666_7130.n2 a_34666_7130.n25 1.883
R14496 a_34666_7130.n1 a_34666_7130.n31 1.13
R14497 a_34666_7130.n6 a_34666_7130.n32 0.967
R14498 a_34666_7130.n7 a_34666_7130.n33 0.943
R14499 a_34666_7130.n8 a_34666_7130.n34 0.92
R14500 a_34666_7130.n39 a_34666_7130.n38 0.78
R14501 a_34666_7130.n38 a_34666_7130.n37 0.625
R14502 a_34666_7130.n38 a_34666_7130.n36 0.576
R14503 a_34666_7130.n9 a_34666_7130.n26 0.377
R14504 a_34666_7130.n0 a_34666_7130.n29 0.377
R14505 a_34666_7130.n0 a_34666_7130.n9 0.359
R14506 a_34666_7130.n1 a_34666_7130.n0 0.359
R14507 a_34666_7130.n2 a_34666_7130.n3 0.359
R14508 a_34666_7130.n4 a_34666_7130.n5 0.359
R14509 a_34666_7130.n3 a_34666_7130.n4 0.359
R14510 a_34666_7130.n5 a_34666_7130.n10 0.359
R14511 a_34666_7130.n15 a_34666_7130.n13 0.295
R14512 a_34666_7130.n8 a_34666_7130.n12 0.295
R14513 a_34666_7130.n7 a_34666_7130.n11 0.295
R14514 a_34666_7130.n35 a_34666_7130.n1 0.286
R14515 a_34666_7130.n12 a_34666_7130.n7 0.273
R14516 a_34666_7130.n11 a_34666_7130.n6 0.272
R14517 a_34666_7130.n13 a_34666_7130.n8 0.271
R14518 a_34666_7130.n14 a_34666_7130.n15 0.269
R14519 a_34666_7130.n1 a_34666_7130.n2 0.21
R14520 a_23698_4566.t0 a_23698_4566.t1 5.053
R14521 a_24364_11382.t0 a_24364_11382.t1 5.031
R14522 a_29758_4670.n1 a_29758_4670.t2 96.409
R14523 a_29758_4670.n0 a_29758_4670.t0 96.409
R14524 a_29758_4670.n6 a_29758_4670.t5 48.936
R14525 a_29758_4670.n6 a_29758_4670.t6 48.67
R14526 a_29758_4670.t4 a_29758_4670.n0 13.11
R14527 a_29758_4670.n5 a_29758_4670.t3 7.141
R14528 a_29758_4670.n2 a_29758_4670.t1 7.141
R14529 a_29758_4670.n1 a_29758_4670.n5 1.198
R14530 a_29758_4670.n0 a_29758_4670.n2 1.198
R14531 a_29758_4670.n1 a_29758_4670.n4 0.942
R14532 a_29758_4670.n0 a_29758_4670.n3 0.939
R14533 a_29758_4670.n1 a_29758_4670.n6 0.491
R14534 a_29758_4670.n0 a_29758_4670.n1 0.482
R14535 DVDD.n12 DVDD.n11 224.905
R14536 DVDD.n28 DVDD.n3 224.769
R14537 DVDD.n22 DVDD.n21 224.769
R14538 DVDD.n17 DVDD.n16 224.752
R14539 DVDD.n73 DVDD.n72 149.458
R14540 DVDD.n63 DVDD.n62 149.458
R14541 DVDD.n58 DVDD.n57 149.458
R14542 DVDD.n47 DVDD.n46 149.458
R14543 DVDD.n42 DVDD.n41 149.458
R14544 DVDD.n32 DVDD.n31 149.458
R14545 DVDD.n27 DVDD.t4 98.99
R14546 DVDD.n27 DVDD.t0 98.99
R14547 DVDD.n9 DVDD.t6 98.99
R14548 DVDD.n9 DVDD.n5 90.999
R14549 DVDD.n0 DVDD.t9 15.654
R14550 DVDD.n49 DVDD.t13 15.596
R14551 DVDD.n0 DVDD.t11 14.998
R14552 DVDD.n23 DVDD.t5 7.141
R14553 DVDD.n23 DVDD.t1 7.141
R14554 DVDD.n4 DVDD.t7 7.141
R14555 DVDD.n4 DVDD.t3 7.141
R14556 DVDD.n5 DVDD.t2 5.221
R14557 DVDD.n27 DVDD.n23 1.681
R14558 DVDD.n13 DVDD.n4 1.681
R14559 DVDD DVDD.n74 0.684
R14560 DVDD.n28 DVDD.n27 0.135
R14561 DVDD.n27 DVDD.n22 0.135
R14562 DVDD.n18 DVDD.n13 0.135
R14563 DVDD.n22 DVDD.n18 0.084
R14564 DVDD.n33 DVDD.n28 0.066
R14565 DVDD.n64 DVDD.n59 0.05
R14566 DVDD.n48 DVDD.n43 0.05
R14567 DVDD.n35 DVDD.n34 0.034
R14568 DVDD.t8 DVDD.n35 0.034
R14569 DVDD.n51 DVDD.n50 0.034
R14570 DVDD.t10 DVDD.n51 0.034
R14571 DVDD.n66 DVDD.n65 0.034
R14572 DVDD.t12 DVDD.n66 0.034
R14573 DVDD.n49 DVDD.n0 0.031
R14574 DVDD.n74 DVDD.n70 0.027
R14575 DVDD.n70 DVDD.n64 0.027
R14576 DVDD.n59 DVDD.n54 0.027
R14577 DVDD.n43 DVDD.n38 0.027
R14578 DVDD.n38 DVDD.n33 0.027
R14579 DVDD.n18 DVDD.n17 0.017
R14580 DVDD.n43 DVDD.n42 0.017
R14581 DVDD.n33 DVDD.n32 0.017
R14582 DVDD.n59 DVDD.n58 0.017
R14583 DVDD.n48 DVDD.n47 0.017
R14584 DVDD.n74 DVDD.n73 0.017
R14585 DVDD.n64 DVDD.n63 0.017
R14586 DVDD.n54 DVDD.n49 0.015
R14587 DVDD.n49 DVDD.n48 0.012
R14588 DVDD.n31 DVDD.n30 0.008
R14589 DVDD.n30 DVDD.n29 0.008
R14590 DVDD.n41 DVDD.n40 0.008
R14591 DVDD.n40 DVDD.n39 0.008
R14592 DVDD.n46 DVDD.n45 0.008
R14593 DVDD.n45 DVDD.n44 0.008
R14594 DVDD.n57 DVDD.n56 0.008
R14595 DVDD.n56 DVDD.n55 0.008
R14596 DVDD.n62 DVDD.n61 0.008
R14597 DVDD.n61 DVDD.n60 0.008
R14598 DVDD.n72 DVDD.n71 0.008
R14599 DVDD.n25 DVDD.n24 0.008
R14600 DVDD.n7 DVDD.n6 0.008
R14601 DVDD.n21 DVDD.n20 0.005
R14602 DVDD.n20 DVDD.n19 0.005
R14603 DVDD.n3 DVDD.n2 0.005
R14604 DVDD.n2 DVDD.n1 0.005
R14605 DVDD.n11 DVDD.n10 0.005
R14606 DVDD.n16 DVDD.n15 0.005
R14607 DVDD.n15 DVDD.n14 0.005
R14608 DVDD.n26 DVDD.n25 0.004
R14609 DVDD.n27 DVDD.n26 0.004
R14610 DVDD.n9 DVDD.n8 0.004
R14611 DVDD.n8 DVDD.n7 0.004
R14612 DVDD.n68 DVDD.n67 0.003
R14613 DVDD.n37 DVDD.n36 0.003
R14614 DVDD.n36 DVDD.t8 0.003
R14615 DVDD.n53 DVDD.n52 0.003
R14616 DVDD.n52 DVDD.t10 0.003
R14617 DVDD.n69 DVDD.n68 0.003
R14618 DVDD.n67 DVDD.t12 0.001
R14619 DVDD.n38 DVDD.n37 0.001
R14620 DVDD.n54 DVDD.n53 0.001
R14621 DVDD.n70 DVDD.n69 0.001
R14622 DVDD.n13 DVDD.n12 0.001
R14623 DVDD.n12 DVDD.n9 0.001
R14624 trim[0].n0 trim[0].t1 38.514
R14625 trim[0].n1 trim[0].t3 37.895
R14626 trim[0].n0 trim[0].t2 37.185
R14627 trim[0].n2 trim[0] 5.806
R14628 trim[0] trim[0].t0 3.65
R14629 trim[0].n2 trim[0].n1 0.6
R14630 trim[0].n1 trim[0].n0 0.432
R14631 trim[0] trim[0].n2 0.013
R14632 trim[2].n0 trim[2].t3 38.514
R14633 trim[2].n1 trim[2].t1 37.895
R14634 trim[2].n0 trim[2].t0 37.185
R14635 trim[2].n2 trim[2] 3.867
R14636 trim[2] trim[2].t2 3.65
R14637 trim[2].n2 trim[2].n1 0.6
R14638 trim[2].n1 trim[2].n0 0.432
R14639 trim[2] trim[2].n2 0.013
R14640 a_32059_n3351.n10 a_32059_n3351.t9 9.321
R14641 a_32059_n3351.n2 a_32059_n3351.t15 9.321
R14642 a_32059_n3351.n4 a_32059_n3351.t13 9.194
R14643 a_32059_n3351.n4 a_32059_n3351.t8 8.266
R14644 a_32059_n3351.n10 a_32059_n3351.t12 8.266
R14645 a_32059_n3351.n3 a_32059_n3351.t10 8.266
R14646 a_32059_n3351.n2 a_32059_n3351.t11 8.266
R14647 a_32059_n3351.t14 a_32059_n3351.n12 8.266
R14648 a_32059_n3351.n8 a_32059_n3351.t6 8.265
R14649 a_32059_n3351.n8 a_32059_n3351.t4 8.265
R14650 a_32059_n3351.n7 a_32059_n3351.t3 8.265
R14651 a_32059_n3351.n7 a_32059_n3351.t7 8.265
R14652 a_32059_n3351.n5 a_32059_n3351.t5 8.265
R14653 a_32059_n3351.n5 a_32059_n3351.t2 8.265
R14654 a_32059_n3351.n6 a_32059_n3351.t0 8.265
R14655 a_32059_n3351.n6 a_32059_n3351.t1 8.265
R14656 a_32059_n3351.n9 a_32059_n3351.n1 5.193
R14657 a_32059_n3351.n11 a_32059_n3351.n9 1.831
R14658 a_32059_n3351.n3 a_32059_n3351.n2 1.705
R14659 a_32059_n3351.n0 a_32059_n3351.n8 1.372
R14660 a_32059_n3351.n1 a_32059_n3351.n6 1.372
R14661 a_32059_n3351.n12 a_32059_n3351.n3 1.055
R14662 a_32059_n3351.n0 a_32059_n3351.n7 0.977
R14663 a_32059_n3351.n1 a_32059_n3351.n5 0.977
R14664 a_32059_n3351.n11 a_32059_n3351.n10 0.957
R14665 a_32059_n3351.n9 a_32059_n3351.n4 0.782
R14666 a_32059_n3351.n12 a_32059_n3351.n11 0.621
R14667 a_32059_n3351.n1 a_32059_n3351.n0 0.394
R14668 en.n1 en.t2 38.514
R14669 en.n2 en.t0 37.894
R14670 en.n1 en.t3 37.185
R14671 en.n0 en 3.955
R14672 en.n0 en.t1 3.683
R14673 en en.n2 0.564
R14674 en.n2 en.n1 0.432
R14675 en en.n0 0.017
R14676 a_12857_n15942.n3 a_12857_n15942.t0 13.851
R14677 a_12857_n15942.n2 a_12857_n15942.t3 13.849
R14678 a_12857_n15942.n2 a_12857_n15942.t5 13.849
R14679 a_12857_n15942.n1 a_12857_n15942.t4 13.849
R14680 a_12857_n15942.n1 a_12857_n15942.t2 13.849
R14681 a_12857_n15942.n0 a_12857_n15942.t1 13.849
R14682 a_12857_n15942.n0 a_12857_n15942.t7 13.849
R14683 a_12857_n15942.t6 a_12857_n15942.n3 13.849
R14684 a_12857_n15942.n3 a_12857_n15942.n0 0.946
R14685 a_12857_n15942.n2 a_12857_n15942.n1 0.795
R14686 a_12857_n15942.n3 a_12857_n15942.n2 0.762
R14687 level_shifter_up_0.x_hv.n6 level_shifter_up_0.x_hv.t6 65.176
R14688 level_shifter_up_0.x_hv.n4 level_shifter_up_0.x_hv.t2 63.759
R14689 level_shifter_up_0.x_hv.n5 level_shifter_up_0.x_hv.t4 63.755
R14690 level_shifter_up_0.x_hv.n5 level_shifter_up_0.x_hv.t8 63.738
R14691 level_shifter_up_0.x_hv.n4 level_shifter_up_0.x_hv.t9 63.734
R14692 level_shifter_up_0.x_hv.n2 level_shifter_up_0.x_hv.t7 63.767
R14693 level_shifter_up_0.x_hv.n1 level_shifter_up_0.x_hv.t3 63.744
R14694 hyst1_hv level_shifter_up_0.x_hv.n0 25.012
R14695 level_shifter_up_0.x_hv level_shifter_up_0.x_hv.t0 17.199
R14696 level_shifter_up_0.x_hv.n6 level_shifter_up_0.x_hv.t1 13.85
R14697 level_shifter_up_0.x_hv.n3 level_shifter_up_0.x_hv.t5 63.708
R14698 level_shifter_up_0.x_hv.t10 level_shifter_up_0.x_hv.n1 63.745
R14699 level_shifter_up_0.x_hv.n1 level_shifter_up_0.x_hv.n0 0.168
R14700 level_shifter_up_0.x_hv hyst1_hv 2.265
R14701 level_shifter_up_0.x_hv level_shifter_up_0.x_hv.n6 0.837
R14702 level_shifter_up_0.x_hv.n2 level_shifter_up_0.x_hv.n5 0.489
R14703 level_shifter_up_0.x_hv.n0 level_shifter_up_0.x_hv.n4 0.366
R14704 level_shifter_up_0.x_hv.n3 level_shifter_up_0.x_hv.n2 0.011
R14705 level_shifter_up_0.x_hv.n0 level_shifter_up_0.x_hv.n3 0.349
R14706 level_shifter_up_3.xb_hv.n0 level_shifter_up_3.xb_hv.t4 193.288
R14707 level_shifter_up_3.xb_hv.n2 level_shifter_up_3.xb_hv.t6 193.286
R14708 level_shifter_up_3.xb_hv.n0 level_shifter_up_3.xb_hv.t10 193.285
R14709 level_shifter_up_3.xb_hv.n1 level_shifter_up_3.xb_hv.t5 193.19
R14710 level_shifter_up_3.xb_hv.n1 level_shifter_up_3.xb_hv.t3 192.83
R14711 level_shifter_up_3.xb_hv.n2 level_shifter_up_3.xb_hv.t2 192.83
R14712 level_shifter_up_3.xb_hv.n0 level_shifter_up_3.xb_hv.t7 192.83
R14713 level_shifter_up_3.xb_hv.n0 level_shifter_up_3.xb_hv.t8 192.83
R14714 level_shifter_up_3.xb_hv.n4 level_shifter_up_3.xb_hv.t9 65.149
R14715 level_shifter_up_3.xb_hv level_shifter_up_3.xb_hv.t1 17.301
R14716 level_shifter_up_3.xb_hv.n4 level_shifter_up_3.xb_hv.t0 13.866
R14717 level_shifter_up_3.xb_hv.n3 level_shifter_up_3.xb_hv.n0 4.981
R14718 level_shifter_up_3.xb_hv.n5 trim5b_hv 1.869
R14719 trim5b_hv level_shifter_up_3.xb_hv.n3 0.961
R14720 level_shifter_up_3.xb_hv.n3 level_shifter_up_3.xb_hv.n1 0.646
R14721 level_shifter_up_3.xb_hv.n5 level_shifter_up_3.xb_hv.n4 0.451
R14722 level_shifter_up_3.xb_hv.n1 level_shifter_up_3.xb_hv.n2 0.367
R14723 level_shifter_up_3.xb_hv level_shifter_up_3.xb_hv.n5 0.262
R14724 Vout.n0 Vout.t0 19.391
R14725 Vout.n0 Vout.t1 17.98
R14726 Vout Vout.n0 0.906
R14727 a_32057_n17742.n11 a_32057_n17742.t4 13.849
R14728 a_32057_n17742.n10 a_32057_n17742.t9 13.849
R14729 a_32057_n17742.n10 a_32057_n17742.t15 13.849
R14730 a_32057_n17742.n9 a_32057_n17742.t3 13.849
R14731 a_32057_n17742.n9 a_32057_n17742.t21 13.849
R14732 a_32057_n17742.n8 a_32057_n17742.t6 13.849
R14733 a_32057_n17742.n8 a_32057_n17742.t12 13.849
R14734 a_32057_n17742.n7 a_32057_n17742.t10 13.849
R14735 a_32057_n17742.n7 a_32057_n17742.t16 13.849
R14736 a_32057_n17742.n6 a_32057_n17742.t0 13.849
R14737 a_32057_n17742.n6 a_32057_n17742.t18 13.849
R14738 a_32057_n17742.n5 a_32057_n17742.t7 13.849
R14739 a_32057_n17742.n5 a_32057_n17742.t13 13.849
R14740 a_32057_n17742.n4 a_32057_n17742.t11 13.849
R14741 a_32057_n17742.n4 a_32057_n17742.t17 13.849
R14742 a_32057_n17742.n3 a_32057_n17742.t1 13.849
R14743 a_32057_n17742.n3 a_32057_n17742.t19 13.849
R14744 a_32057_n17742.n2 a_32057_n17742.t5 13.849
R14745 a_32057_n17742.n2 a_32057_n17742.t23 13.849
R14746 a_32057_n17742.n1 a_32057_n17742.t8 13.849
R14747 a_32057_n17742.n1 a_32057_n17742.t14 13.849
R14748 a_32057_n17742.n0 a_32057_n17742.t2 13.849
R14749 a_32057_n17742.n0 a_32057_n17742.t20 13.849
R14750 a_32057_n17742.t22 a_32057_n17742.n11 13.849
R14751 a_32057_n17742.n11 a_32057_n17742.n10 3.376
R14752 a_32057_n17742.n7 a_32057_n17742.n6 0.868
R14753 a_32057_n17742.n9 a_32057_n17742.n8 0.868
R14754 a_32057_n17742.n2 a_32057_n17742.n1 0.868
R14755 a_32057_n17742.n4 a_32057_n17742.n3 0.868
R14756 a_32057_n17742.n6 a_32057_n17742.n5 0.464
R14757 a_32057_n17742.n8 a_32057_n17742.n7 0.464
R14758 a_32057_n17742.n10 a_32057_n17742.n9 0.464
R14759 a_32057_n17742.n1 a_32057_n17742.n0 0.464
R14760 a_32057_n17742.n3 a_32057_n17742.n2 0.464
R14761 a_32057_n17742.n11 a_32057_n17742.n4 0.464
R14762 a_33659_n2697.n2 a_33659_n2697.t3 8.266
R14763 a_33659_n2697.n1 a_33659_n2697.t1 8.266
R14764 a_33659_n2697.n1 a_33659_n2697.t5 8.266
R14765 a_33659_n2697.n0 a_33659_n2697.t4 8.266
R14766 a_33659_n2697.n0 a_33659_n2697.t0 8.266
R14767 a_33659_n2697.t2 a_33659_n2697.n2 8.266
R14768 a_33659_n2697.n2 a_33659_n2697.n1 0.687
R14769 a_33659_n2697.n1 a_33659_n2697.n0 0.365
R14770 a_12857_n19016.n4 a_12857_n19016.n2 22.014
R14771 a_12857_n19016.n6 a_12857_n19016.t1 14.676
R14772 a_12857_n19016.n5 a_12857_n19016.t3 13.849
R14773 a_12857_n19016.n4 a_12857_n19016.t2 13.849
R14774 a_12857_n19016.t0 a_12857_n19016.n6 13.849
R14775 a_12857_n19016.n2 a_12857_n19016.t6 12.052
R14776 a_12857_n19016.n2 a_12857_n19016.t4 12.05
R14777 a_12857_n19016.n1 a_12857_n19016.t8 12.05
R14778 a_12857_n19016.n1 a_12857_n19016.t12 12.05
R14779 a_12857_n19016.n0 a_12857_n19016.t11 12.05
R14780 a_12857_n19016.n0 a_12857_n19016.t10 12.05
R14781 a_12857_n19016.n3 a_12857_n19016.t9 12.05
R14782 a_12857_n19016.n3 a_12857_n19016.t13 12.05
R14783 a_12857_n19016.n2 a_12857_n19016.t5 8.938
R14784 a_12857_n19016.n2 a_12857_n19016.n1 8.836
R14785 a_12857_n19016.n2 a_12857_n19016.t7 8.652
R14786 a_12857_n19016.n6 a_12857_n19016.n5 1.283
R14787 a_12857_n19016.n5 a_12857_n19016.n4 0.827
R14788 a_12857_n19016.n1 a_12857_n19016.n0 0.703
R14789 a_12857_n19016.n0 a_12857_n19016.n3 0.558
R14790 bias_stg2.n4 bias_stg2.t0 20.406
R14791 bias_stg2.n0 bias_stg2.t4 13.847
R14792 bias_stg2.n0 bias_stg2.t2 13.847
R14793 bias_stg2.n0 bias_stg2.t1 8.601
R14794 bias_stg2.n2 bias_stg2.t3 8.123
R14795 bias_stg2.n3 bias_stg2.t5 8.068
R14796 bias_stg2.n3 bias_stg2.t7 8.068
R14797 bias_stg2.n1 bias_stg2.t8 8.034
R14798 bias_stg2.n1 bias_stg2.t6 8.034
R14799 bias_stg2 bias_stg2.n2 1.942
R14800 bias_stg2.n4 bias_stg2.n1 1.193
R14801 bias_stg2.n2 bias_stg2.n0 0.86
R14802 bias_stg2 bias_stg2.n4 0.847
R14803 bias_stg2.n1 bias_stg2.n3 0.593
R14804 a_2370_7428.n2 a_2370_7428.t9 140.942
R14805 a_2370_7428.n3 a_2370_7428.t11 140.701
R14806 a_2370_7428.n2 a_2370_7428.t10 139.366
R14807 a_2370_7428.n3 a_2370_7428.t8 139.125
R14808 a_2370_7428.n4 a_2370_7428.n3 11.511
R14809 a_2370_7428.n4 a_2370_7428.n2 7.277
R14810 a_2370_7428.n5 a_2370_7428.n4 7.194
R14811 a_2370_7428.n7 a_2370_7428.t0 6.923
R14812 a_2370_7428.n7 a_2370_7428.t2 6.923
R14813 a_2370_7428.n0 a_2370_7428.t5 6.923
R14814 a_2370_7428.n0 a_2370_7428.t4 6.923
R14815 a_2370_7428.n1 a_2370_7428.t7 6.923
R14816 a_2370_7428.n1 a_2370_7428.t6 6.923
R14817 a_2370_7428.n9 a_2370_7428.t1 6.923
R14818 a_2370_7428.t3 a_2370_7428.n9 6.923
R14819 a_2370_7428.n8 a_2370_7428.n7 2.38
R14820 a_2370_7428.n6 a_2370_7428.n0 1.773
R14821 a_2370_7428.n5 a_2370_7428.n1 1.773
R14822 a_2370_7428.n9 a_2370_7428.n8 1.773
R14823 a_2370_7428.n8 a_2370_7428.n6 1.44
R14824 a_2370_7428.n6 a_2370_7428.n5 0.597
R14825 a_12857_n17742.n1 a_12857_n17742.t2 13.851
R14826 a_12857_n17742.n3 a_12857_n17742.t0 13.851
R14827 a_12857_n17742.n2 a_12857_n17742.t1 13.849
R14828 a_12857_n17742.n2 a_12857_n17742.t7 13.849
R14829 a_12857_n17742.n1 a_12857_n17742.t4 13.849
R14830 a_12857_n17742.n0 a_12857_n17742.t3 13.849
R14831 a_12857_n17742.n0 a_12857_n17742.t5 13.849
R14832 a_12857_n17742.t6 a_12857_n17742.n3 13.849
R14833 a_12857_n17742.n1 a_12857_n17742.n0 1.121
R14834 a_12857_n17742.n3 a_12857_n17742.n2 1.121
R14835 a_12857_n17742.n2 a_12857_n17742.n1 0.762
R14836 level_shifter_up_7.x_hv.n0 level_shifter_up_7.x_hv.t6 224.067
R14837 level_shifter_up_7.x_hv.n0 level_shifter_up_7.x_hv.t8 224.061
R14838 level_shifter_up_7.x_hv.n0 level_shifter_up_7.x_hv.t4 223.68
R14839 level_shifter_up_7.x_hv.n0 level_shifter_up_7.x_hv.t7 223.679
R14840 level_shifter_up_7.x_hv.n2 level_shifter_up_7.x_hv.t3 125.496
R14841 level_shifter_up_7.x_hv.n1 level_shifter_up_7.x_hv.t5 125.496
R14842 level_shifter_up_7.x_hv.n5 level_shifter_up_7.x_hv.t2 65.176
R14843 level_shifter_up_7.x_hv.n1 level_shifter_up_7.x_hv.t1 63.646
R14844 level_shifter_up_7.x_hv.n2 level_shifter_up_7.x_hv.t9 63.645
R14845 level_shifter_up_7.x_hv.n4 level_shifter_up_7.x_hv.n3 13.926
R14846 level_shifter_up_7.x_hv.n5 level_shifter_up_7.x_hv.t0 13.85
R14847 level_shifter_up_7.x_hv.n6 level_shifter_up_7.x_hv.n4 4.894
R14848 level_shifter_up_7.x_hv.n3 level_shifter_up_7.x_hv.n2 2.692
R14849 level_shifter_up_7.x_hv.n3 level_shifter_up_7.x_hv.n1 1.694
R14850 level_shifter_up_7.x_hv.n4 level_shifter_up_7.x_hv.n0 0.769
R14851 level_shifter_up_7.x_hv.n6 level_shifter_up_7.x_hv.n5 0.455
R14852 level_shifter_up_7.x_hv level_shifter_up_7.x_hv.n6 0.251
R14853 a_32059_2049.n4 a_32059_2049.t7 8.733
R14854 a_32059_2049.n1 a_32059_2049.t6 8.721
R14855 a_32059_2049.n3 a_32059_2049.t4 8.267
R14856 a_32059_2049.n2 a_32059_2049.t5 8.266
R14857 a_32059_2049.n0 a_32059_2049.t2 8.265
R14858 a_32059_2049.n0 a_32059_2049.t0 8.265
R14859 a_32059_2049.n5 a_32059_2049.t1 8.265
R14860 a_32059_2049.t3 a_32059_2049.n5 8.265
R14861 a_32059_2049.n3 a_32059_2049.n2 1.498
R14862 a_32059_2049.n1 a_32059_2049.n0 1.101
R14863 a_32059_2049.n5 a_32059_2049.n4 1.101
R14864 a_32059_2049.n2 a_32059_2049.n1 0.467
R14865 a_32059_2049.n4 a_32059_2049.n3 0.454
R14866 hyst[1].n1 hyst[1].t1 38.514
R14867 hyst[1].n2 hyst[1].t3 37.894
R14868 hyst[1].n1 hyst[1].t2 37.185
R14869 hyst[1].n0 hyst[1].t0 3.683
R14870 hyst[1].n0 hyst[1] 2.671
R14871 hyst[1] hyst[1].n2 0.564
R14872 hyst[1].n2 hyst[1].n1 0.432
R14873 hyst[1] hyst[1].n0 0.017
R14874 ibias.n2 ibias.t5 51.446
R14875 ibias.n0 ibias.t2 51.437
R14876 ibias.n4 ibias.t6 12.939
R14877 ibias.n0 ibias.t0 12.055
R14878 ibias.n1 ibias.t4 12.05
R14879 ibias.n1 ibias.t3 12.05
R14880 ibias.n0 ibias.t1 8.775
R14881 ibias ibias.n4 3.804
R14882 ibias.n3 ibias.n0 1.371
R14883 ibias.n3 ibias.n2 0.884
R14884 ibias.n4 ibias.n3 0.566
R14885 ibias.n2 ibias.n1 0.002
R14886 a_32059_903.n3 a_32059_903.t5 8.266
R14887 a_32059_903.n2 a_32059_903.t0 8.266
R14888 a_32059_903.n2 a_32059_903.t4 8.266
R14889 a_32059_903.n1 a_32059_903.t7 8.266
R14890 a_32059_903.n1 a_32059_903.t2 8.266
R14891 a_32059_903.n0 a_32059_903.t1 8.266
R14892 a_32059_903.n0 a_32059_903.t6 8.266
R14893 a_32059_903.t3 a_32059_903.n3 8.266
R14894 a_32059_903.n3 a_32059_903.n2 0.687
R14895 a_32059_903.n2 a_32059_903.n1 0.365
R14896 a_32059_903.n3 a_32059_903.n0 0.365
R14897 level_shifter_up_2.xb_hv.n0 level_shifter_up_2.xb_hv.t8 193.288
R14898 level_shifter_up_2.xb_hv.n0 level_shifter_up_2.xb_hv.t9 193.285
R14899 level_shifter_up_2.xb_hv.n0 level_shifter_up_2.xb_hv.t5 192.83
R14900 level_shifter_up_2.xb_hv.n0 level_shifter_up_2.xb_hv.t7 192.83
R14901 level_shifter_up_2.xb_hv.n1 level_shifter_up_2.xb_hv.t6 66.119
R14902 level_shifter_up_2.xb_hv.n3 level_shifter_up_2.xb_hv.t4 66.118
R14903 level_shifter_up_2.xb_hv.n1 level_shifter_up_2.xb_hv.t3 66.116
R14904 level_shifter_up_2.xb_hv.n3 level_shifter_up_2.xb_hv.t2 66.11
R14905 level_shifter_up_2.xb_hv.n2 level_shifter_up_2.xb_hv.t10 64.963
R14906 level_shifter_up_2.xb_hv level_shifter_up_2.xb_hv.t1 17.301
R14907 level_shifter_up_2.xb_hv.n2 level_shifter_up_2.xb_hv.t0 13.976
R14908 trim4b_hv level_shifter_up_2.xb_hv.n4 11.809
R14909 level_shifter_up_2.xb_hv.n4 level_shifter_up_2.xb_hv.n1 7.621
R14910 trim4b_hv level_shifter_up_2.xb_hv.n2 3.32
R14911 level_shifter_up_2.xb_hv.n4 level_shifter_up_2.xb_hv.n0 1.063
R14912 level_shifter_up_2.xb_hv.n2 level_shifter_up_2.xb_hv 0.51
R14913 level_shifter_up_2.xb_hv.n1 level_shifter_up_2.xb_hv.n3 0.381
R14914 a_32057_n22200.n0 a_32057_n22200.t7 14.666
R14915 a_32057_n22200.n1 a_32057_n22200.t4 14.666
R14916 a_32057_n22200.n2 a_32057_n22200.t10 14.666
R14917 a_32057_n22200.n0 a_32057_n22200.t11 13.849
R14918 a_32057_n22200.n1 a_32057_n22200.t8 13.849
R14919 a_32057_n22200.n4 a_32057_n22200.t9 13.849
R14920 a_32057_n22200.n3 a_32057_n22200.t5 13.849
R14921 a_32057_n22200.n2 a_32057_n22200.t6 13.849
R14922 a_32057_n22200.n7 a_32057_n22200.t2 13.847
R14923 a_32057_n22200.n7 a_32057_n22200.t0 13.847
R14924 a_32057_n22200.n9 a_32057_n22200.t1 13.847
R14925 a_32057_n22200.t3 a_32057_n22200.n9 13.847
R14926 a_32057_n22200.n6 a_32057_n22200.n5 2.212
R14927 a_32057_n22200.n8 a_32057_n22200.n7 1.306
R14928 a_32057_n22200.n9 a_32057_n22200.n8 1.306
R14929 a_32057_n22200.n3 a_32057_n22200.n2 1.273
R14930 a_32057_n22200.n4 a_32057_n22200.n3 0.817
R14931 a_32057_n22200.n5 a_32057_n22200.n4 0.775
R14932 a_32057_n22200.n8 a_32057_n22200.n6 0.704
R14933 a_32057_n22200.n6 a_32057_n22200.n0 0.441
R14934 a_32057_n22200.n5 a_32057_n22200.n1 0.427
R14935 trim[4].n0 trim[4].t3 38.514
R14936 trim[4].n1 trim[4].t1 37.895
R14937 trim[4].n0 trim[4].t2 37.185
R14938 trim[4] trim[4].t0 3.676
R14939 trim[4].n2 trim[4] 1.353
R14940 trim[4].n2 trim[4].n1 0.568
R14941 trim[4].n1 trim[4].n0 0.432
R14942 trim[4] trim[4].n2 0.019
R14943 a_12857_n19542.n1 a_12857_n19542.t0 13.851
R14944 a_12857_n19542.n3 a_12857_n19542.t2 13.851
R14945 a_12857_n19542.n2 a_12857_n19542.t1 13.849
R14946 a_12857_n19542.n2 a_12857_n19542.t5 13.849
R14947 a_12857_n19542.n1 a_12857_n19542.t4 13.849
R14948 a_12857_n19542.n0 a_12857_n19542.t3 13.849
R14949 a_12857_n19542.n0 a_12857_n19542.t7 13.849
R14950 a_12857_n19542.t6 a_12857_n19542.n3 13.849
R14951 a_12857_n19542.n2 a_12857_n19542.n1 1.121
R14952 a_12857_n19542.n3 a_12857_n19542.n0 1.121
R14953 a_12857_n19542.n3 a_12857_n19542.n2 0.762
R14954 a_14459_n4755.t0 a_14459_n4755.t1 19.367
R14955 a_32057_n21342.n7 a_32057_n21342.t6 13.849
R14956 a_32057_n21342.n6 a_32057_n21342.t1 13.849
R14957 a_32057_n21342.n6 a_32057_n21342.t11 13.849
R14958 a_32057_n21342.n5 a_32057_n21342.t5 13.849
R14959 a_32057_n21342.n5 a_32057_n21342.t9 13.849
R14960 a_32057_n21342.n4 a_32057_n21342.t2 13.849
R14961 a_32057_n21342.n4 a_32057_n21342.t10 13.849
R14962 a_32057_n21342.n3 a_32057_n21342.t3 13.849
R14963 a_32057_n21342.n3 a_32057_n21342.t12 13.849
R14964 a_32057_n21342.n2 a_32057_n21342.t7 13.849
R14965 a_32057_n21342.n2 a_32057_n21342.t15 13.849
R14966 a_32057_n21342.n1 a_32057_n21342.t0 13.849
R14967 a_32057_n21342.n1 a_32057_n21342.t8 13.849
R14968 a_32057_n21342.n0 a_32057_n21342.t4 13.849
R14969 a_32057_n21342.n0 a_32057_n21342.t13 13.849
R14970 a_32057_n21342.t14 a_32057_n21342.n7 13.849
R14971 a_32057_n21342.n7 a_32057_n21342.n6 4.449
R14972 a_32057_n21342.n2 a_32057_n21342.n1 0.868
R14973 a_32057_n21342.n4 a_32057_n21342.n3 0.868
R14974 a_32057_n21342.n6 a_32057_n21342.n5 0.464
R14975 a_32057_n21342.n1 a_32057_n21342.n0 0.464
R14976 a_32057_n21342.n3 a_32057_n21342.n2 0.464
R14977 a_32057_n21342.n7 a_32057_n21342.n4 0.464
R14978 a_23032_11382.t0 a_23032_11382.t1 5.031
R14979 trim[1].n0 trim[1].t3 38.514
R14980 trim[1].n1 trim[1].t1 37.895
R14981 trim[1].n0 trim[1].t0 37.185
R14982 trim[1].n2 trim[1] 4.866
R14983 trim[1] trim[1].t2 3.65
R14984 trim[1].n2 trim[1].n1 0.6
R14985 trim[1].n1 trim[1].n0 0.432
R14986 trim[1] trim[1].n2 0.013
R14987 level_shifter_up_6.x_hv.n0 level_shifter_up_6.x_hv.t1 224.065
R14988 level_shifter_up_6.x_hv.n1 level_shifter_up_6.x_hv.t3 224.031
R14989 level_shifter_up_6.x_hv.n1 level_shifter_up_6.x_hv.t4 223.689
R14990 level_shifter_up_6.x_hv.n0 level_shifter_up_6.x_hv.t6 223.648
R14991 level_shifter_up_6.x_hv.n2 level_shifter_up_6.x_hv.t7 125.496
R14992 level_shifter_up_6.x_hv.t0 level_shifter_up_6.x_hv.t5 65.176
R14993 level_shifter_up_6.x_hv.n2 level_shifter_up_6.x_hv.t2 63.645
R14994 level_shifter_up_6.x_hv.n4 level_shifter_up_6.x_hv.n2 20.164
R14995 level_shifter_up_6.x_hv.n0 level_shifter_up_6.x_hv.n3 6.4
R14996 level_shifter_up_6.x_hv level_shifter_up_6.x_hv.n4 1.301
R14997 level_shifter_up_6.x_hv level_shifter_up_6.x_hv.t0 0.705
R14998 level_shifter_up_6.x_hv.n4 level_shifter_up_6.x_hv.n1 0.354
R14999 level_shifter_up_6.x_hv.n1 level_shifter_up_6.x_hv.n0 0.344
R15000 a_27926_9740.n1 a_27926_9740.t6 8.967
R15001 a_27926_9740.n2 a_27926_9740.t4 8.37
R15002 a_27926_9740.n3 a_27926_9740.t2 6.923
R15003 a_27926_9740.n3 a_27926_9740.t1 6.923
R15004 a_27926_9740.n0 a_27926_9740.t5 6.923
R15005 a_27926_9740.n0 a_27926_9740.t7 6.923
R15006 a_27926_9740.n5 a_27926_9740.t0 6.923
R15007 a_27926_9740.t3 a_27926_9740.n5 6.923
R15008 a_27926_9740.n4 a_27926_9740.n3 2.044
R15009 a_27926_9740.n1 a_27926_9740.n0 1.447
R15010 a_27926_9740.n5 a_27926_9740.n4 1.447
R15011 a_27926_9740.n4 a_27926_9740.n2 1.117
R15012 a_27926_9740.n2 a_27926_9740.n1 0.607
R15013 level_shifter_up_4.x_hv.n1 level_shifter_up_4.x_hv.t6 223.931
R15014 level_shifter_up_4.x_hv.n3 level_shifter_up_4.x_hv.t2 223.666
R15015 level_shifter_up_4.x_hv.n2 level_shifter_up_4.x_hv.t3 223.666
R15016 level_shifter_up_4.x_hv.n1 level_shifter_up_4.x_hv.t4 223.666
R15017 level_shifter_up_4.x_hv.n0 level_shifter_up_4.x_hv.t5 65.162
R15018 level_shifter_up_4.x_hv level_shifter_up_4.x_hv.t1 17.199
R15019 level_shifter_up_4.x_hv.n0 level_shifter_up_4.x_hv.t0 13.866
R15020 en_hv level_shifter_up_4.x_hv.n3 13.637
R15021 en_hv level_shifter_up_4.x_hv.n0 0.734
R15022 level_shifter_up_4.x_hv.n0 level_shifter_up_4.x_hv 0.706
R15023 level_shifter_up_4.x_hv.n2 level_shifter_up_4.x_hv.n1 0.265
R15024 level_shifter_up_4.x_hv.n3 level_shifter_up_4.x_hv.n2 0.265
R15025 a_33657_n22200.n0 a_33657_n22200.t3 14.666
R15026 a_33657_n22200.n2 a_33657_n22200.t2 14.296
R15027 a_33657_n22200.n1 a_33657_n22200.t4 13.85
R15028 a_33657_n22200.n0 a_33657_n22200.t5 13.849
R15029 a_33657_n22200.t1 a_33657_n22200.n3 13.847
R15030 a_33657_n22200.n3 a_33657_n22200.t0 13.847
R15031 a_33657_n22200.n1 a_33657_n22200.n0 1.274
R15032 a_33657_n22200.n3 a_33657_n22200.n2 1.163
R15033 a_33657_n22200.n2 a_33657_n22200.n1 0.401
R15034 hyst[0].n1 hyst[0].t1 38.514
R15035 hyst[0].n2 hyst[0].t3 37.894
R15036 hyst[0].n1 hyst[0].t2 37.185
R15037 hyst[0].n0 hyst[0].t0 3.683
R15038 hyst[0].n0 hyst[0] 1.434
R15039 hyst[0] hyst[0].n2 0.564
R15040 hyst[0].n2 hyst[0].n1 0.432
R15041 hyst[0] hyst[0].n0 0.017
R15042 a_25030_4566.t0 a_25030_4566.t1 5.053
C0 res_p_bot a_11257_n21342# 0.12fF
C1 AVDD a_31859_n29829# 1.63fF
C2 Vom bias_var_n 17.07fF
C3 level_shifter_up_2.xb_hv level_shifter_up_3.x_hv 0.44fF
C4 Vxm Vfold_bot_m 0.52fF
C5 a_32448_11527# level_shifter_up_7.x_hv 0.42fF
C6 AVDD Vinp 97.46fF
C7 Vxm m2_9760_9570# 0.11fF
C8 Vxp m2_7560_n25770# 0.11fF
C9 Vfold_bot_m m2_10420_n28830# 0.20fF
C10 level_shifter_up_3.x_hv a_32683_n30483# 0.47fF
C11 level_shifter_up_3.xb_hv a_31928_n30483# 0.15fF
C12 Vfold_bot_m Vxp 113.05fF
C13 AVDD level_shifter_up_2.x_hv 1.39fF
C14 Vfold_bot_m m2_11300_n26430# 0.20fF
C15 casc_n bias_p 1.31fF
C16 Vfold_bot_m m2_6900_n30430# 0.20fF
C17 level_shifter_up_5.x_hv a_36699_n29829# 0.39fF
C18 Vfold_bot_m m2_7560_n28030# 0.20fF
C19 a_34648_11527# a_35403_11527# 0.90fF
C20 level_shifter_up_6.x_hv level_shifter_up_4.xb_hv 0.16fF
C21 Vfold_bot_m m2_3820_n29630# 0.20fF
C22 bias_n a_12859_n4755# 0.78fF
C23 level_shifter_up_0.x_hv casc_p 0.27fF
C24 bias_n a_37477_903# 0.17fF
C25 AVDD a_23013_n31913# 1.54fF
C26 Vxp m2_14160_n29770# 0.11fF
C27 Vfold_bot_m level_shifter_up_0.xb_hv 0.29fF
C28 bias_p res_p_bot 9.02fF
C29 level_shifter_up_5.xb_hv level_shifter_up_0.xb_hv 0.83fF
C30 Vfold_bot_m m2_4700_n27230# 0.20fF
C31 level_shifter_up_6.x_hv level_shifter_up_7.x_hv 7.16fF
C32 a_31003_11527# level_shifter_up_6.xb_hv 0.59fF
C33 hyst[1] hyst[0] 0.27fF
C34 Vop casc_p 41.41fF
C35 level_shifter_up_7.x_hv level_shifter_up_4.xb_hv 0.21fF
C36 Vfold_bot_m m2_19220_n25630# 0.20fF
C37 level_shifter_up_0.x_hv a_31859_n29829# 0.11fF
C38 Vfold_bot_m m2_15700_n27230# 0.20fF
C39 a_23013_n31913# a_24345_n31913# 0.30fF
C40 level_shifter_up_1.xb_hv level_shifter_up_3.xb_hv 0.24fF
C41 level_shifter_up_4.x_hv a_31859_n29829# 0.29fF
C42 a_33203_11527# level_shifter_up_7.xb_hv 0.59fF
C43 AVDD a_33203_11527# 1.55fF
C44 Vfold_bot_m m2_11960_n28830# 0.20fF
C45 Vfold_bot_m m2_12620_n26430# 0.20fF
C46 casc_n bias_var_n 8.18fF
C47 level_shifter_up_6.x_hv trim[0] 0.33fF
C48 Vom Vfold_bot_m 28.79fF
C49 level_shifter_up_2.xb_hv a_34883_n30483# 0.64fF
C50 Vfold_bot_m m2_8220_n30430# 0.20fF
C51 AVDD Vinm 100.95fF
C52 Vxp m2_18560_n30570# 0.11fF
C53 Vfold_bot_m m2_9100_n28030# 0.20fF
C54 level_shifter_up_5.xb_hv a_36259_n29829# 0.68fF
C55 a_35403_11527# level_shifter_up_8.x_hv 0.32fF
C56 trim[4] a_34128_n30483# 1.39fF
C57 Vfold_bot_m m2_5360_n29630# 0.20fF
C58 casc_n a_12859_n2697# 0.75fF
C59 level_shifter_up_5.x_hv casc_p 0.58fF
C60 level_shifter_up_4.xb_hv bias_p 3.38fF
C61 bias_n a_11259_n2697# 0.83fF
C62 bias_n a_11877_1191# 0.16fF
C63 Vfold_bot_m m2_6020_n27230# 0.20fF
C64 trim[0] level_shifter_up_7.x_hv 0.18fF
C65 AVDD bias_n 1.87fF
C66 bias_p a_11257_n21342# 0.30fF
C67 Vfold_bot_m m2_16360_n29630# 0.20fF
C68 res_p_bot level_shifter_up_2.xb_hv 0.61fF
C69 level_shifter_up_5.x_hv a_31859_n29829# 0.15fF
C70 Vfold_bot_m m2_17020_n27230# 0.20fF
C71 level_shifter_up_5.xb_hv a_32299_n29829# 0.46fF
C72 a_23679_n25097# a_25011_n25097# 0.30fF
C73 level_shifter_up_6.xb_hv level_shifter_up_8.xb_hv 0.16fF
C74 trim[1] level_shifter_up_8.x_hv 0.17fF
C75 Vxm m2_11960_7170# 0.11fF
C76 AVDD level_shifter_up_7.xb_hv 1.18fF
C77 Vfold_bot_m m2_13500_n28830# 0.20fF
C78 a_36699_n29829# a_36259_n29829# 0.78fF
C79 casc_p Vxp 54.38fF
C80 Vfold_bot_m m2_14160_n26430# 0.20fF
C81 level_shifter_up_1.xb_hv level_shifter_up_2.x_hv 0.19fF
C82 Vfold_bot_m m2_9760_n30430# 0.20fF
C83 level_shifter_up_3.x_hv level_shifter_up_3.xb_hv 4.47fF
C84 Vfold_bot_m m2_10420_n28030# 0.20fF
C85 level_shifter_up_8.x_hv level_shifter_up_8.xb_hv 6.91fF
C86 Vxm m2_5360_6370# 0.11fF
C87 AVDD a_34499_n29829# 1.77fF
C88 Vxm Vinp 78.10fF
C89 AVDD a_24345_n31913# 1.23fF
C90 casc_n Vfold_bot_m 21.77fF
C91 trim[0] trim[2] 0.13fF
C92 Vfold_bot_m m2_3160_n31230# 0.20fF
C93 Vxp Vinp 73.40fF
C94 AVDD a_36328_n30483# 1.62fF
C95 Vxm m2_16360_6370# 0.11fF
C96 bias_n level_shifter_up_0.x_hv 1.15fF
C97 Vfold_bot_m res_p_bot 0.30fF
C98 level_shifter_up_2.xb_hv trim[5] 0.18fF
C99 level_shifter_up_4.xb_hv level_shifter_up_2.xb_hv 0.13fF
C100 Vfold_bot_m m2_17900_n29630# 0.20fF
C101 Vfold_bot_m en 0.12fF
C102 Vop bias_n 0.35fF
C103 level_shifter_up_5.xb_hv en 0.13fF
C104 Vfold_bot_m m2_18560_n27230# 0.20fF
C105 level_shifter_up_0.xb_hv a_31859_n29829# 0.20fF
C106 Vxp m2_11960_n25770# 0.11fF
C107 Vxm m2_14160_9570# 0.11fF
C108 AVDD level_shifter_up_0.x_hv 4.05fF
C109 Vfold_bot_m m2_14820_n28830# 0.20fF
C110 AVDD level_shifter_up_4.x_hv 4.12fF
C111 Vxp m2_7560_n29770# 0.11fF
C112 Vxm m2_9760_5570# 0.11fF
C113 Vom casc_p 41.44fF
C114 AVDD Vop 64.42fF
C115 Vfold_bot_m m2_11300_n30430# 0.20fF
C116 AVDD a_31928_n30483# 1.72fF
C117 Vfold_bot_m m2_11960_n28030# 0.20fF
C118 AVDD hyst[1] 10.10fF
C119 level_shifter_up_0.x_hv a_34499_n29829# 0.38fF
C120 Vxp m2_5360_n26570# 0.11fF
C121 bias_var_n bias_p 0.88fF
C122 a_11877_1191# ibias 0.82fF
C123 bias_n ibias 10.94fF
C124 Vfold_bot_m m2_4700_n31230# 0.20fF
C125 AVDD level_shifter_up_1.x_hv 1.42fF
C126 level_shifter_up_6.x_hv a_31003_11527# 0.52fF
C127 a_34499_n29829# hyst[1] 1.36fF
C128 Vxm Vinm 78.42fF
C129 bias_n a_14459_n2697# 0.89fF
C130 level_shifter_up_4.xb_hv Vfold_bot_m 0.66fF
C131 bias_n level_shifter_up_5.x_hv 1.19fF
C132 level_shifter_up_4.xb_hv level_shifter_up_5.xb_hv 0.11fF
C133 Vxp m2_16360_n26570# 0.11fF
C134 Vfold_bot_m m2_19220_n29630# 0.20fF
C135 AVDD ibias 0.26fF
C136 a_34128_n30483# a_34883_n30483# 0.88fF
C137 Vxp Vinm 73.08fF
C138 Vfold_bot_m m2_15700_n31230# 0.20fF
C139 Vfold_bot_m m2_3160_n25630# 0.20fF
C140 trim[1] a_32448_11527# 1.18fF
C141 a_31003_11527# level_shifter_up_7.x_hv 0.18fF
C142 AVDD level_shifter_up_5.x_hv 5.70fF
C143 AVDD level_shifter_up_1.xb_hv 9.84fF
C144 AVDD a_30248_11527# 1.60fF
C145 level_shifter_up_0.x_hv level_shifter_up_4.x_hv 0.14fF
C146 Vxp m2_9760_n27370# 0.11fF
C147 Vfold_bot_m m2_12620_n30430# 0.20fF
C148 res_p_bot level_shifter_up_3.xb_hv 0.57fF
C149 AVDD trim[4] 3.44fF
C150 a_36328_n30483# level_shifter_up_1.x_hv 0.24fF
C151 Vxm bias_n 22.49fF
C152 a_32299_n29829# a_31859_n29829# 0.81fF
C153 Vfold_bot_m m2_13500_n28030# 0.20fF
C154 level_shifter_up_5.x_hv a_34499_n29829# 0.72fF
C155 casc_n casc_p 0.83fF
C156 AVDD Vom_stg2 1.20fF
C157 AVDD a_34648_11527# 1.62fF
C158 Vfold_bot_m m2_6020_n31230# 0.20fF
C159 Vfold_bot_m m2_6900_n28830# 0.20fF
C160 level_shifter_up_1.xb_hv a_36328_n30483# 0.18fF
C161 AVDD Vxp 325.65fF
C162 Vfold_bot_m bias_p 1.55fF
C163 Vfold_bot_m m2_7560_n26430# 0.20fF
C164 casc_n a_35259_903# 0.71fF
C165 casc_p res_p_bot 1.09fF
C166 a_34883_n30483# level_shifter_up_2.x_hv 0.27fF
C167 Vxm m2_3160_10370# 0.11fF
C168 Vfold_bot_m m2_17020_n31230# 0.20fF
C169 casc_p m2_30910_n8650# 0.21fF
C170 Vfold_bot_m m2_4700_n25630# 0.20fF
C171 trim[1] level_shifter_up_7.x_hv 0.24fF
C172 level_shifter_up_6.x_hv level_shifter_up_8.xb_hv 0.27fF
C173 AVDD level_shifter_up_0.xb_hv 19.94fF
C174 level_shifter_up_0.x_hv level_shifter_up_5.x_hv 8.34fF
C175 AVDD level_shifter_up_6.xb_hv 1.22fF
C176 level_shifter_up_5.x_hv level_shifter_up_4.x_hv 0.23fF
C177 level_shifter_up_0.x_hv level_shifter_up_1.xb_hv 0.17fF
C178 level_shifter_up_4.x_hv level_shifter_up_1.xb_hv 0.12fF
C179 level_shifter_up_3.xb_hv trim[5] 0.17fF
C180 bias_stg2 a_37477_903# 0.21fF
C181 Vfold_bot_m m2_14160_n30430# 0.20fF
C182 Vfold_bot_m m2_14820_n28030# 0.20fF
C183 Vfold_bot_m m2_15700_n25630# 0.20fF
C184 level_shifter_up_5.x_hv hyst[1] 0.36fF
C185 level_shifter_up_5.xb_hv a_34059_n29829# 0.24fF
C186 level_shifter_up_7.xb_hv level_shifter_up_8.x_hv 0.14fF
C187 level_shifter_up_7.x_hv level_shifter_up_8.xb_hv 2.38fF
C188 AVDD level_shifter_up_3.x_hv 1.88fF
C189 AVDD level_shifter_up_8.x_hv 5.66fF
C190 Vom bias_n 1.13fF
C191 Vop Vom_stg2 1.22fF
C192 Vxm m2_7560_9570# 0.11fF
C193 trim[0] trim[1] 2.25fF
C194 Vfold_bot_m m2_8220_n28830# 0.20fF
C195 level_shifter_up_1.xb_hv level_shifter_up_1.x_hv 1.43fF
C196 casc_n a_12859_n4755# 1.08fF
C197 casc_n a_37477_903# 0.32fF
C198 bias_n a_11259_n4497# 0.27fF
C199 level_shifter_up_4.xb_hv casc_p 0.45fF
C200 Vfold_bot_m m2_9100_n26430# 0.20fF
C201 bias_var_n Vfold_bot_m 18.25fF
C202 AVDD Vom 62.24fF
C203 bias_n a_35259_2049# 0.44fF
C204 AVDD a_36259_n29829# 1.60fF
C205 Vfold_bot_m m2_18560_n31230# 0.20fF
C206 Vfold_bot_m m2_6020_n25630# 0.20fF
C207 trim[0] level_shifter_up_8.xb_hv 0.95fF
C208 trim[1] trim[2] 1.32fF
C209 Vxm m2_14160_5570# 0.11fF
C210 casc_p a_11257_n21342# 0.71fF
C211 Vxp m2_11960_n29770# 0.11fF
C212 level_shifter_up_5.x_hv level_shifter_up_1.xb_hv 0.17fF
C213 level_shifter_up_0.x_hv level_shifter_up_0.xb_hv 5.00fF
C214 level_shifter_up_4.x_hv level_shifter_up_0.xb_hv 3.10fF
C215 Vfold_bot_m m2_2500_n27230# 0.20fF
C216 level_shifter_up_4.xb_hv a_31859_n29829# 0.56fF
C217 bias_stg2 bias_n 0.51fF
C218 level_shifter_up_1.xb_hv trim[4] 0.22fF
C219 Vxm ibias 2.09fF
C220 Vfold_bot_m m2_17020_n25630# 0.20fF
C221 trim[2] level_shifter_up_8.xb_hv 0.17fF
C222 AVDD a_32299_n29829# 1.95fF
C223 AVDD bias_stg2 18.06fF
C224 Vxp m2_5360_n30570# 0.11fF
C225 a_32448_11527# a_33203_11527# 0.90fF
C226 Vfold_bot_m m2_9760_n28830# 0.20fF
C227 level_shifter_up_3.x_hv a_31928_n30483# 0.78fF
C228 bias_p casc_p 17.44fF
C229 AVDD a_34883_n30483# 1.55fF
C230 casc_n a_12859_n4497# 0.77fF
C231 Vfold_bot_m m2_10420_n26430# 0.20fF
C232 casc_n a_11259_n2697# 0.75fF
C233 casc_n a_11877_1191# 0.36fF
C234 bias_n casc_n 15.21fF
C235 Vxm m2_5360_7970# 0.11fF
C236 Vom level_shifter_up_0.x_hv 0.36fF
C237 Vxp m2_16360_n30570# 0.11fF
C238 Vfold_bot_m m2_6900_n28030# 0.20fF
C239 Vop Vom 15.00fF
C240 Vfold_bot_m m2_3160_n29630# 0.20fF
C241 AVDD casc_n 0.59fF
C242 AVDD Vop_stg2 0.72fF
C243 bias_n a_36859_903# 0.29fF
C244 level_shifter_up_5.x_hv level_shifter_up_0.xb_hv 0.49fF
C245 level_shifter_up_1.xb_hv level_shifter_up_0.xb_hv 0.57fF
C246 Vfold_bot_m m2_3820_n27230# 0.20fF
C247 Vxm m2_16360_7970# 0.11fF
C248 Vxp m2_14160_n27370# 0.11fF
C249 Vfold_bot_m m2_18560_n25630# 0.20fF
C250 AVDD res_p_bot 17.36fF
C251 AVDD en 12.90fF
C252 level_shifter_up_0.x_hv a_32299_n29829# 0.28fF
C253 level_shifter_up_5.x_hv level_shifter_up_3.x_hv 0.17fF
C254 bias_stg2 level_shifter_up_0.x_hv 0.98fF
C255 level_shifter_up_4.x_hv a_32299_n29829# 0.31fF
C256 level_shifter_up_2.xb_hv level_shifter_up_3.xb_hv 3.11fF
C257 level_shifter_up_1.xb_hv level_shifter_up_3.x_hv 0.32fF
C258 a_33203_11527# level_shifter_up_7.x_hv 0.47fF
C259 Vxm m2_9760_7170# 0.11fF
C260 AVDD m2_30910_n8650# 0.11fF
C261 AVDD a_32448_11527# 1.63fF
C262 Vfold_bot_m m2_11300_n28830# 0.20fF
C263 level_shifter_up_3.xb_hv a_32683_n30483# 0.80fF
C264 AVDD trim[3] 3.43fF
C265 bias_var_n casc_p 3.86fF
C266 Vfold_bot_m m2_11960_n26430# 0.20fF
C267 level_shifter_up_2.xb_hv a_34128_n30483# 0.14fF
C268 Vfold_bot_m m2_7560_n30430# 0.20fF
C269 res_p_bot a_24345_n31913# 0.34fF
C270 level_shifter_up_5.x_hv a_36259_n29829# 0.40fF
C271 Vfold_bot_m m2_8220_n28030# 0.20fF
C272 a_34648_11527# level_shifter_up_8.x_hv 0.36fF
C273 a_12859_n4209# a_12859_n4497# 0.28fF
C274 Vfold_bot_m m2_4700_n29630# 0.20fF
C275 bias_n a_12859_n4209# 0.31fF
C276 AVDD a_23679_n25097# 0.97fF
C277 bias_n a_11259_2049# 0.28fF
C278 level_shifter_up_0.x_hv casc_n 0.23fF
C279 level_shifter_up_4.xb_hv bias_n 2.19fF
C280 Vfold_bot_m m2_5360_n27230# 0.20fF
C281 AVDD level_shifter_up_6.x_hv 4.75fF
C282 Vop casc_n 23.49fF
C283 Vom_stg2 Vom 0.20fF
C284 Vop Vop_stg2 0.16fF
C285 Vxm m2_18560_10370# 0.11fF
C286 level_shifter_up_7.x_hv bias_n 0.39fF
C287 AVDD trim[5] 3.37fF
C288 trim[3] a_36328_n30483# 1.41fF
C289 AVDD level_shifter_up_4.xb_hv 4.72fF
C290 Vfold_bot_m m2_15700_n29630# 0.20fF
C291 level_shifter_up_0.x_hv en 0.24fF
C292 level_shifter_up_5.x_hv a_32299_n29829# 0.57fF
C293 bias_stg2 level_shifter_up_5.x_hv 0.62fF
C294 Vfold_bot_m m2_16360_n27230# 0.20fF
C295 level_shifter_up_6.xb_hv level_shifter_up_8.x_hv 0.11fF
C296 level_shifter_up_7.x_hv level_shifter_up_7.xb_hv 1.14fF
C297 AVDD level_shifter_up_7.x_hv 5.14fF
C298 Vxp m2_9760_n25770# 0.11fF
C299 Vxm m2_11960_9570# 0.11fF
C300 Vfold_bot_m m2_12620_n28830# 0.20fF
C301 AVDD a_11257_n21342# 0.93fF
C302 Vxm m2_7560_5570# 0.11fF
C303 Vop m2_30910_n8650# 0.29fF
C304 casc_n a_14459_n4497# 0.77fF
C305 Vfold_bot_m m2_13500_n26430# 0.20fF
C306 en hyst[1] 1.12fF
C307 level_shifter_up_2.xb_hv level_shifter_up_2.x_hv 1.34fF
C308 Vfold_bot_m m2_9100_n30430# 0.20fF
C309 casc_n ibias 2.43fF
C310 Vfold_bot_m m2_9760_n28030# 0.20fF
C311 bias_stg2 Vom_stg2 0.12fF
C312 a_35403_11527# level_shifter_up_8.xb_hv 0.59fF
C313 Vxm m2_5360_8770# 0.11fF
C314 Vfold_bot_m casc_p 1.57fF
C315 Vfold_bot_m m2_6020_n29630# 0.20fF
C316 casc_n a_14459_n2697# 0.71fF
C317 bias_n bias_p 1.47fF
C318 bias_n a_12859_2049# 0.22fF
C319 level_shifter_up_5.x_hv casc_n 0.23fF
C320 AVDD trim[0] 11.74fF
C321 Vfold_bot_m m2_2500_n31230# 0.20fF
C322 level_shifter_up_6.x_hv level_shifter_up_0.x_hv 0.52fF
C323 level_shifter_up_6.x_hv Vop 0.24fF
C324 AVDD bias_p 212.38fF
C325 level_shifter_up_4.xb_hv level_shifter_up_0.x_hv 0.12fF
C326 Vxm m2_16360_8770# 0.11fF
C327 level_shifter_up_4.xb_hv level_shifter_up_4.x_hv 4.39fF
C328 Vfold_bot_m m2_17020_n29630# 0.20fF
C329 level_shifter_up_5.x_hv en 0.20fF
C330 Vop level_shifter_up_4.xb_hv 1.19fF
C331 Vom_stg2 Vop_stg2 2.85fF
C332 level_shifter_up_0.xb_hv a_32299_n29829# 0.18fF
C333 Vfold_bot_m m2_17900_n27230# 0.20fF
C334 level_shifter_up_5.xb_hv a_31859_n29829# 0.17fF
C335 trim[1] level_shifter_up_8.xb_hv 0.18fF
C336 Vxm casc_n 28.24fF
C337 Vfold_bot_m Vinp 13.28fF
C338 trim[5] a_31928_n30483# 1.33fF
C339 AVDD trim[2] 3.87fF
C340 level_shifter_up_7.x_hv level_shifter_up_0.x_hv 0.22fF
C341 a_36699_n29829# hyst[0] 1.30fF
C342 Vfold_bot_m m2_14160_n28830# 0.20fF
C343 Vfold_bot_m m2_14820_n26430# 0.20fF
C344 level_shifter_up_1.xb_hv trim[3] 0.38fF
C345 Vfold_bot_m m2_10420_n30430# 0.20fF
C346 Vxp m2_7560_n27370# 0.11fF
C347 Vfold_bot_m m2_11300_n28030# 0.20fF
C348 AVDD a_34059_n29829# 1.59fF
C349 bias_n a_14459_n4209# 0.31fF
C350 AVDD a_25011_n25097# 1.32fF
C351 bias_n bias_var_n 0.62fF
C352 Vxp res_p_bot 2.46fF
C353 a_11259_2049# ibias 0.35fF
C354 Vfold_bot_m m2_3820_n31230# 0.20fF
C355 bias_stg2 Vom 0.13fF
C356 level_shifter_up_6.x_hv level_shifter_up_5.x_hv 0.47fF
C357 AVDD a_37083_n30483# 1.59fF
C358 level_shifter_up_6.x_hv a_30248_11527# 0.54fF
C359 a_34499_n29829# a_34059_n29829# 0.78fF
C360 AVDD bias_var_n 5.95fF
C361 level_shifter_up_0.x_hv bias_p 1.38fF
C362 bias_n a_12859_n2697# 0.83fF
C363 bias_p level_shifter_up_4.x_hv 0.54fF
C364 level_shifter_up_4.xb_hv level_shifter_up_5.x_hv 0.20fF
C365 level_shifter_up_1.xb_hv trim[5] 0.18fF
C366 level_shifter_up_4.xb_hv level_shifter_up_1.xb_hv 1.55fF
C367 Vfold_bot_m m2_18560_n29630# 0.20fF
C368 Vop bias_p 13.19fF
C369 Vfold_bot_m m2_19220_n27230# 0.20fF
C370 level_shifter_up_0.xb_hv en 0.55fF
C371 Vxm m2_14160_7170# 0.11fF
C372 Vfold_bot_m m2_2500_n25630# 0.20fF
C373 level_shifter_up_7.x_hv level_shifter_up_5.x_hv 0.12fF
C374 AVDD level_shifter_up_2.xb_hv 7.25fF
C375 Vom casc_n 28.53fF
C376 Vom_stg2 level_shifter_up_4.xb_hv 0.37fF
C377 Vfold_bot_m m2_11960_n30430# 0.20fF
C378 Vom Vop_stg2 1.47fF
C379 res_p_bot level_shifter_up_3.x_hv 0.58fF
C380 AVDD a_32683_n30483# 1.56fF
C381 a_36328_n30483# a_37083_n30483# 0.89fF
C382 Vxm level_shifter_up_4.xb_hv 1.42fF
C383 Vfold_bot_m Vinm 10.70fF
C384 Vfold_bot_m m2_12620_n28030# 0.20fF
C385 Vxp m2_5360_n28970# 0.11fF
C386 level_shifter_up_0.x_hv a_34059_n29829# 0.48fF
C387 casc_n a_11259_n4497# 0.75fF
C388 a_12859_2049# ibias 0.41fF
C389 Vfold_bot_m m2_5360_n31230# 0.20fF
C390 level_shifter_up_6.x_hv level_shifter_up_6.xb_hv 1.12fF
C391 trim[0] a_30248_11527# 1.19fF
C392 Vxp m2_16360_n28970# 0.11fF
C393 level_shifter_up_5.x_hv bias_p 2.53fF
C394 bias_n Vfold_bot_m 1.43fF
C395 Vfold_bot_m m2_6900_n26430# 0.20fF
C396 level_shifter_up_4.xb_hv level_shifter_up_0.xb_hv 0.16fF
C397 a_34128_n30483# level_shifter_up_2.x_hv 0.24fF
C398 Vop bias_var_n 12.46fF
C399 bias_stg2 casc_n 0.49fF
C400 Vfold_bot_m m2_16360_n31230# 0.20fF
C401 Vfold_bot_m m2_3820_n25630# 0.20fF
C402 AVDD Vfold_bot_m 67.60fF
C403 level_shifter_up_6.x_hv level_shifter_up_8.x_hv 0.22fF
C404 level_shifter_up_6.xb_hv level_shifter_up_7.x_hv 0.10fF
C405 Vxp m2_14160_n25770# 0.11fF
C406 AVDD level_shifter_up_5.xb_hv 9.63fF
C407 Vxm m2_11960_5570# 0.11fF
C408 AVDD a_31003_11527# 1.55fF
C409 Vxp m2_9760_n29770# 0.11fF
C410 level_shifter_up_0.x_hv level_shifter_up_2.xb_hv 0.11fF
C411 level_shifter_up_3.x_hv trim[5] 0.34fF
C412 Vfold_bot_m m2_13500_n30430# 0.20fF
C413 a_37083_n30483# level_shifter_up_1.x_hv 0.27fF
C414 a_32299_n29829# en 1.39fF
C415 Vfold_bot_m m2_14160_n28030# 0.20fF
C416 level_shifter_up_6.x_hv Vom 0.27fF
C417 level_shifter_up_5.x_hv a_34059_n29829# 0.22fF
C418 level_shifter_up_5.xb_hv a_34499_n29829# 0.67fF
C419 a_14459_n4209# a_14459_n4497# 0.28fF
C420 bias_p Vxp 0.23fF
C421 trim[2] a_34648_11527# 1.18fF
C422 level_shifter_up_7.x_hv level_shifter_up_8.x_hv 4.10fF
C423 a_31928_n30483# a_32683_n30483# 0.89fF
C424 AVDD a_35403_11527# 1.54fF
C425 Vxp m2_3160_n30570# 0.11fF
C426 Vom level_shifter_up_4.xb_hv 3.04fF
C427 level_shifter_up_6.x_hv a_35259_2049# 0.85fF
C428 Vfold_bot_m m2_7560_n28830# 0.20fF
C429 level_shifter_up_1.xb_hv a_37083_n30483# 0.62fF
C430 level_shifter_up_7.x_hv Vom 0.13fF
C431 casc_n a_36859_903# 0.32fF
C432 Vfold_bot_m m2_8220_n26430# 0.20fF
C433 AVDD a_36699_n29829# 1.89fF
C434 Vfold_bot_m m2_17900_n31230# 0.20fF
C435 Vfold_bot_m m2_5360_n25630# 0.20fF
C436 trim[0] level_shifter_up_8.x_hv 0.18fF
C437 level_shifter_up_6.x_hv bias_stg2 1.11fF
C438 level_shifter_up_0.x_hv Vfold_bot_m 0.24fF
C439 AVDD trim[1] 4.26fF
C440 level_shifter_up_0.x_hv level_shifter_up_5.xb_hv 5.51fF
C441 level_shifter_up_5.x_hv level_shifter_up_2.xb_hv 0.17fF
C442 level_shifter_up_2.xb_hv level_shifter_up_1.xb_hv 7.53fF
C443 level_shifter_up_4.x_hv level_shifter_up_5.xb_hv 0.13fF
C444 Vop Vfold_bot_m 3.41fF
C445 Vxp m2_11960_n27370# 0.11fF
C446 Vfold_bot_m m2_14820_n30430# 0.20fF
C447 bias_stg2 level_shifter_up_4.xb_hv 0.12fF
C448 AVDD DVDD 4.25fF
C449 level_shifter_up_2.xb_hv trim[4] 0.27fF
C450 Vfold_bot_m m2_16360_n25630# 0.20fF
C451 level_shifter_up_0.xb_hv a_34059_n29829# 0.66fF
C452 level_shifter_up_5.xb_hv hyst[1] 0.42fF
C453 trim[2] level_shifter_up_8.x_hv 0.27fF
C454 level_shifter_up_7.x_hv bias_stg2 0.67fF
C455 level_shifter_up_7.xb_hv level_shifter_up_8.xb_hv 0.16fF
C456 AVDD level_shifter_up_3.xb_hv 1.74fF
C457 AVDD level_shifter_up_8.xb_hv 9.00fF
C458 Vom bias_p 8.98fF
C459 Vxm m2_7560_7170# 0.11fF
C460 Vxp m2_5360_n28170# 0.11fF
C461 Vfold_bot_m m2_9100_n28830# 0.20fF
C462 AVDD a_34128_n30483# 1.59fF
C463 Vfold_bot_m m2_9760_n26430# 0.20fF
C464 DVDD Vout 0.62fF
C465 Vinp Vinm 91.58fF
C466 level_shifter_up_4.xb_hv casc_n 0.21fF
C467 Vop_stg2 level_shifter_up_4.xb_hv 0.22fF
C468 AVDD hyst[0] 3.80fF
C469 Vxm m2_5360_10370# 0.11fF
C470 Vxp m2_16360_n28170# 0.11fF
C471 Vfold_bot_m m2_19220_n31230# 0.20fF
C472 AVDD casc_p 236.74fF
C473 trim[0] bias_stg2 0.25fF
C474 Vfold_bot_m m2_2500_n29630# 0.20fF
C475 bias_n a_35259_903# 0.84fF
C476 level_shifter_up_5.x_hv Vfold_bot_m 0.25fF
C477 level_shifter_up_5.x_hv level_shifter_up_5.xb_hv 6.19fF
C478 level_shifter_up_2.xb_hv level_shifter_up_0.xb_hv 1.09fF
C479 level_shifter_up_1.xb_hv level_shifter_up_5.xb_hv 2.08fF
C480 Vfold_bot_m m2_3160_n27230# 0.20fF
C481 a_30248_11527# a_31003_11527# 0.87fF
C482 Vxm m2_16360_10370# 0.11fF
C483 Vfold_bot_m m2_17900_n25630# 0.20fF
C484 ibias DGND 20.87fF
C485 Vout DGND 0.92fF
C486 Vinm DGND 129.23fF
C487 Vinp DGND 157.98fF
C488 DVDD DGND 8.63fF
C489 a_37083_n30483# DGND 1.07fF
C490 a_36328_n30483# DGND 1.86fF
C491 trim[3] DGND 2.58fF
C492 a_34883_n30483# DGND 0.67fF
C493 a_34128_n30483# DGND 1.58fF
C494 trim[4] DGND 2.32fF
C495 a_32683_n30483# DGND 0.34fF
C496 a_31928_n30483# DGND 1.17fF
C497 trim[5] DGND 2.34fF
C498 hyst[0] DGND 2.34fF
C499 a_36699_n29829# DGND 1.60fF
C500 hyst[1] DGND 1.85fF
C501 a_34059_n29829# DGND 0.29fF
C502 a_34499_n29829# DGND 1.53fF
C503 en DGND -1.73fF
C504 a_31859_n29829# DGND 0.60fF
C505 a_32299_n29829# DGND 1.71fF
C506 level_shifter_up_3.xb_hv DGND 2.67fF $ **FLOATING
C507 level_shifter_up_3.x_hv DGND 4.40fF $ **FLOATING
C508 a_25011_n25097# DGND 0.89fF
C509 a_24345_n31913# DGND 0.89fF
C510 a_23679_n25097# DGND 0.89fF
C511 a_23013_n31913# DGND 0.89fF
C512 level_shifter_up_0.xb_hv DGND -9.39fF $ **FLOATING
C513 level_shifter_up_5.xb_hv DGND -4.02fF $ **FLOATING
C514 level_shifter_up_1.xb_hv DGND -3.15fF
C515 level_shifter_up_2.xb_hv DGND 0.15fF $ **FLOATING
C516 level_shifter_up_4.x_hv DGND 2.46fF $ **FLOATING
C517 res_p_bot DGND 4.76fF $ **FLOATING
C518 Vxp DGND -682.67fF $ **FLOATING
C519 a_14459_n4497# DGND 1.73fF
C520 a_14459_n4209# DGND 0.49fF
C521 a_12859_n4497# DGND 1.73fF
C522 a_12859_n4209# DGND 0.49fF
C523 a_12859_n4755# DGND 1.91fF
C524 casc_p DGND -91.55fF $ **FLOATING
C525 a_11259_n4497# DGND 1.46fF
C526 a_14459_n2697# DGND 1.46fF
C527 a_12859_n2697# DGND 1.49fF
C528 bias_p DGND 26.59fF
C529 a_11259_n2697# DGND 1.49fF
C530 a_37477_903# DGND 0.93fF
C531 a_36859_903# DGND 0.68fF
C532 a_35259_903# DGND 1.38fF
C533 Vfold_bot_m DGND 56.46fF $ **FLOATING
C534 bias_var_n DGND 145.27fF
C535 a_12859_2049# DGND 1.10fF
C536 a_11877_1191# DGND 0.94fF
C537 a_11259_2049# DGND 1.08fF
C538 casc_n DGND 93.36fF $ **FLOATING
C539 a_35259_2049# DGND 1.85fF
C540 level_shifter_up_5.x_hv DGND -1.21fF $ **FLOATING
C541 level_shifter_up_0.x_hv DGND 6.06fF $ **FLOATING
C542 bias_n DGND 175.94fF $ **FLOATING
C543 level_shifter_up_4.xb_hv DGND 17.06fF $ **FLOATING
C544 Vop_stg2 DGND 6.72fF
C545 Vom DGND 118.96fF $ **FLOATING
C546 Vom_stg2 DGND 8.88fF
C547 Vop DGND 62.10fF $ **FLOATING
C548 bias_stg2 DGND -2.52fF $ **FLOATING
C549 level_shifter_up_8.xb_hv DGND -2.70fF
C550 level_shifter_up_8.x_hv DGND -1.45fF
C551 a_35403_11527# DGND -0.15fF
C552 a_34648_11527# DGND 1.45fF
C553 trim[2] DGND 3.17fF
C554 level_shifter_up_7.x_hv DGND 2.87fF
C555 a_33203_11527# DGND -0.24fF
C556 a_32448_11527# DGND 1.42fF
C557 trim[1] DGND 2.96fF
C558 a_31003_11527# DGND -0.25fF
C559 a_30248_11527# DGND 1.43fF
C560 trim[0] DGND 0.76fF
C561 level_shifter_up_6.x_hv DGND -0.19fF
C562 Vxm DGND -550.86fF $ **FLOATING
C563 AVDD DGND -73.97fF
C564 a_25030_4566.t1 DGND 0.14fF
C565 a_25030_4566.t0 DGND 2.24fF
C566 hyst[0].t0 DGND 0.33fF
C567 hyst[0].n0 DGND 1.51fF $ **FLOATING
C568 hyst[0].t1 DGND 0.10fF
C569 hyst[0].n1 DGND 0.42fF $ **FLOATING
C570 hyst[0].n2 DGND 0.44fF $ **FLOATING
C571 a_33657_n22200.n0 DGND 1.06fF $ **FLOATING
C572 a_33657_n22200.n1 DGND 0.52fF $ **FLOATING
C573 a_33657_n22200.n2 DGND 1.27fF $ **FLOATING
C574 a_33657_n22200.n3 DGND 0.25fF $ **FLOATING
C575 level_shifter_up_4.x_hv.n0 DGND 2.30fF $ **FLOATING
C576 level_shifter_up_4.x_hv.t5 DGND 0.24fF
C577 level_shifter_up_4.x_hv.t2 DGND 0.52fF
C578 level_shifter_up_4.x_hv.t3 DGND 0.52fF
C579 level_shifter_up_4.x_hv.t4 DGND 0.52fF
C580 level_shifter_up_4.x_hv.t6 DGND 0.52fF
C581 level_shifter_up_4.x_hv.n1 DGND 0.68fF $ **FLOATING
C582 level_shifter_up_4.x_hv.n2 DGND 0.36fF $ **FLOATING
C583 level_shifter_up_4.x_hv.n3 DGND 2.34fF $ **FLOATING
C584 en_hv DGND 2.84fF $ **FLOATING
C585 a_27926_9740.t4 DGND 0.25fF
C586 a_27926_9740.t5 DGND 0.10fF
C587 a_27926_9740.t7 DGND 0.10fF
C588 a_27926_9740.n0 DGND 0.73fF $ **FLOATING
C589 a_27926_9740.t6 DGND 0.30fF
C590 a_27926_9740.n1 DGND 0.94fF $ **FLOATING
C591 a_27926_9740.n2 DGND 0.94fF $ **FLOATING
C592 a_27926_9740.t2 DGND 0.10fF
C593 a_27926_9740.t1 DGND 0.10fF
C594 a_27926_9740.n3 DGND 0.75fF $ **FLOATING
C595 a_27926_9740.n4 DGND 0.28fF $ **FLOATING
C596 a_27926_9740.t0 DGND 0.10fF
C597 a_27926_9740.n5 DGND 0.73fF $ **FLOATING
C598 a_27926_9740.t3 DGND 0.10fF
C599 level_shifter_up_6.x_hv.n0 DGND 0.39fF $ **FLOATING
C600 level_shifter_up_6.x_hv.n1 DGND 0.72fF $ **FLOATING
C601 level_shifter_up_6.x_hv.t7 DGND 0.14fF
C602 level_shifter_up_6.x_hv.n2 DGND 4.49fF $ **FLOATING
C603 level_shifter_up_6.x_hv.t2 DGND 0.14fF
C604 level_shifter_up_6.x_hv.t4 DGND 0.32fF
C605 level_shifter_up_6.x_hv.t3 DGND 0.32fF
C606 level_shifter_up_6.x_hv.t1 DGND 0.32fF
C607 level_shifter_up_6.x_hv.t6 DGND 0.32fF
C608 level_shifter_up_6.x_hv.n4 DGND 2.53fF $ **FLOATING
C609 level_shifter_up_6.x_hv.t5 DGND 0.15fF
C610 level_shifter_up_6.x_hv.t0 DGND 0.96fF
C611 trim[1].t1 DGND 0.11fF
C612 trim[1].t3 DGND 0.11fF
C613 trim[1].t0 DGND 0.10fF
C614 trim[1].n0 DGND 0.47fF $ **FLOATING
C615 trim[1].n1 DGND 0.49fF $ **FLOATING
C616 trim[1].n2 DGND 1.64fF $ **FLOATING
C617 trim[1].t2 DGND 0.36fF
C618 a_23032_11382.t1 DGND 0.15fF
C619 a_23032_11382.t0 DGND 2.41fF
C620 a_32057_n21342.n0 DGND 0.93fF $ **FLOATING
C621 a_32057_n21342.n1 DGND 1.06fF $ **FLOATING
C622 a_32057_n21342.n2 DGND 1.06fF $ **FLOATING
C623 a_32057_n21342.n3 DGND 1.06fF $ **FLOATING
C624 a_32057_n21342.n4 DGND 1.06fF $ **FLOATING
C625 a_32057_n21342.n5 DGND 0.93fF $ **FLOATING
C626 a_32057_n21342.n6 DGND 1.33fF $ **FLOATING
C627 a_32057_n21342.n7 DGND 1.33fF $ **FLOATING
C628 a_14459_n4755.t1 DGND 1.02fF
C629 a_14459_n4755.t0 DGND 1.06fF
C630 a_12857_n19542.n0 DGND 1.06fF $ **FLOATING
C631 a_12857_n19542.n1 DGND 0.97fF $ **FLOATING
C632 a_12857_n19542.n2 DGND 1.23fF $ **FLOATING
C633 a_12857_n19542.n3 DGND 1.14fF $ **FLOATING
C634 trim[4].t3 DGND 0.10fF
C635 trim[4].n0 DGND 0.43fF $ **FLOATING
C636 trim[4].n1 DGND 0.45fF $ **FLOATING
C637 trim[4].n2 DGND 0.56fF $ **FLOATING
C638 trim[4].t0 DGND 0.34fF
C639 a_32057_n22200.n0 DGND 1.32fF $ **FLOATING
C640 a_32057_n22200.n1 DGND 1.31fF $ **FLOATING
C641 a_32057_n22200.n2 DGND 1.54fF $ **FLOATING
C642 a_32057_n22200.n3 DGND 0.90fF $ **FLOATING
C643 a_32057_n22200.n4 DGND 0.76fF $ **FLOATING
C644 a_32057_n22200.n5 DGND 1.29fF $ **FLOATING
C645 a_32057_n22200.n6 DGND 1.14fF $ **FLOATING
C646 a_32057_n22200.n7 DGND 0.40fF $ **FLOATING
C647 a_32057_n22200.n8 DGND 0.88fF $ **FLOATING
C648 a_32057_n22200.n9 DGND 0.40fF $ **FLOATING
C649 level_shifter_up_2.xb_hv.n0 DGND 1.29fF $ **FLOATING
C650 level_shifter_up_2.xb_hv.n1 DGND 2.92fF $ **FLOATING
C651 level_shifter_up_2.xb_hv.t10 DGND 0.20fF
C652 level_shifter_up_2.xb_hv.n2 DGND 2.87fF $ **FLOATING
C653 level_shifter_up_2.xb_hv.t8 DGND 0.41fF
C654 level_shifter_up_2.xb_hv.t7 DGND 0.41fF
C655 level_shifter_up_2.xb_hv.t5 DGND 0.41fF
C656 level_shifter_up_2.xb_hv.t9 DGND 0.41fF
C657 level_shifter_up_2.xb_hv.t2 DGND 0.20fF
C658 level_shifter_up_2.xb_hv.t4 DGND 0.20fF
C659 level_shifter_up_2.xb_hv.n3 DGND 1.19fF $ **FLOATING
C660 level_shifter_up_2.xb_hv.t6 DGND 0.20fF
C661 level_shifter_up_2.xb_hv.t3 DGND 0.20fF
C662 level_shifter_up_2.xb_hv.n4 DGND 3.16fF $ **FLOATING
C663 trim4b_hv DGND 3.15fF $ **FLOATING
C664 a_32059_903.n0 DGND 0.62fF $ **FLOATING
C665 a_32059_903.n1 DGND 0.63fF $ **FLOATING
C666 a_32059_903.n2 DGND 0.76fF $ **FLOATING
C667 a_32059_903.n3 DGND 0.76fF $ **FLOATING
C668 ibias.t0 DGND 2.10fF
C669 ibias.t2 DGND 0.57fF
C670 ibias.n0 DGND 4.82fF $ **FLOATING
C671 ibias.t5 DGND 0.57fF
C672 ibias.t4 DGND 2.10fF
C673 ibias.t3 DGND 2.10fF
C674 ibias.n1 DGND 2.76fF $ **FLOATING
C675 ibias.n2 DGND 3.10fF $ **FLOATING
C676 ibias.n3 DGND 1.95fF $ **FLOATING
C677 ibias.t6 DGND 2.25fF
C678 ibias.n4 DGND 6.61fF $ **FLOATING
C679 hyst[1].t0 DGND 0.64fF
C680 hyst[1].n0 DGND 4.06fF $ **FLOATING
C681 hyst[1].t3 DGND 0.19fF
C682 hyst[1].t1 DGND 0.20fF
C683 hyst[1].t2 DGND 0.18fF
C684 hyst[1].n1 DGND 0.81fF $ **FLOATING
C685 hyst[1].n2 DGND 0.85fF $ **FLOATING
C686 a_32059_2049.n0 DGND 0.29fF $ **FLOATING
C687 a_32059_2049.n1 DGND 1.12fF $ **FLOATING
C688 a_32059_2049.n2 DGND 0.43fF $ **FLOATING
C689 a_32059_2049.n3 DGND 0.42fF $ **FLOATING
C690 a_32059_2049.n4 DGND 1.13fF $ **FLOATING
C691 a_32059_2049.n5 DGND 0.29fF $ **FLOATING
C692 level_shifter_up_7.x_hv.n0 DGND 1.28fF $ **FLOATING
C693 level_shifter_up_7.x_hv.t5 DGND 0.21fF
C694 level_shifter_up_7.x_hv.n1 DGND 1.83fF $ **FLOATING
C695 level_shifter_up_7.x_hv.t8 DGND 0.48fF
C696 level_shifter_up_7.x_hv.t7 DGND 0.48fF
C697 level_shifter_up_7.x_hv.t4 DGND 0.48fF
C698 level_shifter_up_7.x_hv.t6 DGND 0.48fF
C699 level_shifter_up_7.x_hv.t1 DGND 0.22fF
C700 level_shifter_up_7.x_hv.t3 DGND 0.21fF
C701 level_shifter_up_7.x_hv.n2 DGND 2.28fF $ **FLOATING
C702 level_shifter_up_7.x_hv.t9 DGND 0.22fF
C703 level_shifter_up_7.x_hv.n3 DGND 5.00fF $ **FLOATING
C704 level_shifter_up_7.x_hv.n4 DGND 3.14fF $ **FLOATING
C705 level_shifter_up_7.x_hv.t2 DGND 0.22fF
C706 level_shifter_up_7.x_hv.n5 DGND 1.36fF $ **FLOATING
C707 level_shifter_up_7.x_hv.n6 DGND 2.42fF $ **FLOATING
C708 a_12857_n17742.n0 DGND 0.55fF $ **FLOATING
C709 a_12857_n17742.n1 DGND 0.59fF $ **FLOATING
C710 a_12857_n17742.n2 DGND 0.64fF $ **FLOATING
C711 a_12857_n17742.n3 DGND 0.50fF $ **FLOATING
C712 a_2370_7428.n0 DGND 0.66fF $ **FLOATING
C713 a_2370_7428.n1 DGND 0.66fF $ **FLOATING
C714 a_2370_7428.t10 DGND 3.48fF
C715 a_2370_7428.t9 DGND 3.49fF
C716 a_2370_7428.n2 DGND 4.15fF $ **FLOATING
C717 a_2370_7428.t8 DGND 3.32fF
C718 a_2370_7428.t11 DGND 3.34fF
C719 a_2370_7428.n3 DGND 11.59fF $ **FLOATING
C720 a_2370_7428.n4 DGND 38.63fF $ **FLOATING
C721 a_2370_7428.n5 DGND 2.38fF $ **FLOATING
C722 a_2370_7428.n6 DGND 0.32fF $ **FLOATING
C723 a_2370_7428.n7 DGND 0.31fF $ **FLOATING
C724 a_2370_7428.n8 DGND -0.70fF $ **FLOATING
C725 a_2370_7428.n9 DGND 0.66fF $ **FLOATING
C726 bias_stg2.n0 DGND 1.40fF $ **FLOATING
C727 bias_stg2.n1 DGND 3.06fF $ **FLOATING
C728 bias_stg2.t1 DGND 0.74fF
C729 bias_stg2.t3 DGND 0.68fF
C730 bias_stg2.n2 DGND 1.31fF $ **FLOATING
C731 bias_stg2.n3 DGND 2.80fF $ **FLOATING
C732 bias_stg2.t5 DGND 0.67fF
C733 bias_stg2.t7 DGND 0.67fF
C734 bias_stg2.t6 DGND 0.67fF
C735 bias_stg2.t8 DGND 0.67fF
C736 bias_stg2.t0 DGND 1.70fF
C737 bias_stg2.n4 DGND 3.30fF $ **FLOATING
C738 a_12857_n19016.n0 DGND 4.82fF $ **FLOATING
C739 a_12857_n19016.n1 DGND 10.95fF $ **FLOATING
C740 a_12857_n19016.n2 DGND 21.69fF $ **FLOATING
C741 a_12857_n19016.n3 DGND 3.98fF $ **FLOATING
C742 a_12857_n19016.t12 DGND 1.90fF
C743 a_12857_n19016.t8 DGND 1.90fF
C744 a_12857_n19016.t10 DGND 1.90fF
C745 a_12857_n19016.t11 DGND 1.90fF
C746 a_12857_n19016.t13 DGND 1.90fF
C747 a_12857_n19016.t9 DGND 1.90fF
C748 a_12857_n19016.t6 DGND 1.90fF
C749 a_12857_n19016.t4 DGND 1.90fF
C750 a_12857_n19016.n4 DGND 5.32fF $ **FLOATING
C751 a_12857_n19016.n5 DGND 0.55fF $ **FLOATING
C752 a_12857_n19016.n6 DGND 0.94fF $ **FLOATING
C753 a_33659_n2697.n0 DGND 0.58fF $ **FLOATING
C754 a_33659_n2697.n1 DGND 0.71fF $ **FLOATING
C755 a_33659_n2697.n2 DGND 0.67fF $ **FLOATING
C756 a_32057_n17742.n0 DGND 1.19fF $ **FLOATING
C757 a_32057_n17742.n1 DGND 1.36fF $ **FLOATING
C758 a_32057_n17742.n2 DGND 1.36fF $ **FLOATING
C759 a_32057_n17742.n3 DGND 1.36fF $ **FLOATING
C760 a_32057_n17742.n4 DGND 1.36fF $ **FLOATING
C761 a_32057_n17742.n5 DGND 1.19fF $ **FLOATING
C762 a_32057_n17742.n6 DGND 1.36fF $ **FLOATING
C763 a_32057_n17742.n7 DGND 1.36fF $ **FLOATING
C764 a_32057_n17742.n8 DGND 1.36fF $ **FLOATING
C765 a_32057_n17742.n9 DGND 1.36fF $ **FLOATING
C766 a_32057_n17742.n10 DGND 2.11fF $ **FLOATING
C767 a_32057_n17742.n11 DGND 2.15fF $ **FLOATING
C768 level_shifter_up_3.xb_hv.n0 DGND 1.48fF $ **FLOATING
C769 level_shifter_up_3.xb_hv.n1 DGND 0.53fF $ **FLOATING
C770 level_shifter_up_3.xb_hv.t8 DGND 0.34fF
C771 level_shifter_up_3.xb_hv.t7 DGND 0.34fF
C772 level_shifter_up_3.xb_hv.t10 DGND 0.34fF
C773 level_shifter_up_3.xb_hv.t4 DGND 0.34fF
C774 level_shifter_up_3.xb_hv.t3 DGND 0.34fF
C775 level_shifter_up_3.xb_hv.t5 DGND 0.34fF
C776 level_shifter_up_3.xb_hv.t2 DGND 0.34fF
C777 level_shifter_up_3.xb_hv.t6 DGND 0.34fF
C778 level_shifter_up_3.xb_hv.n2 DGND 0.45fF $ **FLOATING
C779 level_shifter_up_3.xb_hv.n3 DGND 1.09fF $ **FLOATING
C780 trim5b_hv DGND 0.89fF $ **FLOATING
C781 level_shifter_up_3.xb_hv.t9 DGND 0.17fF
C782 level_shifter_up_3.xb_hv.n4 DGND 1.03fF $ **FLOATING
C783 level_shifter_up_3.xb_hv.n5 DGND 0.90fF $ **FLOATING
C784 level_shifter_up_0.x_hv.n0 DGND 14.35fF $ **FLOATING
C785 level_shifter_up_0.x_hv.n1 DGND 0.88fF $ **FLOATING
C786 level_shifter_up_0.x_hv.n2 DGND 0.53fF $ **FLOATING
C787 level_shifter_up_0.x_hv.n3 DGND 0.51fF $ **FLOATING
C788 level_shifter_up_0.x_hv.t9 DGND 0.16fF
C789 level_shifter_up_0.x_hv.t2 DGND 0.16fF
C790 level_shifter_up_0.x_hv.n4 DGND 1.01fF $ **FLOATING
C791 level_shifter_up_0.x_hv.t3 DGND 0.16fF
C792 level_shifter_up_0.x_hv.t10 DGND 0.16fF
C793 level_shifter_up_0.x_hv.t7 DGND 0.16fF
C794 level_shifter_up_0.x_hv.t8 DGND 0.16fF
C795 level_shifter_up_0.x_hv.t4 DGND 0.16fF
C796 level_shifter_up_0.x_hv.n5 DGND 1.03fF $ **FLOATING
C797 level_shifter_up_0.x_hv.t5 DGND 0.16fF
C798 hyst1_hv DGND 8.31fF $ **FLOATING
C799 level_shifter_up_0.x_hv.t6 DGND 0.17fF
C800 level_shifter_up_0.x_hv.n6 DGND 1.07fF $ **FLOATING
C801 a_12857_n15942.n0 DGND 0.54fF $ **FLOATING
C802 a_12857_n15942.n1 DGND 0.52fF $ **FLOATING
C803 a_12857_n15942.n2 DGND 0.61fF $ **FLOATING
C804 a_12857_n15942.n3 DGND 0.58fF $ **FLOATING
C805 en.t1 DGND 0.64fF
C806 en.n0 DGND 5.28fF $ **FLOATING
C807 en.t0 DGND 0.19fF
C808 en.t2 DGND 0.20fF
C809 en.t3 DGND 0.18fF
C810 en.n1 DGND 0.82fF $ **FLOATING
C811 en.n2 DGND 0.85fF $ **FLOATING
C812 a_32059_n3351.n0 DGND 0.38fF $ **FLOATING
C813 a_32059_n3351.n1 DGND 3.11fF $ **FLOATING
C814 a_32059_n3351.t15 DGND 0.11fF
C815 a_32059_n3351.n2 DGND 1.20fF $ **FLOATING
C816 a_32059_n3351.n3 DGND 0.72fF $ **FLOATING
C817 a_32059_n3351.t13 DGND 0.11fF
C818 a_32059_n3351.n4 DGND 1.17fF $ **FLOATING
C819 a_32059_n3351.n5 DGND 0.34fF $ **FLOATING
C820 a_32059_n3351.n6 DGND 0.40fF $ **FLOATING
C821 a_32059_n3351.n7 DGND 0.34fF $ **FLOATING
C822 a_32059_n3351.n8 DGND 0.40fF $ **FLOATING
C823 a_32059_n3351.n9 DGND 3.70fF $ **FLOATING
C824 a_32059_n3351.t9 DGND 0.11fF
C825 a_32059_n3351.n10 DGND 1.09fF $ **FLOATING
C826 a_32059_n3351.n11 DGND 1.12fF $ **FLOATING
C827 a_32059_n3351.n12 DGND 0.55fF $ **FLOATING
C828 trim[2].n0 DGND 0.33fF $ **FLOATING
C829 trim[2].n1 DGND 0.35fF $ **FLOATING
C830 trim[2].n2 DGND 0.81fF $ **FLOATING
C831 trim[2].t2 DGND 0.25fF
C832 trim[0].t3 DGND 0.20fF
C833 trim[0].t1 DGND 0.21fF
C834 trim[0].t2 DGND 0.19fF
C835 trim[0].n0 DGND 0.87fF $ **FLOATING
C836 trim[0].n1 DGND 0.91fF $ **FLOATING
C837 trim[0].n2 DGND 4.00fF $ **FLOATING
C838 trim[0].t0 DGND 0.67fF
C839 DVDD.n0 DGND 0.79fF $ **FLOATING
C840 DVDD.n1 DGND 0.72fF $ **FLOATING
C841 DVDD.n2 DGND 0.11fF $ **FLOATING
C842 DVDD.n4 DGND 0.28fF $ **FLOATING
C843 DVDD.t2 DGND 0.79fF
C844 DVDD.n6 DGND 0.11fF $ **FLOATING
C845 DVDD.n7 DGND 0.11fF $ **FLOATING
C846 DVDD.t6 DGND 0.79fF
C847 DVDD.n9 DGND 0.69fF $ **FLOATING
C848 DVDD.n10 DGND 0.85fF $ **FLOATING
C849 DVDD.n12 DGND 0.23fF $ **FLOATING
C850 DVDD.n13 DGND 0.38fF $ **FLOATING
C851 DVDD.n14 DGND 0.72fF $ **FLOATING
C852 DVDD.n15 DGND 0.11fF $ **FLOATING
C853 DVDD.n18 DGND 0.26fF $ **FLOATING
C854 DVDD.n19 DGND 0.72fF $ **FLOATING
C855 DVDD.n20 DGND 0.11fF $ **FLOATING
C856 DVDD.n22 DGND 0.31fF $ **FLOATING
C857 DVDD.n23 DGND 0.28fF $ **FLOATING
C858 DVDD.n24 DGND 0.11fF $ **FLOATING
C859 DVDD.n25 DGND 0.11fF $ **FLOATING
C860 DVDD.t0 DGND 0.79fF
C861 DVDD.t4 DGND 0.79fF
C862 DVDD.n27 DGND 1.05fF $ **FLOATING
C863 DVDD.n28 DGND 0.31fF $ **FLOATING
C864 DVDD.n29 DGND 0.37fF $ **FLOATING
C865 DVDD.n33 DGND 0.26fF $ **FLOATING
C866 DVDD.t8 DGND 0.45fF
C867 DVDD.n38 DGND 0.17fF $ **FLOATING
C868 DVDD.n39 DGND 0.37fF $ **FLOATING
C869 DVDD.n43 DGND 0.26fF $ **FLOATING
C870 DVDD.n44 DGND 0.37fF $ **FLOATING
C871 DVDD.n48 DGND 0.21fF $ **FLOATING
C872 DVDD.n49 DGND 0.55fF $ **FLOATING
C873 DVDD.t10 DGND 0.45fF
C874 DVDD.n54 DGND 0.13fF $ **FLOATING
C875 DVDD.n55 DGND 0.37fF $ **FLOATING
C876 DVDD.n59 DGND 0.26fF $ **FLOATING
C877 DVDD.n60 DGND 0.37fF $ **FLOATING
C878 DVDD.n64 DGND 0.26fF $ **FLOATING
C879 DVDD.t12 DGND 0.45fF
C880 DVDD.n70 DGND 0.17fF $ **FLOATING
C881 DVDD.n71 DGND 0.44fF $ **FLOATING
C882 DVDD.n74 DGND 0.73fF $ **FLOATING
C883 a_29758_4670.n0 DGND 2.15fF $ **FLOATING
C884 a_29758_4670.n1 DGND 0.79fF $ **FLOATING
C885 a_29758_4670.n2 DGND 0.35fF $ **FLOATING
C886 a_29758_4670.n3 DGND 0.56fF $ **FLOATING
C887 a_29758_4670.n4 DGND 0.56fF $ **FLOATING
C888 a_29758_4670.n5 DGND 0.35fF $ **FLOATING
C889 a_29758_4670.t5 DGND 0.34fF
C890 a_29758_4670.t6 DGND 0.34fF
C891 a_29758_4670.n6 DGND 1.79fF $ **FLOATING
C892 a_29758_4670.t2 DGND 0.33fF
C893 a_29758_4670.t0 DGND 0.33fF
C894 a_29758_4670.t4 DGND 1.52fF
C895 a_24364_11382.t1 DGND 0.14fF
C896 a_24364_11382.t0 DGND 2.17fF
C897 a_23698_4566.t1 DGND 0.13fF
C898 a_23698_4566.t0 DGND 1.97fF
C899 a_34666_7130.n0 DGND 1.12fF $ **FLOATING
C900 a_34666_7130.n1 DGND 1.40fF $ **FLOATING
C901 a_34666_7130.n2 DGND 1.14fF $ **FLOATING
C902 a_34666_7130.n3 DGND 1.10fF $ **FLOATING
C903 a_34666_7130.n4 DGND 1.10fF $ **FLOATING
C904 a_34666_7130.n5 DGND 1.12fF $ **FLOATING
C905 a_34666_7130.n6 DGND 1.46fF $ **FLOATING
C906 a_34666_7130.n7 DGND 1.53fF $ **FLOATING
C907 a_34666_7130.n8 DGND 1.53fF $ **FLOATING
C908 a_34666_7130.n9 DGND 1.03fF $ **FLOATING
C909 a_34666_7130.n10 DGND 1.03fF $ **FLOATING
C910 a_34666_7130.n11 DGND 1.51fF $ **FLOATING
C911 a_34666_7130.n12 DGND 1.51fF $ **FLOATING
C912 a_34666_7130.n13 DGND 1.51fF $ **FLOATING
C913 a_34666_7130.n14 DGND 11.61fF $ **FLOATING
C914 a_34666_7130.n15 DGND 1.53fF $ **FLOATING
C915 a_34666_7130.t16 DGND 0.24fF
C916 a_34666_7130.t12 DGND 0.24fF
C917 a_34666_7130.t10 DGND 0.24fF
C918 a_34666_7130.t2 DGND 0.24fF
C919 a_34666_7130.t17 DGND 0.24fF
C920 a_34666_7130.t14 DGND 0.24fF
C921 a_34666_7130.t5 DGND 0.24fF
C922 a_34666_7130.t8 DGND 0.24fF
C923 a_34666_7130.t7 DGND 0.47fF
C924 a_34666_7130.t9 DGND 0.47fF
C925 a_34666_7130.t15 DGND 0.47fF
C926 a_34666_7130.t18 DGND 0.47fF
C927 a_34666_7130.t6 DGND 0.47fF
C928 a_34666_7130.t19 DGND 0.47fF
C929 a_34666_7130.t3 DGND 0.47fF
C930 a_34666_7130.t11 DGND 0.47fF
C931 a_34666_7130.n35 DGND 11.42fF $ **FLOATING
C932 a_34666_7130.n36 DGND 0.44fF $ **FLOATING
C933 a_34666_7130.n37 DGND 0.43fF $ **FLOATING
C934 a_34666_7130.n38 DGND 0.19fF $ **FLOATING
C935 a_34666_7130.n39 DGND 1.79fF $ **FLOATING
C936 a_34666_7130.n40 DGND 0.66fF $ **FLOATING
C937 a_33659_n1551.n0 DGND 0.97fF $ **FLOATING
C938 a_33659_n1551.n1 DGND 2.70fF $ **FLOATING
C939 a_33659_n1551.n2 DGND 2.66fF $ **FLOATING
C940 a_33659_n1551.n3 DGND 0.29fF $ **FLOATING
C941 level_shifter_up_5.x_hv.t5 DGND 0.13fF
C942 level_shifter_up_5.x_hv.n0 DGND 0.85fF $ **FLOATING
C943 level_shifter_up_5.x_hv.t4 DGND 0.13fF
C944 level_shifter_up_5.x_hv.t2 DGND 0.13fF
C945 level_shifter_up_5.x_hv.n1 DGND 0.54fF $ **FLOATING
C946 level_shifter_up_5.x_hv.t3 DGND 0.13fF
C947 level_shifter_up_5.x_hv.n2 DGND 12.23fF $ **FLOATING
C948 hyst0_hv DGND 7.11fF $ **FLOATING
C949 level_shifter_up_5.x_hv.n3 DGND 1.34fF $ **FLOATING
C950 a_9060_4172.n0 DGND 4.23fF $ **FLOATING
C951 a_9060_4172.t1 DGND 0.75fF
C952 a_9060_4172.n1 DGND 7.68fF $ **FLOATING
C953 a_9060_4172.t0 DGND 0.75fF
C954 a_9060_4530.t5 DGND 0.20fF
C955 a_9060_4530.t4 DGND 1.82fF
C956 a_9060_4530.n0 DGND 19.74fF $ **FLOATING
C957 a_9060_4530.n1 DGND 1.54fF $ **FLOATING
C958 a_9060_4530.n2 DGND 14.17fF $ **FLOATING
C959 a_9060_4530.n3 DGND 2.43fF $ **FLOATING
C960 a_9060_4530.n4 DGND 2.16fF $ **FLOATING
C961 a_9060_4530.n5 DGND 2.13fF $ **FLOATING
C962 a_9060_4530.n6 DGND 1.90fF $ **FLOATING
C963 a_11257_n14142.n0 DGND 3.31fF $ **FLOATING
C964 a_25696_11382.t11 DGND 3.64fF
C965 a_25696_11382.t9 DGND 0.18fF
C966 a_25696_11382.n0 DGND 0.41fF $ **FLOATING
C967 a_25696_11382.t0 DGND 0.18fF
C968 a_25696_11382.t12 DGND 0.18fF
C969 a_25696_11382.n1 DGND 0.41fF $ **FLOATING
C970 a_25696_11382.t13 DGND 0.18fF
C971 a_25696_11382.t5 DGND 0.18fF
C972 a_25696_11382.n2 DGND 0.41fF $ **FLOATING
C973 a_25696_11382.t4 DGND 0.18fF
C974 a_25696_11382.t8 DGND 0.21fF
C975 a_25696_11382.t7 DGND 1.77fF
C976 a_25696_11382.n3 DGND 3.45fF $ **FLOATING
C977 a_25696_11382.n4 DGND 1.11fF $ **FLOATING
C978 a_25696_11382.n5 DGND 0.23fF $ **FLOATING
C979 a_25696_11382.n6 DGND 0.57fF $ **FLOATING
C980 a_25696_11382.n7 DGND 0.57fF $ **FLOATING
C981 a_25696_11382.n8 DGND 0.23fF $ **FLOATING
C982 a_25696_11382.n9 DGND 0.71fF $ **FLOATING
C983 a_25696_11382.n10 DGND 0.71fF $ **FLOATING
C984 a_25696_11382.n11 DGND 0.23fF $ **FLOATING
C985 a_25696_11382.n12 DGND 0.77fF $ **FLOATING
C986 a_25696_11382.n13 DGND 10.90fF $ **FLOATING
C987 a_25696_11382.t1 DGND 4.21fF
C988 a_12857_n14142.n0 DGND 0.55fF $ **FLOATING
C989 a_12857_n14142.n1 DGND 0.59fF $ **FLOATING
C990 a_12857_n14142.n2 DGND 0.64fF $ **FLOATING
C991 a_12857_n14142.n3 DGND 0.50fF $ **FLOATING
C992 a_27936_n27260.t0 DGND 0.15fF
C993 a_27936_n27260.t1 DGND 0.15fF
C994 a_27936_n27260.n0 DGND 1.02fF $ **FLOATING
C995 a_27936_n27260.t2 DGND 0.55fF
C996 a_27936_n27260.n1 DGND 1.19fF $ **FLOATING
C997 a_27936_n27260.t4 DGND 0.15fF
C998 a_27936_n27260.t5 DGND 0.15fF
C999 a_27936_n27260.n2 DGND 1.02fF $ **FLOATING
C1000 a_27936_n27260.t7 DGND 0.15fF
C1001 a_27936_n27260.t6 DGND 0.15fF
C1002 a_27936_n27260.n3 DGND 1.07fF $ **FLOATING
C1003 a_27936_n27260.n4 DGND 0.47fF $ **FLOATING
C1004 a_27936_n27260.n5 DGND 1.21fF $ **FLOATING
C1005 a_27936_n27260.t3 DGND 0.45fF
C1006 level_shifter_up_1.xb_hv.n0 DGND 1.45fF $ **FLOATING
C1007 level_shifter_up_1.xb_hv.n1 DGND 3.67fF $ **FLOATING
C1008 level_shifter_up_1.xb_hv.t4 DGND 0.45fF
C1009 level_shifter_up_1.xb_hv.t3 DGND 0.45fF
C1010 level_shifter_up_1.xb_hv.t2 DGND 0.45fF
C1011 level_shifter_up_1.xb_hv.t1 DGND 0.45fF
C1012 level_shifter_up_1.xb_hv.t6 DGND 0.22fF
C1013 level_shifter_up_1.xb_hv.t7 DGND 0.22fF
C1014 level_shifter_up_1.xb_hv.n2 DGND 3.77fF $ **FLOATING
C1015 level_shifter_up_1.xb_hv.n3 DGND 3.65fF $ **FLOATING
C1016 trim3b_hv DGND 3.73fF $ **FLOATING
C1017 level_shifter_up_1.xb_hv.t5 DGND 0.22fF
C1018 a_32059_n4497.n0 DGND 1.16fF $ **FLOATING
C1019 a_32059_n4497.n1 DGND 2.03fF $ **FLOATING
C1020 a_32059_n4497.n2 DGND 1.16fF $ **FLOATING
C1021 a_32059_n4497.n3 DGND 1.42fF $ **FLOATING
C1022 a_32059_n4497.n4 DGND 1.41fF $ **FLOATING
C1023 a_32059_n4497.n5 DGND 1.29fF $ **FLOATING
C1024 a_32059_n4497.n6 DGND 1.30fF $ **FLOATING
C1025 a_32059_n4497.n7 DGND 1.16fF $ **FLOATING
C1026 a_32059_n4497.n8 DGND 1.16fF $ **FLOATING
C1027 a_29757_7018.n0 DGND 1.59fF $ **FLOATING
C1028 a_29757_7018.t1 DGND 0.40fF
C1029 a_29757_7018.n1 DGND 1.41fF $ **FLOATING
C1030 a_29757_7018.n2 DGND 5.95fF $ **FLOATING
C1031 a_29757_7018.t0 DGND 0.28fF
C1032 Vom_stg2.t3 DGND 0.30fF
C1033 Vom_stg2.t4 DGND 0.46fF
C1034 Vom_stg2.n0 DGND 2.36fF $ **FLOATING
C1035 Vom_stg2.t0 DGND 0.43fF
C1036 Vom_stg2.n1 DGND 1.58fF $ **FLOATING
C1037 a_31098_4670.n0 DGND 1.85fF $ **FLOATING
C1038 a_31098_4670.n1 DGND 0.14fF $ **FLOATING
C1039 a_31098_4670.t1 DGND 0.30fF
C1040 a_31098_4670.n2 DGND 0.77fF $ **FLOATING
C1041 a_31098_4670.n3 DGND 0.42fF $ **FLOATING
C1042 a_31098_4670.n4 DGND 0.22fF $ **FLOATING
C1043 a_31098_4670.n5 DGND 0.41fF $ **FLOATING
C1044 a_31098_4670.n6 DGND 0.42fF $ **FLOATING
C1045 a_31098_4670.t2 DGND 1.10fF
C1046 a_31098_4670.n7 DGND 2.04fF $ **FLOATING
C1047 a_31098_4670.n8 DGND 0.23fF $ **FLOATING
C1048 a_31098_4670.n9 DGND 0.24fF $ **FLOATING
C1049 Vop_stg2.n0 DGND 2.11fF $ **FLOATING
C1050 Vop_stg2.t4 DGND 0.30fF
C1051 Vop_stg2.t3 DGND 0.47fF
C1052 Vop_stg2.n1 DGND 2.42fF $ **FLOATING
C1053 Vop_stg2.t0 DGND 0.44fF
C1054 Vop_stg2.n2 DGND 1.51fF $ **FLOATING
C1055 res_p_bot.n0 DGND 0.53fF $ **FLOATING
C1056 res_p_bot.t9 DGND 0.30fF
C1057 res_p_bot.t3 DGND 0.30fF
C1058 res_p_bot.n1 DGND 0.53fF $ **FLOATING
C1059 res_p_bot.t2 DGND 0.30fF
C1060 res_p_bot.n2 DGND 0.67fF $ **FLOATING
C1061 res_p_bot.n3 DGND 0.30fF $ **FLOATING
C1062 res_p_bot.n4 DGND 0.85fF $ **FLOATING
C1063 res_p_bot.n5 DGND 0.85fF $ **FLOATING
C1064 res_p_bot.n6 DGND 0.29fF $ **FLOATING
C1065 res_p_bot.t13 DGND 0.30fF
C1066 res_p_bot.t7 DGND 1.34fF
C1067 res_p_bot.n7 DGND 2.91fF $ **FLOATING
C1068 res_p_bot.n8 DGND 1.08fF $ **FLOATING
C1069 res_p_bot.n9 DGND 6.93fF $ **FLOATING
C1070 res_p_bot.n10 DGND 11.58fF $ **FLOATING
C1071 res_p_bot.t16 DGND 0.30fF
C1072 res_p_bot.n11 DGND 0.53fF $ **FLOATING
C1073 res_p_bot.t5 DGND 0.30fF
C1074 res_p_bot.n12 DGND 0.67fF $ **FLOATING
C1075 res_p_bot.n13 DGND 0.30fF $ **FLOATING
C1076 res_p_bot.n14 DGND 1.06fF $ **FLOATING
C1077 res_p_bot.t6 DGND 5.40fF
C1078 res_p_bot.n15 DGND 2.82fF $ **FLOATING
C1079 a_32059_n4755.n0 DGND 0.56fF $ **FLOATING
C1080 a_32059_n4755.n1 DGND 0.56fF $ **FLOATING
C1081 a_32059_n4755.n2 DGND 0.56fF $ **FLOATING
C1082 a_32059_n4755.n3 DGND 0.65fF $ **FLOATING
C1083 a_32059_n4755.n4 DGND 0.56fF $ **FLOATING
C1084 a_32059_n4755.n5 DGND 0.56fF $ **FLOATING
C1085 a_32059_n4755.n6 DGND 0.56fF $ **FLOATING
C1086 a_32059_n4755.n7 DGND 0.56fF $ **FLOATING
C1087 a_32059_n4755.t6 DGND 0.16fF
C1088 a_32059_n4755.n8 DGND 2.93fF $ **FLOATING
C1089 a_32059_n4755.n9 DGND 1.73fF $ **FLOATING
C1090 a_32059_n4755.n10 DGND 1.73fF $ **FLOATING
C1091 a_32059_n4755.n11 DGND 1.94fF $ **FLOATING
C1092 a_32059_n4755.t15 DGND 0.16fF
C1093 a_32059_n4755.n12 DGND 2.93fF $ **FLOATING
C1094 a_32059_n4755.n13 DGND 1.73fF $ **FLOATING
C1095 a_32059_n4755.n14 DGND 1.73fF $ **FLOATING
C1096 a_32059_n4755.n15 DGND 1.73fF $ **FLOATING
C1097 a_32059_n4755.n16 DGND 2.67fF $ **FLOATING
C1098 a_32059_n4755.n17 DGND 7.09fF $ **FLOATING
C1099 a_32059_n4755.n18 DGND 5.58fF $ **FLOATING
C1100 a_32059_n4755.n19 DGND 0.68fF $ **FLOATING
C1101 a_32059_n4755.n20 DGND 0.68fF $ **FLOATING
C1102 a_32059_n4755.n21 DGND 0.56fF $ **FLOATING
C1103 a_35086_7130.n0 DGND 1.61fF $ **FLOATING
C1104 a_35086_7130.n1 DGND 1.68fF $ **FLOATING
C1105 a_35086_7130.n2 DGND 1.68fF $ **FLOATING
C1106 a_35086_7130.n3 DGND 1.22fF $ **FLOATING
C1107 a_35086_7130.n4 DGND 1.20fF $ **FLOATING
C1108 a_35086_7130.n5 DGND 1.20fF $ **FLOATING
C1109 a_35086_7130.n6 DGND 1.24fF $ **FLOATING
C1110 a_35086_7130.n7 DGND 1.22fF $ **FLOATING
C1111 a_35086_7130.n8 DGND 0.97fF $ **FLOATING
C1112 a_35086_7130.n9 DGND 0.54fF $ **FLOATING
C1113 a_35086_7130.n10 DGND 1.12fF $ **FLOATING
C1114 a_35086_7130.n11 DGND 1.12fF $ **FLOATING
C1115 a_35086_7130.n12 DGND 1.66fF $ **FLOATING
C1116 a_35086_7130.n13 DGND 1.66fF $ **FLOATING
C1117 a_35086_7130.n14 DGND 1.66fF $ **FLOATING
C1118 a_35086_7130.n15 DGND 11.51fF $ **FLOATING
C1119 a_35086_7130.n16 DGND 1.68fF $ **FLOATING
C1120 a_35086_7130.t15 DGND 0.26fF
C1121 a_35086_7130.t8 DGND 0.26fF
C1122 a_35086_7130.t6 DGND 0.26fF
C1123 a_35086_7130.t17 DGND 0.26fF
C1124 a_35086_7130.t16 DGND 0.26fF
C1125 a_35086_7130.t11 DGND 0.26fF
C1126 a_35086_7130.t18 DGND 0.26fF
C1127 a_35086_7130.t2 DGND 0.26fF
C1128 a_35086_7130.t10 DGND 0.52fF
C1129 a_35086_7130.t12 DGND 0.52fF
C1130 a_35086_7130.t19 DGND 0.52fF
C1131 a_35086_7130.t3 DGND 0.52fF
C1132 a_35086_7130.t9 DGND 0.52fF
C1133 a_35086_7130.t4 DGND 0.52fF
C1134 a_35086_7130.t7 DGND 0.52fF
C1135 a_35086_7130.t13 DGND 0.52fF
C1136 a_35086_7130.n36 DGND 11.90fF $ **FLOATING
C1137 a_35086_7130.n37 DGND 0.48fF $ **FLOATING
C1138 a_35086_7130.n38 DGND 0.48fF $ **FLOATING
C1139 a_35086_7130.n39 DGND 0.17fF $ **FLOATING
C1140 a_35086_7130.n40 DGND 1.92fF $ **FLOATING
C1141 a_35086_7130.n41 DGND 0.74fF $ **FLOATING
C1142 level_shifter_up_4.xb_hv.t1 DGND 1.41fF
C1143 level_shifter_up_4.xb_hv.n0 DGND 1.42fF $ **FLOATING
C1144 level_shifter_up_4.xb_hv.t7 DGND 0.16fF
C1145 level_shifter_up_4.xb_hv.t4 DGND 0.15fF
C1146 level_shifter_up_4.xb_hv.t10 DGND 0.15fF
C1147 level_shifter_up_4.xb_hv.t6 DGND 0.15fF
C1148 level_shifter_up_4.xb_hv.t8 DGND 0.15fF
C1149 level_shifter_up_4.xb_hv.n1 DGND 1.53fF $ **FLOATING
C1150 level_shifter_up_4.xb_hv.t2 DGND 0.34fF
C1151 level_shifter_up_4.xb_hv.t9 DGND 0.34fF
C1152 level_shifter_up_4.xb_hv.t5 DGND 0.34fF
C1153 level_shifter_up_4.xb_hv.t3 DGND 0.34fF
C1154 level_shifter_up_4.xb_hv.n2 DGND 0.42fF $ **FLOATING
C1155 level_shifter_up_4.xb_hv.n3 DGND 0.22fF $ **FLOATING
C1156 level_shifter_up_4.xb_hv.n4 DGND 2.89fF $ **FLOATING
C1157 level_shifter_up_4.xb_hv.n5 DGND 20.23fF $ **FLOATING
C1158 enb_hv DGND 6.43fF $ **FLOATING
C1159 Vinm.n0 DGND 6.19fF $ **FLOATING
C1160 Vinm.t21 DGND 2.39fF
C1161 Vinm.t27 DGND 2.56fF
C1162 Vinm.n1 DGND 4.12fF $ **FLOATING
C1163 Vinm.n2 DGND 2.22fF $ **FLOATING
C1164 Vinm.n3 DGND 2.19fF $ **FLOATING
C1165 Vinm.n4 DGND 2.16fF $ **FLOATING
C1166 Vinm.n5 DGND 2.11fF $ **FLOATING
C1167 Vinm.n6 DGND 2.63fF $ **FLOATING
C1168 Vinm.t48 DGND 2.39fF
C1169 Vinm.t19 DGND 2.39fF
C1170 Vinm.t10 DGND 2.39fF
C1171 Vinm.n7 DGND 3.84fF $ **FLOATING
C1172 Vinm.n8 DGND 1.98fF $ **FLOATING
C1173 Vinm.n9 DGND 2.14fF $ **FLOATING
C1174 Vinm.n10 DGND 2.19fF $ **FLOATING
C1175 Vinm.n11 DGND 1.98fF $ **FLOATING
C1176 Vinm.t55 DGND 2.39fF
C1177 Vinm.n12 DGND 2.16fF $ **FLOATING
C1178 Vinm.n13 DGND 2.10fF $ **FLOATING
C1179 Vinm.n14 DGND 2.56fF $ **FLOATING
C1180 Vinm.t17 DGND 2.39fF
C1181 Vinm.t9 DGND 2.39fF
C1182 Vinm.t23 DGND 2.39fF
C1183 Vinm.t18 DGND 2.40fF
C1184 Vinm.n15 DGND 3.80fF $ **FLOATING
C1185 Vinm.n16 DGND 1.98fF $ **FLOATING
C1186 Vinm.n17 DGND 2.16fF $ **FLOATING
C1187 Vinm.n18 DGND 2.22fF $ **FLOATING
C1188 Vinm.n19 DGND 2.40fF $ **FLOATING
C1189 Vinm.n20 DGND 1.98fF $ **FLOATING
C1190 Vinm.n21 DGND 2.16fF $ **FLOATING
C1191 Vinm.n22 DGND 1.86fF $ **FLOATING
C1192 Vinm.n23 DGND 2.56fF $ **FLOATING
C1193 Vinm.t28 DGND 2.39fF
C1194 Vinm.t52 DGND 2.39fF
C1195 Vinm.t4 DGND 2.28fF
C1196 Vinm.n24 DGND 3.96fF $ **FLOATING
C1197 Vinm.n25 DGND 1.98fF $ **FLOATING
C1198 Vinm.t2 DGND 2.39fF
C1199 Vinm.n26 DGND 2.16fF $ **FLOATING
C1200 Vinm.n27 DGND 2.22fF $ **FLOATING
C1201 Vinm.t42 DGND 2.39fF
C1202 Vinm.n28 DGND 2.40fF $ **FLOATING
C1203 Vinm.n29 DGND 1.98fF $ **FLOATING
C1204 Vinm.n30 DGND 2.16fF $ **FLOATING
C1205 Vinm.n31 DGND 1.86fF $ **FLOATING
C1206 Vinm.n32 DGND 2.56fF $ **FLOATING
C1207 Vinm.t35 DGND 2.39fF
C1208 Vinm.t51 DGND 2.39fF
C1209 Vinm.t41 DGND 2.39fF
C1210 Vinm.n33 DGND 4.20fF $ **FLOATING
C1211 Vinm.n34 DGND 2.16fF $ **FLOATING
C1212 Vinm.n35 DGND 2.22fF $ **FLOATING
C1213 Vinm.n36 DGND 2.40fF $ **FLOATING
C1214 Vinm.n37 DGND 1.98fF $ **FLOATING
C1215 Vinm.t31 DGND 2.39fF
C1216 Vinm.n38 DGND 2.16fF $ **FLOATING
C1217 Vinm.n39 DGND 1.86fF $ **FLOATING
C1218 Vinm.n40 DGND 2.56fF $ **FLOATING
C1219 Vinm.t45 DGND 2.39fF
C1220 Vinm.t54 DGND 2.39fF
C1221 Vinm.t15 DGND 2.39fF
C1222 Vinm.t7 DGND 2.41fF
C1223 Vinm.n41 DGND 3.83fF $ **FLOATING
C1224 Vinm.n42 DGND 2.16fF $ **FLOATING
C1225 Vinm.n43 DGND 2.01fF $ **FLOATING
C1226 Vinm.n44 DGND 1.95fF $ **FLOATING
C1227 Vinm.n45 DGND 2.16fF $ **FLOATING
C1228 Vinm.n46 DGND 1.98fF $ **FLOATING
C1229 Vinm.n47 DGND 2.26fF $ **FLOATING
C1230 Vinm.n48 DGND 2.59fF $ **FLOATING
C1231 Vinm.t3 DGND 2.39fF
C1232 Vinm.t29 DGND 2.39fF
C1233 Vinm.t22 DGND 2.39fF
C1234 Vinm.n49 DGND 4.09fF $ **FLOATING
C1235 Vinm.n50 DGND 2.38fF $ **FLOATING
C1236 Vinm.n51 DGND 2.40fF $ **FLOATING
C1237 Vinm.t11 DGND 2.39fF
C1238 Vinm.n52 DGND 2.19fF $ **FLOATING
C1239 Vinm.n53 DGND 2.11fF $ **FLOATING
C1240 Vinm.n54 DGND 2.79fF $ **FLOATING
C1241 Vinm.t46 DGND 2.39fF
C1242 Vinm.t56 DGND 2.56fF
C1243 Vinm.n55 DGND 6.60fF $ **FLOATING
C1244 Vinm.n56 DGND 20.40fF $ **FLOATING
C1245 Vinm.n57 DGND 5.78fF $ **FLOATING
C1246 Vinm.t53 DGND 2.41fF
C1247 Vinm.t33 DGND 2.55fF
C1248 Vinm.n58 DGND 3.49fF $ **FLOATING
C1249 Vinm.n59 DGND 2.39fF $ **FLOATING
C1250 Vinm.n60 DGND 2.41fF $ **FLOATING
C1251 Vinm.n61 DGND 2.20fF $ **FLOATING
C1252 Vinm.n62 DGND 2.03fF $ **FLOATING
C1253 Vinm.n63 DGND 2.00fF $ **FLOATING
C1254 Vinm.t50 DGND 2.41fF
C1255 Vinm.t20 DGND 2.41fF
C1256 Vinm.t12 DGND 2.41fF
C1257 Vinm.n64 DGND 3.24fF $ **FLOATING
C1258 Vinm.n65 DGND 2.18fF $ **FLOATING
C1259 Vinm.n66 DGND 2.02fF $ **FLOATING
C1260 Vinm.n67 DGND 1.96fF $ **FLOATING
C1261 Vinm.n68 DGND 2.18fF $ **FLOATING
C1262 Vinm.t34 DGND 2.41fF
C1263 Vinm.n69 DGND 1.99fF $ **FLOATING
C1264 Vinm.n70 DGND 2.19fF $ **FLOATING
C1265 Vinm.n71 DGND 2.34fF $ **FLOATING
C1266 Vinm.t16 DGND 2.43fF
C1267 Vinm.n72 DGND 3.01fF $ **FLOATING
C1268 Vinm.n73 DGND 2.18fF $ **FLOATING
C1269 Vinm.t24 DGND 2.41fF
C1270 Vinm.n74 DGND 2.23fF $ **FLOATING
C1271 Vinm.n75 DGND 2.41fF $ **FLOATING
C1272 Vinm.t6 DGND 2.41fF
C1273 Vinm.n76 DGND 1.99fF $ **FLOATING
C1274 Vinm.n77 DGND 2.18fF $ **FLOATING
C1275 Vinm.t43 DGND 2.41fF
C1276 Vinm.n78 DGND 1.79fF $ **FLOATING
C1277 Vinm.n79 DGND 2.31fF $ **FLOATING
C1278 Vinm.t26 DGND 2.41fF
C1279 Vinm.t39 DGND 2.41fF
C1280 Vinm.t1 DGND 2.41fF
C1281 Vinm.t49 DGND 2.41fF
C1282 Vinm.n80 DGND 3.01fF $ **FLOATING
C1283 Vinm.n81 DGND 2.18fF $ **FLOATING
C1284 Vinm.n82 DGND 2.23fF $ **FLOATING
C1285 Vinm.n83 DGND 2.41fF $ **FLOATING
C1286 Vinm.n84 DGND 1.99fF $ **FLOATING
C1287 Vinm.n85 DGND 2.18fF $ **FLOATING
C1288 Vinm.n86 DGND 1.79fF $ **FLOATING
C1289 Vinm.n87 DGND 2.31fF $ **FLOATING
C1290 Vinm.t32 DGND 2.41fF
C1291 Vinm.t44 DGND 2.41fF
C1292 Vinm.t36 DGND 2.41fF
C1293 Vinm.n88 DGND 3.01fF $ **FLOATING
C1294 Vinm.n89 DGND 2.18fF $ **FLOATING
C1295 Vinm.n90 DGND 2.23fF $ **FLOATING
C1296 Vinm.n91 DGND 2.41fF $ **FLOATING
C1297 Vinm.n92 DGND 1.99fF $ **FLOATING
C1298 Vinm.n93 DGND 2.18fF $ **FLOATING
C1299 Vinm.t14 DGND 2.41fF
C1300 Vinm.n94 DGND 1.79fF $ **FLOATING
C1301 Vinm.n95 DGND 2.31fF $ **FLOATING
C1302 Vinm.t25 DGND 2.41fF
C1303 Vinm.t38 DGND 2.41fF
C1304 Vinm.t0 DGND 2.41fF
C1305 Vinm.t47 DGND 2.42fF
C1306 Vinm.n96 DGND 3.24fF $ **FLOATING
C1307 Vinm.n97 DGND 1.99fF $ **FLOATING
C1308 Vinm.n98 DGND 2.15fF $ **FLOATING
C1309 Vinm.n99 DGND 2.20fF $ **FLOATING
C1310 Vinm.n100 DGND 1.99fF $ **FLOATING
C1311 Vinm.n101 DGND 2.18fF $ **FLOATING
C1312 Vinm.n102 DGND 2.03fF $ **FLOATING
C1313 Vinm.n103 DGND 2.31fF $ **FLOATING
C1314 Vinm.t40 DGND 2.41fF
C1315 Vinm.t13 DGND 2.41fF
C1316 Vinm.t5 DGND 2.41fF
C1317 Vinm.n104 DGND 3.52fF $ **FLOATING
C1318 Vinm.n105 DGND 2.23fF $ **FLOATING
C1319 Vinm.n106 DGND 2.20fF $ **FLOATING
C1320 Vinm.n107 DGND 2.18fF $ **FLOATING
C1321 Vinm.t30 DGND 2.41fF
C1322 Vinm.n108 DGND 2.03fF $ **FLOATING
C1323 Vinm.n109 DGND 2.55fF $ **FLOATING
C1324 Vinm.t8 DGND 2.41fF
C1325 Vinm.t37 DGND 2.55fF
C1326 Vinm.n110 DGND 5.58fF $ **FLOATING
C1327 Vinm.n111 DGND 26.94fF $ **FLOATING
C1328 a_2370_n28652.n0 DGND 0.50fF $ **FLOATING
C1329 a_2370_n28652.n1 DGND 0.61fF $ **FLOATING
C1330 a_2370_n28652.n2 DGND 0.61fF $ **FLOATING
C1331 a_2370_n28652.t10 DGND 3.08fF
C1332 a_2370_n28652.t8 DGND 3.10fF
C1333 a_2370_n28652.n3 DGND 4.08fF $ **FLOATING
C1334 a_2370_n28652.t11 DGND 3.21fF
C1335 a_2370_n28652.t9 DGND 3.23fF
C1336 a_2370_n28652.n4 DGND 10.29fF $ **FLOATING
C1337 a_2370_n28652.n5 DGND 36.35fF $ **FLOATING
C1338 a_2370_n28652.n6 DGND 2.13fF $ **FLOATING
C1339 a_2370_n28652.n7 DGND 0.29fF $ **FLOATING
C1340 a_2370_n28652.n9 DGND 0.61fF $ **FLOATING
C1341 level_shifter_up_3.x_hv.n0 DGND 1.15fF $ **FLOATING
C1342 level_shifter_up_3.x_hv.n1 DGND 0.79fF $ **FLOATING
C1343 level_shifter_up_3.x_hv.t3 DGND 0.13fF
C1344 level_shifter_up_3.x_hv.n2 DGND 0.84fF $ **FLOATING
C1345 level_shifter_up_3.x_hv.t4 DGND 0.28fF
C1346 level_shifter_up_3.x_hv.t6 DGND 0.28fF
C1347 level_shifter_up_3.x_hv.t5 DGND 0.28fF
C1348 level_shifter_up_3.x_hv.t2 DGND 0.28fF
C1349 level_shifter_up_3.x_hv.t7 DGND 0.28fF
C1350 level_shifter_up_3.x_hv.t10 DGND 0.28fF
C1351 level_shifter_up_3.x_hv.t9 DGND 0.28fF
C1352 level_shifter_up_3.x_hv.t8 DGND 0.28fF
C1353 level_shifter_up_3.x_hv.n3 DGND 0.73fF $ **FLOATING
C1354 trim5_hv DGND 1.03fF $ **FLOATING
C1355 a_32057_n14142.n0 DGND 1.49fF $ **FLOATING
C1356 a_32057_n14142.n1 DGND 1.71fF $ **FLOATING
C1357 a_32057_n14142.n2 DGND 1.71fF $ **FLOATING
C1358 a_32057_n14142.n3 DGND 1.71fF $ **FLOATING
C1359 a_32057_n14142.n4 DGND 1.49fF $ **FLOATING
C1360 a_32057_n14142.n5 DGND 1.71fF $ **FLOATING
C1361 a_32057_n14142.n6 DGND 1.71fF $ **FLOATING
C1362 a_32057_n14142.n7 DGND 1.71fF $ **FLOATING
C1363 a_32057_n14142.n8 DGND 1.71fF $ **FLOATING
C1364 a_32057_n14142.n9 DGND 1.58fF $ **FLOATING
C1365 a_32057_n14142.n10 DGND 1.49fF $ **FLOATING
C1366 a_32057_n14142.n11 DGND 1.71fF $ **FLOATING
C1367 a_32057_n14142.n12 DGND 1.71fF $ **FLOATING
C1368 a_32057_n14142.n13 DGND 1.71fF $ **FLOATING
C1369 a_32057_n14142.n14 DGND 1.71fF $ **FLOATING
C1370 a_32057_n14142.n15 DGND 2.45fF $ **FLOATING
C1371 a_32057_n14142.n16 DGND 2.14fF $ **FLOATING
C1372 a_32057_n14142.n17 DGND 2.45fF $ **FLOATING
C1373 a_32057_n14142.n18 DGND 1.71fF $ **FLOATING
C1374 trim[3].t0 DGND 0.10fF
C1375 trim[3].n0 DGND 0.43fF $ **FLOATING
C1376 trim[3].n1 DGND 0.45fF $ **FLOATING
C1377 trim[3].n2 DGND 0.55fF $ **FLOATING
C1378 trim[3].t1 DGND 0.33fF
C1379 bias_n.n0 DGND 1.88fF $ **FLOATING
C1380 bias_n.n1 DGND 2.05fF $ **FLOATING
C1381 bias_n.n2 DGND 1.88fF $ **FLOATING
C1382 bias_n.n3 DGND 1.88fF $ **FLOATING
C1383 bias_n.n4 DGND 1.88fF $ **FLOATING
C1384 bias_n.n5 DGND 2.05fF $ **FLOATING
C1385 bias_n.n6 DGND 2.05fF $ **FLOATING
C1386 bias_n.n7 DGND 2.05fF $ **FLOATING
C1387 bias_n.n8 DGND 1.88fF $ **FLOATING
C1388 bias_n.n9 DGND 2.05fF $ **FLOATING
C1389 bias_n.n10 DGND 2.05fF $ **FLOATING
C1390 bias_n.n11 DGND 2.05fF $ **FLOATING
C1391 bias_n.n12 DGND 1.88fF $ **FLOATING
C1392 bias_n.n13 DGND 2.05fF $ **FLOATING
C1393 bias_n.n14 DGND 2.05fF $ **FLOATING
C1394 bias_n.n15 DGND 2.05fF $ **FLOATING
C1395 bias_n.n16 DGND 1.88fF $ **FLOATING
C1396 bias_n.n17 DGND 2.05fF $ **FLOATING
C1397 bias_n.n18 DGND 2.05fF $ **FLOATING
C1398 bias_n.n19 DGND 2.05fF $ **FLOATING
C1399 bias_n.n20 DGND 1.88fF $ **FLOATING
C1400 bias_n.n21 DGND 2.05fF $ **FLOATING
C1401 bias_n.n22 DGND 2.05fF $ **FLOATING
C1402 bias_n.n23 DGND 2.05fF $ **FLOATING
C1403 bias_n.n24 DGND 1.88fF $ **FLOATING
C1404 bias_n.n25 DGND 2.44fF $ **FLOATING
C1405 bias_n.n26 DGND 2.05fF $ **FLOATING
C1406 bias_n.n27 DGND 2.05fF $ **FLOATING
C1407 bias_n.n28 DGND 2.44fF $ **FLOATING
C1408 bias_n.n29 DGND 2.05fF $ **FLOATING
C1409 bias_n.n30 DGND 2.05fF $ **FLOATING
C1410 bias_n.n31 DGND 1.89fF $ **FLOATING
C1411 bias_n.n32 DGND 2.24fF $ **FLOATING
C1412 bias_n.n33 DGND 1.89fF $ **FLOATING
C1413 bias_n.n34 DGND 2.25fF $ **FLOATING
C1414 bias_n.n35 DGND 2.08fF $ **FLOATING
C1415 bias_n.n36 DGND 1.89fF $ **FLOATING
C1416 bias_n.n37 DGND 2.08fF $ **FLOATING
C1417 bias_n.n38 DGND 1.89fF $ **FLOATING
C1418 bias_n.n39 DGND 2.08fF $ **FLOATING
C1419 bias_n.n40 DGND 1.92fF $ **FLOATING
C1420 bias_n.t5 DGND 1.70fF
C1421 bias_n.n41 DGND 0.31fF $ **FLOATING
C1422 bias_n.t80 DGND 1.48fF
C1423 bias_n.t57 DGND 1.48fF
C1424 bias_n.n42 DGND 0.31fF $ **FLOATING
C1425 bias_n.t9 DGND 1.48fF
C1426 bias_n.t74 DGND 1.48fF
C1427 bias_n.n43 DGND 1.14fF $ **FLOATING
C1428 bias_n.n44 DGND 0.31fF $ **FLOATING
C1429 bias_n.t73 DGND 1.48fF
C1430 bias_n.t34 DGND 1.48fF
C1431 bias_n.n45 DGND 0.31fF $ **FLOATING
C1432 bias_n.t56 DGND 1.48fF
C1433 bias_n.t19 DGND 1.48fF
C1434 bias_n.n46 DGND 1.66fF $ **FLOATING
C1435 bias_n.n47 DGND 0.31fF $ **FLOATING
C1436 bias_n.t32 DGND 1.48fF
C1437 bias_n.t11 DGND 1.48fF
C1438 bias_n.n48 DGND 0.31fF $ **FLOATING
C1439 bias_n.t18 DGND 1.48fF
C1440 bias_n.t83 DGND 1.48fF
C1441 bias_n.n49 DGND 1.66fF $ **FLOATING
C1442 bias_n.n50 DGND 0.31fF $ **FLOATING
C1443 bias_n.t10 DGND 1.48fF
C1444 bias_n.t77 DGND 1.48fF
C1445 bias_n.n51 DGND 0.31fF $ **FLOATING
C1446 bias_n.t82 DGND 1.48fF
C1447 bias_n.t63 DGND 1.48fF
C1448 bias_n.n52 DGND 1.66fF $ **FLOATING
C1449 bias_n.n53 DGND 0.31fF $ **FLOATING
C1450 bias_n.t76 DGND 1.48fF
C1451 bias_n.t36 DGND 1.48fF
C1452 bias_n.n54 DGND 0.31fF $ **FLOATING
C1453 bias_n.t60 DGND 1.48fF
C1454 bias_n.t22 DGND 1.48fF
C1455 bias_n.n55 DGND 1.66fF $ **FLOATING
C1456 bias_n.n56 DGND 0.31fF $ **FLOATING
C1457 bias_n.t35 DGND 1.48fF
C1458 bias_n.t81 DGND 1.48fF
C1459 bias_n.n57 DGND 0.31fF $ **FLOATING
C1460 bias_n.t21 DGND 1.48fF
C1461 bias_n.t66 DGND 1.48fF
C1462 bias_n.n58 DGND 1.66fF $ **FLOATING
C1463 bias_n.n59 DGND 0.31fF $ **FLOATING
C1464 bias_n.t27 DGND 1.48fF
C1465 bias_n.t8 DGND 1.48fF
C1466 bias_n.n60 DGND 1.52fF $ **FLOATING
C1467 bias_n.n61 DGND 1.79fF $ **FLOATING
C1468 bias_n.n62 DGND 1.35fF $ **FLOATING
C1469 bias_n.n63 DGND 1.35fF $ **FLOATING
C1470 bias_n.n64 DGND 1.35fF $ **FLOATING
C1471 bias_n.n65 DGND 1.35fF $ **FLOATING
C1472 bias_n.n66 DGND 0.25fF $ **FLOATING
C1473 bias_n.n67 DGND 0.31fF $ **FLOATING
C1474 bias_n.t59 DGND 1.48fF
C1475 bias_n.t46 DGND 1.48fF
C1476 bias_n.n68 DGND 0.31fF $ **FLOATING
C1477 bias_n.t31 DGND 1.48fF
C1478 bias_n.t62 DGND 1.48fF
C1479 bias_n.n69 DGND 1.04fF $ **FLOATING
C1480 bias_n.n70 DGND 0.31fF $ **FLOATING
C1481 bias_n.t45 DGND 1.48fF
C1482 bias_n.t87 DGND 1.48fF
C1483 bias_n.n71 DGND 0.31fF $ **FLOATING
C1484 bias_n.t85 DGND 1.48fF
C1485 bias_n.t64 DGND 1.48fF
C1486 bias_n.n72 DGND 1.20fF $ **FLOATING
C1487 bias_n.n73 DGND 0.31fF $ **FLOATING
C1488 bias_n.t24 DGND 1.48fF
C1489 bias_n.t53 DGND 1.48fF
C1490 bias_n.n74 DGND 0.31fF $ **FLOATING
C1491 bias_n.t54 DGND 1.48fF
C1492 bias_n.t17 DGND 1.48fF
C1493 bias_n.n75 DGND 0.31fF $ **FLOATING
C1494 bias_n.t67 DGND 1.48fF
C1495 bias_n.t39 DGND 1.48fF
C1496 bias_n.n76 DGND 0.31fF $ **FLOATING
C1497 bias_n.t28 DGND 1.48fF
C1498 bias_n.t70 DGND 1.48fF
C1499 bias_n.n77 DGND 0.93fF $ **FLOATING
C1500 bias_n.n78 DGND 1.06fF $ **FLOATING
C1501 bias_n.n79 DGND 0.31fF $ **FLOATING
C1502 bias_n.t47 DGND 1.48fF
C1503 bias_n.t14 DGND 1.48fF
C1504 bias_n.t88 DGND 1.55fF
C1505 bias_n.n80 DGND 1.80fF $ **FLOATING
C1506 bias_n.n81 DGND 1.38fF $ **FLOATING
C1507 bias_n.n82 DGND 5.77fF $ **FLOATING
C1508 bias_n.n83 DGND 6.21fF $ **FLOATING
C1509 bias_n.n84 DGND 0.43fF $ **FLOATING
C1510 bias_n.n85 DGND 2.48fF $ **FLOATING
C1511 bias_n.n86 DGND 3.82fF $ **FLOATING
C1512 bias_n.n87 DGND 1.26fF $ **FLOATING
C1513 bias_n.n88 DGND 1.49fF $ **FLOATING
C1514 bias_n.t4 DGND 1.48fF
C1515 bias_n.t6 DGND 1.48fF
C1516 bias_n.n90 DGND 0.31fF $ **FLOATING
C1517 bias_n.t38 DGND 1.48fF
C1518 bias_n.t69 DGND 1.48fF
C1519 bias_n.n91 DGND 0.31fF $ **FLOATING
C1520 bias_n.t79 DGND 1.48fF
C1521 bias_n.t37 DGND 1.48fF
C1522 bias_n.n92 DGND 1.14fF $ **FLOATING
C1523 bias_n.n93 DGND 1.14fF $ **FLOATING
C1524 bias_n.n94 DGND 0.31fF $ **FLOATING
C1525 bias_n.t52 DGND 1.48fF
C1526 bias_n.t26 DGND 1.48fF
C1527 bias_n.n95 DGND 0.31fF $ **FLOATING
C1528 bias_n.t23 DGND 1.48fF
C1529 bias_n.t65 DGND 1.48fF
C1530 bias_n.n96 DGND 1.66fF $ **FLOATING
C1531 bias_n.n97 DGND 1.66fF $ **FLOATING
C1532 bias_n.n98 DGND 0.31fF $ **FLOATING
C1533 bias_n.t13 DGND 1.48fF
C1534 bias_n.t48 DGND 1.48fF
C1535 bias_n.n99 DGND 0.31fF $ **FLOATING
C1536 bias_n.t50 DGND 1.48fF
C1537 bias_n.t12 DGND 1.48fF
C1538 bias_n.n100 DGND 1.66fF $ **FLOATING
C1539 bias_n.n101 DGND 1.66fF $ **FLOATING
C1540 bias_n.n102 DGND 0.31fF $ **FLOATING
C1541 bias_n.t42 DGND 1.48fF
C1542 bias_n.t75 DGND 1.48fF
C1543 bias_n.n103 DGND 0.31fF $ **FLOATING
C1544 bias_n.t84 DGND 1.48fF
C1545 bias_n.t41 DGND 1.48fF
C1546 bias_n.n104 DGND 1.66fF $ **FLOATING
C1547 bias_n.n105 DGND 1.66fF $ **FLOATING
C1548 bias_n.n106 DGND 0.31fF $ **FLOATING
C1549 bias_n.t61 DGND 1.48fF
C1550 bias_n.t33 DGND 1.48fF
C1551 bias_n.n107 DGND 1.66fF $ **FLOATING
C1552 bias_n.n108 DGND 0.31fF $ **FLOATING
C1553 bias_n.t20 DGND 1.48fF
C1554 bias_n.t71 DGND 1.48fF
C1555 bias_n.n109 DGND 0.31fF $ **FLOATING
C1556 bias_n.t58 DGND 1.48fF
C1557 bias_n.t40 DGND 1.48fF
C1558 bias_n.n110 DGND 0.31fF $ **FLOATING
C1559 bias_n.t30 DGND 1.48fF
C1560 bias_n.t72 DGND 1.48fF
C1561 bias_n.n111 DGND 1.66fF $ **FLOATING
C1562 bias_n.n112 DGND 1.66fF $ **FLOATING
C1563 bias_n.n113 DGND 1.66fF $ **FLOATING
C1564 bias_n.n114 DGND 0.31fF $ **FLOATING
C1565 bias_n.t16 DGND 1.48fF
C1566 bias_n.t49 DGND 1.48fF
C1567 bias_n.n115 DGND 0.31fF $ **FLOATING
C1568 bias_n.t86 DGND 1.48fF
C1569 bias_n.t43 DGND 1.48fF
C1570 bias_n.n116 DGND 1.13fF $ **FLOATING
C1571 bias_n.n117 DGND 0.31fF $ **FLOATING
C1572 bias_n.t51 DGND 1.48fF
C1573 bias_n.t15 DGND 1.48fF
C1574 bias_n.n118 DGND 1.66fF $ **FLOATING
C1575 bias_n.n119 DGND 0.31fF $ **FLOATING
C1576 bias_n.t44 DGND 1.48fF
C1577 bias_n.t78 DGND 1.48fF
C1578 bias_n.n120 DGND 2.09fF $ **FLOATING
C1579 bias_n.n121 DGND 0.31fF $ **FLOATING
C1580 bias_n.t55 DGND 1.48fF
C1581 bias_n.t29 DGND 1.48fF
C1582 bias_n.n122 DGND 0.31fF $ **FLOATING
C1583 bias_n.t25 DGND 1.48fF
C1584 bias_n.t68 DGND 1.48fF
C1585 bias_n.n123 DGND 1.66fF $ **FLOATING
C1586 bias_n.n124 DGND 1.46fF $ **FLOATING
C1587 trim[5].t3 DGND 0.10fF
C1588 trim[5].n0 DGND 0.42fF $ **FLOATING
C1589 trim[5].n1 DGND 0.44fF $ **FLOATING
C1590 trim[5].n2 DGND 0.55fF $ **FLOATING
C1591 trim[5].t1 DGND 0.33fF
C1592 a_32057_n9600.n0 DGND 0.45fF $ **FLOATING
C1593 a_32057_n9600.t0 DGND 0.11fF
C1594 a_32057_n9600.n1 DGND 1.69fF $ **FLOATING
C1595 a_32057_n9600.t5 DGND 0.11fF
C1596 a_32057_n9600.n2 DGND 1.89fF $ **FLOATING
C1597 a_32057_n9600.n3 DGND 1.11fF $ **FLOATING
C1598 a_32057_n9600.n4 DGND 0.82fF $ **FLOATING
C1599 a_32057_n9600.n5 DGND 8.22fF $ **FLOATING
C1600 a_32057_n9600.n6 DGND 0.45fF $ **FLOATING
C1601 a_32057_n9600.t6 DGND 0.13fF
C1602 a_32057_n9600.n7 DGND 0.81fF $ **FLOATING
C1603 a_32057_n9600.n8 DGND 7.82fF $ **FLOATING
C1604 a_32057_n9600.n9 DGND 0.81fF $ **FLOATING
C1605 a_32057_n9600.t10 DGND 0.13fF
C1606 level_shifter_up_5.xb_hv.n0 DGND 0.87fF $ **FLOATING
C1607 level_shifter_up_5.xb_hv.n1 DGND 2.07fF $ **FLOATING
C1608 level_shifter_up_5.xb_hv.n2 DGND 0.91fF $ **FLOATING
C1609 level_shifter_up_5.xb_hv.t4 DGND 0.35fF
C1610 level_shifter_up_5.xb_hv.n3 DGND 2.29fF $ **FLOATING
C1611 level_shifter_up_5.xb_hv.t3 DGND 0.36fF
C1612 level_shifter_up_5.xb_hv.t2 DGND 0.35fF
C1613 level_shifter_up_5.xb_hv.n4 DGND 2.00fF $ **FLOATING
C1614 level_shifter_up_5.xb_hv.t5 DGND 0.35fF
C1615 level_shifter_up_5.xb_hv.t8 DGND 0.36fF
C1616 level_shifter_up_5.xb_hv.t7 DGND 0.35fF
C1617 level_shifter_up_5.xb_hv.t6 DGND 0.35fF
C1618 level_shifter_up_5.xb_hv.n5 DGND 5.10fF $ **FLOATING
C1619 hyst0b_hv DGND 6.14fF $ **FLOATING
C1620 level_shifter_up_5.xb_hv.t1 DGND 3.49fF
C1621 a_23032_4566.n0 DGND 1.53fF $ **FLOATING
C1622 a_23032_4566.n1 DGND 0.91fF $ **FLOATING
C1623 a_23032_4566.n2 DGND 0.91fF $ **FLOATING
C1624 a_23032_4566.n3 DGND 0.91fF $ **FLOATING
C1625 a_23032_4566.n4 DGND 6.17fF $ **FLOATING
C1626 a_23032_4566.t4 DGND 0.26fF
C1627 a_23032_4566.n5 DGND 0.61fF $ **FLOATING
C1628 a_23032_4566.t7 DGND 0.26fF
C1629 a_23032_4566.t17 DGND 0.26fF
C1630 a_23032_4566.n6 DGND 0.61fF $ **FLOATING
C1631 a_23032_4566.t16 DGND 0.26fF
C1632 a_23032_4566.n7 DGND 0.61fF $ **FLOATING
C1633 a_23032_4566.n8 DGND 0.57fF $ **FLOATING
C1634 a_23032_4566.n9 DGND 0.60fF $ **FLOATING
C1635 a_23032_4566.n10 DGND 1.29fF $ **FLOATING
C1636 a_23032_4566.n11 DGND 0.30fF $ **FLOATING
C1637 a_23032_4566.n12 DGND 0.83fF $ **FLOATING
C1638 a_23032_4566.n13 DGND 0.83fF $ **FLOATING
C1639 a_23032_4566.n14 DGND 0.30fF $ **FLOATING
C1640 a_23032_4566.n15 DGND 2.22fF $ **FLOATING
C1641 a_23032_4566.t3 DGND 22.39fF
C1642 a_2370_6628.n0 DGND 0.66fF $ **FLOATING
C1643 a_2370_6628.t8 DGND 3.36fF
C1644 a_2370_6628.t11 DGND 3.43fF
C1645 a_2370_6628.n1 DGND 4.61fF $ **FLOATING
C1646 a_2370_6628.t10 DGND 3.22fF
C1647 a_2370_6628.t9 DGND 3.30fF
C1648 a_2370_6628.n2 DGND 13.73fF $ **FLOATING
C1649 a_2370_6628.n3 DGND 33.48fF $ **FLOATING
C1650 a_2370_6628.n4 DGND 3.06fF $ **FLOATING
C1651 a_2370_6628.n5 DGND 0.66fF $ **FLOATING
C1652 a_2370_6628.n6 DGND 0.49fF $ **FLOATING
C1653 a_2370_6628.n7 DGND 0.23fF $ **FLOATING
C1654 a_2370_6628.n8 DGND 0.85fF $ **FLOATING
C1655 a_2370_6628.n9 DGND 0.66fF $ **FLOATING
C1656 level_shifter_up_8.xb_hv.n0 DGND 1.42fF $ **FLOATING
C1657 level_shifter_up_8.xb_hv.n1 DGND 2.16fF $ **FLOATING
C1658 level_shifter_up_8.xb_hv.n2 DGND 6.15fF $ **FLOATING
C1659 level_shifter_up_8.xb_hv.t8 DGND 0.56fF
C1660 level_shifter_up_8.xb_hv.t5 DGND 0.56fF
C1661 level_shifter_up_8.xb_hv.t6 DGND 0.56fF
C1662 level_shifter_up_8.xb_hv.t4 DGND 0.56fF
C1663 level_shifter_up_8.xb_hv.t1 DGND 0.56fF
C1664 level_shifter_up_8.xb_hv.t2 DGND 0.56fF
C1665 level_shifter_up_8.xb_hv.t3 DGND 0.56fF
C1666 level_shifter_up_8.xb_hv.t9 DGND 0.56fF
C1667 level_shifter_up_8.xb_hv.n3 DGND 2.94fF $ **FLOATING
C1668 level_shifter_up_8.xb_hv.t7 DGND 0.26fF
C1669 a_11257_n8742.n0 DGND 0.71fF $ **FLOATING
C1670 a_11257_n8742.n1 DGND 0.80fF $ **FLOATING
C1671 a_11257_n8742.n2 DGND 0.79fF $ **FLOATING
C1672 a_11257_n8742.n3 DGND 0.70fF $ **FLOATING
C1673 a_11257_n8742.t10 DGND 0.11fF
C1674 a_11257_n8742.n4 DGND 1.51fF $ **FLOATING
C1675 a_11257_n8742.n5 DGND 0.88fF $ **FLOATING
C1676 a_11257_n8742.n6 DGND 1.36fF $ **FLOATING
C1677 a_11257_n8742.n7 DGND 2.06fF $ **FLOATING
C1678 a_11257_n8742.n8 DGND 0.65fF $ **FLOATING
C1679 a_11257_n8742.n9 DGND 0.83fF $ **FLOATING
C1680 a_11257_n8742.n10 DGND 1.42fF $ **FLOATING
C1681 a_11257_n8742.t5 DGND 0.11fF
C1682 a_11160_n9542.n0 DGND 4.52fF $ **FLOATING
C1683 a_11160_n9542.n1 DGND 2.21fF $ **FLOATING
C1684 a_11160_n9542.n2 DGND 1.90fF $ **FLOATING
C1685 a_11160_n9542.n3 DGND 0.83fF $ **FLOATING
C1686 a_11160_n9542.n4 DGND 0.76fF $ **FLOATING
C1687 a_11160_n9542.t6 DGND 0.17fF
C1688 a_11160_n9542.n5 DGND 0.40fF $ **FLOATING
C1689 a_11160_n9542.t2 DGND 0.17fF
C1690 a_11160_n9542.n6 DGND 1.59fF $ **FLOATING
C1691 a_11160_n9542.t4 DGND 0.17fF
C1692 a_11160_n9542.t10 DGND 0.17fF
C1693 a_11160_n9542.t0 DGND 0.17fF
C1694 a_11160_n9542.t14 DGND 1.61fF
C1695 a_11160_n9542.t13 DGND 1.61fF
C1696 a_11160_n9542.n8 DGND 0.12fF $ **FLOATING
C1697 a_11160_n9542.n9 DGND 0.12fF $ **FLOATING
C1698 a_11160_n9542.t12 DGND 0.77fF
C1699 a_11160_n9542.t8 DGND 0.17fF
C1700 a_11160_n9542.n10 DGND 0.40fF $ **FLOATING
C1701 a_32057_n13616.t13 DGND 0.10fF
C1702 a_32057_n13616.n0 DGND 0.84fF $ **FLOATING
C1703 a_32057_n13616.n1 DGND 1.14fF $ **FLOATING
C1704 a_32057_n13616.n2 DGND 1.14fF $ **FLOATING
C1705 a_32057_n13616.n3 DGND 0.84fF $ **FLOATING
C1706 a_32057_n13616.t25 DGND 0.10fF
C1707 a_32057_n13616.n4 DGND 1.75fF $ **FLOATING
C1708 a_32057_n13616.n5 DGND 0.84fF $ **FLOATING
C1709 a_32057_n13616.n6 DGND 1.14fF $ **FLOATING
C1710 a_32057_n13616.n7 DGND 1.14fF $ **FLOATING
C1711 a_32057_n13616.n8 DGND 0.84fF $ **FLOATING
C1712 a_32057_n13616.t29 DGND 0.10fF
C1713 a_32057_n13616.n9 DGND 1.75fF $ **FLOATING
C1714 a_32057_n13616.t35 DGND 0.11fF
C1715 a_32057_n13616.t7 DGND 0.11fF
C1716 a_32057_n13616.n10 DGND 0.82fF $ **FLOATING
C1717 a_32057_n13616.t39 DGND 0.11fF
C1718 a_32057_n13616.t0 DGND 0.11fF
C1719 a_32057_n13616.n11 DGND 0.82fF $ **FLOATING
C1720 a_32057_n13616.t33 DGND 0.11fF
C1721 a_32057_n13616.t3 DGND 0.11fF
C1722 a_32057_n13616.n12 DGND 0.82fF $ **FLOATING
C1723 a_32057_n13616.t2 DGND 0.11fF
C1724 a_32057_n13616.t5 DGND 0.11fF
C1725 a_32057_n13616.n13 DGND 0.82fF $ **FLOATING
C1726 a_32057_n13616.t32 DGND 0.11fF
C1727 a_32057_n13616.t37 DGND 0.11fF
C1728 a_32057_n13616.n14 DGND 0.82fF $ **FLOATING
C1729 a_32057_n13616.t1 DGND 0.11fF
C1730 a_32057_n13616.t36 DGND 0.11fF
C1731 a_32057_n13616.n15 DGND 0.82fF $ **FLOATING
C1732 a_32057_n13616.t34 DGND 0.11fF
C1733 a_32057_n13616.t4 DGND 0.11fF
C1734 a_32057_n13616.n16 DGND 0.82fF $ **FLOATING
C1735 a_32057_n13616.t38 DGND 0.11fF
C1736 a_32057_n13616.t6 DGND 0.11fF
C1737 a_32057_n13616.n17 DGND 0.82fF $ **FLOATING
C1738 a_32057_n13616.n18 DGND 1.11fF $ **FLOATING
C1739 a_32057_n13616.n19 DGND 1.11fF $ **FLOATING
C1740 a_32057_n13616.n20 DGND 1.11fF $ **FLOATING
C1741 a_32057_n13616.n21 DGND 7.56fF $ **FLOATING
C1742 a_32057_n13616.t19 DGND 0.10fF
C1743 a_32057_n13616.n22 DGND 1.75fF $ **FLOATING
C1744 a_32057_n13616.n23 DGND 1.96fF $ **FLOATING
C1745 a_32057_n13616.n24 DGND 1.14fF $ **FLOATING
C1746 a_32057_n13616.n25 DGND 1.14fF $ **FLOATING
C1747 a_32057_n13616.n26 DGND 0.84fF $ **FLOATING
C1748 a_32057_n13616.n27 DGND 7.76fF $ **FLOATING
C1749 a_32057_n13616.n28 DGND 2.38fF $ **FLOATING
C1750 a_32057_n13616.n29 DGND 2.38fF $ **FLOATING
C1751 a_32057_n13616.n30 DGND 2.36fF $ **FLOATING
C1752 a_32057_n13616.n31 DGND 2.36fF $ **FLOATING
C1753 a_32057_n13616.n32 DGND 1.96fF $ **FLOATING
C1754 a_32057_n13616.n33 DGND 1.14fF $ **FLOATING
C1755 a_32057_n13616.n34 DGND 1.14fF $ **FLOATING
C1756 a_32057_n13616.n35 DGND 0.84fF $ **FLOATING
C1757 a_32057_n13616.n36 DGND 1.53fF $ **FLOATING
C1758 a_32057_n13616.n37 DGND 1.75fF $ **FLOATING
C1759 a_32057_n8742.n0 DGND 0.92fF $ **FLOATING
C1760 a_32057_n8742.n1 DGND 1.05fF $ **FLOATING
C1761 a_32057_n8742.n2 DGND 1.05fF $ **FLOATING
C1762 a_32057_n8742.n3 DGND 0.92fF $ **FLOATING
C1763 a_32057_n8742.n4 DGND 1.05fF $ **FLOATING
C1764 a_32057_n8742.n5 DGND 1.05fF $ **FLOATING
C1765 bias_var_n.n0 DGND 3.85fF $ **FLOATING
C1766 bias_var_n.n1 DGND 3.85fF $ **FLOATING
C1767 bias_var_n.n2 DGND 1.34fF $ **FLOATING
C1768 bias_var_n.n3 DGND 3.85fF $ **FLOATING
C1769 bias_var_n.n4 DGND 3.85fF $ **FLOATING
C1770 bias_var_n.n5 DGND 3.92fF $ **FLOATING
C1771 bias_var_n.n6 DGND 1.93fF $ **FLOATING
C1772 bias_var_n.n7 DGND 3.85fF $ **FLOATING
C1773 bias_var_n.n8 DGND 3.24fF $ **FLOATING
C1774 bias_var_n.n9 DGND 7.20fF $ **FLOATING
C1775 bias_var_n.n10 DGND 2.73fF $ **FLOATING
C1776 bias_var_n.n11 DGND 2.73fF $ **FLOATING
C1777 bias_var_n.n12 DGND 2.54fF $ **FLOATING
C1778 bias_var_n.n13 DGND 5.39fF $ **FLOATING
C1779 bias_var_n.n14 DGND 2.73fF $ **FLOATING
C1780 bias_var_n.n15 DGND 2.54fF $ **FLOATING
C1781 bias_var_n.n16 DGND 2.54fF $ **FLOATING
C1782 bias_var_n.n17 DGND 2.73fF $ **FLOATING
C1783 bias_var_n.n18 DGND 2.73fF $ **FLOATING
C1784 bias_var_n.n19 DGND 2.73fF $ **FLOATING
C1785 bias_var_n.n20 DGND 2.54fF $ **FLOATING
C1786 bias_var_n.n21 DGND 2.73fF $ **FLOATING
C1787 bias_var_n.n22 DGND 2.73fF $ **FLOATING
C1788 bias_var_n.n23 DGND 2.73fF $ **FLOATING
C1789 bias_var_n.n24 DGND 2.54fF $ **FLOATING
C1790 bias_var_n.n25 DGND 2.73fF $ **FLOATING
C1791 bias_var_n.n26 DGND 2.73fF $ **FLOATING
C1792 bias_var_n.n27 DGND 2.73fF $ **FLOATING
C1793 bias_var_n.n28 DGND 2.54fF $ **FLOATING
C1794 bias_var_n.n29 DGND 2.73fF $ **FLOATING
C1795 bias_var_n.n30 DGND 2.73fF $ **FLOATING
C1796 bias_var_n.n31 DGND 3.19fF $ **FLOATING
C1797 bias_var_n.n32 DGND 2.73fF $ **FLOATING
C1798 bias_var_n.n33 DGND 2.73fF $ **FLOATING
C1799 bias_var_n.n34 DGND 2.73fF $ **FLOATING
C1800 bias_var_n.n35 DGND 2.73fF $ **FLOATING
C1801 bias_var_n.n36 DGND 4.12fF $ **FLOATING
C1802 bias_var_n.t39 DGND 1.72fF
C1803 bias_var_n.t10 DGND 1.72fF
C1804 bias_var_n.t42 DGND 1.72fF
C1805 bias_var_n.t11 DGND 1.72fF
C1806 bias_var_n.t22 DGND 1.72fF
C1807 bias_var_n.t49 DGND 1.72fF
C1808 bias_var_n.t58 DGND 1.72fF
C1809 bias_var_n.t29 DGND 1.72fF
C1810 bias_var_n.t7 DGND 1.72fF
C1811 bias_var_n.t46 DGND 1.72fF
C1812 bias_var_n.t8 DGND 1.72fF
C1813 bias_var_n.t40 DGND 1.72fF
C1814 bias_var_n.t27 DGND 1.72fF
C1815 bias_var_n.t13 DGND 1.72fF
C1816 bias_var_n.t41 DGND 1.72fF
C1817 bias_var_n.t28 DGND 1.72fF
C1818 bias_var_n.t19 DGND 1.72fF
C1819 bias_var_n.t48 DGND 1.72fF
C1820 bias_var_n.t35 DGND 1.72fF
C1821 bias_var_n.t21 DGND 1.72fF
C1822 bias_var_n.t44 DGND 1.72fF
C1823 bias_var_n.t31 DGND 1.72fF
C1824 bias_var_n.n37 DGND 1.31fF $ **FLOATING
C1825 bias_var_n.t37 DGND 1.72fF
C1826 bias_var_n.t57 DGND 1.72fF
C1827 bias_var_n.t61 DGND 1.72fF
C1828 bias_var_n.t36 DGND 1.72fF
C1829 bias_var_n.n38 DGND 1.31fF $ **FLOATING
C1830 bias_var_n.t60 DGND 1.72fF
C1831 bias_var_n.t38 DGND 1.72fF
C1832 bias_var_n.t12 DGND 1.72fF
C1833 bias_var_n.t45 DGND 1.72fF
C1834 bias_var_n.n39 DGND 2.07fF $ **FLOATING
C1835 bias_var_n.n40 DGND 1.93fF $ **FLOATING
C1836 bias_var_n.t63 DGND 1.72fF
C1837 bias_var_n.t43 DGND 1.72fF
C1838 bias_var_n.t17 DGND 1.72fF
C1839 bias_var_n.t62 DGND 1.72fF
C1840 bias_var_n.t50 DGND 1.72fF
C1841 bias_var_n.t14 DGND 1.72fF
C1842 bias_var_n.t32 DGND 1.72fF
C1843 bias_var_n.t18 DGND 1.72fF
C1844 bias_var_n.t30 DGND 1.72fF
C1845 bias_var_n.t53 DGND 1.72fF
C1846 bias_var_n.t23 DGND 1.72fF
C1847 bias_var_n.t9 DGND 1.72fF
C1848 bias_var_n.t16 DGND 1.72fF
C1849 bias_var_n.t47 DGND 1.72fF
C1850 bias_var_n.t51 DGND 1.72fF
C1851 bias_var_n.t15 DGND 1.72fF
C1852 bias_var_n.n41 DGND 1.93fF $ **FLOATING
C1853 bias_var_n.t54 DGND 1.72fF
C1854 bias_var_n.t24 DGND 1.72fF
C1855 bias_var_n.t33 DGND 1.72fF
C1856 bias_var_n.t20 DGND 1.72fF
C1857 bias_var_n.t59 DGND 1.72fF
C1858 bias_var_n.t34 DGND 1.72fF
C1859 bias_var_n.n42 DGND 3.19fF $ **FLOATING
C1860 bias_var_n.t52 DGND 1.72fF
C1861 bias_var_n.t26 DGND 1.72fF
C1862 bias_var_n.t25 DGND 1.72fF
C1863 bias_var_n.t56 DGND 1.72fF
C1864 bias_var_n.n43 DGND 0.86fF $ **FLOATING
C1865 bias_var_n.n44 DGND 0.50fF $ **FLOATING
C1866 bias_var_n.n45 DGND 4.43fF $ **FLOATING
C1867 bias_var_n.n46 DGND 1.31fF $ **FLOATING
C1868 Vinp.n0 DGND 6.35fF $ **FLOATING
C1869 Vinp.t44 DGND 2.53fF
C1870 Vinp.t51 DGND 2.77fF
C1871 Vinp.n1 DGND 3.85fF $ **FLOATING
C1872 Vinp.n2 DGND 2.86fF $ **FLOATING
C1873 Vinp.n3 DGND 2.83fF $ **FLOATING
C1874 Vinp.n4 DGND 2.28fF $ **FLOATING
C1875 Vinp.n5 DGND 1.89fF $ **FLOATING
C1876 Vinp.n6 DGND 1.85fF $ **FLOATING
C1877 Vinp.t19 DGND 2.53fF
C1878 Vinp.t41 DGND 2.53fF
C1879 Vinp.t32 DGND 2.55fF
C1880 Vinp.n7 DGND 4.05fF $ **FLOATING
C1881 Vinp.n8 DGND 2.28fF $ **FLOATING
C1882 Vinp.n9 DGND 2.13fF $ **FLOATING
C1883 Vinp.n10 DGND 2.07fF $ **FLOATING
C1884 Vinp.n11 DGND 2.28fF $ **FLOATING
C1885 Vinp.n12 DGND 2.10fF $ **FLOATING
C1886 Vinp.t0 DGND 2.53fF
C1887 Vinp.n13 DGND 2.30fF $ **FLOATING
C1888 Vinp.n14 DGND 2.47fF $ **FLOATING
C1889 Vinp.t38 DGND 2.53fF
C1890 Vinp.t29 DGND 2.53fF
C1891 Vinp.t55 DGND 2.53fF
C1892 Vinp.t45 DGND 2.53fF
C1893 Vinp.n15 DGND 4.95fF $ **FLOATING
C1894 Vinp.n16 DGND 2.28fF $ **FLOATING
C1895 Vinp.n17 DGND 1.85fF $ **FLOATING
C1896 Vinp.n18 DGND 2.03fF $ **FLOATING
C1897 Vinp.n19 DGND 2.10fF $ **FLOATING
C1898 Vinp.n20 DGND 2.28fF $ **FLOATING
C1899 Vinp.n21 DGND 2.14fF $ **FLOATING
C1900 Vinp.n22 DGND 2.69fF $ **FLOATING
C1901 Vinp.t9 DGND 2.53fF
C1902 Vinp.t34 DGND 2.53fF
C1903 Vinp.t23 DGND 2.53fF
C1904 Vinp.n23 DGND 4.50fF $ **FLOATING
C1905 Vinp.n24 DGND 2.10fF $ **FLOATING
C1906 Vinp.n25 DGND 2.28fF $ **FLOATING
C1907 Vinp.n26 DGND 1.85fF $ **FLOATING
C1908 Vinp.n27 DGND 2.03fF $ **FLOATING
C1909 Vinp.n28 DGND 2.10fF $ **FLOATING
C1910 Vinp.t14 DGND 2.53fF
C1911 Vinp.n29 DGND 2.28fF $ **FLOATING
C1912 Vinp.n30 DGND 2.14fF $ **FLOATING
C1913 Vinp.n31 DGND 2.69fF $ **FLOATING
C1914 Vinp.t8 DGND 2.53fF
C1915 Vinp.t2 DGND 2.53fF
C1916 Vinp.t24 DGND 2.53fF
C1917 Vinp.t13 DGND 2.53fF
C1918 Vinp.t52 DGND 2.47fF
C1919 Vinp.n32 DGND 4.65fF $ **FLOATING
C1920 Vinp.n33 DGND 2.10fF $ **FLOATING
C1921 Vinp.n34 DGND 2.28fF $ **FLOATING
C1922 Vinp.n35 DGND 1.85fF $ **FLOATING
C1923 Vinp.n36 DGND 2.03fF $ **FLOATING
C1924 Vinp.n37 DGND 2.10fF $ **FLOATING
C1925 Vinp.n38 DGND 2.28fF $ **FLOATING
C1926 Vinp.n39 DGND 2.14fF $ **FLOATING
C1927 Vinp.n40 DGND 2.69fF $ **FLOATING
C1928 Vinp.t17 DGND 2.53fF
C1929 Vinp.t46 DGND 2.53fF
C1930 Vinp.t37 DGND 2.53fF
C1931 Vinp.n41 DGND 4.06fF $ **FLOATING
C1932 Vinp.n42 DGND 2.10fF $ **FLOATING
C1933 Vinp.n43 DGND 2.25fF $ **FLOATING
C1934 Vinp.n44 DGND 2.31fF $ **FLOATING
C1935 Vinp.n45 DGND 2.10fF $ **FLOATING
C1936 Vinp.t25 DGND 2.53fF
C1937 Vinp.n46 DGND 2.28fF $ **FLOATING
C1938 Vinp.n47 DGND 2.14fF $ **FLOATING
C1939 Vinp.n48 DGND 2.44fF $ **FLOATING
C1940 Vinp.t3 DGND 2.53fF
C1941 Vinp.t36 DGND 2.53fF
C1942 Vinp.t50 DGND 2.53fF
C1943 Vinp.t43 DGND 2.55fF
C1944 Vinp.n49 DGND 3.82fF $ **FLOATING
C1945 Vinp.n50 DGND 3.01fF $ **FLOATING
C1946 Vinp.n51 DGND 3.04fF $ **FLOATING
C1947 Vinp.n52 DGND 2.31fF $ **FLOATING
C1948 Vinp.n53 DGND 1.89fF $ **FLOATING
C1949 Vinp.n54 DGND 2.44fF $ **FLOATING
C1950 Vinp.t20 DGND 2.78fF
C1951 Vinp.t12 DGND 2.53fF
C1952 Vinp.n55 DGND 7.06fF $ **FLOATING
C1953 Vinp.n56 DGND 20.62fF $ **FLOATING
C1954 Vinp.n57 DGND 6.41fF $ **FLOATING
C1955 Vinp.t28 DGND 2.55fF
C1956 Vinp.t56 DGND 2.76fF
C1957 Vinp.n58 DGND 3.18fF $ **FLOATING
C1958 Vinp.n59 DGND 3.03fF $ **FLOATING
C1959 Vinp.n60 DGND 3.06fF $ **FLOATING
C1960 Vinp.n61 DGND 2.32fF $ **FLOATING
C1961 Vinp.n62 DGND 1.99fF $ **FLOATING
C1962 Vinp.n63 DGND 2.34fF $ **FLOATING
C1963 Vinp.t22 DGND 2.55fF
C1964 Vinp.t42 DGND 2.55fF
C1965 Vinp.t33 DGND 2.56fF
C1966 Vinp.n64 DGND 3.43fF $ **FLOATING
C1967 Vinp.n65 DGND 2.11fF $ **FLOATING
C1968 Vinp.n66 DGND 2.27fF $ **FLOATING
C1969 Vinp.n67 DGND 2.32fF $ **FLOATING
C1970 Vinp.n68 DGND 2.11fF $ **FLOATING
C1971 Vinp.n69 DGND 2.30fF $ **FLOATING
C1972 Vinp.t7 DGND 2.55fF
C1973 Vinp.n70 DGND 2.24fF $ **FLOATING
C1974 Vinp.n71 DGND 2.71fF $ **FLOATING
C1975 Vinp.t10 DGND 2.55fF
C1976 Vinp.t27 DGND 2.55fF
C1977 Vinp.t54 DGND 2.55fF
C1978 Vinp.t47 DGND 2.55fF
C1979 Vinp.n72 DGND 3.69fF $ **FLOATING
C1980 Vinp.n73 DGND 2.30fF $ **FLOATING
C1981 Vinp.n74 DGND 1.86fF $ **FLOATING
C1982 Vinp.n75 DGND 2.04fF $ **FLOATING
C1983 Vinp.n76 DGND 2.11fF $ **FLOATING
C1984 Vinp.n77 DGND 2.30fF $ **FLOATING
C1985 Vinp.n78 DGND 2.25fF $ **FLOATING
C1986 Vinp.n79 DGND 2.95fF $ **FLOATING
C1987 Vinp.t6 DGND 2.55fF
C1988 Vinp.t31 DGND 2.55fF
C1989 Vinp.t21 DGND 2.55fF
C1990 Vinp.n80 DGND 3.69fF $ **FLOATING
C1991 Vinp.n81 DGND 2.30fF $ **FLOATING
C1992 Vinp.n82 DGND 1.86fF $ **FLOATING
C1993 Vinp.n83 DGND 2.04fF $ **FLOATING
C1994 Vinp.n84 DGND 2.11fF $ **FLOATING
C1995 Vinp.n85 DGND 2.30fF $ **FLOATING
C1996 Vinp.t49 DGND 2.55fF
C1997 Vinp.n86 DGND 2.25fF $ **FLOATING
C1998 Vinp.n87 DGND 2.95fF $ **FLOATING
C1999 Vinp.t35 DGND 2.55fF
C2000 Vinp.t53 DGND 2.55fF
C2001 Vinp.t15 DGND 2.55fF
C2002 Vinp.t11 DGND 2.55fF
C2003 Vinp.n88 DGND 3.69fF $ **FLOATING
C2004 Vinp.n89 DGND 2.30fF $ **FLOATING
C2005 Vinp.n90 DGND 1.86fF $ **FLOATING
C2006 Vinp.n91 DGND 2.04fF $ **FLOATING
C2007 Vinp.n92 DGND 2.11fF $ **FLOATING
C2008 Vinp.n93 DGND 2.30fF $ **FLOATING
C2009 Vinp.n94 DGND 2.25fF $ **FLOATING
C2010 Vinp.n95 DGND 2.95fF $ **FLOATING
C2011 Vinp.t5 DGND 2.55fF
C2012 Vinp.t30 DGND 2.55fF
C2013 Vinp.t18 DGND 2.55fF
C2014 Vinp.n96 DGND 3.42fF $ **FLOATING
C2015 Vinp.n97 DGND 2.30fF $ **FLOATING
C2016 Vinp.n98 DGND 2.14fF $ **FLOATING
C2017 Vinp.n99 DGND 2.08fF $ **FLOATING
C2018 Vinp.n100 DGND 2.30fF $ **FLOATING
C2019 Vinp.t48 DGND 2.55fF
C2020 Vinp.n101 DGND 2.11fF $ **FLOATING
C2021 Vinp.n102 DGND 2.40fF $ **FLOATING
C2022 Vinp.n103 DGND 2.73fF $ **FLOATING
C2023 Vinp.t26 DGND 2.57fF
C2024 Vinp.n104 DGND 3.21fF $ **FLOATING
C2025 Vinp.t39 DGND 2.55fF
C2026 Vinp.n105 DGND 2.87fF $ **FLOATING
C2027 Vinp.t16 DGND 2.55fF
C2028 Vinp.n106 DGND 2.84fF $ **FLOATING
C2029 Vinp.n107 DGND 2.30fF $ **FLOATING
C2030 Vinp.t1 DGND 2.55fF
C2031 Vinp.n108 DGND 1.99fF $ **FLOATING
C2032 Vinp.n109 DGND 2.71fF $ **FLOATING
C2033 Vinp.t40 DGND 2.55fF
C2034 Vinp.t4 DGND 2.75fF
C2035 Vinp.n110 DGND 6.19fF $ **FLOATING
C2036 Vinp.n111 DGND 28.03fF $ **FLOATING
C2037 a_32059_n897.n0 DGND 1.00fF $ **FLOATING
C2038 a_32059_n897.n1 DGND 1.22fF $ **FLOATING
C2039 a_32059_n897.n2 DGND 1.22fF $ **FLOATING
C2040 a_32059_n897.n3 DGND 1.22fF $ **FLOATING
C2041 a_32059_n897.n4 DGND 1.22fF $ **FLOATING
C2042 a_32059_n897.n5 DGND 1.00fF $ **FLOATING
C2043 a_2458_6570.t5 DGND 1.68fF
C2044 a_2458_6570.t12 DGND 1.68fF
C2045 a_2458_6570.t1 DGND 1.68fF
C2046 a_2458_6570.t13 DGND 1.68fF
C2047 a_2458_6570.t4 DGND 1.68fF
C2048 a_2458_6570.t3 DGND 1.68fF
C2049 a_2458_6570.t2 DGND 1.81fF
C2050 a_2458_6570.n0 DGND 7.68fF $ **FLOATING
C2051 a_2458_6570.n1 DGND 2.60fF $ **FLOATING
C2052 a_2458_6570.n2 DGND 4.01fF $ **FLOATING
C2053 a_2458_6570.n3 DGND 1.51fF $ **FLOATING
C2054 a_2458_6570.n4 DGND 0.90fF $ **FLOATING
C2055 a_2458_6570.n5 DGND 0.90fF $ **FLOATING
C2056 a_2458_6570.n6 DGND 0.90fF $ **FLOATING
C2057 a_2458_6570.n7 DGND 4.91fF $ **FLOATING
C2058 a_2458_6570.n8 DGND 31.58fF $ **FLOATING
C2059 a_2458_6570.n9 DGND 19.10fF $ **FLOATING
C2060 a_2458_6570.n10 DGND 2.60fF $ **FLOATING
C2061 a_2458_6570.n11 DGND 7.68fF $ **FLOATING
C2062 a_2458_6570.t0 DGND 1.82fF
C2063 a_32057_n15000.n0 DGND 0.46fF $ **FLOATING
C2064 a_32057_n15000.n1 DGND 0.46fF $ **FLOATING
C2065 a_32057_n15000.n2 DGND 0.46fF $ **FLOATING
C2066 a_32057_n15000.n3 DGND 0.46fF $ **FLOATING
C2067 a_32057_n15000.t9 DGND 0.11fF
C2068 a_32057_n15000.n4 DGND 1.92fF $ **FLOATING
C2069 a_32057_n15000.n5 DGND 1.12fF $ **FLOATING
C2070 a_32057_n15000.n6 DGND 0.93fF $ **FLOATING
C2071 a_32057_n15000.t16 DGND 0.11fF
C2072 a_32057_n15000.n7 DGND 1.63fF $ **FLOATING
C2073 a_32057_n15000.t1 DGND 0.11fF
C2074 a_32057_n15000.n8 DGND 1.92fF $ **FLOATING
C2075 a_32057_n15000.n9 DGND 1.12fF $ **FLOATING
C2076 a_32057_n15000.n10 DGND 0.93fF $ **FLOATING
C2077 a_32057_n15000.t8 DGND 0.11fF
C2078 a_32057_n15000.n11 DGND 1.63fF $ **FLOATING
C2079 a_32057_n15000.t4 DGND 0.11fF
C2080 a_32057_n15000.n12 DGND 1.92fF $ **FLOATING
C2081 a_32057_n15000.n13 DGND 1.12fF $ **FLOATING
C2082 a_32057_n15000.n14 DGND 0.93fF $ **FLOATING
C2083 a_32057_n15000.t10 DGND 0.11fF
C2084 a_32057_n15000.n15 DGND 1.63fF $ **FLOATING
C2085 a_32057_n15000.n16 DGND 1.67fF $ **FLOATING
C2086 a_32057_n15000.n17 DGND 2.56fF $ **FLOATING
C2087 a_32057_n15000.n18 DGND 6.82fF $ **FLOATING
C2088 a_32057_n15000.n19 DGND 0.46fF $ **FLOATING
C2089 a_32057_n15000.n20 DGND 0.46fF $ **FLOATING
C2090 a_32057_n15000.n21 DGND 0.55fF $ **FLOATING
C2091 a_32057_n15000.n22 DGND 0.52fF $ **FLOATING
C2092 a_32057_n15000.n23 DGND 0.32fF $ **FLOATING
C2093 a_32057_n15000.n24 DGND 5.85fF $ **FLOATING
C2094 a_32057_n15000.n25 DGND 0.21fF $ **FLOATING
C2095 a_32057_n15000.n26 DGND 0.33fF $ **FLOATING
C2096 a_32057_n15000.n27 DGND 0.33fF $ **FLOATING
C2097 a_32057_n15000.n28 DGND 0.52fF $ **FLOATING
C2098 a_32057_n15000.n29 DGND 0.55fF $ **FLOATING
C2099 level_shifter_up_0.xb_hv.n0 DGND 3.51fF $ **FLOATING
C2100 level_shifter_up_0.xb_hv.n1 DGND 3.76fF $ **FLOATING
C2101 level_shifter_up_0.xb_hv.n2 DGND 3.58fF $ **FLOATING
C2102 level_shifter_up_0.xb_hv.t4 DGND 0.31fF
C2103 level_shifter_up_0.xb_hv.n3 DGND 1.64fF $ **FLOATING
C2104 level_shifter_up_0.xb_hv.n7 DGND 0.19fF $ **FLOATING
C2105 level_shifter_up_0.xb_hv.t2 DGND 0.31fF
C2106 level_shifter_up_0.xb_hv.n8 DGND 0.19fF $ **FLOATING
C2107 level_shifter_up_0.xb_hv.n9 DGND 0.19fF $ **FLOATING
C2108 level_shifter_up_0.xb_hv.t14 DGND 0.31fF
C2109 level_shifter_up_0.xb_hv.t6 DGND 0.30fF
C2110 level_shifter_up_0.xb_hv.t5 DGND 0.30fF
C2111 level_shifter_up_0.xb_hv.n10 DGND 1.86fF $ **FLOATING
C2112 level_shifter_up_0.xb_hv.n11 DGND 1.65fF $ **FLOATING
C2113 level_shifter_up_0.xb_hv.t13 DGND 0.30fF
C2114 level_shifter_up_0.xb_hv.t10 DGND 0.30fF
C2115 level_shifter_up_0.xb_hv.t15 DGND 0.30fF
C2116 level_shifter_up_0.xb_hv.t12 DGND 0.30fF
C2117 level_shifter_up_0.xb_hv.t16 DGND 0.30fF
C2118 level_shifter_up_0.xb_hv.t8 DGND 0.30fF
C2119 level_shifter_up_0.xb_hv.t18 DGND 0.30fF
C2120 level_shifter_up_0.xb_hv.t9 DGND 0.30fF
C2121 level_shifter_up_0.xb_hv.t11 DGND 0.30fF
C2122 level_shifter_up_0.xb_hv.t17 DGND 0.31fF
C2123 level_shifter_up_0.xb_hv.t3 DGND 0.31fF
C2124 level_shifter_up_0.xb_hv.t7 DGND 0.30fF
C2125 level_shifter_up_0.xb_hv.n18 DGND 6.46fF $ **FLOATING
C2126 hyst1b_hv DGND 4.66fF $ **FLOATING
C2127 a_2467_n30310.n0 DGND 1.53fF $ **FLOATING
C2128 a_2467_n30310.n1 DGND 1.53fF $ **FLOATING
C2129 a_2467_n30310.n2 DGND 1.70fF $ **FLOATING
C2130 a_2467_n30310.n3 DGND 1.53fF $ **FLOATING
C2131 a_2467_n30310.n4 DGND 1.70fF $ **FLOATING
C2132 a_2467_n30310.n5 DGND 1.53fF $ **FLOATING
C2133 a_2467_n30310.n6 DGND 1.70fF $ **FLOATING
C2134 a_2467_n30310.n7 DGND 1.53fF $ **FLOATING
C2135 a_2467_n30310.n8 DGND 1.70fF $ **FLOATING
C2136 a_2467_n30310.n9 DGND 1.53fF $ **FLOATING
C2137 a_2467_n30310.n10 DGND 2.55fF $ **FLOATING
C2138 a_2467_n30310.n11 DGND 1.95fF $ **FLOATING
C2139 a_2467_n30310.n12 DGND 1.78fF $ **FLOATING
C2140 a_2467_n30310.n13 DGND 2.21fF $ **FLOATING
C2141 a_2467_n30310.t58 DGND 0.18fF
C2142 a_2467_n30310.n14 DGND 5.29fF $ **FLOATING
C2143 a_2467_n30310.t6 DGND 0.18fF
C2144 a_2467_n30310.n15 DGND 4.14fF $ **FLOATING
C2145 a_2467_n30310.t64 DGND 0.18fF
C2146 a_2467_n30310.n16 DGND 4.14fF $ **FLOATING
C2147 a_2467_n30310.t29 DGND 0.18fF
C2148 a_2467_n30310.n17 DGND 5.18fF $ **FLOATING
C2149 a_2467_n30310.t38 DGND 0.18fF
C2150 a_2467_n30310.t11 DGND 0.18fF
C2151 a_2467_n30310.t27 DGND 0.18fF
C2152 a_2467_n30310.t10 DGND 0.18fF
C2153 a_2467_n30310.n18 DGND 5.38fF $ **FLOATING
C2154 a_2467_n30310.n19 DGND 4.14fF $ **FLOATING
C2155 a_2467_n30310.n20 DGND 4.14fF $ **FLOATING
C2156 a_2467_n30310.n21 DGND 5.26fF $ **FLOATING
C2157 a_2467_n30310.t2 DGND 0.18fF
C2158 a_2467_n30310.t45 DGND 0.18fF
C2159 a_2467_n30310.n22 DGND 6.37fF $ **FLOATING
C2160 a_2467_n30310.n23 DGND 3.93fF $ **FLOATING
C2161 a_2467_n30310.n24 DGND 3.19fF $ **FLOATING
C2162 a_2467_n30310.t66 DGND 0.18fF
C2163 a_2467_n30310.t118 DGND 0.18fF
C2164 a_2467_n30310.t33 DGND 0.18fF
C2165 a_2467_n30310.t8 DGND 0.18fF
C2166 a_2467_n30310.n25 DGND 5.29fF $ **FLOATING
C2167 a_2467_n30310.n26 DGND 4.14fF $ **FLOATING
C2168 a_2467_n30310.n27 DGND 4.14fF $ **FLOATING
C2169 a_2467_n30310.n28 DGND 5.18fF $ **FLOATING
C2170 a_2467_n30310.n29 DGND 2.25fF $ **FLOATING
C2171 a_2467_n30310.t68 DGND 0.18fF
C2172 a_2467_n30310.t65 DGND 0.18fF
C2173 a_2467_n30310.n30 DGND 6.37fF $ **FLOATING
C2174 a_2467_n30310.n31 DGND 3.93fF $ **FLOATING
C2175 a_2467_n30310.n32 DGND 1.28fF $ **FLOATING
C2176 a_2467_n30310.t18 DGND 0.18fF
C2177 a_2467_n30310.t12 DGND 0.18fF
C2178 a_2467_n30310.n33 DGND 6.37fF $ **FLOATING
C2179 a_2467_n30310.n34 DGND 3.93fF $ **FLOATING
C2180 a_2467_n30310.n35 DGND 1.28fF $ **FLOATING
C2181 a_2467_n30310.t9 DGND 0.18fF
C2182 a_2467_n30310.t1 DGND 0.18fF
C2183 a_2467_n30310.t39 DGND 0.18fF
C2184 a_2467_n30310.t0 DGND 0.18fF
C2185 a_2467_n30310.n36 DGND 5.29fF $ **FLOATING
C2186 a_2467_n30310.n37 DGND 4.14fF $ **FLOATING
C2187 a_2467_n30310.n38 DGND 4.14fF $ **FLOATING
C2188 a_2467_n30310.n39 DGND 5.18fF $ **FLOATING
C2189 a_2467_n30310.n40 DGND 2.25fF $ **FLOATING
C2190 a_2467_n30310.t44 DGND 0.18fF
C2191 a_2467_n30310.t25 DGND 0.18fF
C2192 a_2467_n30310.n41 DGND 6.37fF $ **FLOATING
C2193 a_2467_n30310.n42 DGND 3.93fF $ **FLOATING
C2194 a_2467_n30310.n43 DGND 1.28fF $ **FLOATING
C2195 a_2467_n30310.n44 DGND 15.81fF $ **FLOATING
C2196 a_2467_n30310.n45 DGND 1.53fF $ **FLOATING
C2197 a_2467_n30310.n46 DGND 1.70fF $ **FLOATING
C2198 a_2467_n30310.n47 DGND 1.53fF $ **FLOATING
C2199 a_2467_n30310.n48 DGND 1.70fF $ **FLOATING
C2200 a_2467_n30310.n49 DGND 1.53fF $ **FLOATING
C2201 a_2467_n30310.n50 DGND 1.70fF $ **FLOATING
C2202 a_2467_n30310.n51 DGND 1.53fF $ **FLOATING
C2203 a_2467_n30310.n52 DGND 2.55fF $ **FLOATING
C2204 a_2467_n30310.n53 DGND 1.95fF $ **FLOATING
C2205 a_2467_n30310.n54 DGND 1.78fF $ **FLOATING
C2206 a_2467_n30310.n55 DGND 2.21fF $ **FLOATING
C2207 a_2467_n30310.n56 DGND 1.53fF $ **FLOATING
C2208 a_2467_n30310.n57 DGND 1.70fF $ **FLOATING
C2209 a_2467_n30310.n58 DGND 1.53fF $ **FLOATING
C2210 a_2467_n30310.n59 DGND 1.70fF $ **FLOATING
C2211 a_2467_n30310.n60 DGND 1.53fF $ **FLOATING
C2212 a_2467_n30310.n61 DGND 1.70fF $ **FLOATING
C2213 a_2467_n30310.n62 DGND 1.53fF $ **FLOATING
C2214 a_2467_n30310.n63 DGND 2.55fF $ **FLOATING
C2215 a_2467_n30310.n64 DGND 1.95fF $ **FLOATING
C2216 a_2467_n30310.n65 DGND 1.78fF $ **FLOATING
C2217 a_2467_n30310.n66 DGND 2.21fF $ **FLOATING
C2218 a_2467_n30310.t7 DGND 0.18fF
C2219 a_2467_n30310.t21 DGND 0.18fF
C2220 a_2467_n30310.n67 DGND 6.37fF $ **FLOATING
C2221 a_2467_n30310.n68 DGND 4.06fF $ **FLOATING
C2222 a_2467_n30310.t110 DGND 0.18fF
C2223 a_2467_n30310.t26 DGND 0.18fF
C2224 a_2467_n30310.n69 DGND 6.37fF $ **FLOATING
C2225 a_2467_n30310.n70 DGND 4.06fF $ **FLOATING
C2226 a_2467_n30310.t17 DGND 0.18fF
C2227 a_2467_n30310.t119 DGND 0.18fF
C2228 a_2467_n30310.n71 DGND 6.37fF $ **FLOATING
C2229 a_2467_n30310.n72 DGND 4.06fF $ **FLOATING
C2230 a_2467_n30310.t67 DGND 0.18fF
C2231 a_2467_n30310.t32 DGND 0.18fF
C2232 a_2467_n30310.n73 DGND 6.37fF $ **FLOATING
C2233 a_2467_n30310.n74 DGND 4.06fF $ **FLOATING
C2234 a_2467_n30310.n75 DGND 3.66fF $ **FLOATING
C2235 a_2467_n30310.n76 DGND 2.50fF $ **FLOATING
C2236 a_2467_n30310.n77 DGND 1.51fF $ **FLOATING
C2237 a_2467_n30310.n78 DGND 1.51fF $ **FLOATING
C2238 a_2467_n30310.n79 DGND 2.50fF $ **FLOATING
C2239 a_2467_n30310.n80 DGND 1.51fF $ **FLOATING
C2240 a_2467_n30310.n81 DGND 29.37fF $ **FLOATING
C2241 a_2467_n30310.n82 DGND 31.13fF $ **FLOATING
C2242 a_2467_n30310.n83 DGND 3.95fF $ **FLOATING
C2243 a_2467_n30310.n84 DGND 16.81fF $ **FLOATING
C2244 a_2467_n30310.n85 DGND 6.18fF $ **FLOATING
C2245 a_2467_n30310.n86 DGND 1.53fF $ **FLOATING
C2246 a_2467_n30310.n87 DGND 1.70fF $ **FLOATING
C2247 a_2467_n30310.n88 DGND 1.53fF $ **FLOATING
C2248 a_2467_n30310.n89 DGND 2.64fF $ **FLOATING
C2249 a_2467_n30310.n90 DGND 2.40fF $ **FLOATING
C2250 a_2467_n30310.t60 DGND 0.25fF
C2251 a_2467_n30310.n91 DGND 0.65fF $ **FLOATING
C2252 a_2467_n30310.n92 DGND 0.65fF $ **FLOATING
C2253 a_2467_n30310.n93 DGND 0.65fF $ **FLOATING
C2254 a_2467_n30310.t117 DGND 0.32fF
C2255 a_2467_n30310.n94 DGND 1.37fF $ **FLOATING
C2256 a_2467_n30310.n95 DGND 0.48fF $ **FLOATING
C2257 a_2467_n30310.n96 DGND 0.48fF $ **FLOATING
C2258 a_2467_n30310.n97 DGND 12.07fF $ **FLOATING
C2259 a_2467_n30310.n98 DGND 22.39fF $ **FLOATING
C2260 a_2467_n30310.n99 DGND 6.30fF $ **FLOATING
C2261 a_2467_n30310.n100 DGND 2.21fF $ **FLOATING
C2262 a_2467_n30310.n101 DGND 1.51fF $ **FLOATING
C2263 a_2467_n30310.n102 DGND 1.54fF $ **FLOATING
C2264 a_2467_n30310.n103 DGND 1.53fF $ **FLOATING
C2265 a_2467_n30310.n104 DGND 1.70fF $ **FLOATING
C2266 a_2467_n30310.n105 DGND 1.51fF $ **FLOATING
C2267 a_2467_n30310.n106 DGND 1.54fF $ **FLOATING
C2268 a_2467_n30310.n107 DGND 1.53fF $ **FLOATING
C2269 a_2467_n30310.n108 DGND 1.70fF $ **FLOATING
C2270 a_2467_n30310.n109 DGND 1.15fF $ **FLOATING
C2271 a_2467_n30310.n110 DGND 1.91fF $ **FLOATING
C2272 a_2467_n30310.n111 DGND 1.77fF $ **FLOATING
C2273 a_2467_n30310.n112 DGND 1.70fF $ **FLOATING
C2274 bias_p.n0 DGND 2.83fF $ **FLOATING
C2275 bias_p.n1 DGND 2.61fF $ **FLOATING
C2276 bias_p.n2 DGND 2.61fF $ **FLOATING
C2277 bias_p.n3 DGND 2.61fF $ **FLOATING
C2278 bias_p.n4 DGND 2.61fF $ **FLOATING
C2279 bias_p.n5 DGND 2.61fF $ **FLOATING
C2280 bias_p.n6 DGND 2.61fF $ **FLOATING
C2281 bias_p.n7 DGND 2.09fF $ **FLOATING
C2282 bias_p.n8 DGND 2.26fF $ **FLOATING
C2283 bias_p.n9 DGND 2.26fF $ **FLOATING
C2284 bias_p.n10 DGND 2.26fF $ **FLOATING
C2285 bias_p.n11 DGND 2.26fF $ **FLOATING
C2286 bias_p.n12 DGND 2.26fF $ **FLOATING
C2287 bias_p.n13 DGND 2.26fF $ **FLOATING
C2288 bias_p.n14 DGND 2.26fF $ **FLOATING
C2289 bias_p.n15 DGND 2.09fF $ **FLOATING
C2290 bias_p.n16 DGND 2.26fF $ **FLOATING
C2291 bias_p.n17 DGND 2.26fF $ **FLOATING
C2292 bias_p.n18 DGND 2.26fF $ **FLOATING
C2293 bias_p.n19 DGND 2.26fF $ **FLOATING
C2294 bias_p.n20 DGND 2.26fF $ **FLOATING
C2295 bias_p.n21 DGND 2.26fF $ **FLOATING
C2296 bias_p.n22 DGND 2.26fF $ **FLOATING
C2297 bias_p.n23 DGND 2.09fF $ **FLOATING
C2298 bias_p.n24 DGND 2.26fF $ **FLOATING
C2299 bias_p.n25 DGND 2.26fF $ **FLOATING
C2300 bias_p.n26 DGND 2.26fF $ **FLOATING
C2301 bias_p.n27 DGND 2.26fF $ **FLOATING
C2302 bias_p.n28 DGND 2.26fF $ **FLOATING
C2303 bias_p.n29 DGND 2.26fF $ **FLOATING
C2304 bias_p.n30 DGND 2.09fF $ **FLOATING
C2305 bias_p.n31 DGND 2.32fF $ **FLOATING
C2306 bias_p.n32 DGND 2.09fF $ **FLOATING
C2307 bias_p.n33 DGND 2.32fF $ **FLOATING
C2308 bias_p.n34 DGND 2.09fF $ **FLOATING
C2309 bias_p.n35 DGND 2.32fF $ **FLOATING
C2310 bias_p.n36 DGND 2.71fF $ **FLOATING
C2311 bias_p.n37 DGND 2.30fF $ **FLOATING
C2312 bias_p.n38 DGND 2.45fF $ **FLOATING
C2313 bias_p.n39 DGND 3.16fF $ **FLOATING
C2314 bias_p.t1 DGND 5.88fF
C2315 bias_p.t65 DGND 1.69fF
C2316 bias_p.t24 DGND 1.69fF
C2317 bias_p.t18 DGND 1.69fF
C2318 bias_p.t70 DGND 1.69fF
C2319 bias_p.n41 DGND 0.12fF $ **FLOATING
C2320 bias_p.n42 DGND 0.12fF $ **FLOATING
C2321 bias_p.n43 DGND 0.11fF $ **FLOATING
C2322 bias_p.n44 DGND 2.65fF $ **FLOATING
C2323 bias_p.t89 DGND 1.69fF
C2324 bias_p.t42 DGND 1.69fF
C2325 bias_p.n46 DGND 0.12fF $ **FLOATING
C2326 bias_p.n47 DGND 0.12fF $ **FLOATING
C2327 bias_p.n48 DGND 0.12fF $ **FLOATING
C2328 bias_p.n49 DGND 0.29fF $ **FLOATING
C2329 bias_p.t37 DGND 1.69fF
C2330 bias_p.t44 DGND 1.69fF
C2331 bias_p.n51 DGND 0.12fF $ **FLOATING
C2332 bias_p.n52 DGND 0.12fF $ **FLOATING
C2333 bias_p.n53 DGND 0.12fF $ **FLOATING
C2334 bias_p.t41 DGND 1.69fF
C2335 bias_p.t91 DGND 1.69fF
C2336 bias_p.n55 DGND 0.12fF $ **FLOATING
C2337 bias_p.n56 DGND 0.12fF $ **FLOATING
C2338 bias_p.n57 DGND 0.12fF $ **FLOATING
C2339 bias_p.t87 DGND 1.69fF
C2340 bias_p.t40 DGND 1.69fF
C2341 bias_p.n59 DGND 0.12fF $ **FLOATING
C2342 bias_p.n60 DGND 0.12fF $ **FLOATING
C2343 bias_p.n61 DGND 0.12fF $ **FLOATING
C2344 bias_p.t90 DGND 1.69fF
C2345 bias_p.t96 DGND 1.69fF
C2346 bias_p.n63 DGND 0.12fF $ **FLOATING
C2347 bias_p.n64 DGND 0.12fF $ **FLOATING
C2348 bias_p.n65 DGND 0.12fF $ **FLOATING
C2349 bias_p.t39 DGND 1.69fF
C2350 bias_p.t47 DGND 1.69fF
C2351 bias_p.n67 DGND 0.12fF $ **FLOATING
C2352 bias_p.n68 DGND 0.12fF $ **FLOATING
C2353 bias_p.n69 DGND 0.12fF $ **FLOATING
C2354 bias_p.t94 DGND 1.69fF
C2355 bias_p.t49 DGND 1.69fF
C2356 bias_p.n71 DGND 0.12fF $ **FLOATING
C2357 bias_p.n72 DGND 0.12fF $ **FLOATING
C2358 bias_p.n73 DGND 0.12fF $ **FLOATING
C2359 bias_p.t43 DGND 1.69fF
C2360 bias_p.t93 DGND 1.69fF
C2361 bias_p.n75 DGND 0.12fF $ **FLOATING
C2362 bias_p.n76 DGND 0.12fF $ **FLOATING
C2363 bias_p.n77 DGND 0.12fF $ **FLOATING
C2364 bias_p.n78 DGND 1.26fF $ **FLOATING
C2365 bias_p.n79 DGND 1.84fF $ **FLOATING
C2366 bias_p.n80 DGND 1.84fF $ **FLOATING
C2367 bias_p.t84 DGND 1.69fF
C2368 bias_p.t88 DGND 1.69fF
C2369 bias_p.n82 DGND 0.12fF $ **FLOATING
C2370 bias_p.n83 DGND 0.12fF $ **FLOATING
C2371 bias_p.n84 DGND 0.12fF $ **FLOATING
C2372 bias_p.t71 DGND 1.69fF
C2373 bias_p.t86 DGND 1.69fF
C2374 bias_p.n86 DGND 0.12fF $ **FLOATING
C2375 bias_p.n87 DGND 0.12fF $ **FLOATING
C2376 bias_p.n88 DGND 0.12fF $ **FLOATING
C2377 bias_p.t15 DGND 1.69fF
C2378 bias_p.t32 DGND 1.69fF
C2379 bias_p.n90 DGND 0.12fF $ **FLOATING
C2380 bias_p.n91 DGND 0.12fF $ **FLOATING
C2381 bias_p.n92 DGND 0.12fF $ **FLOATING
C2382 bias_p.t59 DGND 1.69fF
C2383 bias_p.t73 DGND 1.69fF
C2384 bias_p.n94 DGND 0.12fF $ **FLOATING
C2385 bias_p.n95 DGND 0.12fF $ **FLOATING
C2386 bias_p.n96 DGND 0.12fF $ **FLOATING
C2387 bias_p.t36 DGND 1.69fF
C2388 bias_p.t79 DGND 1.69fF
C2389 bias_p.t82 DGND 1.69fF
C2390 bias_p.t30 DGND 1.69fF
C2391 bias_p.n97 DGND 2.63fF $ **FLOATING
C2392 bias_p.n98 DGND 1.32fF $ **FLOATING
C2393 bias_p.t83 DGND 1.69fF
C2394 bias_p.t67 DGND 1.69fF
C2395 bias_p.t35 DGND 1.69fF
C2396 bias_p.t19 DGND 1.69fF
C2397 bias_p.n99 DGND 2.63fF $ **FLOATING
C2398 bias_p.n100 DGND 1.90fF $ **FLOATING
C2399 bias_p.t74 DGND 1.69fF
C2400 bias_p.t21 DGND 1.69fF
C2401 bias_p.t26 DGND 1.69fF
C2402 bias_p.t66 DGND 1.69fF
C2403 bias_p.n101 DGND 2.63fF $ **FLOATING
C2404 bias_p.n102 DGND 1.90fF $ **FLOATING
C2405 bias_p.t12 DGND 1.69fF
C2406 bias_p.t27 DGND 1.69fF
C2407 bias_p.n104 DGND 0.12fF $ **FLOATING
C2408 bias_p.n105 DGND 0.12fF $ **FLOATING
C2409 bias_p.n106 DGND 0.12fF $ **FLOATING
C2410 bias_p.t17 DGND 1.69fF
C2411 bias_p.t62 DGND 1.69fF
C2412 bias_p.t28 DGND 1.69fF
C2413 bias_p.t14 DGND 1.69fF
C2414 bias_p.t77 DGND 1.69fF
C2415 bias_p.t25 DGND 1.69fF
C2416 bias_p.n107 DGND 1.25fF $ **FLOATING
C2417 bias_p.n108 DGND 1.84fF $ **FLOATING
C2418 bias_p.n109 DGND 1.84fF $ **FLOATING
C2419 bias_p.t56 DGND 1.69fF
C2420 bias_p.t64 DGND 1.69fF
C2421 bias_p.n111 DGND 0.12fF $ **FLOATING
C2422 bias_p.n112 DGND 0.12fF $ **FLOATING
C2423 bias_p.n113 DGND 0.12fF $ **FLOATING
C2424 bias_p.t50 DGND 1.69fF
C2425 bias_p.t20 DGND 1.69fF
C2426 bias_p.n114 DGND 2.37fF $ **FLOATING
C2427 bias_p.n115 DGND 1.32fF $ **FLOATING
C2428 bias_p.t22 DGND 1.69fF
C2429 bias_p.t80 DGND 1.69fF
C2430 bias_p.n116 DGND 2.37fF $ **FLOATING
C2431 bias_p.n117 DGND 1.90fF $ **FLOATING
C2432 bias_p.t81 DGND 1.69fF
C2433 bias_p.t45 DGND 1.69fF
C2434 bias_p.n118 DGND 2.37fF $ **FLOATING
C2435 bias_p.n119 DGND 1.90fF $ **FLOATING
C2436 bias_p.t97 DGND 1.69fF
C2437 bias_p.t46 DGND 1.69fF
C2438 bias_p.n121 DGND 0.12fF $ **FLOATING
C2439 bias_p.n122 DGND 0.12fF $ **FLOATING
C2440 bias_p.n123 DGND 0.12fF $ **FLOATING
C2441 bias_p.n124 DGND 1.84fF $ **FLOATING
C2442 bias_p.n125 DGND 1.84fF $ **FLOATING
C2443 bias_p.n126 DGND 1.84fF $ **FLOATING
C2444 bias_p.n127 DGND 1.25fF $ **FLOATING
C2445 bias_p.n128 DGND 1.25fF $ **FLOATING
C2446 bias_p.n129 DGND 1.25fF $ **FLOATING
C2447 bias_p.n130 DGND 1.84fF $ **FLOATING
C2448 bias_p.t29 DGND 1.69fF
C2449 bias_p.t38 DGND 1.69fF
C2450 bias_p.n132 DGND 0.12fF $ **FLOATING
C2451 bias_p.n133 DGND 0.12fF $ **FLOATING
C2452 bias_p.n134 DGND 0.12fF $ **FLOATING
C2453 bias_p.t69 DGND 1.69fF
C2454 bias_p.t85 DGND 1.69fF
C2455 bias_p.n136 DGND 0.12fF $ **FLOATING
C2456 bias_p.n137 DGND 0.12fF $ **FLOATING
C2457 bias_p.n138 DGND 0.12fF $ **FLOATING
C2458 bias_p.t58 DGND 1.69fF
C2459 bias_p.t72 DGND 1.69fF
C2460 bias_p.n140 DGND 0.12fF $ **FLOATING
C2461 bias_p.n141 DGND 0.12fF $ **FLOATING
C2462 bias_p.n142 DGND 0.12fF $ **FLOATING
C2463 bias_p.t101 DGND 1.69fF
C2464 bias_p.t16 DGND 1.69fF
C2465 bias_p.n144 DGND 0.12fF $ **FLOATING
C2466 bias_p.n145 DGND 0.12fF $ **FLOATING
C2467 bias_p.n146 DGND 0.12fF $ **FLOATING
C2468 bias_p.t52 DGND 1.69fF
C2469 bias_p.t60 DGND 1.69fF
C2470 bias_p.n148 DGND 0.12fF $ **FLOATING
C2471 bias_p.n149 DGND 0.12fF $ **FLOATING
C2472 bias_p.n150 DGND 0.12fF $ **FLOATING
C2473 bias_p.t99 DGND 1.69fF
C2474 bias_p.t13 DGND 1.69fF
C2475 bias_p.n152 DGND 0.12fF $ **FLOATING
C2476 bias_p.n153 DGND 0.12fF $ **FLOATING
C2477 bias_p.n154 DGND 0.12fF $ **FLOATING
C2478 bias_p.t48 DGND 1.69fF
C2479 bias_p.t57 DGND 1.69fF
C2480 bias_p.n156 DGND 0.12fF $ **FLOATING
C2481 bias_p.n157 DGND 0.12fF $ **FLOATING
C2482 bias_p.n158 DGND 0.12fF $ **FLOATING
C2483 bias_p.t31 DGND 1.69fF
C2484 bias_p.t68 DGND 1.69fF
C2485 bias_p.n160 DGND 0.12fF $ **FLOATING
C2486 bias_p.n161 DGND 0.12fF $ **FLOATING
C2487 bias_p.n162 DGND 0.12fF $ **FLOATING
C2488 bias_p.n163 DGND 1.84fF $ **FLOATING
C2489 bias_p.n164 DGND 1.84fF $ **FLOATING
C2490 bias_p.n165 DGND 1.84fF $ **FLOATING
C2491 bias_p.n166 DGND 1.84fF $ **FLOATING
C2492 bias_p.n167 DGND 1.84fF $ **FLOATING
C2493 bias_p.n168 DGND 1.84fF $ **FLOATING
C2494 bias_p.n169 DGND 1.84fF $ **FLOATING
C2495 bias_p.n170 DGND 1.79fF $ **FLOATING
C2496 bias_p.n171 DGND 0.47fF $ **FLOATING
C2497 bias_p.n172 DGND 1.04fF $ **FLOATING
C2498 bias_p.t78 DGND 1.69fF
C2499 bias_p.t34 DGND 1.69fF
C2500 bias_p.n174 DGND 0.12fF $ **FLOATING
C2501 bias_p.n175 DGND 0.12fF $ **FLOATING
C2502 bias_p.n176 DGND 0.12fF $ **FLOATING
C2503 bias_p.t23 DGND 1.69fF
C2504 bias_p.t75 DGND 1.69fF
C2505 bias_p.n178 DGND 0.12fF $ **FLOATING
C2506 bias_p.n179 DGND 0.12fF $ **FLOATING
C2507 bias_p.n180 DGND 0.12fF $ **FLOATING
C2508 bias_p.t11 DGND 1.69fF
C2509 bias_p.t63 DGND 1.69fF
C2510 bias_p.n182 DGND 0.12fF $ **FLOATING
C2511 bias_p.n183 DGND 0.12fF $ **FLOATING
C2512 bias_p.n184 DGND 0.12fF $ **FLOATING
C2513 bias_p.t55 DGND 1.69fF
C2514 bias_p.t102 DGND 1.69fF
C2515 bias_p.n186 DGND 0.12fF $ **FLOATING
C2516 bias_p.n187 DGND 0.12fF $ **FLOATING
C2517 bias_p.n188 DGND 0.12fF $ **FLOATING
C2518 bias_p.t98 DGND 1.69fF
C2519 bias_p.t54 DGND 1.69fF
C2520 bias_p.n190 DGND 0.12fF $ **FLOATING
C2521 bias_p.n191 DGND 0.12fF $ **FLOATING
C2522 bias_p.n192 DGND 0.12fF $ **FLOATING
C2523 bias_p.t53 DGND 1.69fF
C2524 bias_p.t100 DGND 1.69fF
C2525 bias_p.n194 DGND 0.12fF $ **FLOATING
C2526 bias_p.n195 DGND 0.12fF $ **FLOATING
C2527 bias_p.n196 DGND 0.12fF $ **FLOATING
C2528 bias_p.t95 DGND 1.69fF
C2529 bias_p.t51 DGND 1.69fF
C2530 bias_p.n198 DGND 0.12fF $ **FLOATING
C2531 bias_p.n199 DGND 0.12fF $ **FLOATING
C2532 bias_p.n200 DGND 0.12fF $ **FLOATING
C2533 bias_p.t92 DGND 1.69fF
C2534 bias_p.t33 DGND 1.69fF
C2535 bias_p.n202 DGND 0.12fF $ **FLOATING
C2536 bias_p.n203 DGND 0.12fF $ **FLOATING
C2537 bias_p.n204 DGND 0.12fF $ **FLOATING
C2538 bias_p.n205 DGND 1.25fF $ **FLOATING
C2539 bias_p.n206 DGND 1.25fF $ **FLOATING
C2540 bias_p.n207 DGND 1.25fF $ **FLOATING
C2541 bias_p.n208 DGND 1.25fF $ **FLOATING
C2542 bias_p.n209 DGND 1.25fF $ **FLOATING
C2543 bias_p.n210 DGND 1.25fF $ **FLOATING
C2544 bias_p.n211 DGND 1.25fF $ **FLOATING
C2545 bias_p.n212 DGND 1.03fF $ **FLOATING
C2546 bias_p.n213 DGND 5.00fF $ **FLOATING
C2547 bias_p.n214 DGND 8.22fF $ **FLOATING
C2548 bias_p.n215 DGND 4.81fF $ **FLOATING
C2549 bias_p.n216 DGND 0.32fF $ **FLOATING
C2550 a_23013_n25097.n0 DGND 1.45fF $ **FLOATING
C2551 a_23013_n25097.n1 DGND 0.85fF $ **FLOATING
C2552 a_23013_n25097.n2 DGND 0.85fF $ **FLOATING
C2553 a_23013_n25097.n3 DGND 0.85fF $ **FLOATING
C2554 a_23013_n25097.n4 DGND 0.71fF $ **FLOATING
C2555 a_23013_n25097.n5 DGND 1.45fF $ **FLOATING
C2556 a_23013_n25097.n6 DGND 0.85fF $ **FLOATING
C2557 a_23013_n25097.n7 DGND 0.85fF $ **FLOATING
C2558 a_23013_n25097.n8 DGND 0.85fF $ **FLOATING
C2559 a_23013_n25097.n9 DGND 1.53fF $ **FLOATING
C2560 a_23013_n25097.n10 DGND 5.81fF $ **FLOATING
C2561 a_23013_n25097.n11 DGND 0.66fF $ **FLOATING
C2562 a_23013_n25097.n12 DGND 0.66fF $ **FLOATING
C2563 a_23013_n25097.t21 DGND 0.36fF
C2564 a_23013_n25097.n13 DGND 0.66fF $ **FLOATING
C2565 a_23013_n25097.t1 DGND 0.36fF
C2566 a_23013_n25097.t6 DGND 0.36fF
C2567 a_23013_n25097.n14 DGND 0.66fF $ **FLOATING
C2568 a_23013_n25097.t7 DGND 0.42fF
C2569 a_23013_n25097.n15 DGND 0.96fF $ **FLOATING
C2570 a_23013_n25097.n16 DGND 0.82fF $ **FLOATING
C2571 a_23013_n25097.n17 DGND 0.82fF $ **FLOATING
C2572 a_23013_n25097.n18 DGND 0.33fF $ **FLOATING
C2573 a_23013_n25097.n19 DGND 1.32fF $ **FLOATING
C2574 a_23013_n25097.n20 DGND 0.85fF $ **FLOATING
C2575 a_23013_n25097.n21 DGND 1.42fF $ **FLOATING
C2576 a_23013_n25097.t22 DGND 21.68fF
C2577 a_33657_n21342.n0 DGND 0.51fF $ **FLOATING
C2578 a_33657_n21342.n1 DGND 0.51fF $ **FLOATING
C2579 a_33657_n21342.n2 DGND 0.59fF $ **FLOATING
C2580 a_33657_n21342.n3 DGND 0.59fF $ **FLOATING
C2581 level_shifter_up_8.x_hv.n0 DGND 1.96fF $ **FLOATING
C2582 level_shifter_up_8.x_hv.n1 DGND 0.61fF $ **FLOATING
C2583 level_shifter_up_8.x_hv.n2 DGND 3.37fF $ **FLOATING
C2584 level_shifter_up_8.x_hv.n3 DGND 5.38fF $ **FLOATING
C2585 level_shifter_up_8.x_hv.t8 DGND 0.25fF
C2586 level_shifter_up_8.x_hv.t9 DGND 0.54fF
C2587 level_shifter_up_8.x_hv.t1 DGND 0.54fF
C2588 level_shifter_up_8.x_hv.t6 DGND 0.54fF
C2589 level_shifter_up_8.x_hv.t7 DGND 0.54fF
C2590 level_shifter_up_8.x_hv.t4 DGND 0.54fF
C2591 level_shifter_up_8.x_hv.t5 DGND 0.54fF
C2592 level_shifter_up_8.x_hv.t2 DGND 0.54fF
C2593 level_shifter_up_8.x_hv.t3 DGND 0.54fF
C2594 Vxp.t146 DGND 0.30fF
C2595 Vxp.t2 DGND 0.30fF
C2596 Vxp.t28 DGND 0.30fF
C2597 Vxp.n0 DGND 7.33fF $ **FLOATING
C2598 Vxp.n1 DGND 7.33fF $ **FLOATING
C2599 Vxp.n2 DGND 7.06fF $ **FLOATING
C2600 Vxp.t36 DGND 0.30fF
C2601 Vxp.t25 DGND 0.30fF
C2602 Vxp.t22 DGND 0.30fF
C2603 Vxp.n3 DGND 7.33fF $ **FLOATING
C2604 Vxp.n4 DGND 7.33fF $ **FLOATING
C2605 Vxp.n5 DGND 7.06fF $ **FLOATING
C2606 Vxp.t149 DGND 0.30fF
C2607 Vxp.t13 DGND 0.30fF
C2608 Vxp.n6 DGND 7.33fF $ **FLOATING
C2609 Vxp.n7 DGND 7.98fF $ **FLOATING
C2610 Vxp.t16 DGND 0.30fF
C2611 Vxp.t18 DGND 0.30fF
C2612 Vxp.n8 DGND 7.33fF $ **FLOATING
C2613 Vxp.n9 DGND 7.98fF $ **FLOATING
C2614 Vxp.t40 DGND 0.30fF
C2615 Vxp.t6 DGND 0.30fF
C2616 Vxp.n10 DGND 7.33fF $ **FLOATING
C2617 Vxp.n11 DGND 7.98fF $ **FLOATING
C2618 Vxp.t138 DGND 0.30fF
C2619 Vxp.t139 DGND 0.30fF
C2620 Vxp.n12 DGND 7.33fF $ **FLOATING
C2621 Vxp.n13 DGND 7.98fF $ **FLOATING
C2622 Vxp.t7 DGND 0.30fF
C2623 Vxp.t20 DGND 0.30fF
C2624 Vxp.t34 DGND 0.30fF
C2625 Vxp.n14 DGND 7.33fF $ **FLOATING
C2626 Vxp.n15 DGND 7.33fF $ **FLOATING
C2627 Vxp.n16 DGND 7.68fF $ **FLOATING
C2628 Vxp.t5 DGND 0.30fF
C2629 Vxp.t37 DGND 0.30fF
C2630 Vxp.t21 DGND 0.30fF
C2631 Vxp.n17 DGND 7.33fF $ **FLOATING
C2632 Vxp.n18 DGND 7.33fF $ **FLOATING
C2633 Vxp.n19 DGND 7.06fF $ **FLOATING
C2634 Vxp.n20 DGND 5.91fF $ **FLOATING
C2635 Vxp.n21 DGND 3.59fF $ **FLOATING
C2636 Vxp.n22 DGND 3.59fF $ **FLOATING
C2637 Vxp.n23 DGND 3.59fF $ **FLOATING
C2638 Vxp.n24 DGND 3.59fF $ **FLOATING
C2639 Vxp.n25 DGND 2.82fF $ **FLOATING
C2640 Vxp.n26 DGND 18.43fF $ **FLOATING
C2641 Vxp.t42 DGND 0.13fF
C2642 Vxp.n27 DGND 2.49fF $ **FLOATING
C2643 Vxp.n28 DGND 1.19fF $ **FLOATING
C2644 Vxp.n29 DGND 2.00fF $ **FLOATING
C2645 Vxp.t87 DGND 0.13fF
C2646 Vxp.n30 DGND 2.49fF $ **FLOATING
C2647 Vxp.n31 DGND 1.19fF $ **FLOATING
C2648 Vxp.n32 DGND 3.08fF $ **FLOATING
C2649 Vxp.t132 DGND 0.13fF
C2650 Vxp.n33 DGND 2.49fF $ **FLOATING
C2651 Vxp.n34 DGND 1.19fF $ **FLOATING
C2652 Vxp.n35 DGND 3.08fF $ **FLOATING
C2653 Vxp.t85 DGND 0.13fF
C2654 Vxp.n36 DGND 2.49fF $ **FLOATING
C2655 Vxp.n37 DGND 1.19fF $ **FLOATING
C2656 Vxp.n38 DGND 3.08fF $ **FLOATING
C2657 Vxp.t128 DGND 0.13fF
C2658 Vxp.n39 DGND 2.49fF $ **FLOATING
C2659 Vxp.n40 DGND 1.19fF $ **FLOATING
C2660 Vxp.n41 DGND 3.08fF $ **FLOATING
C2661 Vxp.t75 DGND 0.13fF
C2662 Vxp.n42 DGND 2.49fF $ **FLOATING
C2663 Vxp.n43 DGND 1.19fF $ **FLOATING
C2664 Vxp.n44 DGND 3.08fF $ **FLOATING
C2665 Vxp.t116 DGND 0.13fF
C2666 Vxp.n45 DGND 2.49fF $ **FLOATING
C2667 Vxp.n46 DGND 1.19fF $ **FLOATING
C2668 Vxp.n47 DGND 3.08fF $ **FLOATING
C2669 Vxp.t105 DGND 0.13fF
C2670 Vxp.n48 DGND 2.49fF $ **FLOATING
C2671 Vxp.n49 DGND 1.19fF $ **FLOATING
C2672 Vxp.n50 DGND 3.60fF $ **FLOATING
C2673 Vxp.n51 DGND 20.33fF $ **FLOATING
C2674 Vxp.n52 DGND 1.19fF $ **FLOATING
C2675 Vxp.n53 DGND 1.34fF $ **FLOATING
C2676 Vxp.n54 DGND 1.34fF $ **FLOATING
C2677 Vxp.n55 DGND 1.19fF $ **FLOATING
C2678 Vxp.n56 DGND 2.00fF $ **FLOATING
C2679 Vxp.n57 DGND 3.08fF $ **FLOATING
C2680 Vxp.n58 DGND 1.34fF $ **FLOATING
C2681 Vxp.n59 DGND 1.19fF $ **FLOATING
C2682 Vxp.n60 DGND 3.08fF $ **FLOATING
C2683 Vxp.n61 DGND 1.34fF $ **FLOATING
C2684 Vxp.n62 DGND 1.19fF $ **FLOATING
C2685 Vxp.n63 DGND 3.08fF $ **FLOATING
C2686 Vxp.n64 DGND 1.34fF $ **FLOATING
C2687 Vxp.n65 DGND 1.19fF $ **FLOATING
C2688 Vxp.n66 DGND 3.08fF $ **FLOATING
C2689 Vxp.n67 DGND 1.34fF $ **FLOATING
C2690 Vxp.n68 DGND 1.19fF $ **FLOATING
C2691 Vxp.n69 DGND 3.08fF $ **FLOATING
C2692 Vxp.n70 DGND 1.34fF $ **FLOATING
C2693 Vxp.n71 DGND 1.19fF $ **FLOATING
C2694 Vxp.n72 DGND 3.08fF $ **FLOATING
C2695 Vxp.n73 DGND 1.34fF $ **FLOATING
C2696 Vxp.n74 DGND 1.19fF $ **FLOATING
C2697 Vxp.n75 DGND 3.60fF $ **FLOATING
C2698 Vxp.n76 DGND 6.13fF $ **FLOATING
C2699 Vxp.n77 DGND 1.19fF $ **FLOATING
C2700 Vxp.n78 DGND 1.34fF $ **FLOATING
C2701 Vxp.n79 DGND 1.34fF $ **FLOATING
C2702 Vxp.n80 DGND 1.19fF $ **FLOATING
C2703 Vxp.n81 DGND 2.00fF $ **FLOATING
C2704 Vxp.n82 DGND 1.34fF $ **FLOATING
C2705 Vxp.n83 DGND 1.19fF $ **FLOATING
C2706 Vxp.n84 DGND 3.08fF $ **FLOATING
C2707 Vxp.n85 DGND 1.34fF $ **FLOATING
C2708 Vxp.n86 DGND 1.19fF $ **FLOATING
C2709 Vxp.n87 DGND 3.08fF $ **FLOATING
C2710 Vxp.n88 DGND 1.34fF $ **FLOATING
C2711 Vxp.n89 DGND 1.19fF $ **FLOATING
C2712 Vxp.n90 DGND 3.08fF $ **FLOATING
C2713 Vxp.n91 DGND 1.34fF $ **FLOATING
C2714 Vxp.n92 DGND 1.19fF $ **FLOATING
C2715 Vxp.n93 DGND 3.08fF $ **FLOATING
C2716 Vxp.n94 DGND 1.34fF $ **FLOATING
C2717 Vxp.n95 DGND 1.19fF $ **FLOATING
C2718 Vxp.n96 DGND 3.08fF $ **FLOATING
C2719 Vxp.n97 DGND 1.34fF $ **FLOATING
C2720 Vxp.n98 DGND 1.19fF $ **FLOATING
C2721 Vxp.n99 DGND 3.08fF $ **FLOATING
C2722 Vxp.n100 DGND 3.60fF $ **FLOATING
C2723 Vxp.n101 DGND 5.15fF $ **FLOATING
C2724 Vxp.t140 DGND 0.30fF
C2725 Vxp.t29 DGND 0.30fF
C2726 Vxp.t23 DGND 0.30fF
C2727 Vxp.t12 DGND 0.30fF
C2728 Vxp.t24 DGND 0.30fF
C2729 Vxp.n102 DGND 7.33fF $ **FLOATING
C2730 Vxp.n103 DGND 7.33fF $ **FLOATING
C2731 Vxp.n104 DGND 7.33fF $ **FLOATING
C2732 Vxp.n105 DGND 7.33fF $ **FLOATING
C2733 Vxp.n106 DGND 7.06fF $ **FLOATING
C2734 Vxp.t148 DGND 0.30fF
C2735 Vxp.t0 DGND 0.30fF
C2736 Vxp.t14 DGND 0.30fF
C2737 Vxp.t27 DGND 0.30fF
C2738 Vxp.t15 DGND 0.30fF
C2739 Vxp.n107 DGND 7.33fF $ **FLOATING
C2740 Vxp.n108 DGND 7.33fF $ **FLOATING
C2741 Vxp.n109 DGND 7.33fF $ **FLOATING
C2742 Vxp.n110 DGND 7.33fF $ **FLOATING
C2743 Vxp.n111 DGND 7.68fF $ **FLOATING
C2744 Vxp.n112 DGND 5.91fF $ **FLOATING
C2745 Vxp.t32 DGND 0.30fF
C2746 Vxp.t11 DGND 0.30fF
C2747 Vxp.t30 DGND 0.30fF
C2748 Vxp.t150 DGND 0.30fF
C2749 Vxp.n113 DGND 7.33fF $ **FLOATING
C2750 Vxp.n114 DGND 7.33fF $ **FLOATING
C2751 Vxp.n115 DGND 7.33fF $ **FLOATING
C2752 Vxp.n116 DGND 7.98fF $ **FLOATING
C2753 Vxp.n117 DGND 3.59fF $ **FLOATING
C2754 Vxp.t151 DGND 0.30fF
C2755 Vxp.t142 DGND 0.30fF
C2756 Vxp.t17 DGND 0.30fF
C2757 Vxp.t143 DGND 0.30fF
C2758 Vxp.n118 DGND 7.33fF $ **FLOATING
C2759 Vxp.n119 DGND 7.33fF $ **FLOATING
C2760 Vxp.n120 DGND 7.33fF $ **FLOATING
C2761 Vxp.n121 DGND 7.98fF $ **FLOATING
C2762 Vxp.n122 DGND 3.59fF $ **FLOATING
C2763 Vxp.t26 DGND 0.30fF
C2764 Vxp.t8 DGND 0.30fF
C2765 Vxp.t31 DGND 0.30fF
C2766 Vxp.t1 DGND 0.30fF
C2767 Vxp.n123 DGND 7.33fF $ **FLOATING
C2768 Vxp.n124 DGND 7.33fF $ **FLOATING
C2769 Vxp.n125 DGND 7.33fF $ **FLOATING
C2770 Vxp.n126 DGND 7.98fF $ **FLOATING
C2771 Vxp.n127 DGND 3.59fF $ **FLOATING
C2772 Vxp.t147 DGND 0.30fF
C2773 Vxp.t3 DGND 0.30fF
C2774 Vxp.t35 DGND 0.30fF
C2775 Vxp.t4 DGND 0.30fF
C2776 Vxp.n128 DGND 7.33fF $ **FLOATING
C2777 Vxp.n129 DGND 7.33fF $ **FLOATING
C2778 Vxp.n130 DGND 7.33fF $ **FLOATING
C2779 Vxp.n131 DGND 7.98fF $ **FLOATING
C2780 Vxp.n132 DGND 3.59fF $ **FLOATING
C2781 Vxp.t10 DGND 0.30fF
C2782 Vxp.t19 DGND 0.30fF
C2783 Vxp.t33 DGND 0.30fF
C2784 Vxp.t145 DGND 0.30fF
C2785 Vxp.t137 DGND 0.30fF
C2786 Vxp.n133 DGND 7.33fF $ **FLOATING
C2787 Vxp.n134 DGND 7.33fF $ **FLOATING
C2788 Vxp.n135 DGND 7.33fF $ **FLOATING
C2789 Vxp.n136 DGND 7.33fF $ **FLOATING
C2790 Vxp.n137 DGND 7.06fF $ **FLOATING
C2791 Vxp.n138 DGND 2.82fF $ **FLOATING
C2792 Vxp.t141 DGND 0.30fF
C2793 Vxp.t144 DGND 0.30fF
C2794 Vxp.t38 DGND 0.30fF
C2795 Vxp.t9 DGND 0.30fF
C2796 Vxp.t39 DGND 0.30fF
C2797 Vxp.n139 DGND 7.33fF $ **FLOATING
C2798 Vxp.n140 DGND 7.33fF $ **FLOATING
C2799 Vxp.n141 DGND 7.33fF $ **FLOATING
C2800 Vxp.n142 DGND 7.33fF $ **FLOATING
C2801 Vxp.n143 DGND 7.06fF $ **FLOATING
C2802 Vxp.n144 DGND 3.99fF $ **FLOATING
C2803 Vxp.n145 DGND 2.76fF $ **FLOATING
C2804 Vxp.n146 DGND 1.34fF $ **FLOATING
C2805 Vxp.n147 DGND 3.33fF $ **FLOATING
C2806 Vxp.n148 DGND 1.34fF $ **FLOATING
C2807 Vxp.n149 DGND 2.91fF $ **FLOATING
C2808 Vxp.n150 DGND 1.34fF $ **FLOATING
C2809 Vxp.n151 DGND 2.91fF $ **FLOATING
C2810 Vxp.n152 DGND 1.34fF $ **FLOATING
C2811 Vxp.n153 DGND 2.91fF $ **FLOATING
C2812 Vxp.n154 DGND 1.34fF $ **FLOATING
C2813 Vxp.n155 DGND 2.91fF $ **FLOATING
C2814 Vxp.n156 DGND 1.34fF $ **FLOATING
C2815 Vxp.n157 DGND 2.91fF $ **FLOATING
C2816 Vxp.n158 DGND 1.34fF $ **FLOATING
C2817 Vxp.n159 DGND 3.64fF $ **FLOATING
C2818 Vxp.n160 DGND 10.91fF $ **FLOATING
C2819 Vxp.n161 DGND 1.19fF $ **FLOATING
C2820 Vxp.n162 DGND 1.34fF $ **FLOATING
C2821 Vxp.n163 DGND 1.34fF $ **FLOATING
C2822 Vxp.n164 DGND 1.19fF $ **FLOATING
C2823 Vxp.n165 DGND 2.00fF $ **FLOATING
C2824 Vxp.n166 DGND 1.34fF $ **FLOATING
C2825 Vxp.n167 DGND 1.19fF $ **FLOATING
C2826 Vxp.n168 DGND 3.08fF $ **FLOATING
C2827 Vxp.n169 DGND 1.34fF $ **FLOATING
C2828 Vxp.n170 DGND 1.19fF $ **FLOATING
C2829 Vxp.n171 DGND 3.08fF $ **FLOATING
C2830 Vxp.n172 DGND 1.34fF $ **FLOATING
C2831 Vxp.n173 DGND 1.19fF $ **FLOATING
C2832 Vxp.n174 DGND 3.08fF $ **FLOATING
C2833 Vxp.n175 DGND 1.34fF $ **FLOATING
C2834 Vxp.n176 DGND 1.19fF $ **FLOATING
C2835 Vxp.n177 DGND 3.08fF $ **FLOATING
C2836 Vxp.n178 DGND 1.34fF $ **FLOATING
C2837 Vxp.n179 DGND 1.19fF $ **FLOATING
C2838 Vxp.n180 DGND 3.08fF $ **FLOATING
C2839 Vxp.n181 DGND 1.34fF $ **FLOATING
C2840 Vxp.n182 DGND 1.19fF $ **FLOATING
C2841 Vxp.n183 DGND 3.08fF $ **FLOATING
C2842 Vxp.n184 DGND 3.60fF $ **FLOATING
C2843 Vxp.n185 DGND 5.55fF $ **FLOATING
C2844 Vxp.n186 DGND 1.19fF $ **FLOATING
C2845 Vxp.n187 DGND 1.34fF $ **FLOATING
C2846 Vxp.n188 DGND 1.19fF $ **FLOATING
C2847 Vxp.n189 DGND 1.34fF $ **FLOATING
C2848 Vxp.n190 DGND 1.19fF $ **FLOATING
C2849 Vxp.n191 DGND 1.34fF $ **FLOATING
C2850 Vxp.n192 DGND 1.19fF $ **FLOATING
C2851 Vxp.n193 DGND 1.34fF $ **FLOATING
C2852 Vxp.n194 DGND 1.19fF $ **FLOATING
C2853 Vxp.n195 DGND 1.34fF $ **FLOATING
C2854 Vxp.n196 DGND 1.34fF $ **FLOATING
C2855 Vxp.n197 DGND 1.19fF $ **FLOATING
C2856 Vxp.n198 DGND 2.00fF $ **FLOATING
C2857 Vxp.n199 DGND 1.34fF $ **FLOATING
C2858 Vxp.n200 DGND 1.19fF $ **FLOATING
C2859 Vxp.n201 DGND 3.08fF $ **FLOATING
C2860 Vxp.n202 DGND 3.08fF $ **FLOATING
C2861 Vxp.n203 DGND 3.08fF $ **FLOATING
C2862 Vxp.n204 DGND 3.08fF $ **FLOATING
C2863 Vxp.n205 DGND 3.08fF $ **FLOATING
C2864 Vxp.n206 DGND 3.08fF $ **FLOATING
C2865 Vxp.n207 DGND 1.34fF $ **FLOATING
C2866 Vxp.n208 DGND 1.19fF $ **FLOATING
C2867 Vxp.n209 DGND 3.60fF $ **FLOATING
C2868 Vxp.n210 DGND 5.06fF $ **FLOATING
C2869 Vop.t39 DGND 0.12fF
C2870 Vop.n0 DGND 1.95fF $ **FLOATING
C2871 Vop.t35 DGND 0.12fF
C2872 Vop.n1 DGND 1.95fF $ **FLOATING
C2873 Vop.t74 DGND 0.12fF
C2874 Vop.n2 DGND 1.95fF $ **FLOATING
C2875 Vop.t29 DGND 0.12fF
C2876 Vop.n3 DGND 1.95fF $ **FLOATING
C2877 Vop.t64 DGND 0.12fF
C2878 Vop.n4 DGND 2.09fF $ **FLOATING
C2879 Vop.t67 DGND 0.12fF
C2880 Vop.n5 DGND 1.95fF $ **FLOATING
C2881 Vop.t20 DGND 0.12fF
C2882 Vop.n6 DGND 2.09fF $ **FLOATING
C2883 Vop.t22 DGND 0.12fF
C2884 Vop.n7 DGND 1.95fF $ **FLOATING
C2885 Vop.t53 DGND 0.12fF
C2886 Vop.n8 DGND 2.09fF $ **FLOATING
C2887 Vop.t58 DGND 0.12fF
C2888 Vop.n9 DGND 1.95fF $ **FLOATING
C2889 Vop.t47 DGND 0.12fF
C2890 Vop.n10 DGND 2.09fF $ **FLOATING
C2891 Vop.t48 DGND 0.12fF
C2892 Vop.n11 DGND 1.95fF $ **FLOATING
C2893 Vop.n12 DGND 1.18fF $ **FLOATING
C2894 Vop.n13 DGND 2.81fF $ **FLOATING
C2895 Vop.n14 DGND 2.81fF $ **FLOATING
C2896 Vop.n15 DGND 2.81fF $ **FLOATING
C2897 Vop.n16 DGND 2.54fF $ **FLOATING
C2898 Vop.n17 DGND 2.54fF $ **FLOATING
C2899 Vop.n18 DGND 2.54fF $ **FLOATING
C2900 Vop.n19 DGND 2.22fF $ **FLOATING
C2901 Vop.t106 DGND 0.14fF
C2902 Vop.n20 DGND 2.17fF $ **FLOATING
C2903 Vop.t115 DGND 0.14fF
C2904 Vop.n21 DGND 2.17fF $ **FLOATING
C2905 Vop.t85 DGND 0.14fF
C2906 Vop.n22 DGND 2.32fF $ **FLOATING
C2907 Vop.t107 DGND 0.14fF
C2908 Vop.n23 DGND 2.36fF $ **FLOATING
C2909 Vop.t102 DGND 0.14fF
C2910 Vop.n24 DGND 2.33fF $ **FLOATING
C2911 Vop.t94 DGND 0.14fF
C2912 Vop.n25 DGND 2.17fF $ **FLOATING
C2913 Vop.n26 DGND 1.10fF $ **FLOATING
C2914 Vop.n27 DGND 2.88fF $ **FLOATING
C2915 Vop.n28 DGND 2.46fF $ **FLOATING
C2916 Vop.n29 DGND 2.61fF $ **FLOATING
C2917 Vop.t97 DGND 0.14fF
C2918 Vop.n30 DGND 2.17fF $ **FLOATING
C2919 Vop.t111 DGND 0.14fF
C2920 Vop.n31 DGND 3.50fF $ **FLOATING
C2921 Vop.n32 DGND 2.83fF $ **FLOATING
C2922 Vop.t31 DGND 0.12fF
C2923 Vop.n33 DGND 1.95fF $ **FLOATING
C2924 Vop.t66 DGND 0.12fF
C2925 Vop.n34 DGND 1.95fF $ **FLOATING
C2926 Vop.t21 DGND 0.12fF
C2927 Vop.n35 DGND 1.95fF $ **FLOATING
C2928 Vop.t62 DGND 0.12fF
C2929 Vop.n36 DGND -4.38fF $ **FLOATING
C2930 Vop.n37 DGND 1.36fF $ **FLOATING
C2931 Vop.n38 DGND 2.54fF $ **FLOATING
C2932 Vop.n39 DGND 2.22fF $ **FLOATING
C2933 Vop.t120 DGND 2.26fF
C2934 Vop.n40 DGND 41.65fF $ **FLOATING
C2935 Vop.n41 DGND 7.06fF $ **FLOATING
C2936 Vop.t5 DGND 0.12fF
C2937 Vop.n42 DGND 1.95fF $ **FLOATING
C2938 Vop.t43 DGND 0.12fF
C2939 Vop.n43 DGND 1.95fF $ **FLOATING
C2940 Vop.t7 DGND 0.12fF
C2941 Vop.n44 DGND 1.95fF $ **FLOATING
C2942 Vop.t41 DGND 0.12fF
C2943 Vop.n45 DGND 1.95fF $ **FLOATING
C2944 Vop.t3 DGND 0.12fF
C2945 Vop.n46 DGND 1.95fF $ **FLOATING
C2946 Vop.t34 DGND 0.12fF
C2947 Vop.n47 DGND 1.95fF $ **FLOATING
C2948 Vop.t73 DGND 0.12fF
C2949 Vop.n48 DGND 1.95fF $ **FLOATING
C2950 Vop.t63 DGND 0.12fF
C2951 Vop.n49 DGND 2.71fF $ **FLOATING
C2952 Vop.n50 DGND 2.68fF $ **FLOATING
C2953 Vop.n51 DGND 2.54fF $ **FLOATING
C2954 Vop.n52 DGND 2.54fF $ **FLOATING
C2955 Vop.n53 DGND 2.54fF $ **FLOATING
C2956 Vop.n54 DGND 2.54fF $ **FLOATING
C2957 Vop.n55 DGND 2.54fF $ **FLOATING
C2958 Vop.n56 DGND 2.22fF $ **FLOATING
C2959 Vop.t113 DGND 0.14fF
C2960 Vop.n57 DGND 2.17fF $ **FLOATING
C2961 Vop.t108 DGND 0.14fF
C2962 Vop.n58 DGND 2.17fF $ **FLOATING
C2963 Vop.t114 DGND 0.14fF
C2964 Vop.n59 DGND 2.17fF $ **FLOATING
C2965 Vop.t119 DGND 0.14fF
C2966 Vop.n60 DGND 2.83fF $ **FLOATING
C2967 Vop.n61 DGND 2.58fF $ **FLOATING
C2968 Vop.n62 DGND 2.46fF $ **FLOATING
C2969 Vop.n63 DGND 2.61fF $ **FLOATING
C2970 Vop.t14 DGND 0.12fF
C2971 Vop.n64 DGND 1.86fF $ **FLOATING
C2972 Vop.t55 DGND 0.12fF
C2973 Vop.n65 DGND 1.86fF $ **FLOATING
C2974 Vop.t15 DGND 0.12fF
C2975 Vop.n66 DGND 1.86fF $ **FLOATING
C2976 Vop.t49 DGND 0.12fF
C2977 Vop.n67 DGND 1.86fF $ **FLOATING
C2978 Vop.t11 DGND 0.12fF
C2979 Vop.n68 DGND 1.86fF $ **FLOATING
C2980 Vop.t45 DGND 0.12fF
C2981 Vop.n69 DGND 1.86fF $ **FLOATING
C2982 Vop.t9 DGND 0.12fF
C2983 Vop.n70 DGND 1.86fF $ **FLOATING
C2984 Vop.t2 DGND 0.12fF
C2985 Vop.n71 DGND 2.61fF $ **FLOATING
C2986 Vop.n72 DGND 2.68fF $ **FLOATING
C2987 Vop.n73 DGND 2.54fF $ **FLOATING
C2988 Vop.n74 DGND 2.54fF $ **FLOATING
C2989 Vop.n75 DGND 2.54fF $ **FLOATING
C2990 Vop.n76 DGND 2.54fF $ **FLOATING
C2991 Vop.n77 DGND 2.54fF $ **FLOATING
C2992 Vop.n78 DGND 2.21fF $ **FLOATING
C2993 Vop.t88 DGND 0.14fF
C2994 Vop.n79 DGND 2.17fF $ **FLOATING
C2995 Vop.t92 DGND 0.14fF
C2996 Vop.n80 DGND 2.17fF $ **FLOATING
C2997 Vop.t81 DGND 0.14fF
C2998 Vop.n81 DGND 2.17fF $ **FLOATING
C2999 Vop.t86 DGND 0.14fF
C3000 Vop.n82 DGND 2.83fF $ **FLOATING
C3001 Vop.n83 DGND 2.58fF $ **FLOATING
C3002 Vop.n84 DGND 2.46fF $ **FLOATING
C3003 Vop.n85 DGND 2.61fF $ **FLOATING
C3004 Vop.n86 DGND 6.12fF $ **FLOATING
C3005 Vop.n87 DGND 9.65fF $ **FLOATING
C3006 Vop.t82 DGND 0.14fF
C3007 Vop.n88 DGND 2.17fF $ **FLOATING
C3008 Vop.t101 DGND 0.14fF
C3009 Vop.n89 DGND 2.17fF $ **FLOATING
C3010 Vop.t83 DGND 0.14fF
C3011 Vop.n90 DGND 2.17fF $ **FLOATING
C3012 Vop.t98 DGND 0.14fF
C3013 Vop.n91 DGND 2.83fF $ **FLOATING
C3014 Vop.n92 DGND 2.58fF $ **FLOATING
C3015 Vop.n93 DGND 2.46fF $ **FLOATING
C3016 Vop.n94 DGND 2.61fF $ **FLOATING
C3017 Vop.t18 DGND 0.12fF
C3018 Vop.n95 DGND 1.95fF $ **FLOATING
C3019 Vop.t6 DGND 0.12fF
C3020 Vop.n96 DGND 1.95fF $ **FLOATING
C3021 Vop.t1 DGND 0.12fF
C3022 Vop.n97 DGND 1.95fF $ **FLOATING
C3023 Vop.t30 DGND 0.12fF
C3024 Vop.n98 DGND 1.95fF $ **FLOATING
C3025 Vop.t69 DGND 0.12fF
C3026 Vop.n99 DGND 1.95fF $ **FLOATING
C3027 Vop.t24 DGND 0.12fF
C3028 Vop.n100 DGND 1.95fF $ **FLOATING
C3029 Vop.t19 DGND 0.12fF
C3030 Vop.n101 DGND 2.71fF $ **FLOATING
C3031 Vop.n102 DGND 2.68fF $ **FLOATING
C3032 Vop.n103 DGND 2.54fF $ **FLOATING
C3033 Vop.n104 DGND 2.54fF $ **FLOATING
C3034 Vop.n105 DGND 2.54fF $ **FLOATING
C3035 Vop.t36 DGND 0.12fF
C3036 Vop.n106 DGND 1.95fF $ **FLOATING
C3037 Vop.n107 DGND 2.54fF $ **FLOATING
C3038 Vop.n108 DGND 2.54fF $ **FLOATING
C3039 Vop.n109 DGND 2.22fF $ **FLOATING
C3040 Vop.n110 DGND 8.33fF $ **FLOATING
C3041 a_2458_6128.n0 DGND 1.57fF $ **FLOATING
C3042 a_2458_6128.n1 DGND 1.55fF $ **FLOATING
C3043 a_2458_6128.n2 DGND 1.57fF $ **FLOATING
C3044 a_2458_6128.n3 DGND 1.66fF $ **FLOATING
C3045 a_2458_6128.n4 DGND 1.15fF $ **FLOATING
C3046 a_2458_6128.n5 DGND 1.57fF $ **FLOATING
C3047 a_2458_6128.n6 DGND 1.55fF $ **FLOATING
C3048 a_2458_6128.n7 DGND 1.57fF $ **FLOATING
C3049 a_2458_6128.n8 DGND 1.66fF $ **FLOATING
C3050 a_2458_6128.n9 DGND 1.57fF $ **FLOATING
C3051 a_2458_6128.n10 DGND 1.55fF $ **FLOATING
C3052 a_2458_6128.n11 DGND 1.57fF $ **FLOATING
C3053 a_2458_6128.n12 DGND 1.66fF $ **FLOATING
C3054 a_2458_6128.n13 DGND 1.57fF $ **FLOATING
C3055 a_2458_6128.n14 DGND 1.66fF $ **FLOATING
C3056 a_2458_6128.n15 DGND 1.57fF $ **FLOATING
C3057 a_2458_6128.n16 DGND 1.66fF $ **FLOATING
C3058 a_2458_6128.n17 DGND 1.57fF $ **FLOATING
C3059 a_2458_6128.n18 DGND 1.66fF $ **FLOATING
C3060 a_2458_6128.n19 DGND 1.57fF $ **FLOATING
C3061 a_2458_6128.n20 DGND 1.66fF $ **FLOATING
C3062 a_2458_6128.n21 DGND 1.57fF $ **FLOATING
C3063 a_2458_6128.n22 DGND 1.66fF $ **FLOATING
C3064 a_2458_6128.n23 DGND 1.57fF $ **FLOATING
C3065 a_2458_6128.n24 DGND 1.66fF $ **FLOATING
C3066 a_2458_6128.n25 DGND 1.57fF $ **FLOATING
C3067 a_2458_6128.n26 DGND 1.66fF $ **FLOATING
C3068 a_2458_6128.n27 DGND 1.57fF $ **FLOATING
C3069 a_2458_6128.n28 DGND 1.66fF $ **FLOATING
C3070 a_2458_6128.n29 DGND 1.57fF $ **FLOATING
C3071 a_2458_6128.n30 DGND 1.66fF $ **FLOATING
C3072 a_2458_6128.n31 DGND 1.57fF $ **FLOATING
C3073 a_2458_6128.n32 DGND 1.66fF $ **FLOATING
C3074 a_2458_6128.n33 DGND 1.57fF $ **FLOATING
C3075 a_2458_6128.n34 DGND 1.66fF $ **FLOATING
C3076 a_2458_6128.n35 DGND 1.57fF $ **FLOATING
C3077 a_2458_6128.n36 DGND 2.49fF $ **FLOATING
C3078 a_2458_6128.n37 DGND 2.00fF $ **FLOATING
C3079 a_2458_6128.n38 DGND 1.80fF $ **FLOATING
C3080 a_2458_6128.n39 DGND 1.80fF $ **FLOATING
C3081 a_2458_6128.n40 DGND 1.80fF $ **FLOATING
C3082 a_2458_6128.n41 DGND 1.80fF $ **FLOATING
C3083 a_2458_6128.n42 DGND 1.80fF $ **FLOATING
C3084 a_2458_6128.n43 DGND 1.44fF $ **FLOATING
C3085 a_2458_6128.t174 DGND 0.19fF
C3086 a_2458_6128.t83 DGND 0.19fF
C3087 a_2458_6128.n44 DGND 6.59fF $ **FLOATING
C3088 a_2458_6128.n45 DGND 4.20fF $ **FLOATING
C3089 a_2458_6128.t75 DGND 0.19fF
C3090 a_2458_6128.t5 DGND 0.19fF
C3091 a_2458_6128.t62 DGND 0.19fF
C3092 a_2458_6128.t78 DGND 0.19fF
C3093 a_2458_6128.n46 DGND 5.36fF $ **FLOATING
C3094 a_2458_6128.n47 DGND 4.29fF $ **FLOATING
C3095 a_2458_6128.n48 DGND 4.29fF $ **FLOATING
C3096 a_2458_6128.n49 DGND 5.47fF $ **FLOATING
C3097 a_2458_6128.t182 DGND 0.19fF
C3098 a_2458_6128.t68 DGND 0.19fF
C3099 a_2458_6128.n50 DGND 6.59fF $ **FLOATING
C3100 a_2458_6128.n51 DGND 4.20fF $ **FLOATING
C3101 a_2458_6128.t181 DGND 0.19fF
C3102 a_2458_6128.t93 DGND 0.19fF
C3103 a_2458_6128.n52 DGND 6.59fF $ **FLOATING
C3104 a_2458_6128.n53 DGND 4.20fF $ **FLOATING
C3105 a_2458_6128.t82 DGND 0.19fF
C3106 a_2458_6128.t85 DGND 0.19fF
C3107 a_2458_6128.t88 DGND 0.19fF
C3108 a_2458_6128.t70 DGND 0.19fF
C3109 a_2458_6128.n54 DGND 5.36fF $ **FLOATING
C3110 a_2458_6128.n55 DGND 4.29fF $ **FLOATING
C3111 a_2458_6128.n56 DGND 4.29fF $ **FLOATING
C3112 a_2458_6128.n57 DGND 5.47fF $ **FLOATING
C3113 a_2458_6128.t73 DGND 0.19fF
C3114 a_2458_6128.t71 DGND 0.19fF
C3115 a_2458_6128.n58 DGND 6.59fF $ **FLOATING
C3116 a_2458_6128.n59 DGND 4.20fF $ **FLOATING
C3117 a_2458_6128.t79 DGND 0.19fF
C3118 a_2458_6128.t175 DGND 0.19fF
C3119 a_2458_6128.t80 DGND 0.19fF
C3120 a_2458_6128.t89 DGND 0.19fF
C3121 a_2458_6128.n60 DGND 5.44fF $ **FLOATING
C3122 a_2458_6128.n61 DGND 4.29fF $ **FLOATING
C3123 a_2458_6128.n62 DGND 4.29fF $ **FLOATING
C3124 a_2458_6128.n63 DGND 5.56fF $ **FLOATING
C3125 a_2458_6128.n64 DGND 3.77fF $ **FLOATING
C3126 a_2458_6128.n65 DGND 2.58fF $ **FLOATING
C3127 a_2458_6128.n66 DGND 1.55fF $ **FLOATING
C3128 a_2458_6128.n67 DGND 1.55fF $ **FLOATING
C3129 a_2458_6128.n68 DGND 2.58fF $ **FLOATING
C3130 a_2458_6128.n69 DGND 1.55fF $ **FLOATING
C3131 a_2458_6128.t67 DGND 0.19fF
C3132 a_2458_6128.t63 DGND 0.19fF
C3133 a_2458_6128.t199 DGND 0.19fF
C3134 a_2458_6128.t188 DGND 0.19fF
C3135 a_2458_6128.n70 DGND 5.36fF $ **FLOATING
C3136 a_2458_6128.n71 DGND 4.29fF $ **FLOATING
C3137 a_2458_6128.n72 DGND 4.29fF $ **FLOATING
C3138 a_2458_6128.n73 DGND 5.47fF $ **FLOATING
C3139 a_2458_6128.n74 DGND 13.43fF $ **FLOATING
C3140 a_2458_6128.n75 DGND 1.57fF $ **FLOATING
C3141 a_2458_6128.n76 DGND 1.66fF $ **FLOATING
C3142 a_2458_6128.n77 DGND 1.57fF $ **FLOATING
C3143 a_2458_6128.n78 DGND 1.66fF $ **FLOATING
C3144 a_2458_6128.n79 DGND 1.57fF $ **FLOATING
C3145 a_2458_6128.n80 DGND 1.66fF $ **FLOATING
C3146 a_2458_6128.n81 DGND 1.57fF $ **FLOATING
C3147 a_2458_6128.n82 DGND 1.66fF $ **FLOATING
C3148 a_2458_6128.n83 DGND 1.57fF $ **FLOATING
C3149 a_2458_6128.n84 DGND 1.66fF $ **FLOATING
C3150 a_2458_6128.n85 DGND 1.57fF $ **FLOATING
C3151 a_2458_6128.n86 DGND 1.66fF $ **FLOATING
C3152 a_2458_6128.n87 DGND 1.57fF $ **FLOATING
C3153 a_2458_6128.n88 DGND 1.66fF $ **FLOATING
C3154 a_2458_6128.n89 DGND 1.57fF $ **FLOATING
C3155 a_2458_6128.n90 DGND 2.49fF $ **FLOATING
C3156 a_2458_6128.n91 DGND 2.00fF $ **FLOATING
C3157 a_2458_6128.n92 DGND 1.80fF $ **FLOATING
C3158 a_2458_6128.n93 DGND 1.80fF $ **FLOATING
C3159 a_2458_6128.n94 DGND 1.80fF $ **FLOATING
C3160 a_2458_6128.n95 DGND 1.80fF $ **FLOATING
C3161 a_2458_6128.n96 DGND 1.80fF $ **FLOATING
C3162 a_2458_6128.n97 DGND 1.44fF $ **FLOATING
C3163 a_2458_6128.n98 DGND 1.57fF $ **FLOATING
C3164 a_2458_6128.n99 DGND 1.66fF $ **FLOATING
C3165 a_2458_6128.n100 DGND 1.57fF $ **FLOATING
C3166 a_2458_6128.n101 DGND 1.66fF $ **FLOATING
C3167 a_2458_6128.n102 DGND 1.57fF $ **FLOATING
C3168 a_2458_6128.n103 DGND 1.66fF $ **FLOATING
C3169 a_2458_6128.n104 DGND 1.57fF $ **FLOATING
C3170 a_2458_6128.n105 DGND 1.66fF $ **FLOATING
C3171 a_2458_6128.n106 DGND 1.57fF $ **FLOATING
C3172 a_2458_6128.n107 DGND 1.66fF $ **FLOATING
C3173 a_2458_6128.n108 DGND 1.57fF $ **FLOATING
C3174 a_2458_6128.n109 DGND 1.66fF $ **FLOATING
C3175 a_2458_6128.n110 DGND 1.57fF $ **FLOATING
C3176 a_2458_6128.n111 DGND 1.66fF $ **FLOATING
C3177 a_2458_6128.n112 DGND 1.57fF $ **FLOATING
C3178 a_2458_6128.n113 DGND 2.49fF $ **FLOATING
C3179 a_2458_6128.n114 DGND 2.00fF $ **FLOATING
C3180 a_2458_6128.n115 DGND 1.80fF $ **FLOATING
C3181 a_2458_6128.n116 DGND 1.80fF $ **FLOATING
C3182 a_2458_6128.n117 DGND 1.80fF $ **FLOATING
C3183 a_2458_6128.n118 DGND 1.80fF $ **FLOATING
C3184 a_2458_6128.n119 DGND 1.80fF $ **FLOATING
C3185 a_2458_6128.n120 DGND 1.44fF $ **FLOATING
C3186 a_2458_6128.t90 DGND 0.19fF
C3187 a_2458_6128.t84 DGND 0.19fF
C3188 a_2458_6128.n121 DGND 6.59fF $ **FLOATING
C3189 a_2458_6128.n122 DGND 4.07fF $ **FLOATING
C3190 a_2458_6128.n123 DGND 3.30fF $ **FLOATING
C3191 a_2458_6128.n124 DGND 2.33fF $ **FLOATING
C3192 a_2458_6128.t183 DGND 0.19fF
C3193 a_2458_6128.t69 DGND 0.19fF
C3194 a_2458_6128.n125 DGND 6.59fF $ **FLOATING
C3195 a_2458_6128.n126 DGND 4.07fF $ **FLOATING
C3196 a_2458_6128.n127 DGND 1.33fF $ **FLOATING
C3197 a_2458_6128.t192 DGND 0.19fF
C3198 a_2458_6128.t176 DGND 0.19fF
C3199 a_2458_6128.n128 DGND 6.59fF $ **FLOATING
C3200 a_2458_6128.n129 DGND 4.07fF $ **FLOATING
C3201 a_2458_6128.n130 DGND 1.33fF $ **FLOATING
C3202 a_2458_6128.n131 DGND 2.33fF $ **FLOATING
C3203 a_2458_6128.t72 DGND 0.19fF
C3204 a_2458_6128.t74 DGND 0.19fF
C3205 a_2458_6128.n132 DGND 6.59fF $ **FLOATING
C3206 a_2458_6128.n133 DGND 4.07fF $ **FLOATING
C3207 a_2458_6128.n134 DGND 1.33fF $ **FLOATING
C3208 a_2458_6128.n135 DGND 26.30fF $ **FLOATING
C3209 a_2458_6128.n136 DGND 27.38fF $ **FLOATING
C3210 a_2458_6128.n137 DGND 4.49fF $ **FLOATING
C3211 a_2458_6128.n138 DGND 14.00fF $ **FLOATING
C3212 a_2458_6128.n139 DGND 4.32fF $ **FLOATING
C3213 a_2458_6128.n140 DGND 1.57fF $ **FLOATING
C3214 a_2458_6128.n141 DGND 1.66fF $ **FLOATING
C3215 a_2458_6128.n142 DGND 1.57fF $ **FLOATING
C3216 a_2458_6128.n143 DGND 1.66fF $ **FLOATING
C3217 a_2458_6128.n144 DGND 1.57fF $ **FLOATING
C3218 a_2458_6128.n145 DGND 1.66fF $ **FLOATING
C3219 a_2458_6128.n146 DGND 1.57fF $ **FLOATING
C3220 a_2458_6128.n147 DGND -2.11fF $ **FLOATING
C3221 a_2458_6128.n148 DGND 0.87fF $ **FLOATING
C3222 a_2458_6128.n149 DGND 1.80fF $ **FLOATING
C3223 a_2458_6128.n150 DGND 1.44fF $ **FLOATING
C3224 a_2458_6128.n151 DGND 0.36fF $ **FLOATING
C3225 a_2458_6128.n152 DGND 0.36fF $ **FLOATING
C3226 a_2458_6128.n153 DGND 0.36fF $ **FLOATING
C3227 a_2458_6128.t196 DGND 0.16fF
C3228 a_2458_6128.n154 DGND 0.94fF $ **FLOATING
C3229 a_2458_6128.n155 DGND 0.39fF $ **FLOATING
C3230 a_2458_6128.n156 DGND 0.57fF $ **FLOATING
C3231 a_2458_6128.n157 DGND 10.21fF $ **FLOATING
C3232 a_2458_6128.n158 DGND 19.78fF $ **FLOATING
C3233 a_2458_6128.n159 DGND 5.68fF $ **FLOATING
C3234 a_2458_6128.n160 DGND 1.44fF $ **FLOATING
C3235 a_2458_6128.n161 DGND 1.80fF $ **FLOATING
C3236 a_2458_6128.n162 DGND 1.80fF $ **FLOATING
C3237 a_2458_6128.n163 DGND 1.80fF $ **FLOATING
C3238 a_2458_6128.n164 DGND 1.90fF $ **FLOATING
C3239 a_2458_6128.n165 DGND 1.90fF $ **FLOATING
C3240 a_2458_6128.n166 DGND 1.57fF $ **FLOATING
C3241 a_2458_6128.n167 DGND 1.66fF $ **FLOATING
C3242 a_2458_6128.n168 DGND 1.90fF $ **FLOATING
C3243 a_2458_6128.n169 DGND 1.57fF $ **FLOATING
C3244 a_2458_6128.n170 DGND 1.55fF $ **FLOATING
C3245 a_2467_n29152.t0 DGND 2.42fF
C3246 a_2467_n29152.t19 DGND 2.42fF
C3247 a_2467_n29152.t3 DGND 2.42fF
C3248 a_2467_n29152.t4 DGND 2.43fF
C3249 a_2467_n29152.t1 DGND 2.43fF
C3250 a_2467_n29152.t18 DGND 2.43fF
C3251 a_2467_n29152.t2 DGND 2.63fF
C3252 a_2467_n29152.n0 DGND 13.82fF $ **FLOATING
C3253 a_2467_n29152.n1 DGND 4.82fF $ **FLOATING
C3254 a_2467_n29152.n2 DGND 7.19fF $ **FLOATING
C3255 a_2467_n29152.t7 DGND 0.12fF
C3256 a_2467_n29152.n3 DGND 2.22fF $ **FLOATING
C3257 a_2467_n29152.n4 DGND 1.30fF $ **FLOATING
C3258 a_2467_n29152.n5 DGND 1.30fF $ **FLOATING
C3259 a_2467_n29152.n6 DGND 1.30fF $ **FLOATING
C3260 a_2467_n29152.n7 DGND 0.94fF $ **FLOATING
C3261 a_2467_n29152.t14 DGND 0.12fF
C3262 a_2467_n29152.n8 DGND 2.22fF $ **FLOATING
C3263 a_2467_n29152.n9 DGND 1.30fF $ **FLOATING
C3264 a_2467_n29152.n10 DGND 1.30fF $ **FLOATING
C3265 a_2467_n29152.n11 DGND 1.30fF $ **FLOATING
C3266 a_2467_n29152.n12 DGND 2.21fF $ **FLOATING
C3267 a_2467_n29152.n13 DGND 9.08fF $ **FLOATING
C3268 a_2467_n29152.n14 DGND 54.65fF $ **FLOATING
C3269 a_2467_n29152.n15 DGND 32.46fF $ **FLOATING
C3270 a_2467_n29152.n16 DGND 4.81fF $ **FLOATING
C3271 a_2467_n29152.n17 DGND 13.80fF $ **FLOATING
C3272 a_2467_n29152.t5 DGND 2.62fF
C3273 Vfold_bot_m.t54 DGND 0.29fF
C3274 Vfold_bot_m.n0 DGND 0.72fF $ **FLOATING
C3275 Vfold_bot_m.n1 DGND 0.72fF $ **FLOATING
C3276 Vfold_bot_m.n2 DGND 0.72fF $ **FLOATING
C3277 Vfold_bot_m.t109 DGND 0.36fF
C3278 Vfold_bot_m.n3 DGND 1.52fF $ **FLOATING
C3279 Vfold_bot_m.n4 DGND 0.53fF $ **FLOATING
C3280 Vfold_bot_m.n5 DGND 0.53fF $ **FLOATING
C3281 Vfold_bot_m.n6 DGND 12.55fF $ **FLOATING
C3282 Vfold_bot_m.n7 DGND 1.69fF $ **FLOATING
C3283 Vfold_bot_m.n8 DGND 1.88fF $ **FLOATING
C3284 Vfold_bot_m.n9 DGND 1.69fF $ **FLOATING
C3285 Vfold_bot_m.n10 DGND 1.88fF $ **FLOATING
C3286 Vfold_bot_m.n11 DGND 1.69fF $ **FLOATING
C3287 Vfold_bot_m.n12 DGND 2.07fF $ **FLOATING
C3288 Vfold_bot_m.n13 DGND 2.06fF $ **FLOATING
C3289 Vfold_bot_m.n14 DGND 1.88fF $ **FLOATING
C3290 Vfold_bot_m.n15 DGND 1.69fF $ **FLOATING
C3291 Vfold_bot_m.n16 DGND 2.07fF $ **FLOATING
C3292 Vfold_bot_m.n17 DGND 2.06fF $ **FLOATING
C3293 Vfold_bot_m.n18 DGND 2.82fF $ **FLOATING
C3294 Vfold_bot_m.n19 DGND 2.16fF $ **FLOATING
C3295 Vfold_bot_m.n20 DGND 1.97fF $ **FLOATING
C3296 Vfold_bot_m.n21 DGND 1.59fF $ **FLOATING
C3297 Vfold_bot_m.n22 DGND 1.69fF $ **FLOATING
C3298 Vfold_bot_m.n23 DGND 1.88fF $ **FLOATING
C3299 Vfold_bot_m.n24 DGND 1.69fF $ **FLOATING
C3300 Vfold_bot_m.n25 DGND 0.26fF $ **FLOATING
C3301 Vfold_bot_m.n26 DGND 1.26fF $ **FLOATING
C3302 Vfold_bot_m.n27 DGND 1.69fF $ **FLOATING
C3303 Vfold_bot_m.n28 DGND 1.88fF $ **FLOATING
C3304 Vfold_bot_m.n29 DGND 1.69fF $ **FLOATING
C3305 Vfold_bot_m.n30 DGND 1.88fF $ **FLOATING
C3306 Vfold_bot_m.n31 DGND 1.69fF $ **FLOATING
C3307 Vfold_bot_m.n32 DGND 1.88fF $ **FLOATING
C3308 Vfold_bot_m.n33 DGND 1.69fF $ **FLOATING
C3309 Vfold_bot_m.n34 DGND 2.82fF $ **FLOATING
C3310 Vfold_bot_m.n35 DGND 2.16fF $ **FLOATING
C3311 Vfold_bot_m.n36 DGND 1.97fF $ **FLOATING
C3312 Vfold_bot_m.n37 DGND 1.59fF $ **FLOATING
C3313 Vfold_bot_m.t2 DGND 0.24fF
C3314 Vfold_bot_m.n38 DGND 7.08fF $ **FLOATING
C3315 Vfold_bot_m.t115 DGND 0.24fF
C3316 Vfold_bot_m.n39 DGND 4.48fF $ **FLOATING
C3317 Vfold_bot_m.t32 DGND 0.24fF
C3318 Vfold_bot_m.n40 DGND 5.75fF $ **FLOATING
C3319 Vfold_bot_m.t111 DGND 0.24fF
C3320 Vfold_bot_m.n41 DGND 4.61fF $ **FLOATING
C3321 Vfold_bot_m.t61 DGND 0.24fF
C3322 Vfold_bot_m.n42 DGND 4.61fF $ **FLOATING
C3323 Vfold_bot_m.t22 DGND 0.24fF
C3324 Vfold_bot_m.n43 DGND 5.86fF $ **FLOATING
C3325 Vfold_bot_m.t118 DGND 0.24fF
C3326 Vfold_bot_m.n44 DGND 7.08fF $ **FLOATING
C3327 Vfold_bot_m.t16 DGND 0.24fF
C3328 Vfold_bot_m.n45 DGND 4.48fF $ **FLOATING
C3329 Vfold_bot_m.t7 DGND 0.23fF
C3330 Vfold_bot_m.n46 DGND 5.71fF $ **FLOATING
C3331 Vfold_bot_m.t30 DGND 0.23fF
C3332 Vfold_bot_m.n47 DGND 4.56fF $ **FLOATING
C3333 Vfold_bot_m.t1 DGND 0.23fF
C3334 Vfold_bot_m.n48 DGND 4.56fF $ **FLOATING
C3335 Vfold_bot_m.t10 DGND 0.23fF
C3336 Vfold_bot_m.n49 DGND 5.82fF $ **FLOATING
C3337 Vfold_bot_m.t106 DGND 0.23fF
C3338 Vfold_bot_m.n50 DGND 5.71fF $ **FLOATING
C3339 Vfold_bot_m.t9 DGND 0.23fF
C3340 Vfold_bot_m.n51 DGND 4.56fF $ **FLOATING
C3341 Vfold_bot_m.t107 DGND 0.23fF
C3342 Vfold_bot_m.n52 DGND 4.56fF $ **FLOATING
C3343 Vfold_bot_m.t5 DGND 0.23fF
C3344 Vfold_bot_m.n53 DGND 5.82fF $ **FLOATING
C3345 Vfold_bot_m.t62 DGND 0.23fF
C3346 Vfold_bot_m.n54 DGND 7.03fF $ **FLOATING
C3347 Vfold_bot_m.t19 DGND 0.23fF
C3348 Vfold_bot_m.n55 DGND 4.46fF $ **FLOATING
C3349 Vfold_bot_m.t20 DGND 0.23fF
C3350 Vfold_bot_m.n56 DGND 7.03fF $ **FLOATING
C3351 Vfold_bot_m.t6 DGND 0.23fF
C3352 Vfold_bot_m.n57 DGND 4.58fF $ **FLOATING
C3353 Vfold_bot_m.t21 DGND 0.23fF
C3354 Vfold_bot_m.t24 DGND 0.23fF
C3355 Vfold_bot_m.t8 DGND 0.23fF
C3356 Vfold_bot_m.t23 DGND 0.23fF
C3357 Vfold_bot_m.n58 DGND 5.71fF $ **FLOATING
C3358 Vfold_bot_m.n59 DGND 4.56fF $ **FLOATING
C3359 Vfold_bot_m.n60 DGND 4.56fF $ **FLOATING
C3360 Vfold_bot_m.n61 DGND 5.82fF $ **FLOATING
C3361 Vfold_bot_m.n62 DGND 3.84fF $ **FLOATING
C3362 Vfold_bot_m.n63 DGND 1.69fF $ **FLOATING
C3363 Vfold_bot_m.n64 DGND 2.79fF $ **FLOATING
C3364 Vfold_bot_m.n65 DGND 2.79fF $ **FLOATING
C3365 Vfold_bot_m.n66 DGND 1.72fF $ **FLOATING
C3366 Vfold_bot_m.n67 DGND 2.81fF $ **FLOATING
C3367 Vfold_bot_m.n68 DGND 19.00fF $ **FLOATING
C3368 Vfold_bot_m.n69 DGND 1.69fF $ **FLOATING
C3369 Vfold_bot_m.n70 DGND 1.88fF $ **FLOATING
C3370 Vfold_bot_m.n71 DGND 1.69fF $ **FLOATING
C3371 Vfold_bot_m.n72 DGND 1.88fF $ **FLOATING
C3372 Vfold_bot_m.n73 DGND 1.69fF $ **FLOATING
C3373 Vfold_bot_m.n74 DGND 1.88fF $ **FLOATING
C3374 Vfold_bot_m.n75 DGND 1.69fF $ **FLOATING
C3375 Vfold_bot_m.n76 DGND 2.82fF $ **FLOATING
C3376 Vfold_bot_m.n77 DGND 2.16fF $ **FLOATING
C3377 Vfold_bot_m.n78 DGND 1.97fF $ **FLOATING
C3378 Vfold_bot_m.n79 DGND 1.59fF $ **FLOATING
C3379 Vfold_bot_m.t117 DGND 0.23fF
C3380 Vfold_bot_m.t0 DGND 0.23fF
C3381 Vfold_bot_m.n80 DGND 7.02fF $ **FLOATING
C3382 Vfold_bot_m.n81 DGND 4.42fF $ **FLOATING
C3383 Vfold_bot_m.n82 DGND 3.25fF $ **FLOATING
C3384 Vfold_bot_m.t18 DGND 0.23fF
C3385 Vfold_bot_m.t31 DGND 0.23fF
C3386 Vfold_bot_m.n83 DGND 7.02fF $ **FLOATING
C3387 Vfold_bot_m.n84 DGND 4.31fF $ **FLOATING
C3388 Vfold_bot_m.n85 DGND 1.41fF $ **FLOATING
C3389 Vfold_bot_m.n86 DGND 2.48fF $ **FLOATING
C3390 Vfold_bot_m.n87 DGND 2.48fF $ **FLOATING
C3391 Vfold_bot_m.t17 DGND 0.24fF
C3392 Vfold_bot_m.t116 DGND 0.24fF
C3393 Vfold_bot_m.n88 DGND 7.08fF $ **FLOATING
C3394 Vfold_bot_m.n89 DGND 4.34fF $ **FLOATING
C3395 Vfold_bot_m.n90 DGND 1.44fF $ **FLOATING
C3396 Vfold_bot_m.n91 DGND 2.50fF $ **FLOATING
C3397 Vfold_bot_m.t105 DGND 0.24fF
C3398 Vfold_bot_m.t110 DGND 0.24fF
C3399 Vfold_bot_m.n92 DGND 7.08fF $ **FLOATING
C3400 Vfold_bot_m.n93 DGND 4.34fF $ **FLOATING
C3401 Vfold_bot_m.n94 DGND 32.16fF $ **FLOATING
C3402 Vfold_bot_m.n95 DGND 1.69fF $ **FLOATING
C3403 Vfold_bot_m.n96 DGND 1.88fF $ **FLOATING
C3404 Vfold_bot_m.n97 DGND 1.69fF $ **FLOATING
C3405 Vfold_bot_m.n98 DGND 1.88fF $ **FLOATING
C3406 Vfold_bot_m.n99 DGND 1.69fF $ **FLOATING
C3407 Vfold_bot_m.n100 DGND 2.82fF $ **FLOATING
C3408 Vfold_bot_m.n101 DGND 2.16fF $ **FLOATING
C3409 Vfold_bot_m.n102 DGND 1.69fF $ **FLOATING
C3410 Vfold_bot_m.n103 DGND 1.88fF $ **FLOATING
C3411 Vfold_bot_m.n104 DGND 1.97fF $ **FLOATING
C3412 Vfold_bot_m.n105 DGND 1.59fF $ **FLOATING
C3413 Vfold_bot_m.n106 DGND 35.55fF $ **FLOATING
C3414 Vfold_bot_m.n107 DGND 5.54fF $ **FLOATING
C3415 Vfold_bot_m.n108 DGND 20.64fF $ **FLOATING
C3416 Vfold_bot_m.n109 DGND 3.96fF $ **FLOATING
C3417 Vfold_bot_m.n110 DGND 6.12fF $ **FLOATING
C3418 Vfold_bot_m.n111 DGND 8.18fF $ **FLOATING
C3419 a_2370_n29452.t4 DGND 0.11fF
C3420 a_2370_n29452.t3 DGND 0.11fF
C3421 a_2370_n29452.n0 DGND 0.85fF $ **FLOATING
C3422 a_2370_n29452.t2 DGND 0.11fF
C3423 a_2370_n29452.t1 DGND 0.11fF
C3424 a_2370_n29452.n1 DGND 0.85fF $ **FLOATING
C3425 a_2370_n29452.t7 DGND 0.11fF
C3426 a_2370_n29452.t6 DGND 0.11fF
C3427 a_2370_n29452.n2 DGND 0.85fF $ **FLOATING
C3428 a_2370_n29452.t9 DGND 4.17fF
C3429 a_2370_n29452.t11 DGND 4.27fF
C3430 a_2370_n29452.n3 DGND 6.29fF $ **FLOATING
C3431 a_2370_n29452.t10 DGND 4.37fF
C3432 a_2370_n29452.t8 DGND 4.46fF
C3433 a_2370_n29452.n4 DGND 17.13fF $ **FLOATING
C3434 a_2370_n29452.n5 DGND 45.32fF $ **FLOATING
C3435 a_2370_n29452.n6 DGND 2.99fF $ **FLOATING
C3436 a_2370_n29452.n7 DGND 1.09fF $ **FLOATING
C3437 a_2370_n29452.n8 DGND 1.18fF $ **FLOATING
C3438 a_2370_n29452.t5 DGND 0.11fF
C3439 a_2370_n29452.n9 DGND 0.88fF $ **FLOATING
C3440 a_2370_n29452.t0 DGND 0.11fF
C3441 a_12760_n20342.n0 DGND 3.69fF $ **FLOATING
C3442 a_12760_n20342.n1 DGND 3.69fF $ **FLOATING
C3443 a_12760_n20342.n2 DGND 3.10fF $ **FLOATING
C3444 a_12760_n20342.n3 DGND 1.84fF $ **FLOATING
C3445 a_12760_n20342.n4 DGND 3.69fF $ **FLOATING
C3446 a_12760_n20342.n5 DGND 3.10fF $ **FLOATING
C3447 a_12760_n20342.n6 DGND 3.69fF $ **FLOATING
C3448 a_12760_n20342.n7 DGND 3.10fF $ **FLOATING
C3449 a_12760_n20342.n8 DGND 1.26fF $ **FLOATING
C3450 a_12760_n20342.n9 DGND 3.69fF $ **FLOATING
C3451 a_12760_n20342.n10 DGND 3.69fF $ **FLOATING
C3452 a_12760_n20342.n11 DGND 3.68fF $ **FLOATING
C3453 a_12760_n20342.n12 DGND 1.84fF $ **FLOATING
C3454 a_12760_n20342.n13 DGND 3.69fF $ **FLOATING
C3455 a_12760_n20342.n14 DGND 3.10fF $ **FLOATING
C3456 a_12760_n20342.n15 DGND 3.69fF $ **FLOATING
C3457 a_12760_n20342.n16 DGND 3.69fF $ **FLOATING
C3458 a_12760_n20342.n17 DGND 4.06fF $ **FLOATING
C3459 a_12760_n20342.n18 DGND 3.36fF $ **FLOATING
C3460 a_12760_n20342.n19 DGND 5.85fF $ **FLOATING
C3461 a_12760_n20342.n20 DGND 1.32fF $ **FLOATING
C3462 a_12760_n20342.n21 DGND 2.39fF $ **FLOATING
C3463 a_12760_n20342.n22 DGND 2.39fF $ **FLOATING
C3464 a_12760_n20342.n23 DGND 2.39fF $ **FLOATING
C3465 a_12760_n20342.n24 DGND 2.39fF $ **FLOATING
C3466 a_12760_n20342.n25 DGND 2.22fF $ **FLOATING
C3467 a_12760_n20342.n26 DGND 2.39fF $ **FLOATING
C3468 a_12760_n20342.n27 DGND 2.39fF $ **FLOATING
C3469 a_12760_n20342.n28 DGND 2.39fF $ **FLOATING
C3470 a_12760_n20342.n29 DGND 2.22fF $ **FLOATING
C3471 a_12760_n20342.n30 DGND 2.39fF $ **FLOATING
C3472 a_12760_n20342.n31 DGND 2.39fF $ **FLOATING
C3473 a_12760_n20342.n32 DGND 2.39fF $ **FLOATING
C3474 a_12760_n20342.n33 DGND 2.39fF $ **FLOATING
C3475 a_12760_n20342.n34 DGND 2.39fF $ **FLOATING
C3476 a_12760_n20342.n35 DGND 2.39fF $ **FLOATING
C3477 a_12760_n20342.n36 DGND 2.39fF $ **FLOATING
C3478 a_12760_n20342.n37 DGND 2.39fF $ **FLOATING
C3479 a_12760_n20342.n38 DGND 2.39fF $ **FLOATING
C3480 a_12760_n20342.n39 DGND 2.22fF $ **FLOATING
C3481 a_12760_n20342.n40 DGND 2.22fF $ **FLOATING
C3482 a_12760_n20342.n41 DGND 2.22fF $ **FLOATING
C3483 a_12760_n20342.n42 DGND 2.39fF $ **FLOATING
C3484 a_12760_n20342.n43 DGND 2.39fF $ **FLOATING
C3485 a_12760_n20342.n44 DGND 2.39fF $ **FLOATING
C3486 a_12760_n20342.n45 DGND 2.22fF $ **FLOATING
C3487 a_12760_n20342.n46 DGND 2.39fF $ **FLOATING
C3488 a_12760_n20342.n47 DGND 2.22fF $ **FLOATING
C3489 a_12760_n20342.n48 DGND 2.39fF $ **FLOATING
C3490 a_12760_n20342.n49 DGND 2.39fF $ **FLOATING
C3491 a_12760_n20342.n50 DGND 2.39fF $ **FLOATING
C3492 a_12760_n20342.n51 DGND 2.39fF $ **FLOATING
C3493 a_12760_n20342.n52 DGND 2.39fF $ **FLOATING
C3494 a_12760_n20342.n53 DGND 2.39fF $ **FLOATING
C3495 a_12760_n20342.n54 DGND 2.82fF $ **FLOATING
C3496 a_12760_n20342.n55 DGND 2.39fF $ **FLOATING
C3497 a_12760_n20342.n56 DGND 2.39fF $ **FLOATING
C3498 a_12760_n20342.n57 DGND 2.39fF $ **FLOATING
C3499 a_12760_n20342.n58 DGND 2.82fF $ **FLOATING
C3500 a_12760_n20342.n59 DGND 2.39fF $ **FLOATING
C3501 a_12760_n20342.n60 DGND 2.39fF $ **FLOATING
C3502 a_12760_n20342.n61 DGND 2.39fF $ **FLOATING
C3503 a_12760_n20342.n62 DGND 2.39fF $ **FLOATING
C3504 a_12760_n20342.n63 DGND 2.39fF $ **FLOATING
C3505 a_12760_n20342.n64 DGND 2.39fF $ **FLOATING
C3506 a_12760_n20342.n65 DGND 2.39fF $ **FLOATING
C3507 a_12760_n20342.n66 DGND 2.39fF $ **FLOATING
C3508 a_12760_n20342.n67 DGND 2.39fF $ **FLOATING
C3509 a_12760_n20342.n68 DGND 2.39fF $ **FLOATING
C3510 a_12760_n20342.n69 DGND 2.39fF $ **FLOATING
C3511 a_12760_n20342.n70 DGND 2.39fF $ **FLOATING
C3512 a_12760_n20342.n71 DGND 2.39fF $ **FLOATING
C3513 a_12760_n20342.n72 DGND 2.39fF $ **FLOATING
C3514 a_12760_n20342.n73 DGND 2.39fF $ **FLOATING
C3515 a_12760_n20342.n74 DGND 2.39fF $ **FLOATING
C3516 a_12760_n20342.n75 DGND 2.39fF $ **FLOATING
C3517 a_12760_n20342.n76 DGND 2.39fF $ **FLOATING
C3518 a_12760_n20342.n77 DGND 2.41fF $ **FLOATING
C3519 a_12760_n20342.n78 DGND 2.47fF $ **FLOATING
C3520 a_12760_n20342.n79 DGND 2.28fF $ **FLOATING
C3521 a_12760_n20342.n80 DGND 2.36fF $ **FLOATING
C3522 a_12760_n20342.n81 DGND 2.19fF $ **FLOATING
C3523 a_12760_n20342.n82 DGND 2.83fF $ **FLOATING
C3524 a_12760_n20342.t32 DGND 1.70fF
C3525 a_12760_n20342.t42 DGND 1.70fF
C3526 a_12760_n20342.n84 DGND 0.12fF $ **FLOATING
C3527 a_12760_n20342.n85 DGND 0.12fF $ **FLOATING
C3528 a_12760_n20342.t92 DGND 1.70fF
C3529 a_12760_n20342.t107 DGND 1.70fF
C3530 a_12760_n20342.n87 DGND 0.12fF $ **FLOATING
C3531 a_12760_n20342.n88 DGND 0.12fF $ **FLOATING
C3532 a_12760_n20342.n89 DGND 2.43fF $ **FLOATING
C3533 a_12760_n20342.t4 DGND 1.34fF
C3534 a_12760_n20342.t11 DGND 1.70fF
C3535 a_12760_n20342.t24 DGND 1.70fF
C3536 a_12760_n20342.n91 DGND 0.12fF $ **FLOATING
C3537 a_12760_n20342.n92 DGND 0.12fF $ **FLOATING
C3538 a_12760_n20342.t10 DGND 1.70fF
C3539 a_12760_n20342.t22 DGND 1.70fF
C3540 a_12760_n20342.n94 DGND 0.12fF $ **FLOATING
C3541 a_12760_n20342.n95 DGND 0.12fF $ **FLOATING
C3542 a_12760_n20342.t70 DGND 1.70fF
C3543 a_12760_n20342.t84 DGND 1.70fF
C3544 a_12760_n20342.n97 DGND 0.12fF $ **FLOATING
C3545 a_12760_n20342.n98 DGND 0.12fF $ **FLOATING
C3546 a_12760_n20342.t78 DGND 1.70fF
C3547 a_12760_n20342.t90 DGND 1.70fF
C3548 a_12760_n20342.n100 DGND 0.12fF $ **FLOATING
C3549 a_12760_n20342.n101 DGND 0.12fF $ **FLOATING
C3550 a_12760_n20342.t19 DGND 1.70fF
C3551 a_12760_n20342.t31 DGND 1.70fF
C3552 a_12760_n20342.n103 DGND 0.12fF $ **FLOATING
C3553 a_12760_n20342.n104 DGND 0.12fF $ **FLOATING
C3554 a_12760_n20342.t47 DGND 1.70fF
C3555 a_12760_n20342.t62 DGND 1.70fF
C3556 a_12760_n20342.n106 DGND 0.12fF $ **FLOATING
C3557 a_12760_n20342.n107 DGND 0.12fF $ **FLOATING
C3558 a_12760_n20342.t101 DGND 1.70fF
C3559 a_12760_n20342.t121 DGND 1.70fF
C3560 a_12760_n20342.n109 DGND 0.12fF $ **FLOATING
C3561 a_12760_n20342.n110 DGND 0.12fF $ **FLOATING
C3562 a_12760_n20342.t55 DGND 1.70fF
C3563 a_12760_n20342.t106 DGND 1.70fF
C3564 a_12760_n20342.n112 DGND 0.12fF $ **FLOATING
C3565 a_12760_n20342.n113 DGND 0.12fF $ **FLOATING
C3566 a_12760_n20342.n114 DGND 1.26fF $ **FLOATING
C3567 a_12760_n20342.n115 DGND 1.26fF $ **FLOATING
C3568 a_12760_n20342.t111 DGND 1.70fF
C3569 a_12760_n20342.t125 DGND 1.70fF
C3570 a_12760_n20342.n117 DGND 0.12fF $ **FLOATING
C3571 a_12760_n20342.n118 DGND 0.12fF $ **FLOATING
C3572 a_12760_n20342.t112 DGND 1.70fF
C3573 a_12760_n20342.t51 DGND 1.70fF
C3574 a_12760_n20342.n120 DGND 0.12fF $ **FLOATING
C3575 a_12760_n20342.n121 DGND 0.12fF $ **FLOATING
C3576 a_12760_n20342.t39 DGND 1.70fF
C3577 a_12760_n20342.t108 DGND 1.70fF
C3578 a_12760_n20342.n123 DGND 0.12fF $ **FLOATING
C3579 a_12760_n20342.n124 DGND 0.12fF $ **FLOATING
C3580 a_12760_n20342.t13 DGND 1.70fF
C3581 a_12760_n20342.t56 DGND 1.70fF
C3582 a_12760_n20342.n126 DGND 0.12fF $ **FLOATING
C3583 a_12760_n20342.n127 DGND 0.12fF $ **FLOATING
C3584 a_12760_n20342.n128 DGND 1.84fF $ **FLOATING
C3585 a_12760_n20342.n129 DGND 1.84fF $ **FLOATING
C3586 a_12760_n20342.t46 DGND 1.70fF
C3587 a_12760_n20342.t115 DGND 1.70fF
C3588 a_12760_n20342.n131 DGND 0.12fF $ **FLOATING
C3589 a_12760_n20342.n132 DGND 0.12fF $ **FLOATING
C3590 a_12760_n20342.t99 DGND 1.70fF
C3591 a_12760_n20342.t117 DGND 1.70fF
C3592 a_12760_n20342.n134 DGND 0.12fF $ **FLOATING
C3593 a_12760_n20342.n135 DGND 0.12fF $ **FLOATING
C3594 a_12760_n20342.t36 DGND 1.70fF
C3595 a_12760_n20342.t50 DGND 1.70fF
C3596 a_12760_n20342.n137 DGND 0.12fF $ **FLOATING
C3597 a_12760_n20342.n138 DGND 0.12fF $ **FLOATING
C3598 a_12760_n20342.t37 DGND 1.70fF
C3599 a_12760_n20342.t52 DGND 1.70fF
C3600 a_12760_n20342.n140 DGND 0.12fF $ **FLOATING
C3601 a_12760_n20342.n141 DGND 0.12fF $ **FLOATING
C3602 a_12760_n20342.t98 DGND 1.70fF
C3603 a_12760_n20342.t116 DGND 1.70fF
C3604 a_12760_n20342.n143 DGND 0.12fF $ **FLOATING
C3605 a_12760_n20342.n144 DGND 0.12fF $ **FLOATING
C3606 a_12760_n20342.t27 DGND 1.70fF
C3607 a_12760_n20342.t91 DGND 1.70fF
C3608 a_12760_n20342.n146 DGND 0.12fF $ **FLOATING
C3609 a_12760_n20342.n147 DGND 0.12fF $ **FLOATING
C3610 a_12760_n20342.t93 DGND 1.70fF
C3611 a_12760_n20342.t109 DGND 1.70fF
C3612 a_12760_n20342.n149 DGND 0.12fF $ **FLOATING
C3613 a_12760_n20342.n150 DGND 0.12fF $ **FLOATING
C3614 a_12760_n20342.t34 DGND 1.70fF
C3615 a_12760_n20342.t44 DGND 1.70fF
C3616 a_12760_n20342.n152 DGND 0.12fF $ **FLOATING
C3617 a_12760_n20342.n153 DGND 0.12fF $ **FLOATING
C3618 a_12760_n20342.t81 DGND 1.70fF
C3619 a_12760_n20342.t26 DGND 1.70fF
C3620 a_12760_n20342.n155 DGND 0.12fF $ **FLOATING
C3621 a_12760_n20342.n156 DGND 0.12fF $ **FLOATING
C3622 a_12760_n20342.t80 DGND 1.70fF
C3623 a_12760_n20342.t14 DGND 1.70fF
C3624 a_12760_n20342.n158 DGND 0.12fF $ **FLOATING
C3625 a_12760_n20342.n159 DGND 0.12fF $ **FLOATING
C3626 a_12760_n20342.t41 DGND 1.70fF
C3627 a_12760_n20342.t95 DGND 1.70fF
C3628 a_12760_n20342.n161 DGND 0.12fF $ **FLOATING
C3629 a_12760_n20342.n162 DGND 0.12fF $ **FLOATING
C3630 a_12760_n20342.t72 DGND 1.70fF
C3631 a_12760_n20342.t120 DGND 1.70fF
C3632 a_12760_n20342.n164 DGND 0.12fF $ **FLOATING
C3633 a_12760_n20342.n165 DGND 0.12fF $ **FLOATING
C3634 a_12760_n20342.t88 DGND 1.70fF
C3635 a_12760_n20342.t30 DGND 1.70fF
C3636 a_12760_n20342.n167 DGND 0.12fF $ **FLOATING
C3637 a_12760_n20342.n168 DGND 0.12fF $ **FLOATING
C3638 a_12760_n20342.t79 DGND 1.70fF
C3639 a_12760_n20342.t23 DGND 1.70fF
C3640 a_12760_n20342.n170 DGND 0.12fF $ **FLOATING
C3641 a_12760_n20342.n171 DGND 0.12fF $ **FLOATING
C3642 a_12760_n20342.t73 DGND 1.70fF
C3643 a_12760_n20342.t87 DGND 1.70fF
C3644 a_12760_n20342.n173 DGND 0.12fF $ **FLOATING
C3645 a_12760_n20342.n174 DGND 0.12fF $ **FLOATING
C3646 a_12760_n20342.t20 DGND 1.70fF
C3647 a_12760_n20342.t74 DGND 1.70fF
C3648 a_12760_n20342.n176 DGND 0.12fF $ **FLOATING
C3649 a_12760_n20342.n177 DGND 0.12fF $ **FLOATING
C3650 a_12760_n20342.n178 DGND 1.84fF $ **FLOATING
C3651 a_12760_n20342.t15 DGND 1.70fF
C3652 a_12760_n20342.t77 DGND 1.70fF
C3653 a_12760_n20342.n180 DGND 0.12fF $ **FLOATING
C3654 a_12760_n20342.n181 DGND 0.12fF $ **FLOATING
C3655 a_12760_n20342.t105 DGND 1.70fF
C3656 a_12760_n20342.t21 DGND 1.70fF
C3657 a_12760_n20342.n183 DGND 0.12fF $ **FLOATING
C3658 a_12760_n20342.n184 DGND 0.12fF $ **FLOATING
C3659 a_12760_n20342.n185 DGND 1.26fF $ **FLOATING
C3660 a_12760_n20342.t18 DGND 1.70fF
C3661 a_12760_n20342.t82 DGND 1.70fF
C3662 a_12760_n20342.n187 DGND 0.12fF $ **FLOATING
C3663 a_12760_n20342.n188 DGND 0.12fF $ **FLOATING
C3664 a_12760_n20342.t69 DGND 1.70fF
C3665 a_12760_n20342.t83 DGND 1.70fF
C3666 a_12760_n20342.n190 DGND 0.12fF $ **FLOATING
C3667 a_12760_n20342.n191 DGND 0.12fF $ **FLOATING
C3668 a_12760_n20342.t86 DGND 1.70fF
C3669 a_12760_n20342.t28 DGND 1.70fF
C3670 a_12760_n20342.n193 DGND 0.12fF $ **FLOATING
C3671 a_12760_n20342.n194 DGND 0.12fF $ **FLOATING
C3672 a_12760_n20342.t29 DGND 1.70fF
C3673 a_12760_n20342.t94 DGND 1.70fF
C3674 a_12760_n20342.n196 DGND 0.12fF $ **FLOATING
C3675 a_12760_n20342.n197 DGND 0.12fF $ **FLOATING
C3676 a_12760_n20342.t100 DGND 1.70fF
C3677 a_12760_n20342.t118 DGND 1.70fF
C3678 a_12760_n20342.n199 DGND 0.12fF $ **FLOATING
C3679 a_12760_n20342.n200 DGND 0.12fF $ **FLOATING
C3680 a_12760_n20342.t38 DGND 1.70fF
C3681 a_12760_n20342.t103 DGND 1.70fF
C3682 a_12760_n20342.n202 DGND 0.12fF $ **FLOATING
C3683 a_12760_n20342.n203 DGND 0.12fF $ **FLOATING
C3684 a_12760_n20342.t45 DGND 1.70fF
C3685 a_12760_n20342.t60 DGND 1.70fF
C3686 a_12760_n20342.n205 DGND 0.12fF $ **FLOATING
C3687 a_12760_n20342.n206 DGND 0.12fF $ **FLOATING
C3688 a_12760_n20342.n207 DGND 2.01fF $ **FLOATING
C3689 a_12760_n20342.t110 DGND 1.70fF
C3690 a_12760_n20342.t48 DGND 1.70fF
C3691 a_12760_n20342.n209 DGND 0.12fF $ **FLOATING
C3692 a_12760_n20342.n210 DGND 0.12fF $ **FLOATING
C3693 a_12760_n20342.n211 DGND 1.26fF $ **FLOATING
C3694 a_12760_n20342.t54 DGND 1.70fF
C3695 a_12760_n20342.t65 DGND 1.70fF
C3696 a_12760_n20342.n213 DGND 0.12fF $ **FLOATING
C3697 a_12760_n20342.n214 DGND 0.12fF $ **FLOATING
C3698 a_12760_n20342.t124 DGND 1.70fF
C3699 a_12760_n20342.t7 DGND 1.70fF
C3700 a_12760_n20342.n216 DGND 0.12fF $ **FLOATING
C3701 a_12760_n20342.n217 DGND 0.12fF $ **FLOATING
C3702 a_12760_n20342.t6 DGND 1.70fF
C3703 a_12760_n20342.t17 DGND 1.70fF
C3704 a_12760_n20342.n219 DGND 0.12fF $ **FLOATING
C3705 a_12760_n20342.n220 DGND 0.12fF $ **FLOATING
C3706 a_12760_n20342.t71 DGND 1.70fF
C3707 a_12760_n20342.t85 DGND 1.70fF
C3708 a_12760_n20342.n222 DGND 0.12fF $ **FLOATING
C3709 a_12760_n20342.n223 DGND 0.12fF $ **FLOATING
C3710 a_12760_n20342.n224 DGND 1.26fF $ **FLOATING
C3711 a_12760_n20342.n225 DGND 1.26fF $ **FLOATING
C3712 a_12760_n20342.n226 DGND 1.26fF $ **FLOATING
C3713 a_12760_n20342.t119 DGND 1.70fF
C3714 a_12760_n20342.t58 DGND 1.70fF
C3715 a_12760_n20342.n228 DGND 0.12fF $ **FLOATING
C3716 a_12760_n20342.n229 DGND 0.12fF $ **FLOATING
C3717 a_12760_n20342.t61 DGND 1.70fF
C3718 a_12760_n20342.t127 DGND 1.70fF
C3719 a_12760_n20342.n231 DGND 0.12fF $ **FLOATING
C3720 a_12760_n20342.n232 DGND 0.12fF $ **FLOATING
C3721 a_12760_n20342.t67 DGND 1.70fF
C3722 a_12760_n20342.t8 DGND 1.70fF
C3723 a_12760_n20342.n234 DGND 0.12fF $ **FLOATING
C3724 a_12760_n20342.n235 DGND 0.12fF $ **FLOATING
C3725 a_12760_n20342.n236 DGND 1.84fF $ **FLOATING
C3726 a_12760_n20342.n237 DGND 1.84fF $ **FLOATING
C3727 a_12760_n20342.t104 DGND 1.70fF
C3728 a_12760_n20342.t122 DGND 1.70fF
C3729 a_12760_n20342.n239 DGND 0.12fF $ **FLOATING
C3730 a_12760_n20342.n240 DGND 0.12fF $ **FLOATING
C3731 a_12760_n20342.t49 DGND 1.70fF
C3732 a_12760_n20342.t64 DGND 1.70fF
C3733 a_12760_n20342.n242 DGND 0.12fF $ **FLOATING
C3734 a_12760_n20342.n243 DGND 0.12fF $ **FLOATING
C3735 a_12760_n20342.t63 DGND 1.70fF
C3736 a_12760_n20342.t68 DGND 1.70fF
C3737 a_12760_n20342.n245 DGND 0.12fF $ **FLOATING
C3738 a_12760_n20342.n246 DGND 0.12fF $ **FLOATING
C3739 a_12760_n20342.t12 DGND 1.70fF
C3740 a_12760_n20342.t75 DGND 1.70fF
C3741 a_12760_n20342.n248 DGND 0.12fF $ **FLOATING
C3742 a_12760_n20342.n249 DGND 0.12fF $ **FLOATING
C3743 a_12760_n20342.n250 DGND 2.01fF $ **FLOATING
C3744 a_12760_n20342.t5 DGND 1.70fF
C3745 a_12760_n20342.t16 DGND 1.70fF
C3746 a_12760_n20342.n252 DGND 0.12fF $ **FLOATING
C3747 a_12760_n20342.n253 DGND 0.12fF $ **FLOATING
C3748 a_12760_n20342.n254 DGND 1.52fF $ **FLOATING
C3749 a_12760_n20342.n255 DGND 1.84fF $ **FLOATING
C3750 a_12760_n20342.n256 DGND 1.84fF $ **FLOATING
C3751 a_12760_n20342.t43 DGND 1.70fF
C3752 a_12760_n20342.t59 DGND 1.70fF
C3753 a_12760_n20342.n258 DGND 0.12fF $ **FLOATING
C3754 a_12760_n20342.n259 DGND 0.12fF $ **FLOATING
C3755 a_12760_n20342.t33 DGND 1.70fF
C3756 a_12760_n20342.t96 DGND 1.70fF
C3757 a_12760_n20342.n261 DGND 0.12fF $ **FLOATING
C3758 a_12760_n20342.n262 DGND 0.12fF $ **FLOATING
C3759 a_12760_n20342.t114 DGND 1.70fF
C3760 a_12760_n20342.t128 DGND 1.70fF
C3761 a_12760_n20342.n264 DGND 0.12fF $ **FLOATING
C3762 a_12760_n20342.n265 DGND 0.12fF $ **FLOATING
C3763 a_12760_n20342.t97 DGND 1.70fF
C3764 a_12760_n20342.t40 DGND 1.70fF
C3765 a_12760_n20342.n267 DGND 0.12fF $ **FLOATING
C3766 a_12760_n20342.n268 DGND 0.12fF $ **FLOATING
C3767 a_12760_n20342.t126 DGND 1.70fF
C3768 a_12760_n20342.t9 DGND 1.70fF
C3769 a_12760_n20342.n270 DGND 0.12fF $ **FLOATING
C3770 a_12760_n20342.n271 DGND 0.12fF $ **FLOATING
C3771 a_12760_n20342.t66 DGND 1.70fF
C3772 a_12760_n20342.t76 DGND 1.70fF
C3773 a_12760_n20342.n273 DGND 0.12fF $ **FLOATING
C3774 a_12760_n20342.n274 DGND 0.12fF $ **FLOATING
C3775 a_12760_n20342.n275 DGND 1.52fF $ **FLOATING
C3776 a_12760_n20342.n276 DGND 1.84fF $ **FLOATING
C3777 a_12760_n20342.t113 DGND 1.70fF
C3778 a_12760_n20342.t53 DGND 1.70fF
C3779 a_12760_n20342.n278 DGND 0.12fF $ **FLOATING
C3780 a_12760_n20342.n279 DGND 0.12fF $ **FLOATING
C3781 a_12760_n20342.t57 DGND 1.70fF
C3782 a_12760_n20342.t123 DGND 1.70fF
C3783 a_12760_n20342.n281 DGND 0.12fF $ **FLOATING
C3784 a_12760_n20342.n282 DGND 0.12fF $ **FLOATING
C3785 a_12760_n20342.n283 DGND 1.52fF $ **FLOATING
C3786 a_12760_n20342.n284 DGND 1.84fF $ **FLOATING
C3787 a_12760_n20342.t25 DGND 1.70fF
C3788 a_12760_n20342.t35 DGND 1.70fF
C3789 a_12760_n20342.n286 DGND 0.12fF $ **FLOATING
C3790 a_12760_n20342.n287 DGND 0.12fF $ **FLOATING
C3791 a_12760_n20342.t89 DGND 1.70fF
C3792 a_12760_n20342.t102 DGND 1.70fF
C3793 a_12760_n20342.n289 DGND 0.12fF $ **FLOATING
C3794 a_12760_n20342.n290 DGND 0.12fF $ **FLOATING
C3795 a_12760_n20342.n291 DGND 1.84fF $ **FLOATING
C3796 Vom.n0 DGND 4.83fF $ **FLOATING
C3797 Vom.n1 DGND 5.09fF $ **FLOATING
C3798 Vom.n2 DGND 4.25fF $ **FLOATING
C3799 Vom.n3 DGND 5.09fF $ **FLOATING
C3800 Vom.n4 DGND 4.25fF $ **FLOATING
C3801 Vom.n5 DGND 4.25fF $ **FLOATING
C3802 Vom.n6 DGND 4.83fF $ **FLOATING
C3803 Vom.n7 DGND 4.25fF $ **FLOATING
C3804 Vom.n8 DGND 4.25fF $ **FLOATING
C3805 Vom.n9 DGND 4.25fF $ **FLOATING
C3806 Vom.n10 DGND 4.83fF $ **FLOATING
C3807 Vom.n11 DGND 4.25fF $ **FLOATING
C3808 Vom.n12 DGND 1.39fF $ **FLOATING
C3809 Vom.n13 DGND 1.39fF $ **FLOATING
C3810 Vom.n14 DGND 1.39fF $ **FLOATING
C3811 Vom.n15 DGND 1.39fF $ **FLOATING
C3812 Vom.n16 DGND 1.64fF $ **FLOATING
C3813 Vom.n17 DGND 0.96fF $ **FLOATING
C3814 Vom.n18 DGND 0.70fF $ **FLOATING
C3815 Vom.n19 DGND 1.64fF $ **FLOATING
C3816 Vom.n20 DGND 0.96fF $ **FLOATING
C3817 Vom.n21 DGND 0.70fF $ **FLOATING
C3818 Vom.n22 DGND 1.64fF $ **FLOATING
C3819 Vom.n23 DGND 0.96fF $ **FLOATING
C3820 Vom.n24 DGND 0.70fF $ **FLOATING
C3821 Vom.n25 DGND 1.64fF $ **FLOATING
C3822 Vom.n26 DGND 0.96fF $ **FLOATING
C3823 Vom.n27 DGND 1.25fF $ **FLOATING
C3824 Vom.n28 DGND 1.91fF $ **FLOATING
C3825 Vom.n29 DGND 1.81fF $ **FLOATING
C3826 Vom.n30 DGND 1.81fF $ **FLOATING
C3827 Vom.n31 DGND 1.81fF $ **FLOATING
C3828 Vom.n32 DGND 1.81fF $ **FLOATING
C3829 Vom.n33 DGND 1.81fF $ **FLOATING
C3830 Vom.n34 DGND 1.91fF $ **FLOATING
C3831 Vom.t105 DGND 0.10fF
C3832 Vom.n35 DGND 1.55fF $ **FLOATING
C3833 Vom.t109 DGND 0.10fF
C3834 Vom.n36 DGND 1.69fF $ **FLOATING
C3835 Vom.n37 DGND 1.99fF $ **FLOATING
C3836 Vom.n38 DGND 1.21fF $ **FLOATING
C3837 Vom.n39 DGND 0.87fF $ **FLOATING
C3838 Vom.n40 DGND 1.99fF $ **FLOATING
C3839 Vom.n41 DGND 1.21fF $ **FLOATING
C3840 Vom.n42 DGND 1.40fF $ **FLOATING
C3841 Vom.n43 DGND 1.90fF $ **FLOATING
C3842 Vom.n44 DGND 1.82fF $ **FLOATING
C3843 Vom.n45 DGND 1.53fF $ **FLOATING
C3844 Vom.n46 DGND 0.64fF $ **FLOATING
C3845 Vom.t132 DGND 3.08fF
C3846 Vom.t143 DGND 3.08fF
C3847 Vom.n47 DGND 0.64fF $ **FLOATING
C3848 Vom.t144 DGND 3.08fF
C3849 Vom.t130 DGND 3.08fF
C3850 Vom.n48 DGND 2.50fF $ **FLOATING
C3851 Vom.t124 DGND 1.64fF
C3852 Vom.n49 DGND 25.96fF $ **FLOATING
C3853 Vom.n50 DGND 0.64fF $ **FLOATING
C3854 Vom.t138 DGND 3.08fF
C3855 Vom.t121 DGND 3.08fF
C3856 Vom.n51 DGND 0.64fF $ **FLOATING
C3857 Vom.t122 DGND 3.08fF
C3858 Vom.t135 DGND 3.08fF
C3859 Vom.n52 DGND 0.64fF $ **FLOATING
C3860 Vom.t128 DGND 3.08fF
C3861 Vom.t120 DGND 3.08fF
C3862 Vom.n53 DGND 0.64fF $ **FLOATING
C3863 Vom.t133 DGND 3.08fF
C3864 Vom.t125 DGND 3.08fF
C3865 Vom.n54 DGND 2.50fF $ **FLOATING
C3866 Vom.n55 DGND 2.50fF $ **FLOATING
C3867 Vom.n56 DGND 0.64fF $ **FLOATING
C3868 Vom.t136 DGND 3.08fF
C3869 Vom.t131 DGND 3.08fF
C3870 Vom.n57 DGND 0.64fF $ **FLOATING
C3871 Vom.t140 DGND 3.08fF
C3872 Vom.t134 DGND 3.08fF
C3873 Vom.n58 DGND 5.11fF $ **FLOATING
C3874 Vom.n59 DGND 3.71fF $ **FLOATING
C3875 Vom.n60 DGND 3.71fF $ **FLOATING
C3876 Vom.n61 DGND 3.71fF $ **FLOATING
C3877 Vom.n62 DGND 3.45fF $ **FLOATING
C3878 Vom.n63 DGND 2.88fF $ **FLOATING
C3879 Vom.n64 DGND 0.64fF $ **FLOATING
C3880 Vom.t126 DGND 3.08fF
C3881 Vom.t142 DGND 3.08fF
C3882 Vom.n65 DGND 0.64fF $ **FLOATING
C3883 Vom.t139 DGND 3.08fF
C3884 Vom.t127 DGND 3.08fF
C3885 Vom.n66 DGND 0.64fF $ **FLOATING
C3886 Vom.t123 DGND 3.08fF
C3887 Vom.t137 DGND 3.08fF
C3888 Vom.n67 DGND 0.64fF $ **FLOATING
C3889 Vom.t129 DGND 3.08fF
C3890 Vom.t141 DGND 3.08fF
C3891 Vom.n68 DGND 2.50fF $ **FLOATING
C3892 Vom.n69 DGND 2.50fF $ **FLOATING
C3893 Vom.n70 DGND 2.50fF $ **FLOATING
C3894 Vom.n71 DGND 3.84fF $ **FLOATING
C3895 Vom.n72 DGND 1.37fF $ **FLOATING
C3896 Vom.n73 DGND 1.37fF $ **FLOATING
C3897 Vom.n74 DGND 1.37fF $ **FLOATING
C3898 Vom.n75 DGND 1.18fF $ **FLOATING
C3899 Vom.n76 DGND 1.77fF $ **FLOATING
C3900 Vom.n77 DGND 1.81fF $ **FLOATING
C3901 Vom.n78 DGND 1.91fF $ **FLOATING
C3902 Vom.t116 DGND 0.10fF
C3903 Vom.n79 DGND 1.55fF $ **FLOATING
C3904 Vom.t87 DGND 0.10fF
C3905 Vom.n80 DGND -0.54fF $ **FLOATING
C3906 Vom.n81 DGND 1.17fF $ **FLOATING
C3907 Vom.n82 DGND 1.39fF $ **FLOATING
C3908 Vom.n83 DGND 1.39fF $ **FLOATING
C3909 Vom.n84 DGND 1.39fF $ **FLOATING
C3910 Vom.n85 DGND 1.39fF $ **FLOATING
C3911 Vom.n86 DGND 1.39fF $ **FLOATING
C3912 Vom.n87 DGND 1.39fF $ **FLOATING
C3913 Vom.n88 DGND 1.39fF $ **FLOATING
C3914 Vom.n89 DGND 1.93fF $ **FLOATING
C3915 Vom.n90 DGND 1.91fF $ **FLOATING
C3916 Vom.n91 DGND 1.81fF $ **FLOATING
C3917 Vom.n92 DGND 1.81fF $ **FLOATING
C3918 Vom.n93 DGND 1.81fF $ **FLOATING
C3919 Vom.n94 DGND 1.81fF $ **FLOATING
C3920 Vom.n95 DGND 1.81fF $ **FLOATING
C3921 Vom.n96 DGND 1.91fF $ **FLOATING
C3922 Vom.t110 DGND 0.10fF
C3923 Vom.n97 DGND 1.55fF $ **FLOATING
C3924 Vom.t81 DGND 0.10fF
C3925 Vom.n98 DGND 1.55fF $ **FLOATING
C3926 Vom.t111 DGND 0.10fF
C3927 Vom.n99 DGND 1.55fF $ **FLOATING
C3928 Vom.t101 DGND 0.10fF
C3929 Vom.n100 DGND 2.02fF $ **FLOATING
C3930 Vom.n101 DGND 1.83fF $ **FLOATING
C3931 Vom.n102 DGND 1.76fF $ **FLOATING
C3932 Vom.n103 DGND 1.53fF $ **FLOATING
C3933 Vom.n104 DGND 1.32fF $ **FLOATING
C3934 Vom.n105 DGND 1.32fF $ **FLOATING
C3935 Vom.n106 DGND 1.32fF $ **FLOATING
C3936 Vom.n107 DGND 1.32fF $ **FLOATING
C3937 Vom.n108 DGND 1.32fF $ **FLOATING
C3938 Vom.n109 DGND 1.32fF $ **FLOATING
C3939 Vom.n110 DGND 1.32fF $ **FLOATING
C3940 Vom.n111 DGND 1.86fF $ **FLOATING
C3941 Vom.n112 DGND 1.91fF $ **FLOATING
C3942 Vom.n113 DGND 1.81fF $ **FLOATING
C3943 Vom.n114 DGND 1.81fF $ **FLOATING
C3944 Vom.n115 DGND 1.81fF $ **FLOATING
C3945 Vom.n116 DGND 1.81fF $ **FLOATING
C3946 Vom.n117 DGND 1.81fF $ **FLOATING
C3947 Vom.n118 DGND 1.91fF $ **FLOATING
C3948 Vom.t90 DGND 0.10fF
C3949 Vom.n119 DGND 1.55fF $ **FLOATING
C3950 Vom.t118 DGND 0.10fF
C3951 Vom.n120 DGND 1.55fF $ **FLOATING
C3952 Vom.t91 DGND 0.10fF
C3953 Vom.n121 DGND 1.55fF $ **FLOATING
C3954 Vom.t112 DGND 0.10fF
C3955 Vom.n122 DGND 2.02fF $ **FLOATING
C3956 Vom.n123 DGND 1.83fF $ **FLOATING
C3957 Vom.n124 DGND 1.76fF $ **FLOATING
C3958 Vom.n125 DGND 1.53fF $ **FLOATING
C3959 Vom.n126 DGND 4.36fF $ **FLOATING
C3960 Vom.n127 DGND 6.87fF $ **FLOATING
C3961 Vom.t107 DGND 0.10fF
C3962 Vom.n128 DGND 1.55fF $ **FLOATING
C3963 Vom.t80 DGND 0.10fF
C3964 Vom.n129 DGND 1.55fF $ **FLOATING
C3965 Vom.t108 DGND 0.10fF
C3966 Vom.n130 DGND 1.55fF $ **FLOATING
C3967 Vom.t85 DGND 0.10fF
C3968 Vom.n131 DGND 2.02fF $ **FLOATING
C3969 Vom.n132 DGND 1.83fF $ **FLOATING
C3970 Vom.n133 DGND 1.76fF $ **FLOATING
C3971 Vom.n134 DGND 1.53fF $ **FLOATING
C3972 Vom.n135 DGND 1.39fF $ **FLOATING
C3973 Vom.n136 DGND 1.39fF $ **FLOATING
C3974 Vom.n137 DGND 1.39fF $ **FLOATING
C3975 Vom.n138 DGND 1.39fF $ **FLOATING
C3976 Vom.n139 DGND 1.39fF $ **FLOATING
C3977 Vom.n140 DGND 1.39fF $ **FLOATING
C3978 Vom.n141 DGND 1.93fF $ **FLOATING
C3979 Vom.n142 DGND 1.91fF $ **FLOATING
C3980 Vom.n143 DGND 1.39fF $ **FLOATING
C3981 Vom.n144 DGND 1.81fF $ **FLOATING
C3982 Vom.n145 DGND 1.81fF $ **FLOATING
C3983 Vom.n146 DGND 1.81fF $ **FLOATING
C3984 Vom.n147 DGND 1.81fF $ **FLOATING
C3985 Vom.n148 DGND 1.81fF $ **FLOATING
C3986 Vom.n149 DGND 1.91fF $ **FLOATING
C3987 Vom.n150 DGND 6.87fF $ **FLOATING
C3988 Vom.n151 DGND 4.57fF $ **FLOATING
C3989 a_2458_5328.t18 DGND 0.25fF
C3990 a_2458_5328.t15 DGND 0.25fF
C3991 a_2458_5328.t192 DGND 0.25fF
C3992 a_2458_5328.t40 DGND 0.25fF
C3993 a_2458_5328.t189 DGND 0.25fF
C3994 a_2458_5328.n0 DGND 5.82fF $ **FLOATING
C3995 a_2458_5328.n1 DGND 4.56fF $ **FLOATING
C3996 a_2458_5328.n2 DGND 4.56fF $ **FLOATING
C3997 a_2458_5328.n3 DGND 5.70fF $ **FLOATING
C3998 a_2458_5328.n4 DGND 1.68fF $ **FLOATING
C3999 a_2458_5328.n5 DGND 1.78fF $ **FLOATING
C4000 a_2458_5328.n6 DGND 1.68fF $ **FLOATING
C4001 a_2458_5328.n7 DGND 1.78fF $ **FLOATING
C4002 a_2458_5328.n8 DGND 1.68fF $ **FLOATING
C4003 a_2458_5328.n9 DGND 1.78fF $ **FLOATING
C4004 a_2458_5328.n10 DGND 1.68fF $ **FLOATING
C4005 a_2458_5328.n11 DGND 1.78fF $ **FLOATING
C4006 a_2458_5328.n12 DGND 1.68fF $ **FLOATING
C4007 a_2458_5328.n13 DGND 1.78fF $ **FLOATING
C4008 a_2458_5328.n14 DGND 1.68fF $ **FLOATING
C4009 a_2458_5328.n15 DGND 1.78fF $ **FLOATING
C4010 a_2458_5328.n16 DGND 1.68fF $ **FLOATING
C4011 a_2458_5328.n17 DGND 1.78fF $ **FLOATING
C4012 a_2458_5328.n18 DGND 1.68fF $ **FLOATING
C4013 a_2458_5328.n19 DGND 2.68fF $ **FLOATING
C4014 a_2458_5328.n20 DGND 2.15fF $ **FLOATING
C4015 a_2458_5328.n21 DGND 1.93fF $ **FLOATING
C4016 a_2458_5328.n22 DGND 1.93fF $ **FLOATING
C4017 a_2458_5328.n23 DGND 1.93fF $ **FLOATING
C4018 a_2458_5328.n24 DGND 1.93fF $ **FLOATING
C4019 a_2458_5328.n25 DGND 1.93fF $ **FLOATING
C4020 a_2458_5328.n26 DGND 2.40fF $ **FLOATING
C4021 a_2458_5328.n27 DGND 1.68fF $ **FLOATING
C4022 a_2458_5328.n28 DGND 1.78fF $ **FLOATING
C4023 a_2458_5328.n29 DGND 1.68fF $ **FLOATING
C4024 a_2458_5328.n30 DGND 1.78fF $ **FLOATING
C4025 a_2458_5328.n31 DGND 1.68fF $ **FLOATING
C4026 a_2458_5328.n32 DGND 1.78fF $ **FLOATING
C4027 a_2458_5328.n33 DGND 1.68fF $ **FLOATING
C4028 a_2458_5328.n34 DGND 1.96fF $ **FLOATING
C4029 a_2458_5328.n35 DGND 1.97fF $ **FLOATING
C4030 a_2458_5328.n36 DGND 1.93fF $ **FLOATING
C4031 a_2458_5328.n37 DGND 2.40fF $ **FLOATING
C4032 a_2458_5328.n38 DGND 1.68fF $ **FLOATING
C4033 a_2458_5328.n39 DGND 1.78fF $ **FLOATING
C4034 a_2458_5328.n40 DGND 1.68fF $ **FLOATING
C4035 a_2458_5328.n41 DGND 1.78fF $ **FLOATING
C4036 a_2458_5328.n42 DGND 1.68fF $ **FLOATING
C4037 a_2458_5328.n43 DGND 1.78fF $ **FLOATING
C4038 a_2458_5328.n44 DGND 1.68fF $ **FLOATING
C4039 a_2458_5328.n45 DGND 1.78fF $ **FLOATING
C4040 a_2458_5328.n46 DGND 1.68fF $ **FLOATING
C4041 a_2458_5328.n47 DGND 1.93fF $ **FLOATING
C4042 a_2458_5328.n48 DGND 1.93fF $ **FLOATING
C4043 a_2458_5328.n49 DGND 1.78fF $ **FLOATING
C4044 a_2458_5328.n50 DGND 1.68fF $ **FLOATING
C4045 a_2458_5328.n51 DGND 1.93fF $ **FLOATING
C4046 a_2458_5328.n52 DGND 1.93fF $ **FLOATING
C4047 a_2458_5328.n53 DGND 1.78fF $ **FLOATING
C4048 a_2458_5328.n54 DGND 1.68fF $ **FLOATING
C4049 a_2458_5328.n55 DGND 1.93fF $ **FLOATING
C4050 a_2458_5328.n56 DGND 1.93fF $ **FLOATING
C4051 a_2458_5328.n57 DGND 1.78fF $ **FLOATING
C4052 a_2458_5328.n58 DGND 1.68fF $ **FLOATING
C4053 a_2458_5328.n59 DGND 1.93fF $ **FLOATING
C4054 a_2458_5328.n60 DGND 1.93fF $ **FLOATING
C4055 a_2458_5328.n61 DGND 2.68fF $ **FLOATING
C4056 a_2458_5328.n62 DGND 2.15fF $ **FLOATING
C4057 a_2458_5328.n63 DGND 1.93fF $ **FLOATING
C4058 a_2458_5328.n64 DGND 1.93fF $ **FLOATING
C4059 a_2458_5328.n65 DGND 1.93fF $ **FLOATING
C4060 a_2458_5328.n66 DGND 1.93fF $ **FLOATING
C4061 a_2458_5328.n67 DGND 1.93fF $ **FLOATING
C4062 a_2458_5328.n68 DGND 2.40fF $ **FLOATING
C4063 a_2458_5328.n69 DGND 0.39fF $ **FLOATING
C4064 a_2458_5328.n70 DGND 0.39fF $ **FLOATING
C4065 a_2458_5328.n71 DGND 0.39fF $ **FLOATING
C4066 a_2458_5328.t198 DGND 0.18fF
C4067 a_2458_5328.n72 DGND 1.01fF $ **FLOATING
C4068 a_2458_5328.n73 DGND 0.42fF $ **FLOATING
C4069 a_2458_5328.n74 DGND 0.47fF $ **FLOATING
C4070 a_2458_5328.n75 DGND 10.76fF $ **FLOATING
C4071 a_2458_5328.n76 DGND 21.84fF $ **FLOATING
C4072 a_2458_5328.n77 DGND 6.96fF $ **FLOATING
C4073 a_2458_5328.n78 DGND 5.46fF $ **FLOATING
C4074 a_2458_5328.n79 DGND 1.68fF $ **FLOATING
C4075 a_2458_5328.n80 DGND 1.78fF $ **FLOATING
C4076 a_2458_5328.n81 DGND 1.68fF $ **FLOATING
C4077 a_2458_5328.n82 DGND 1.78fF $ **FLOATING
C4078 a_2458_5328.n83 DGND 1.68fF $ **FLOATING
C4079 a_2458_5328.n84 DGND 1.78fF $ **FLOATING
C4080 a_2458_5328.n85 DGND 1.68fF $ **FLOATING
C4081 a_2458_5328.n86 DGND 1.78fF $ **FLOATING
C4082 a_2458_5328.n87 DGND 1.68fF $ **FLOATING
C4083 a_2458_5328.n88 DGND 1.78fF $ **FLOATING
C4084 a_2458_5328.n89 DGND 1.68fF $ **FLOATING
C4085 a_2458_5328.n90 DGND 1.78fF $ **FLOATING
C4086 a_2458_5328.n91 DGND 1.68fF $ **FLOATING
C4087 a_2458_5328.n92 DGND 1.78fF $ **FLOATING
C4088 a_2458_5328.n93 DGND 1.68fF $ **FLOATING
C4089 a_2458_5328.n94 DGND 2.68fF $ **FLOATING
C4090 a_2458_5328.n95 DGND 2.15fF $ **FLOATING
C4091 a_2458_5328.n96 DGND 1.93fF $ **FLOATING
C4092 a_2458_5328.n97 DGND 1.93fF $ **FLOATING
C4093 a_2458_5328.n98 DGND 1.93fF $ **FLOATING
C4094 a_2458_5328.n99 DGND 1.93fF $ **FLOATING
C4095 a_2458_5328.n100 DGND 1.93fF $ **FLOATING
C4096 a_2458_5328.n101 DGND 2.40fF $ **FLOATING
C4097 a_2458_5328.n102 DGND 1.68fF $ **FLOATING
C4098 a_2458_5328.n103 DGND 1.78fF $ **FLOATING
C4099 a_2458_5328.n104 DGND 1.68fF $ **FLOATING
C4100 a_2458_5328.n105 DGND 1.78fF $ **FLOATING
C4101 a_2458_5328.n106 DGND 1.68fF $ **FLOATING
C4102 a_2458_5328.n107 DGND 1.78fF $ **FLOATING
C4103 a_2458_5328.n108 DGND 1.68fF $ **FLOATING
C4104 a_2458_5328.n109 DGND 1.78fF $ **FLOATING
C4105 a_2458_5328.n110 DGND 1.68fF $ **FLOATING
C4106 a_2458_5328.n111 DGND 1.78fF $ **FLOATING
C4107 a_2458_5328.n112 DGND 1.68fF $ **FLOATING
C4108 a_2458_5328.n113 DGND 1.78fF $ **FLOATING
C4109 a_2458_5328.n114 DGND 1.68fF $ **FLOATING
C4110 a_2458_5328.n115 DGND 1.78fF $ **FLOATING
C4111 a_2458_5328.n116 DGND 1.68fF $ **FLOATING
C4112 a_2458_5328.n117 DGND 2.68fF $ **FLOATING
C4113 a_2458_5328.n118 DGND 2.15fF $ **FLOATING
C4114 a_2458_5328.n119 DGND 1.93fF $ **FLOATING
C4115 a_2458_5328.n120 DGND 1.93fF $ **FLOATING
C4116 a_2458_5328.n121 DGND 1.93fF $ **FLOATING
C4117 a_2458_5328.n122 DGND 1.93fF $ **FLOATING
C4118 a_2458_5328.n123 DGND 1.93fF $ **FLOATING
C4119 a_2458_5328.n124 DGND 2.40fF $ **FLOATING
C4120 a_2458_5328.n125 DGND 26.96fF $ **FLOATING
C4121 a_2458_5328.n126 DGND 5.72fF $ **FLOATING
C4122 a_2458_5328.n127 DGND 12.56fF $ **FLOATING
C4123 a_2458_5328.t16 DGND 0.26fF
C4124 a_2458_5328.t6 DGND 0.26fF
C4125 a_2458_5328.t17 DGND 0.26fF
C4126 a_2458_5328.n128 DGND 7.08fF $ **FLOATING
C4127 a_2458_5328.n129 DGND 7.08fF $ **FLOATING
C4128 a_2458_5328.n130 DGND 4.34fF $ **FLOATING
C4129 a_2458_5328.n131 DGND 10.40fF $ **FLOATING
C4130 a_2458_5328.t19 DGND 0.25fF
C4131 a_2458_5328.t187 DGND 0.25fF
C4132 a_2458_5328.t191 DGND 0.25fF
C4133 a_2458_5328.t14 DGND 0.25fF
C4134 a_2458_5328.n132 DGND 5.82fF $ **FLOATING
C4135 a_2458_5328.n133 DGND 4.56fF $ **FLOATING
C4136 a_2458_5328.n134 DGND 4.56fF $ **FLOATING
C4137 a_2458_5328.n135 DGND 5.70fF $ **FLOATING
C4138 a_2458_5328.n136 DGND 2.48fF $ **FLOATING
C4139 a_2458_5328.t197 DGND 0.25fF
C4140 a_2458_5328.t195 DGND 0.25fF
C4141 a_2458_5328.t42 DGND 0.25fF
C4142 a_2458_5328.n137 DGND 7.02fF $ **FLOATING
C4143 a_2458_5328.n138 DGND 7.02fF $ **FLOATING
C4144 a_2458_5328.n139 DGND 4.30fF $ **FLOATING
C4145 a_2458_5328.n140 DGND 1.41fF $ **FLOATING
C4146 a_2458_5328.t194 DGND 0.25fF
C4147 a_2458_5328.t7 DGND 0.25fF
C4148 a_2458_5328.t188 DGND 0.25fF
C4149 a_2458_5328.t20 DGND 0.25fF
C4150 a_2458_5328.n141 DGND 5.82fF $ **FLOATING
C4151 a_2458_5328.n142 DGND 4.56fF $ **FLOATING
C4152 a_2458_5328.n143 DGND 4.56fF $ **FLOATING
C4153 a_2458_5328.n144 DGND 5.70fF $ **FLOATING
C4154 a_2458_5328.n145 DGND 2.48fF $ **FLOATING
C4155 a_2458_5328.t11 DGND 0.25fF
C4156 a_2458_5328.t41 DGND 0.25fF
C4157 a_2458_5328.t1 DGND 0.25fF
C4158 a_2458_5328.t51 DGND 0.25fF
C4159 a_2458_5328.n146 DGND 5.82fF $ **FLOATING
C4160 a_2458_5328.n147 DGND 4.56fF $ **FLOATING
C4161 a_2458_5328.n148 DGND 4.56fF $ **FLOATING
C4162 a_2458_5328.n149 DGND 5.70fF $ **FLOATING
C4163 a_2458_5328.n150 DGND 2.48fF $ **FLOATING
C4164 a_2458_5328.t10 DGND 0.25fF
C4165 a_2458_5328.t178 DGND 0.25fF
C4166 a_2458_5328.t13 DGND 0.25fF
C4167 a_2458_5328.n151 DGND 7.02fF $ **FLOATING
C4168 a_2458_5328.n152 DGND 7.02fF $ **FLOATING
C4169 a_2458_5328.n153 DGND 4.30fF $ **FLOATING
C4170 a_2458_5328.n154 DGND 1.41fF $ **FLOATING
C4171 a_2458_5328.n155 DGND 3.25fF $ **FLOATING
C4172 a_2458_5328.n156 DGND 4.42fF $ **FLOATING
C4173 a_2458_5328.t185 DGND 0.25fF
C4174 a_2458_5328.t190 DGND 0.25fF
C4175 a_2458_5328.t8 DGND 0.25fF
C4176 a_2458_5328.n157 DGND 4.45fF $ **FLOATING
C4177 a_2458_5328.t9 DGND 0.25fF
C4178 a_2458_5328.n158 DGND 4.45fF $ **FLOATING
C4179 a_2458_5328.t179 DGND 0.26fF
C4180 a_2458_5328.n159 DGND 4.48fF $ **FLOATING
C4181 a_2458_5328.n160 DGND 24.16fF $ **FLOATING
C4182 a_2458_5328.n161 DGND 2.79fF $ **FLOATING
C4183 a_2458_5328.n162 DGND 1.70fF $ **FLOATING
C4184 a_2458_5328.n163 DGND 2.79fF $ **FLOATING
C4185 a_2458_5328.n164 DGND 2.79fF $ **FLOATING
C4186 a_2458_5328.n165 DGND 1.70fF $ **FLOATING
C4187 a_2458_5328.n166 DGND 3.84fF $ **FLOATING
C4188 a_2458_5328.n167 DGND 4.57fF $ **FLOATING
C4189 a_2458_5328.n168 DGND 7.02fF $ **FLOATING
C4190 a_2458_5328.n169 DGND 7.02fF $ **FLOATING
C4191 a_2458_5328.t0 DGND 0.25fF
C4192 casc_p.n0 DGND 3.62fF $ **FLOATING
C4193 casc_p.n1 DGND 0.36fF $ **FLOATING
C4194 casc_p.n2 DGND 0.36fF $ **FLOATING
C4195 casc_p.t283 DGND 0.33fF
C4196 casc_p.t79 DGND 0.30fF
C4197 casc_p.n3 DGND 2.59fF $ **FLOATING
C4198 casc_p.t152 DGND 0.30fF
C4199 casc_p.n4 DGND 1.40fF $ **FLOATING
C4200 casc_p.t286 DGND 0.30fF
C4201 casc_p.n5 DGND 1.40fF $ **FLOATING
C4202 casc_p.t381 DGND 0.30fF
C4203 casc_p.n6 DGND 1.40fF $ **FLOATING
C4204 casc_p.t155 DGND 0.30fF
C4205 casc_p.n7 DGND 1.40fF $ **FLOATING
C4206 casc_p.t240 DGND 0.30fF
C4207 casc_p.n8 DGND 1.39fF $ **FLOATING
C4208 casc_p.t384 DGND 0.30fF
C4209 casc_p.n9 DGND 1.39fF $ **FLOATING
C4210 casc_p.t313 DGND 0.30fF
C4211 casc_p.n10 DGND 1.40fF $ **FLOATING
C4212 casc_p.t127 DGND 0.30fF
C4213 casc_p.n11 DGND 1.40fF $ **FLOATING
C4214 casc_p.t221 DGND 0.30fF
C4215 casc_p.n12 DGND 1.40fF $ **FLOATING
C4216 casc_p.t318 DGND 0.30fF
C4217 casc_p.n13 DGND 1.40fF $ **FLOATING
C4218 casc_p.t78 DGND 0.30fF
C4219 casc_p.n14 DGND 1.40fF $ **FLOATING
C4220 casc_p.t223 DGND 0.30fF
C4221 casc_p.n15 DGND 1.40fF $ **FLOATING
C4222 casc_p.t285 DGND 0.30fF
C4223 casc_p.n16 DGND 1.40fF $ **FLOATING
C4224 casc_p.t80 DGND 0.30fF
C4225 casc_p.n17 DGND 1.40fF $ **FLOATING
C4226 casc_p.t154 DGND 0.30fF
C4227 casc_p.n18 DGND 1.40fF $ **FLOATING
C4228 casc_p.t287 DGND 0.30fF
C4229 casc_p.n19 DGND 1.40fF $ **FLOATING
C4230 casc_p.t382 DGND 0.30fF
C4231 casc_p.n20 DGND 1.40fF $ **FLOATING
C4232 casc_p.t198 DGND 0.30fF
C4233 casc_p.n21 DGND 1.40fF $ **FLOATING
C4234 casc_p.t125 DGND 0.30fF
C4235 casc_p.n22 DGND 1.40fF $ **FLOATING
C4236 casc_p.t242 DGND 0.30fF
C4237 casc_p.n23 DGND 1.40fF $ **FLOATING
C4238 casc_p.t314 DGND 0.30fF
C4239 casc_p.n24 DGND 1.40fF $ **FLOATING
C4240 casc_p.t128 DGND 0.30fF
C4241 casc_p.n25 DGND 1.11fF $ **FLOATING
C4242 casc_p.n26 DGND 1.02fF $ **FLOATING
C4243 casc_p.t319 DGND 0.31fF
C4244 casc_p.n28 DGND 0.82fF $ **FLOATING
C4245 casc_p.t2 DGND 2.84fF
C4246 casc_p.t66 DGND 2.84fF
C4247 casc_p.t64 DGND 2.84fF
C4248 casc_p.t0 DGND 2.84fF
C4249 casc_p.n30 DGND 3.36fF $ **FLOATING
C4250 casc_p.n31 DGND 1.01fF $ **FLOATING
C4251 casc_p.n32 DGND 0.73fF $ **FLOATING
C4252 casc_p.n33 DGND 0.73fF $ **FLOATING
C4253 casc_p.n34 DGND 0.82fF $ **FLOATING
C4254 casc_p.n35 DGND 0.21fF $ **FLOATING
C4255 casc_p.n36 DGND 0.21fF $ **FLOATING
C4256 casc_p.n37 DGND 0.21fF $ **FLOATING
C4257 casc_p.n38 DGND 3.67fF $ **FLOATING
C4258 casc_p.t195 DGND 0.33fF
C4259 casc_p.t378 DGND 0.30fF
C4260 casc_p.n39 DGND 2.60fF $ **FLOATING
C4261 casc_p.t277 DGND 0.30fF
C4262 casc_p.n40 DGND 1.40fF $ **FLOATING
C4263 casc_p.t193 DGND 0.30fF
C4264 casc_p.n41 DGND 1.40fF $ **FLOATING
C4265 casc_p.t99 DGND 0.30fF
C4266 casc_p.n42 DGND 1.40fF $ **FLOATING
C4267 casc_p.t275 DGND 0.30fF
C4268 casc_p.n43 DGND 1.40fF $ **FLOATING
C4269 casc_p.t217 DGND 0.30fF
C4270 casc_p.n44 DGND 1.40fF $ **FLOATING
C4271 casc_p.t73 DGND 0.30fF
C4272 casc_p.n45 DGND 1.40fF $ **FLOATING
C4273 casc_p.t308 DGND 0.30fF
C4274 casc_p.n46 DGND 1.40fF $ **FLOATING
C4275 casc_p.t215 DGND 0.30fF
C4276 casc_p.n47 DGND 1.40fF $ **FLOATING
C4277 casc_p.t119 DGND 0.30fF
C4278 casc_p.n48 DGND 1.39fF $ **FLOATING
C4279 casc_p.t385 DGND 0.30fF
C4280 casc_p.n49 DGND 0.81fF $ **FLOATING
C4281 casc_p.t118 DGND 0.33fF
C4282 casc_p.t94 DGND 0.30fF
C4283 casc_p.n50 DGND 2.60fF $ **FLOATING
C4284 casc_p.t276 DGND 0.30fF
C4285 casc_p.n51 DGND 1.40fF $ **FLOATING
C4286 casc_p.t111 DGND 0.30fF
C4287 casc_p.n52 DGND 1.40fF $ **FLOATING
C4288 casc_p.t307 DGND 0.30fF
C4289 casc_p.n53 DGND 1.40fF $ **FLOATING
C4290 casc_p.t267 DGND 0.30fF
C4291 casc_p.n54 DGND 1.40fF $ **FLOATING
C4292 casc_p.t146 DGND 0.30fF
C4293 casc_p.n55 DGND 1.40fF $ **FLOATING
C4294 casc_p.t108 DGND 0.30fF
C4295 casc_p.n56 DGND 1.40fF $ **FLOATING
C4296 casc_p.t302 DGND 0.30fF
C4297 casc_p.n57 DGND 1.40fF $ **FLOATING
C4298 casc_p.t132 DGND 0.30fF
C4299 casc_p.n58 DGND 1.40fF $ **FLOATING
C4300 casc_p.t336 DGND 0.30fF
C4301 casc_p.n59 DGND 1.39fF $ **FLOATING
C4302 casc_p.t252 DGND 0.30fF
C4303 casc_p.n60 DGND 0.81fF $ **FLOATING
C4304 casc_p.t292 DGND 0.33fF
C4305 casc_p.t145 DGND 0.30fF
C4306 casc_p.n61 DGND 2.59fF $ **FLOATING
C4307 casc_p.t266 DGND 0.30fF
C4308 casc_p.n62 DGND 1.40fF $ **FLOATING
C4309 casc_p.t304 DGND 0.30fF
C4310 casc_p.n63 DGND 1.40fF $ **FLOATING
C4311 casc_p.t109 DGND 0.30fF
C4312 casc_p.n64 DGND 1.40fF $ **FLOATING
C4313 casc_p.t274 DGND 0.30fF
C4314 casc_p.n65 DGND 1.40fF $ **FLOATING
C4315 casc_p.t93 DGND 0.30fF
C4316 casc_p.n66 DGND 1.39fF $ **FLOATING
C4317 casc_p.t116 DGND 0.30fF
C4318 casc_p.n67 DGND 1.39fF $ **FLOATING
C4319 casc_p.t394 DGND 0.30fF
C4320 casc_p.n68 DGND 1.40fF $ **FLOATING
C4321 casc_p.t95 DGND 0.30fF
C4322 casc_p.n69 DGND 1.40fF $ **FLOATING
C4323 casc_p.t232 DGND 0.30fF
C4324 casc_p.n70 DGND 1.40fF $ **FLOATING
C4325 casc_p.t81 DGND 0.30fF
C4326 casc_p.n71 DGND 1.40fF $ **FLOATING
C4327 casc_p.t212 DGND 0.30fF
C4328 casc_p.n72 DGND 1.40fF $ **FLOATING
C4329 casc_p.t243 DGND 0.30fF
C4330 casc_p.n73 DGND 1.40fF $ **FLOATING
C4331 casc_p.t375 DGND 0.30fF
C4332 casc_p.n74 DGND 1.40fF $ **FLOATING
C4333 casc_p.t224 DGND 0.30fF
C4334 casc_p.n75 DGND 1.40fF $ **FLOATING
C4335 casc_p.t356 DGND 0.30fF
C4336 casc_p.n76 DGND 1.40fF $ **FLOATING
C4337 casc_p.t388 DGND 0.30fF
C4338 casc_p.n77 DGND 1.40fF $ **FLOATING
C4339 casc_p.t192 DGND 0.30fF
C4340 casc_p.n78 DGND 1.40fF $ **FLOATING
C4341 casc_p.t225 DGND 0.30fF
C4342 casc_p.n79 DGND 1.40fF $ **FLOATING
C4343 casc_p.t157 DGND 0.30fF
C4344 casc_p.n80 DGND 1.40fF $ **FLOATING
C4345 casc_p.t333 DGND 0.30fF
C4346 casc_p.n81 DGND 1.40fF $ **FLOATING
C4347 casc_p.t126 DGND 0.30fF
C4348 casc_p.n82 DGND 1.40fF $ **FLOATING
C4349 casc_p.t172 DGND 0.30fF
C4350 casc_p.n83 DGND 1.40fF $ **FLOATING
C4351 casc_p.t290 DGND 0.30fF
C4352 casc_p.n84 DGND 1.40fF $ **FLOATING
C4353 casc_p.t141 DGND 0.30fF
C4354 casc_p.n85 DGND 1.11fF $ **FLOATING
C4355 casc_p.n86 DGND 0.94fF $ **FLOATING
C4356 casc_p.n87 DGND 0.68fF $ **FLOATING
C4357 casc_p.t28 DGND 0.30fF
C4358 casc_p.n88 DGND 0.51fF $ **FLOATING
C4359 casc_p.n89 DGND 0.51fF $ **FLOATING
C4360 casc_p.n90 DGND 0.68fF $ **FLOATING
C4361 casc_p.t16 DGND 0.30fF
C4362 casc_p.n91 DGND 0.66fF $ **FLOATING
C4363 casc_p.n92 DGND 0.65fF $ **FLOATING
C4364 casc_p.n93 DGND 0.68fF $ **FLOATING
C4365 casc_p.t58 DGND 0.30fF
C4366 casc_p.n94 DGND 0.51fF $ **FLOATING
C4367 casc_p.n95 DGND 0.51fF $ **FLOATING
C4368 casc_p.n96 DGND 0.68fF $ **FLOATING
C4369 casc_p.t43 DGND 0.30fF
C4370 casc_p.n97 DGND 0.66fF $ **FLOATING
C4371 casc_p.n98 DGND 0.65fF $ **FLOATING
C4372 casc_p.n99 DGND 0.68fF $ **FLOATING
C4373 casc_p.t25 DGND 0.30fF
C4374 casc_p.n100 DGND 0.51fF $ **FLOATING
C4375 casc_p.n101 DGND 0.51fF $ **FLOATING
C4376 casc_p.n102 DGND 0.68fF $ **FLOATING
C4377 casc_p.t55 DGND 0.30fF
C4378 casc_p.n103 DGND 0.60fF $ **FLOATING
C4379 casc_p.t298 DGND 0.33fF
C4380 casc_p.t263 DGND 0.30fF
C4381 casc_p.n104 DGND 2.60fF $ **FLOATING
C4382 casc_p.t140 DGND 0.30fF
C4383 casc_p.n105 DGND 1.40fF $ **FLOATING
C4384 casc_p.t289 DGND 0.30fF
C4385 casc_p.n106 DGND 1.40fF $ **FLOATING
C4386 casc_p.t171 DGND 0.30fF
C4387 casc_p.n107 DGND 1.40fF $ **FLOATING
C4388 casc_p.t124 DGND 0.30fF
C4389 casc_p.n108 DGND 1.40fF $ **FLOATING
C4390 casc_p.t332 DGND 0.30fF
C4391 casc_p.n109 DGND 1.40fF $ **FLOATING
C4392 casc_p.t282 DGND 0.30fF
C4393 casc_p.n110 DGND 1.40fF $ **FLOATING
C4394 casc_p.t168 DGND 0.30fF
C4395 casc_p.n111 DGND 1.40fF $ **FLOATING
C4396 casc_p.t311 DGND 0.30fF
C4397 casc_p.n112 DGND 1.40fF $ **FLOATING
C4398 casc_p.t190 DGND 0.30fF
C4399 casc_p.n113 DGND 1.39fF $ **FLOATING
C4400 casc_p.t100 DGND 0.30fF
C4401 casc_p.n114 DGND 0.81fF $ **FLOATING
C4402 casc_p.t151 DGND 0.33fF
C4403 casc_p.t330 DGND 0.30fF
C4404 casc_p.n115 DGND 2.59fF $ **FLOATING
C4405 casc_p.t122 DGND 0.30fF
C4406 casc_p.n116 DGND 1.40fF $ **FLOATING
C4407 casc_p.t170 DGND 0.30fF
C4408 casc_p.n117 DGND 1.40fF $ **FLOATING
C4409 casc_p.t284 DGND 0.30fF
C4410 casc_p.n118 DGND 1.40fF $ **FLOATING
C4411 casc_p.t138 DGND 0.30fF
C4412 casc_p.n119 DGND 1.40fF $ **FLOATING
C4413 casc_p.t262 DGND 0.30fF
C4414 casc_p.n120 DGND 1.39fF $ **FLOATING
C4415 casc_p.t297 DGND 0.30fF
C4416 casc_p.n121 DGND 1.39fF $ **FLOATING
C4417 casc_p.t245 DGND 0.30fF
C4418 casc_p.n122 DGND 1.40fF $ **FLOATING
C4419 casc_p.t264 DGND 0.30fF
C4420 casc_p.n123 DGND 1.40fF $ **FLOATING
C4421 casc_p.t84 DGND 0.30fF
C4422 casc_p.n124 DGND 1.40fF $ **FLOATING
C4423 casc_p.t251 DGND 0.30fF
C4424 casc_p.n125 DGND 1.40fF $ **FLOATING
C4425 casc_p.t391 DGND 0.30fF
C4426 casc_p.n126 DGND 1.40fF $ **FLOATING
C4427 casc_p.t91 DGND 0.30fF
C4428 casc_p.n127 DGND 1.40fF $ **FLOATING
C4429 casc_p.t228 DGND 0.30fF
C4430 casc_p.n128 DGND 1.40fF $ **FLOATING
C4431 casc_p.t72 DGND 0.30fF
C4432 casc_p.n129 DGND 1.40fF $ **FLOATING
C4433 casc_p.t207 DGND 0.30fF
C4434 casc_p.n130 DGND 1.40fF $ **FLOATING
C4435 casc_p.t236 DGND 0.30fF
C4436 casc_p.n131 DGND 1.40fF $ **FLOATING
C4437 casc_p.t367 DGND 0.30fF
C4438 casc_p.n132 DGND 1.40fF $ **FLOATING
C4439 casc_p.t75 DGND 0.30fF
C4440 casc_p.n133 DGND 1.40fF $ **FLOATING
C4441 casc_p.t338 DGND 0.30fF
C4442 casc_p.n134 DGND 1.40fF $ **FLOATING
C4443 casc_p.t187 DGND 0.30fF
C4444 casc_p.n135 DGND 1.40fF $ **FLOATING
C4445 casc_p.t305 DGND 0.30fF
C4446 casc_p.n136 DGND 1.40fF $ **FLOATING
C4447 casc_p.t350 DGND 0.30fF
C4448 casc_p.n137 DGND 1.40fF $ **FLOATING
C4449 casc_p.t147 DGND 0.30fF
C4450 casc_p.n138 DGND 1.40fF $ **FLOATING
C4451 casc_p.t322 DGND 0.30fF
C4452 casc_p.n139 DGND 1.40fF $ **FLOATING
C4453 casc_p.t115 DGND 0.30fF
C4454 casc_p.n140 DGND 1.40fF $ **FLOATING
C4455 casc_p.t161 DGND 0.30fF
C4456 casc_p.n141 DGND 1.40fF $ **FLOATING
C4457 casc_p.t278 DGND 0.30fF
C4458 casc_p.n142 DGND 1.40fF $ **FLOATING
C4459 casc_p.t325 DGND 0.30fF
C4460 casc_p.n143 DGND 1.11fF $ **FLOATING
C4461 casc_p.n144 DGND 0.94fF $ **FLOATING
C4462 casc_p.n145 DGND 0.68fF $ **FLOATING
C4463 casc_p.t52 DGND 0.30fF
C4464 casc_p.n146 DGND 0.51fF $ **FLOATING
C4465 casc_p.n147 DGND 0.51fF $ **FLOATING
C4466 casc_p.n148 DGND 0.68fF $ **FLOATING
C4467 casc_p.t19 DGND 0.30fF
C4468 casc_p.n149 DGND 0.60fF $ **FLOATING
C4469 casc_p.t139 DGND 0.33fF
C4470 casc_p.t104 DGND 0.30fF
C4471 casc_p.n150 DGND 2.60fF $ **FLOATING
C4472 casc_p.t295 DGND 0.30fF
C4473 casc_p.n151 DGND 1.40fF $ **FLOATING
C4474 casc_p.t123 DGND 0.30fF
C4475 casc_p.n152 DGND 1.40fF $ **FLOATING
C4476 casc_p.t331 DGND 0.30fF
C4477 casc_p.n153 DGND 1.40fF $ **FLOATING
C4478 casc_p.t281 DGND 0.30fF
C4479 casc_p.n154 DGND 1.40fF $ **FLOATING
C4480 casc_p.t167 DGND 0.30fF
C4481 casc_p.n155 DGND 1.40fF $ **FLOATING
C4482 casc_p.t120 DGND 0.30fF
C4483 casc_p.n156 DGND 1.40fF $ **FLOATING
C4484 casc_p.t327 DGND 0.30fF
C4485 casc_p.n157 DGND 1.40fF $ **FLOATING
C4486 casc_p.t150 DGND 0.30fF
C4487 casc_p.n158 DGND 1.40fF $ **FLOATING
C4488 casc_p.t354 DGND 0.30fF
C4489 casc_p.n159 DGND 1.39fF $ **FLOATING
C4490 casc_p.t259 DGND 0.30fF
C4491 casc_p.n160 DGND 0.81fF $ **FLOATING
C4492 casc_p.t309 DGND 0.33fF
C4493 casc_p.t165 DGND 0.30fF
C4494 casc_p.n161 DGND 2.59fF $ **FLOATING
C4495 casc_p.t280 DGND 0.30fF
C4496 casc_p.n162 DGND 1.40fF $ **FLOATING
C4497 casc_p.t328 DGND 0.30fF
C4498 casc_p.n163 DGND 1.40fF $ **FLOATING
C4499 casc_p.t121 DGND 0.30fF
C4500 casc_p.n164 DGND 1.40fF $ **FLOATING
C4501 casc_p.t294 DGND 0.30fF
C4502 casc_p.n165 DGND 1.40fF $ **FLOATING
C4503 casc_p.t103 DGND 0.30fF
C4504 casc_p.n166 DGND 1.39fF $ **FLOATING
C4505 casc_p.t136 DGND 0.30fF
C4506 casc_p.n167 DGND 1.39fF $ **FLOATING
C4507 casc_p.t83 DGND 0.30fF
C4508 casc_p.n168 DGND 1.40fF $ **FLOATING
C4509 casc_p.t105 DGND 0.30fF
C4510 casc_p.n169 DGND 1.40fF $ **FLOATING
C4511 casc_p.t244 DGND 0.30fF
C4512 casc_p.n170 DGND 1.40fF $ **FLOATING
C4513 casc_p.t90 DGND 0.30fF
C4514 casc_p.n171 DGND 1.40fF $ **FLOATING
C4515 casc_p.t227 DGND 0.30fF
C4516 casc_p.n172 DGND 1.40fF $ **FLOATING
C4517 casc_p.t250 DGND 0.30fF
C4518 casc_p.n173 DGND 1.40fF $ **FLOATING
C4519 casc_p.t390 DGND 0.30fF
C4520 casc_p.n174 DGND 1.40fF $ **FLOATING
C4521 casc_p.t234 DGND 0.30fF
C4522 casc_p.n175 DGND 1.40fF $ **FLOATING
C4523 casc_p.t366 DGND 0.30fF
C4524 casc_p.n176 DGND 1.40fF $ **FLOATING
C4525 casc_p.t71 DGND 0.30fF
C4526 casc_p.n177 DGND 1.40fF $ **FLOATING
C4527 casc_p.t206 DGND 0.30fF
C4528 casc_p.n178 DGND 1.40fF $ **FLOATING
C4529 casc_p.t235 DGND 0.30fF
C4530 casc_p.n179 DGND 1.40fF $ **FLOATING
C4531 casc_p.t174 DGND 0.30fF
C4532 casc_p.n180 DGND 1.40fF $ **FLOATING
C4533 casc_p.t348 DGND 0.30fF
C4534 casc_p.n181 DGND 1.40fF $ **FLOATING
C4535 casc_p.t144 DGND 0.30fF
C4536 casc_p.n182 DGND 1.40fF $ **FLOATING
C4537 casc_p.t186 DGND 0.30fF
C4538 casc_p.n183 DGND 1.40fF $ **FLOATING
C4539 casc_p.t303 DGND 0.30fF
C4540 casc_p.n184 DGND 1.40fF $ **FLOATING
C4541 casc_p.t159 DGND 0.30fF
C4542 casc_p.n185 DGND 1.40fF $ **FLOATING
C4543 casc_p.t273 DGND 0.30fF
C4544 casc_p.n186 DGND 1.40fF $ **FLOATING
C4545 casc_p.t321 DGND 0.30fF
C4546 casc_p.n187 DGND 1.40fF $ **FLOATING
C4547 casc_p.t114 DGND 0.30fF
C4548 casc_p.n188 DGND 1.40fF $ **FLOATING
C4549 casc_p.t160 DGND 0.30fF
C4550 casc_p.n189 DGND 1.11fF $ **FLOATING
C4551 casc_p.n190 DGND 0.94fF $ **FLOATING
C4552 casc_p.n191 DGND 0.68fF $ **FLOATING
C4553 casc_p.t22 DGND 0.30fF
C4554 casc_p.n192 DGND 0.51fF $ **FLOATING
C4555 casc_p.n193 DGND 0.51fF $ **FLOATING
C4556 casc_p.n194 DGND 0.68fF $ **FLOATING
C4557 casc_p.t49 DGND 0.30fF
C4558 casc_p.n195 DGND 0.60fF $ **FLOATING
C4559 casc_p.t320 DGND 0.33fF
C4560 casc_p.t271 DGND 0.30fF
C4561 casc_p.n196 DGND 2.60fF $ **FLOATING
C4562 casc_p.t156 DGND 0.30fF
C4563 casc_p.n197 DGND 1.40fF $ **FLOATING
C4564 casc_p.t301 DGND 0.30fF
C4565 casc_p.n198 DGND 1.40fF $ **FLOATING
C4566 casc_p.t185 DGND 0.30fF
C4567 casc_p.n199 DGND 1.40fF $ **FLOATING
C4568 casc_p.t143 DGND 0.30fF
C4569 casc_p.n200 DGND 1.40fF $ **FLOATING
C4570 casc_p.t346 DGND 0.30fF
C4571 casc_p.n201 DGND 1.40fF $ **FLOATING
C4572 casc_p.t299 DGND 0.30fF
C4573 casc_p.n202 DGND 1.40fF $ **FLOATING
C4574 casc_p.t181 DGND 0.30fF
C4575 casc_p.n203 DGND 1.40fF $ **FLOATING
C4576 casc_p.t334 DGND 0.30fF
C4577 casc_p.n204 DGND 1.40fF $ **FLOATING
C4578 casc_p.t203 DGND 0.30fF
C4579 casc_p.n205 DGND 1.39fF $ **FLOATING
C4580 casc_p.t112 DGND 0.30fF
C4581 casc_p.n206 DGND 0.81fF $ **FLOATING
C4582 casc_p.t173 DGND 0.33fF
C4583 casc_p.t344 DGND 0.30fF
C4584 casc_p.n207 DGND 2.59fF $ **FLOATING
C4585 casc_p.t142 DGND 0.30fF
C4586 casc_p.n208 DGND 1.40fF $ **FLOATING
C4587 casc_p.t183 DGND 0.30fF
C4588 casc_p.n209 DGND 1.40fF $ **FLOATING
C4589 casc_p.t300 DGND 0.30fF
C4590 casc_p.n210 DGND 1.40fF $ **FLOATING
C4591 casc_p.t153 DGND 0.30fF
C4592 casc_p.n211 DGND 1.40fF $ **FLOATING
C4593 casc_p.t270 DGND 0.30fF
C4594 casc_p.n212 DGND 1.40fF $ **FLOATING
C4595 casc_p.t316 DGND 0.30fF
C4596 casc_p.n213 DGND 1.40fF $ **FLOATING
C4597 casc_p.t254 DGND 0.30fF
C4598 casc_p.n214 DGND 1.40fF $ **FLOATING
C4599 casc_p.t272 DGND 0.30fF
C4600 casc_p.n215 DGND 1.40fF $ **FLOATING
C4601 casc_p.t92 DGND 0.30fF
C4602 casc_p.n216 DGND 1.40fF $ **FLOATING
C4603 casc_p.t258 DGND 0.30fF
C4604 casc_p.n217 DGND 1.40fF $ **FLOATING
C4605 casc_p.t77 DGND 0.30fF
C4606 casc_p.n218 DGND 1.40fF $ **FLOATING
C4607 casc_p.t98 DGND 0.30fF
C4608 casc_p.n219 DGND 1.40fF $ **FLOATING
C4609 casc_p.t241 DGND 0.30fF
C4610 casc_p.n220 DGND 1.40fF $ **FLOATING
C4611 casc_p.t86 DGND 0.30fF
C4612 casc_p.n221 DGND 1.40fF $ **FLOATING
C4613 casc_p.t220 DGND 0.30fF
C4614 casc_p.n222 DGND 1.40fF $ **FLOATING
C4615 casc_p.t247 DGND 0.30fF
C4616 casc_p.n223 DGND 1.40fF $ **FLOATING
C4617 casc_p.t387 DGND 0.30fF
C4618 casc_p.n224 DGND 1.40fF $ **FLOATING
C4619 casc_p.t87 DGND 0.30fF
C4620 casc_p.n225 DGND 1.40fF $ **FLOATING
C4621 casc_p.t355 DGND 0.30fF
C4622 casc_p.n226 DGND 1.40fF $ **FLOATING
C4623 casc_p.t201 DGND 0.30fF
C4624 casc_p.n227 DGND 1.40fF $ **FLOATING
C4625 casc_p.t329 DGND 0.30fF
C4626 casc_p.n228 DGND 1.40fF $ **FLOATING
C4627 casc_p.t364 DGND 0.30fF
C4628 casc_p.n229 DGND 1.40fF $ **FLOATING
C4629 casc_p.t169 DGND 0.30fF
C4630 casc_p.n230 DGND 1.40fF $ **FLOATING
C4631 casc_p.t340 DGND 0.30fF
C4632 casc_p.n231 DGND 1.40fF $ **FLOATING
C4633 casc_p.t137 DGND 0.30fF
C4634 casc_p.n232 DGND 1.40fF $ **FLOATING
C4635 casc_p.t178 DGND 0.30fF
C4636 casc_p.n233 DGND 1.40fF $ **FLOATING
C4637 casc_p.t296 DGND 0.30fF
C4638 casc_p.n234 DGND 1.40fF $ **FLOATING
C4639 casc_p.t341 DGND 0.30fF
C4640 casc_p.n235 DGND 1.11fF $ **FLOATING
C4641 casc_p.n236 DGND 0.94fF $ **FLOATING
C4642 casc_p.n237 DGND 0.68fF $ **FLOATING
C4643 casc_p.t46 DGND 0.30fF
C4644 casc_p.n238 DGND 0.51fF $ **FLOATING
C4645 casc_p.n239 DGND 0.51fF $ **FLOATING
C4646 casc_p.n240 DGND 0.68fF $ **FLOATING
C4647 casc_p.t13 DGND 0.30fF
C4648 casc_p.n241 DGND 0.60fF $ **FLOATING
C4649 casc_p.t177 DGND 0.33fF
C4650 casc_p.t133 DGND 0.30fF
C4651 casc_p.n242 DGND 2.60fF $ **FLOATING
C4652 casc_p.t337 DGND 0.30fF
C4653 casc_p.n243 DGND 1.40fF $ **FLOATING
C4654 casc_p.t166 DGND 0.30fF
C4655 casc_p.n244 DGND 1.40fF $ **FLOATING
C4656 casc_p.t363 DGND 0.30fF
C4657 casc_p.n245 DGND 1.40fF $ **FLOATING
C4658 casc_p.t326 DGND 0.30fF
C4659 casc_p.n246 DGND 1.40fF $ **FLOATING
C4660 casc_p.t199 DGND 0.30fF
C4661 casc_p.n247 DGND 1.40fF $ **FLOATING
C4662 casc_p.t162 DGND 0.30fF
C4663 casc_p.n248 DGND 1.40fF $ **FLOATING
C4664 casc_p.t360 DGND 0.30fF
C4665 casc_p.n249 DGND 1.40fF $ **FLOATING
C4666 casc_p.t188 DGND 0.30fF
C4667 casc_p.n250 DGND 1.40fF $ **FLOATING
C4668 casc_p.t383 DGND 0.30fF
C4669 casc_p.n251 DGND 1.39fF $ **FLOATING
C4670 casc_p.t291 DGND 0.30fF
C4671 casc_p.n252 DGND 0.81fF $ **FLOATING
C4672 casc_p.t353 DGND 0.33fF
C4673 casc_p.t197 DGND 0.30fF
C4674 casc_p.n253 DGND 2.59fF $ **FLOATING
C4675 casc_p.t324 DGND 0.30fF
C4676 casc_p.n254 DGND 1.40fF $ **FLOATING
C4677 casc_p.t361 DGND 0.30fF
C4678 casc_p.n255 DGND 1.40fF $ **FLOATING
C4679 casc_p.t164 DGND 0.30fF
C4680 casc_p.n256 DGND 1.40fF $ **FLOATING
C4681 casc_p.t335 DGND 0.30fF
C4682 casc_p.n257 DGND 1.40fF $ **FLOATING
C4683 casc_p.t131 DGND 0.30fF
C4684 casc_p.n258 DGND 1.40fF $ **FLOATING
C4685 casc_p.t176 DGND 0.30fF
C4686 casc_p.n259 DGND 1.40fF $ **FLOATING
C4687 casc_p.t102 DGND 0.30fF
C4688 casc_p.n260 DGND 1.40fF $ **FLOATING
C4689 casc_p.t135 DGND 0.30fF
C4690 casc_p.n261 DGND 1.40fF $ **FLOATING
C4691 casc_p.t261 DGND 0.30fF
C4692 casc_p.n262 DGND 1.40fF $ **FLOATING
C4693 casc_p.t110 DGND 0.30fF
C4694 casc_p.n263 DGND 1.40fF $ **FLOATING
C4695 casc_p.t249 DGND 0.30fF
C4696 casc_p.n264 DGND 1.40fF $ **FLOATING
C4697 casc_p.t268 DGND 0.30fF
C4698 casc_p.n265 DGND 1.40fF $ **FLOATING
C4699 casc_p.t89 DGND 0.30fF
C4700 casc_p.n266 DGND 1.40fF $ **FLOATING
C4701 casc_p.t255 DGND 0.30fF
C4702 casc_p.n267 DGND 1.40fF $ **FLOATING
C4703 casc_p.t70 DGND 0.30fF
C4704 casc_p.n268 DGND 1.40fF $ **FLOATING
C4705 casc_p.t96 DGND 0.30fF
C4706 casc_p.n269 DGND 1.40fF $ **FLOATING
C4707 casc_p.t233 DGND 0.30fF
C4708 casc_p.n270 DGND 1.40fF $ **FLOATING
C4709 casc_p.t256 DGND 0.30fF
C4710 casc_p.n271 DGND 1.40fF $ **FLOATING
C4711 casc_p.t205 DGND 0.30fF
C4712 casc_p.n272 DGND 1.40fF $ **FLOATING
C4713 casc_p.t377 DGND 0.30fF
C4714 casc_p.n273 DGND 1.40fF $ **FLOATING
C4715 casc_p.t184 DGND 0.30fF
C4716 casc_p.n274 DGND 1.40fF $ **FLOATING
C4717 casc_p.t216 DGND 0.30fF
C4718 casc_p.n275 DGND 1.40fF $ **FLOATING
C4719 casc_p.t347 DGND 0.30fF
C4720 casc_p.n276 DGND 1.40fF $ **FLOATING
C4721 casc_p.t194 DGND 0.30fF
C4722 casc_p.n277 DGND 1.40fF $ **FLOATING
C4723 casc_p.t317 DGND 0.30fF
C4724 casc_p.n278 DGND 1.40fF $ **FLOATING
C4725 casc_p.t359 DGND 0.30fF
C4726 casc_p.n279 DGND 1.40fF $ **FLOATING
C4727 casc_p.t158 DGND 0.30fF
C4728 casc_p.n280 DGND 1.40fF $ **FLOATING
C4729 casc_p.t196 DGND 0.30fF
C4730 casc_p.n281 DGND 1.11fF $ **FLOATING
C4731 casc_p.n282 DGND 0.94fF $ **FLOATING
C4732 casc_p.n283 DGND 0.68fF $ **FLOATING
C4733 casc_p.t10 DGND 0.30fF
C4734 casc_p.n284 DGND 0.51fF $ **FLOATING
C4735 casc_p.n285 DGND 0.51fF $ **FLOATING
C4736 casc_p.n286 DGND 0.68fF $ **FLOATING
C4737 casc_p.t40 DGND 0.30fF
C4738 casc_p.n287 DGND 0.59fF $ **FLOATING
C4739 casc_p.t358 DGND 0.33fF
C4740 casc_p.t312 DGND 0.30fF
C4741 casc_p.n288 DGND 2.60fF $ **FLOATING
C4742 casc_p.t191 DGND 0.30fF
C4743 casc_p.n289 DGND 1.40fF $ **FLOATING
C4744 casc_p.t345 DGND 0.30fF
C4745 casc_p.n290 DGND 1.40fF $ **FLOATING
C4746 casc_p.t214 DGND 0.30fF
C4747 casc_p.n291 DGND 1.40fF $ **FLOATING
C4748 casc_p.t180 DGND 0.30fF
C4749 casc_p.n292 DGND 1.40fF $ **FLOATING
C4750 casc_p.t374 DGND 0.30fF
C4751 casc_p.n293 DGND 1.40fF $ **FLOATING
C4752 casc_p.t342 DGND 0.30fF
C4753 casc_p.n294 DGND 1.40fF $ **FLOATING
C4754 casc_p.t211 DGND 0.30fF
C4755 casc_p.n295 DGND 1.40fF $ **FLOATING
C4756 casc_p.t365 DGND 0.30fF
C4757 casc_p.n296 DGND 1.40fF $ **FLOATING
C4758 casc_p.t231 DGND 0.30fF
C4759 casc_p.n297 DGND 1.39fF $ **FLOATING
C4760 casc_p.t148 DGND 0.30fF
C4761 casc_p.n298 DGND 0.81fF $ **FLOATING
C4762 casc_p.t202 DGND 0.33fF
C4763 casc_p.t373 DGND 0.30fF
C4764 casc_p.n299 DGND 2.59fF $ **FLOATING
C4765 casc_p.t179 DGND 0.30fF
C4766 casc_p.n300 DGND 1.40fF $ **FLOATING
C4767 casc_p.t213 DGND 0.30fF
C4768 casc_p.n301 DGND 1.40fF $ **FLOATING
C4769 casc_p.t343 DGND 0.30fF
C4770 casc_p.n302 DGND 1.40fF $ **FLOATING
C4771 casc_p.t189 DGND 0.30fF
C4772 casc_p.n303 DGND 1.40fF $ **FLOATING
C4773 casc_p.t310 DGND 0.30fF
C4774 casc_p.n304 DGND 1.40fF $ **FLOATING
C4775 casc_p.t357 DGND 0.30fF
C4776 casc_p.n305 DGND 1.40fF $ **FLOATING
C4777 casc_p.t269 DGND 0.30fF
C4778 casc_p.n306 DGND 1.40fF $ **FLOATING
C4779 casc_p.t315 DGND 0.30fF
C4780 casc_p.n307 DGND 1.40fF $ **FLOATING
C4781 casc_p.t113 DGND 0.30fF
C4782 casc_p.n308 DGND 1.40fF $ **FLOATING
C4783 casc_p.t288 DGND 0.30fF
C4784 casc_p.n309 DGND 1.40fF $ **FLOATING
C4785 casc_p.t97 DGND 0.30fF
C4786 casc_p.n310 DGND 1.40fF $ **FLOATING
C4787 casc_p.t129 DGND 0.30fF
C4788 casc_p.n311 DGND 1.40fF $ **FLOATING
C4789 casc_p.t257 DGND 0.30fF
C4790 casc_p.n312 DGND 1.40fF $ **FLOATING
C4791 casc_p.t106 DGND 0.30fF
C4792 casc_p.n313 DGND 1.40fF $ **FLOATING
C4793 casc_p.t246 DGND 0.30fF
C4794 casc_p.n314 DGND 1.40fF $ **FLOATING
C4795 casc_p.t265 DGND 0.30fF
C4796 casc_p.n315 DGND 1.40fF $ **FLOATING
C4797 casc_p.t85 DGND 0.30fF
C4798 casc_p.n316 DGND 1.40fF $ **FLOATING
C4799 casc_p.t107 DGND 0.30fF
C4800 casc_p.n317 DGND 1.40fF $ **FLOATING
C4801 casc_p.t386 DGND 0.30fF
C4802 casc_p.n318 DGND 1.40fF $ **FLOATING
C4803 casc_p.t229 DGND 0.30fF
C4804 casc_p.n319 DGND 1.40fF $ **FLOATING
C4805 casc_p.t362 DGND 0.30fF
C4806 casc_p.n320 DGND 1.40fF $ **FLOATING
C4807 casc_p.t393 DGND 0.30fF
C4808 casc_p.n321 DGND 1.40fF $ **FLOATING
C4809 casc_p.t200 DGND 0.30fF
C4810 casc_p.n322 DGND 1.40fF $ **FLOATING
C4811 casc_p.t369 DGND 0.30fF
C4812 casc_p.n323 DGND 1.40fF $ **FLOATING
C4813 casc_p.t175 DGND 0.30fF
C4814 casc_p.n324 DGND 1.40fF $ **FLOATING
C4815 casc_p.t210 DGND 0.30fF
C4816 casc_p.n325 DGND 1.40fF $ **FLOATING
C4817 casc_p.t339 DGND 0.30fF
C4818 casc_p.n326 DGND 1.40fF $ **FLOATING
C4819 casc_p.t372 DGND 0.30fF
C4820 casc_p.n327 DGND 1.11fF $ **FLOATING
C4821 casc_p.n328 DGND 0.94fF $ **FLOATING
C4822 casc_p.n329 DGND 0.68fF $ **FLOATING
C4823 casc_p.t37 DGND 0.30fF
C4824 casc_p.n330 DGND 0.51fF $ **FLOATING
C4825 casc_p.n331 DGND 0.51fF $ **FLOATING
C4826 casc_p.n332 DGND 0.68fF $ **FLOATING
C4827 casc_p.t7 DGND 0.30fF
C4828 casc_p.n333 DGND 0.60fF $ **FLOATING
C4829 casc_p.t230 DGND 0.33fF
C4830 casc_p.t74 DGND 0.30fF
C4831 casc_p.n334 DGND 2.59fF $ **FLOATING
C4832 casc_p.t208 DGND 0.30fF
C4833 casc_p.n335 DGND 1.40fF $ **FLOATING
C4834 casc_p.t238 DGND 0.30fF
C4835 casc_p.n336 DGND 1.40fF $ **FLOATING
C4836 casc_p.t370 DGND 0.30fF
C4837 casc_p.n337 DGND 1.40fF $ **FLOATING
C4838 casc_p.t218 DGND 0.30fF
C4839 casc_p.n338 DGND 1.40fF $ **FLOATING
C4840 casc_p.t349 DGND 0.30fF
C4841 casc_p.n339 DGND 1.40fF $ **FLOATING
C4842 casc_p.t379 DGND 0.30fF
C4843 casc_p.n340 DGND 1.40fF $ **FLOATING
C4844 casc_p.t306 DGND 0.30fF
C4845 casc_p.n341 DGND 1.40fF $ **FLOATING
C4846 casc_p.t352 DGND 0.30fF
C4847 casc_p.n342 DGND 1.40fF $ **FLOATING
C4848 casc_p.t149 DGND 0.30fF
C4849 casc_p.n343 DGND 1.40fF $ **FLOATING
C4850 casc_p.t323 DGND 0.30fF
C4851 casc_p.n344 DGND 1.40fF $ **FLOATING
C4852 casc_p.t117 DGND 0.30fF
C4853 casc_p.n345 DGND 1.40fF $ **FLOATING
C4854 casc_p.t163 DGND 0.30fF
C4855 casc_p.n346 DGND 1.40fF $ **FLOATING
C4856 casc_p.t279 DGND 0.30fF
C4857 casc_p.n347 DGND 1.40fF $ **FLOATING
C4858 casc_p.t130 DGND 0.30fF
C4859 casc_p.n348 DGND 1.40fF $ **FLOATING
C4860 casc_p.t260 DGND 0.30fF
C4861 casc_p.n349 DGND 1.40fF $ **FLOATING
C4862 casc_p.t293 DGND 0.30fF
C4863 casc_p.n350 DGND 1.40fF $ **FLOATING
C4864 casc_p.t101 DGND 0.30fF
C4865 casc_p.n351 DGND 1.40fF $ **FLOATING
C4866 casc_p.t134 DGND 0.30fF
C4867 casc_p.n352 DGND 1.40fF $ **FLOATING
C4868 casc_p.t82 DGND 0.30fF
C4869 casc_p.n353 DGND 1.40fF $ **FLOATING
C4870 casc_p.t248 DGND 0.30fF
C4871 casc_p.n354 DGND 1.40fF $ **FLOATING
C4872 casc_p.t389 DGND 0.30fF
C4873 casc_p.n355 DGND 1.40fF $ **FLOATING
C4874 casc_p.t88 DGND 0.30fF
C4875 casc_p.n356 DGND 1.40fF $ **FLOATING
C4876 casc_p.t226 DGND 0.30fF
C4877 casc_p.n357 DGND 1.40fF $ **FLOATING
C4878 casc_p.t395 DGND 0.30fF
C4879 casc_p.n358 DGND 1.11fF $ **FLOATING
C4880 casc_p.n359 DGND 0.94fF $ **FLOATING
C4881 casc_p.n360 DGND 0.68fF $ **FLOATING
C4882 casc_p.t34 DGND 0.30fF
C4883 casc_p.n361 DGND 0.51fF $ **FLOATING
C4884 casc_p.n362 DGND 0.51fF $ **FLOATING
C4885 casc_p.n363 DGND 0.68fF $ **FLOATING
C4886 casc_p.t31 DGND 0.30fF
C4887 casc_p.n364 DGND 0.66fF $ **FLOATING
C4888 casc_p.n365 DGND 0.65fF $ **FLOATING
C4889 casc_p.n366 DGND 0.68fF $ **FLOATING
C4890 casc_p.t4 DGND 0.30fF
C4891 casc_p.n367 DGND 0.51fF $ **FLOATING
C4892 casc_p.n368 DGND 0.51fF $ **FLOATING
C4893 casc_p.n369 DGND 0.68fF $ **FLOATING
C4894 casc_p.t61 DGND 0.30fF
C4895 casc_p.n370 DGND 0.95fF $ **FLOATING
C4896 casc_p.t204 DGND 0.30fF
C4897 casc_p.n371 DGND 1.11fF $ **FLOATING
C4898 casc_p.t376 DGND 0.30fF
C4899 casc_p.n372 DGND 1.02fF $ **FLOATING
C4900 casc_p.t380 DGND 0.33fF
C4901 casc_p.t351 DGND 0.30fF
C4902 casc_p.n373 DGND 2.60fF $ **FLOATING
C4903 casc_p.t219 DGND 0.30fF
C4904 casc_p.n374 DGND 1.40fF $ **FLOATING
C4905 casc_p.t371 DGND 0.30fF
C4906 casc_p.n375 DGND 1.40fF $ **FLOATING
C4907 casc_p.t239 DGND 0.30fF
C4908 casc_p.n376 DGND 1.40fF $ **FLOATING
C4909 casc_p.t209 DGND 0.30fF
C4910 casc_p.n377 DGND 1.40fF $ **FLOATING
C4911 casc_p.t76 DGND 0.30fF
C4912 casc_p.n378 DGND 1.40fF $ **FLOATING
C4913 casc_p.t368 DGND 0.30fF
C4914 casc_p.n379 DGND 1.40fF $ **FLOATING
C4915 casc_p.t237 DGND 0.30fF
C4916 casc_p.n380 DGND 1.40fF $ **FLOATING
C4917 casc_p.t392 DGND 0.30fF
C4918 casc_p.n381 DGND 1.40fF $ **FLOATING
C4919 casc_p.t253 DGND 0.30fF
C4920 casc_p.n382 DGND 1.39fF $ **FLOATING
C4921 casc_p.t182 DGND 0.30fF
C4922 casc_p.n383 DGND 0.81fF $ **FLOATING
C4923 casc_p.n384 DGND 0.89fF $ **FLOATING
C4924 casc_p.n385 DGND 2.09fF $ **FLOATING
C4925 casc_p.n386 DGND 2.09fF $ **FLOATING
C4926 casc_p.n387 DGND 2.09fF $ **FLOATING
C4927 casc_p.n388 DGND 2.09fF $ **FLOATING
C4928 casc_p.n389 DGND 2.09fF $ **FLOATING
C4929 casc_p.n390 DGND 2.09fF $ **FLOATING
C4930 casc_p.n391 DGND 2.60fF $ **FLOATING
C4931 casc_p.n392 DGND 6.00fF $ **FLOATING
C4932 casc_p.n393 DGND 1.97fF $ **FLOATING
C4933 casc_p.t222 DGND 0.30fF
C4934 a_1657_n21342.n0 DGND 1.91fF $ **FLOATING
C4935 a_1657_n21342.n1 DGND 1.72fF $ **FLOATING
C4936 a_1657_n21342.n2 DGND 1.72fF $ **FLOATING
C4937 a_1657_n21342.n3 DGND 2.02fF $ **FLOATING
C4938 a_1657_n21342.n4 DGND 1.42fF $ **FLOATING
C4939 a_1657_n21342.n5 DGND 1.72fF $ **FLOATING
C4940 a_1657_n21342.n6 DGND 2.02fF $ **FLOATING
C4941 a_1657_n21342.n7 DGND 1.42fF $ **FLOATING
C4942 a_1657_n21342.n8 DGND 1.91fF $ **FLOATING
C4943 a_1657_n21342.n9 DGND 1.72fF $ **FLOATING
C4944 a_1657_n21342.n10 DGND 1.72fF $ **FLOATING
C4945 a_1657_n21342.n11 DGND 2.02fF $ **FLOATING
C4946 a_1657_n21342.n12 DGND 2.17fF $ **FLOATING
C4947 a_1657_n21342.n13 DGND 1.91fF $ **FLOATING
C4948 a_1657_n21342.n14 DGND 1.72fF $ **FLOATING
C4949 a_1657_n21342.n15 DGND 2.81fF $ **FLOATING
C4950 a_1657_n21342.n16 DGND 2.02fF $ **FLOATING
C4951 a_1657_n21342.n17 DGND 1.42fF $ **FLOATING
C4952 a_1657_n21342.n18 DGND 1.72fF $ **FLOATING
C4953 a_1657_n21342.n19 DGND 2.02fF $ **FLOATING
C4954 a_1657_n21342.n20 DGND 1.42fF $ **FLOATING
C4955 a_1657_n21342.n21 DGND 1.72fF $ **FLOATING
C4956 a_1657_n21342.n22 DGND 2.02fF $ **FLOATING
C4957 a_1657_n21342.n23 DGND 1.42fF $ **FLOATING
C4958 a_1657_n21342.n24 DGND 1.72fF $ **FLOATING
C4959 a_1657_n21342.n25 DGND 2.02fF $ **FLOATING
C4960 a_1657_n21342.n26 DGND 2.17fF $ **FLOATING
C4961 a_1657_n21342.n27 DGND 1.72fF $ **FLOATING
C4962 a_1657_n21342.n28 DGND 2.02fF $ **FLOATING
C4963 a_1657_n21342.n29 DGND 2.17fF $ **FLOATING
C4964 a_1657_n21342.n30 DGND 1.72fF $ **FLOATING
C4965 a_1657_n21342.n31 DGND 2.02fF $ **FLOATING
C4966 a_1657_n21342.n32 DGND 2.17fF $ **FLOATING
C4967 a_1657_n21342.n33 DGND 1.72fF $ **FLOATING
C4968 a_1657_n21342.n34 DGND 2.02fF $ **FLOATING
C4969 a_1657_n21342.n35 DGND 2.17fF $ **FLOATING
C4970 a_1657_n21342.n36 DGND 1.72fF $ **FLOATING
C4971 a_1657_n21342.n37 DGND 2.02fF $ **FLOATING
C4972 a_1657_n21342.n38 DGND 2.17fF $ **FLOATING
C4973 a_1657_n21342.n39 DGND 1.91fF $ **FLOATING
C4974 a_1657_n21342.n40 DGND 1.72fF $ **FLOATING
C4975 a_1657_n21342.n41 DGND 1.72fF $ **FLOATING
C4976 a_1657_n21342.n42 DGND 2.02fF $ **FLOATING
C4977 a_1657_n21342.n43 DGND 2.17fF $ **FLOATING
C4978 a_1657_n21342.n44 DGND 1.72fF $ **FLOATING
C4979 a_1657_n21342.n45 DGND 2.02fF $ **FLOATING
C4980 a_1657_n21342.n46 DGND 1.91fF $ **FLOATING
C4981 a_1657_n21342.n47 DGND 1.72fF $ **FLOATING
C4982 a_1657_n21342.n48 DGND 1.01fF $ **FLOATING
C4983 a_1657_n21342.n49 DGND 1.91fF $ **FLOATING
C4984 a_1657_n21342.n50 DGND 1.72fF $ **FLOATING
C4985 a_1657_n21342.n51 DGND 1.72fF $ **FLOATING
C4986 a_1657_n21342.n52 DGND 2.02fF $ **FLOATING
C4987 a_1657_n21342.n53 DGND 1.16fF $ **FLOATING
C4988 a_1657_n21342.n54 DGND 1.72fF $ **FLOATING
C4989 a_1657_n21342.n55 DGND 2.02fF $ **FLOATING
C4990 a_1657_n21342.n56 DGND 2.17fF $ **FLOATING
C4991 a_1657_n21342.n57 DGND 1.72fF $ **FLOATING
C4992 a_1657_n21342.n58 DGND 2.02fF $ **FLOATING
C4993 a_1657_n21342.n59 DGND 2.17fF $ **FLOATING
C4994 a_1657_n21342.n60 DGND 1.91fF $ **FLOATING
C4995 a_1657_n21342.n61 DGND 1.72fF $ **FLOATING
C4996 a_1657_n21342.n62 DGND 1.72fF $ **FLOATING
C4997 a_1657_n21342.n63 DGND 2.02fF $ **FLOATING
C4998 a_1657_n21342.n64 DGND 2.17fF $ **FLOATING
C4999 a_1657_n21342.n65 DGND 1.72fF $ **FLOATING
C5000 a_1657_n21342.n66 DGND 2.02fF $ **FLOATING
C5001 a_1657_n21342.n67 DGND 2.17fF $ **FLOATING
C5002 a_1657_n21342.n68 DGND 1.72fF $ **FLOATING
C5003 a_1657_n21342.n69 DGND 2.02fF $ **FLOATING
C5004 a_1657_n21342.n70 DGND 2.17fF $ **FLOATING
C5005 a_1657_n21342.n71 DGND 1.72fF $ **FLOATING
C5006 a_1657_n21342.n72 DGND 2.02fF $ **FLOATING
C5007 a_1657_n21342.n73 DGND 2.17fF $ **FLOATING
C5008 a_1657_n21342.n74 DGND 1.72fF $ **FLOATING
C5009 a_1657_n21342.n75 DGND 2.02fF $ **FLOATING
C5010 a_1657_n21342.n76 DGND 2.17fF $ **FLOATING
C5011 a_1657_n21342.n77 DGND 1.72fF $ **FLOATING
C5012 a_1657_n21342.n78 DGND 2.02fF $ **FLOATING
C5013 a_1657_n21342.n79 DGND 2.17fF $ **FLOATING
C5014 a_1657_n21342.n80 DGND 1.72fF $ **FLOATING
C5015 a_1657_n21342.n81 DGND 2.02fF $ **FLOATING
C5016 a_1657_n21342.n82 DGND 2.17fF $ **FLOATING
C5017 a_1657_n21342.n83 DGND 2.45fF $ **FLOATING
C5018 a_1657_n21342.n84 DGND 2.02fF $ **FLOATING
C5019 a_1657_n21342.n85 DGND 1.01fF $ **FLOATING
C5020 a_1657_n21342.n86 DGND 1.72fF $ **FLOATING
C5021 a_1657_n21342.n87 DGND 2.02fF $ **FLOATING
C5022 a_1657_n21342.n88 DGND 1.01fF $ **FLOATING
C5023 a_1657_n21342.n89 DGND 1.72fF $ **FLOATING
C5024 a_1657_n21342.n90 DGND 2.02fF $ **FLOATING
C5025 a_1657_n21342.n91 DGND 1.01fF $ **FLOATING
C5026 a_1657_n21342.n92 DGND 1.72fF $ **FLOATING
C5027 a_1657_n21342.n93 DGND 2.02fF $ **FLOATING
C5028 a_1657_n21342.n94 DGND 2.17fF $ **FLOATING
C5029 a_1657_n21342.n95 DGND 1.72fF $ **FLOATING
C5030 a_1657_n21342.n96 DGND 2.02fF $ **FLOATING
C5031 a_1657_n21342.n97 DGND 2.17fF $ **FLOATING
C5032 a_1657_n21342.n98 DGND 1.72fF $ **FLOATING
C5033 a_1657_n21342.n99 DGND 2.02fF $ **FLOATING
C5034 a_1657_n21342.n100 DGND 2.17fF $ **FLOATING
C5035 a_1657_n21342.n101 DGND 1.72fF $ **FLOATING
C5036 a_1657_n21342.n102 DGND 2.02fF $ **FLOATING
C5037 a_1657_n21342.n103 DGND 2.17fF $ **FLOATING
C5038 a_1657_n21342.n104 DGND 1.72fF $ **FLOATING
C5039 a_1657_n21342.n105 DGND 2.02fF $ **FLOATING
C5040 a_1657_n21342.n106 DGND 2.17fF $ **FLOATING
C5041 a_1657_n21342.n107 DGND 1.72fF $ **FLOATING
C5042 a_1657_n21342.n108 DGND 2.02fF $ **FLOATING
C5043 a_1657_n21342.n109 DGND 2.17fF $ **FLOATING
C5044 a_1657_n21342.n110 DGND 1.72fF $ **FLOATING
C5045 a_1657_n21342.n111 DGND 2.02fF $ **FLOATING
C5046 a_1657_n21342.n112 DGND 2.17fF $ **FLOATING
C5047 a_1657_n21342.n113 DGND 1.72fF $ **FLOATING
C5048 a_1657_n21342.n114 DGND 2.02fF $ **FLOATING
C5049 a_1657_n21342.n115 DGND 2.17fF $ **FLOATING
C5050 a_1657_n21342.n116 DGND 1.72fF $ **FLOATING
C5051 a_1657_n21342.n117 DGND 2.02fF $ **FLOATING
C5052 a_1657_n21342.n118 DGND 2.17fF $ **FLOATING
C5053 a_1657_n21342.n119 DGND 2.12fF $ **FLOATING
C5054 a_1657_n21342.n120 DGND 1.98fF $ **FLOATING
C5055 a_1657_n21342.n121 DGND 1.98fF $ **FLOATING
C5056 a_1657_n21342.n122 DGND 2.07fF $ **FLOATING
C5057 a_1657_n21342.n123 DGND 1.98fF $ **FLOATING
C5058 a_1657_n21342.n124 DGND 1.98fF $ **FLOATING
C5059 a_1657_n21342.n125 DGND 1.72fF $ **FLOATING
C5060 a_1657_n21342.n126 DGND 2.02fF $ **FLOATING
C5061 a_1657_n21342.n127 DGND 2.17fF $ **FLOATING
C5062 a_1657_n21342.n128 DGND 1.72fF $ **FLOATING
C5063 a_1657_n21342.n129 DGND 2.02fF $ **FLOATING
C5064 a_1657_n21342.n130 DGND 2.17fF $ **FLOATING
C5065 a_1657_n21342.n131 DGND 1.72fF $ **FLOATING
C5066 a_1657_n21342.n132 DGND 2.02fF $ **FLOATING
C5067 a_1657_n21342.n133 DGND 2.17fF $ **FLOATING
C5068 a_1657_n21342.n134 DGND 1.72fF $ **FLOATING
C5069 a_1657_n21342.n135 DGND 2.02fF $ **FLOATING
C5070 a_1657_n21342.n136 DGND 2.17fF $ **FLOATING
C5071 a_1657_n21342.n137 DGND 1.72fF $ **FLOATING
C5072 a_1657_n21342.n138 DGND 2.02fF $ **FLOATING
C5073 a_1657_n21342.n139 DGND 2.17fF $ **FLOATING
C5074 a_1657_n21342.n140 DGND 1.72fF $ **FLOATING
C5075 a_1657_n21342.n141 DGND 1.91fF $ **FLOATING
C5076 a_1560_n22142.n0 DGND 1.46fF $ **FLOATING
C5077 a_1560_n22142.n1 DGND 11.66fF $ **FLOATING
C5078 a_1560_n22142.n2 DGND 2.71fF $ **FLOATING
C5079 a_1560_n22142.n3 DGND 2.20fF $ **FLOATING
C5080 a_1560_n22142.n4 DGND 2.12fF $ **FLOATING
C5081 a_1560_n22142.n5 DGND 2.35fF $ **FLOATING
C5082 a_1560_n22142.n6 DGND 2.12fF $ **FLOATING
C5083 a_1560_n22142.n7 DGND 2.35fF $ **FLOATING
C5084 a_1560_n22142.n8 DGND 2.12fF $ **FLOATING
C5085 a_1560_n22142.n9 DGND 2.35fF $ **FLOATING
C5086 a_1560_n22142.n10 DGND 2.24fF $ **FLOATING
C5087 a_1560_n22142.n11 DGND 2.24fF $ **FLOATING
C5088 a_1560_n22142.n12 DGND 2.24fF $ **FLOATING
C5089 a_1560_n22142.n13 DGND 2.24fF $ **FLOATING
C5090 a_1560_n22142.n14 DGND 2.24fF $ **FLOATING
C5091 a_1560_n22142.n15 DGND 2.24fF $ **FLOATING
C5092 a_1560_n22142.n16 DGND 2.24fF $ **FLOATING
C5093 a_1560_n22142.n17 DGND 2.62fF $ **FLOATING
C5094 a_1560_n22142.n18 DGND 2.26fF $ **FLOATING
C5095 a_1560_n22142.n19 DGND 2.24fF $ **FLOATING
C5096 a_1560_n22142.n20 DGND 2.09fF $ **FLOATING
C5097 a_1560_n22142.n21 DGND 2.24fF $ **FLOATING
C5098 a_1560_n22142.n22 DGND 2.09fF $ **FLOATING
C5099 a_1560_n22142.n23 DGND 2.24fF $ **FLOATING
C5100 a_1560_n22142.n24 DGND 2.24fF $ **FLOATING
C5101 a_1560_n22142.n25 DGND 2.24fF $ **FLOATING
C5102 a_1560_n22142.n26 DGND 2.24fF $ **FLOATING
C5103 a_1560_n22142.n27 DGND 2.24fF $ **FLOATING
C5104 a_1560_n22142.n28 DGND 2.24fF $ **FLOATING
C5105 a_1560_n22142.n29 DGND 2.24fF $ **FLOATING
C5106 a_1560_n22142.n30 DGND 2.24fF $ **FLOATING
C5107 a_1560_n22142.n31 DGND 2.24fF $ **FLOATING
C5108 a_1560_n22142.n32 DGND 2.09fF $ **FLOATING
C5109 a_1560_n22142.n33 DGND 2.24fF $ **FLOATING
C5110 a_1560_n22142.n34 DGND 2.24fF $ **FLOATING
C5111 a_1560_n22142.n35 DGND 2.24fF $ **FLOATING
C5112 a_1560_n22142.n36 DGND 2.09fF $ **FLOATING
C5113 a_1560_n22142.n37 DGND 2.24fF $ **FLOATING
C5114 a_1560_n22142.n38 DGND 2.24fF $ **FLOATING
C5115 a_1560_n22142.n39 DGND 2.09fF $ **FLOATING
C5116 a_1560_n22142.n40 DGND 2.24fF $ **FLOATING
C5117 a_1560_n22142.n41 DGND 2.24fF $ **FLOATING
C5118 a_1560_n22142.n42 DGND 2.09fF $ **FLOATING
C5119 a_1560_n22142.n43 DGND 2.24fF $ **FLOATING
C5120 a_1560_n22142.n44 DGND 2.24fF $ **FLOATING
C5121 a_1560_n22142.n45 DGND 2.24fF $ **FLOATING
C5122 a_1560_n22142.n46 DGND 2.24fF $ **FLOATING
C5123 a_1560_n22142.n47 DGND 2.24fF $ **FLOATING
C5124 a_1560_n22142.n48 DGND 2.24fF $ **FLOATING
C5125 a_1560_n22142.n49 DGND 2.24fF $ **FLOATING
C5126 a_1560_n22142.n50 DGND 2.24fF $ **FLOATING
C5127 a_1560_n22142.n51 DGND 2.24fF $ **FLOATING
C5128 a_1560_n22142.n52 DGND 2.24fF $ **FLOATING
C5129 a_1560_n22142.n53 DGND 2.24fF $ **FLOATING
C5130 a_1560_n22142.n54 DGND 2.24fF $ **FLOATING
C5131 a_1560_n22142.n55 DGND 2.20fF $ **FLOATING
C5132 a_1560_n22142.n56 DGND 2.64fF $ **FLOATING
C5133 a_1560_n22142.n57 DGND 2.64fF $ **FLOATING
C5134 a_1560_n22142.n58 DGND 2.64fF $ **FLOATING
C5135 a_1560_n22142.n59 DGND 2.64fF $ **FLOATING
C5136 a_1560_n22142.n60 DGND 0.66fF $ **FLOATING
C5137 a_1560_n22142.n61 DGND 0.70fF $ **FLOATING
C5138 a_1560_n22142.t22 DGND 1.72fF
C5139 a_1560_n22142.t43 DGND 1.72fF
C5140 a_1560_n22142.n63 DGND 0.13fF $ **FLOATING
C5141 a_1560_n22142.n64 DGND 0.13fF $ **FLOATING
C5142 a_1560_n22142.n65 DGND 0.11fF $ **FLOATING
C5143 a_1560_n22142.t93 DGND 1.72fF
C5144 a_1560_n22142.t42 DGND 1.72fF
C5145 a_1560_n22142.n67 DGND 0.13fF $ **FLOATING
C5146 a_1560_n22142.n68 DGND 0.13fF $ **FLOATING
C5147 a_1560_n22142.n69 DGND 0.11fF $ **FLOATING
C5148 a_1560_n22142.t26 DGND 1.72fF
C5149 a_1560_n22142.t89 DGND 1.72fF
C5150 a_1560_n22142.n71 DGND 0.13fF $ **FLOATING
C5151 a_1560_n22142.n72 DGND 0.13fF $ **FLOATING
C5152 a_1560_n22142.n73 DGND 0.11fF $ **FLOATING
C5153 a_1560_n22142.t13 DGND 1.72fF
C5154 a_1560_n22142.t32 DGND 1.72fF
C5155 a_1560_n22142.n75 DGND 0.13fF $ **FLOATING
C5156 a_1560_n22142.n76 DGND 0.13fF $ **FLOATING
C5157 a_1560_n22142.n77 DGND 0.11fF $ **FLOATING
C5158 a_1560_n22142.t70 DGND 1.72fF
C5159 a_1560_n22142.t82 DGND 1.72fF
C5160 a_1560_n22142.n79 DGND 0.13fF $ **FLOATING
C5161 a_1560_n22142.n80 DGND 0.13fF $ **FLOATING
C5162 a_1560_n22142.n81 DGND 0.11fF $ **FLOATING
C5163 a_1560_n22142.n82 DGND 1.19fF $ **FLOATING
C5164 a_1560_n22142.t80 DGND 1.72fF
C5165 a_1560_n22142.t99 DGND 1.72fF
C5166 a_1560_n22142.n84 DGND 0.13fF $ **FLOATING
C5167 a_1560_n22142.n85 DGND 0.13fF $ **FLOATING
C5168 a_1560_n22142.n86 DGND 0.11fF $ **FLOATING
C5169 a_1560_n22142.n87 DGND 1.19fF $ **FLOATING
C5170 a_1560_n22142.n88 DGND 1.80fF $ **FLOATING
C5171 a_1560_n22142.t85 DGND 1.72fF
C5172 a_1560_n22142.t104 DGND 1.72fF
C5173 a_1560_n22142.n90 DGND 0.13fF $ **FLOATING
C5174 a_1560_n22142.n91 DGND 0.13fF $ **FLOATING
C5175 a_1560_n22142.n92 DGND 0.11fF $ **FLOATING
C5176 a_1560_n22142.t34 DGND 1.72fF
C5177 a_1560_n22142.t53 DGND 1.72fF
C5178 a_1560_n22142.n94 DGND 0.13fF $ **FLOATING
C5179 a_1560_n22142.n95 DGND 0.13fF $ **FLOATING
C5180 a_1560_n22142.n96 DGND 0.11fF $ **FLOATING
C5181 a_1560_n22142.n97 DGND 1.80fF $ **FLOATING
C5182 a_1560_n22142.t24 DGND 1.72fF
C5183 a_1560_n22142.t45 DGND 1.72fF
C5184 a_1560_n22142.n99 DGND 0.13fF $ **FLOATING
C5185 a_1560_n22142.n100 DGND 0.13fF $ **FLOATING
C5186 a_1560_n22142.n101 DGND 0.11fF $ **FLOATING
C5187 a_1560_n22142.t77 DGND 1.72fF
C5188 a_1560_n22142.t21 DGND 1.72fF
C5189 a_1560_n22142.n103 DGND 0.13fF $ **FLOATING
C5190 a_1560_n22142.n104 DGND 0.13fF $ **FLOATING
C5191 a_1560_n22142.n105 DGND 0.11fF $ **FLOATING
C5192 a_1560_n22142.n106 DGND 1.80fF $ **FLOATING
C5193 a_1560_n22142.t17 DGND 1.72fF
C5194 a_1560_n22142.t37 DGND 1.72fF
C5195 a_1560_n22142.n108 DGND 0.13fF $ **FLOATING
C5196 a_1560_n22142.n109 DGND 0.13fF $ **FLOATING
C5197 a_1560_n22142.n110 DGND 0.11fF $ **FLOATING
C5198 a_1560_n22142.t11 DGND 1.72fF
C5199 a_1560_n22142.t23 DGND 1.72fF
C5200 a_1560_n22142.n112 DGND 0.13fF $ **FLOATING
C5201 a_1560_n22142.n113 DGND 0.13fF $ **FLOATING
C5202 a_1560_n22142.n114 DGND 0.11fF $ **FLOATING
C5203 a_1560_n22142.t67 DGND 1.72fF
C5204 a_1560_n22142.t74 DGND 1.72fF
C5205 a_1560_n22142.n116 DGND 0.13fF $ **FLOATING
C5206 a_1560_n22142.n117 DGND 0.13fF $ **FLOATING
C5207 a_1560_n22142.n118 DGND 0.11fF $ **FLOATING
C5208 a_1560_n22142.t57 DGND 1.72fF
C5209 a_1560_n22142.t109 DGND 1.72fF
C5210 a_1560_n22142.n120 DGND 0.13fF $ **FLOATING
C5211 a_1560_n22142.n121 DGND 0.13fF $ **FLOATING
C5212 a_1560_n22142.n122 DGND 0.11fF $ **FLOATING
C5213 a_1560_n22142.n123 DGND 1.19fF $ **FLOATING
C5214 a_1560_n22142.n124 DGND 1.19fF $ **FLOATING
C5215 a_1560_n22142.n125 DGND 1.19fF $ **FLOATING
C5216 a_1560_n22142.t19 DGND 1.72fF
C5217 a_1560_n22142.t83 DGND 1.72fF
C5218 a_1560_n22142.n127 DGND 0.13fF $ **FLOATING
C5219 a_1560_n22142.n128 DGND 0.13fF $ **FLOATING
C5220 a_1560_n22142.n129 DGND 0.11fF $ **FLOATING
C5221 a_1560_n22142.t72 DGND 1.72fF
C5222 a_1560_n22142.t14 DGND 1.72fF
C5223 a_1560_n22142.n131 DGND 0.13fF $ **FLOATING
C5224 a_1560_n22142.n132 DGND 0.13fF $ **FLOATING
C5225 a_1560_n22142.n133 DGND 0.11fF $ **FLOATING
C5226 a_1560_n22142.t108 DGND 1.72fF
C5227 a_1560_n22142.t16 DGND 1.72fF
C5228 a_1560_n22142.n135 DGND 0.13fF $ **FLOATING
C5229 a_1560_n22142.n136 DGND 0.13fF $ **FLOATING
C5230 a_1560_n22142.n137 DGND 0.11fF $ **FLOATING
C5231 a_1560_n22142.n138 DGND 1.80fF $ **FLOATING
C5232 a_1560_n22142.n139 DGND 1.80fF $ **FLOATING
C5233 a_1560_n22142.n140 DGND 1.80fF $ **FLOATING
C5234 a_1560_n22142.t78 DGND 1.72fF
C5235 a_1560_n22142.t96 DGND 1.72fF
C5236 a_1560_n22142.n142 DGND 0.13fF $ **FLOATING
C5237 a_1560_n22142.n143 DGND 0.13fF $ **FLOATING
C5238 a_1560_n22142.n144 DGND 0.11fF $ **FLOATING
C5239 a_1560_n22142.t12 DGND 1.72fF
C5240 a_1560_n22142.t28 DGND 1.72fF
C5241 a_1560_n22142.n146 DGND 0.13fF $ **FLOATING
C5242 a_1560_n22142.n147 DGND 0.13fF $ **FLOATING
C5243 a_1560_n22142.n148 DGND 0.11fF $ **FLOATING
C5244 a_1560_n22142.t15 DGND 1.72fF
C5245 a_1560_n22142.t68 DGND 1.72fF
C5246 a_1560_n22142.n150 DGND 0.13fF $ **FLOATING
C5247 a_1560_n22142.n151 DGND 0.13fF $ **FLOATING
C5248 a_1560_n22142.n152 DGND 0.11fF $ **FLOATING
C5249 a_1560_n22142.n153 DGND 1.80fF $ **FLOATING
C5250 a_1560_n22142.n154 DGND 1.80fF $ **FLOATING
C5251 a_1560_n22142.n155 DGND 1.80fF $ **FLOATING
C5252 a_1560_n22142.n156 DGND 1.80fF $ **FLOATING
C5253 a_1560_n22142.t76 DGND 1.72fF
C5254 a_1560_n22142.t94 DGND 1.72fF
C5255 a_1560_n22142.n158 DGND 0.13fF $ **FLOATING
C5256 a_1560_n22142.n159 DGND 0.13fF $ **FLOATING
C5257 a_1560_n22142.n160 DGND 0.11fF $ **FLOATING
C5258 a_1560_n22142.t18 DGND 1.72fF
C5259 a_1560_n22142.t38 DGND 1.72fF
C5260 a_1560_n22142.n162 DGND 0.13fF $ **FLOATING
C5261 a_1560_n22142.n163 DGND 0.13fF $ **FLOATING
C5262 a_1560_n22142.n164 DGND 0.11fF $ **FLOATING
C5263 a_1560_n22142.t71 DGND 1.72fF
C5264 a_1560_n22142.t86 DGND 1.72fF
C5265 a_1560_n22142.n166 DGND 0.13fF $ **FLOATING
C5266 a_1560_n22142.n167 DGND 0.13fF $ **FLOATING
C5267 a_1560_n22142.n168 DGND 0.11fF $ **FLOATING
C5268 a_1560_n22142.t64 DGND 1.72fF
C5269 a_1560_n22142.t119 DGND 1.72fF
C5270 a_1560_n22142.n170 DGND 0.13fF $ **FLOATING
C5271 a_1560_n22142.n171 DGND 0.13fF $ **FLOATING
C5272 a_1560_n22142.n172 DGND 0.11fF $ **FLOATING
C5273 a_1560_n22142.n173 DGND 1.80fF $ **FLOATING
C5274 a_1560_n22142.n174 DGND 1.80fF $ **FLOATING
C5275 a_1560_n22142.n175 DGND 1.80fF $ **FLOATING
C5276 a_1560_n22142.n176 DGND 1.80fF $ **FLOATING
C5277 a_1560_n22142.t91 DGND 1.72fF
C5278 a_1560_n22142.t113 DGND 1.72fF
C5279 a_1560_n22142.n178 DGND 0.13fF $ **FLOATING
C5280 a_1560_n22142.n179 DGND 0.13fF $ **FLOATING
C5281 a_1560_n22142.n180 DGND 0.11fF $ **FLOATING
C5282 a_1560_n22142.n181 DGND 1.80fF $ **FLOATING
C5283 a_1560_n22142.t39 DGND 1.72fF
C5284 a_1560_n22142.t101 DGND 1.72fF
C5285 a_1560_n22142.n183 DGND 0.13fF $ **FLOATING
C5286 a_1560_n22142.n184 DGND 0.13fF $ **FLOATING
C5287 a_1560_n22142.n185 DGND 0.11fF $ **FLOATING
C5288 a_1560_n22142.t87 DGND 1.72fF
C5289 a_1560_n22142.t35 DGND 1.72fF
C5290 a_1560_n22142.n187 DGND 0.13fF $ **FLOATING
C5291 a_1560_n22142.n188 DGND 0.13fF $ **FLOATING
C5292 a_1560_n22142.n189 DGND 0.11fF $ **FLOATING
C5293 a_1560_n22142.t30 DGND 1.72fF
C5294 a_1560_n22142.t95 DGND 1.72fF
C5295 a_1560_n22142.n191 DGND 0.13fF $ **FLOATING
C5296 a_1560_n22142.n192 DGND 0.13fF $ **FLOATING
C5297 a_1560_n22142.n193 DGND 0.11fF $ **FLOATING
C5298 a_1560_n22142.n194 DGND 1.80fF $ **FLOATING
C5299 a_1560_n22142.n195 DGND 1.80fF $ **FLOATING
C5300 a_1560_n22142.t105 DGND 1.72fF
C5301 a_1560_n22142.t51 DGND 1.72fF
C5302 a_1560_n22142.n197 DGND 0.13fF $ **FLOATING
C5303 a_1560_n22142.n198 DGND 0.13fF $ **FLOATING
C5304 a_1560_n22142.n199 DGND 0.11fF $ **FLOATING
C5305 a_1560_n22142.n200 DGND 1.80fF $ **FLOATING
C5306 a_1560_n22142.t73 DGND 1.72fF
C5307 a_1560_n22142.t115 DGND 1.72fF
C5308 a_1560_n22142.n202 DGND 0.13fF $ **FLOATING
C5309 a_1560_n22142.n203 DGND 0.13fF $ **FLOATING
C5310 a_1560_n22142.n204 DGND 0.11fF $ **FLOATING
C5311 a_1560_n22142.t10 DGND 1.72fF
C5312 a_1560_n22142.t48 DGND 1.72fF
C5313 a_1560_n22142.n206 DGND 0.13fF $ **FLOATING
C5314 a_1560_n22142.n207 DGND 0.13fF $ **FLOATING
C5315 a_1560_n22142.n208 DGND 0.11fF $ **FLOATING
C5316 a_1560_n22142.t69 DGND 1.72fF
C5317 a_1560_n22142.t106 DGND 1.72fF
C5318 a_1560_n22142.n210 DGND 0.13fF $ **FLOATING
C5319 a_1560_n22142.n211 DGND 0.13fF $ **FLOATING
C5320 a_1560_n22142.n212 DGND 0.11fF $ **FLOATING
C5321 a_1560_n22142.t79 DGND 1.72fF
C5322 a_1560_n22142.t27 DGND 1.72fF
C5323 a_1560_n22142.n214 DGND 0.13fF $ **FLOATING
C5324 a_1560_n22142.n215 DGND 0.13fF $ **FLOATING
C5325 a_1560_n22142.n216 DGND 0.11fF $ **FLOATING
C5326 a_1560_n22142.t118 DGND 1.72fF
C5327 a_1560_n22142.t29 DGND 1.72fF
C5328 a_1560_n22142.n218 DGND 0.13fF $ **FLOATING
C5329 a_1560_n22142.n219 DGND 0.13fF $ **FLOATING
C5330 a_1560_n22142.n220 DGND 0.11fF $ **FLOATING
C5331 a_1560_n22142.n221 DGND 1.80fF $ **FLOATING
C5332 a_1560_n22142.n222 DGND 1.80fF $ **FLOATING
C5333 a_1560_n22142.t125 DGND 1.72fF
C5334 a_1560_n22142.t41 DGND 1.72fF
C5335 a_1560_n22142.n224 DGND 0.13fF $ **FLOATING
C5336 a_1560_n22142.n225 DGND 0.13fF $ **FLOATING
C5337 a_1560_n22142.n226 DGND 0.11fF $ **FLOATING
C5338 a_1560_n22142.t60 DGND 1.72fF
C5339 a_1560_n22142.t75 DGND 1.72fF
C5340 a_1560_n22142.n228 DGND 0.13fF $ **FLOATING
C5341 a_1560_n22142.n229 DGND 0.13fF $ **FLOATING
C5342 a_1560_n22142.n230 DGND 0.11fF $ **FLOATING
C5343 a_1560_n22142.n231 DGND 1.19fF $ **FLOATING
C5344 a_1560_n22142.n232 DGND 1.19fF $ **FLOATING
C5345 a_1560_n22142.n233 DGND 1.19fF $ **FLOATING
C5346 a_1560_n22142.n234 DGND 1.19fF $ **FLOATING
C5347 a_1560_n22142.t20 DGND 1.72fF
C5348 a_1560_n22142.t59 DGND 1.72fF
C5349 a_1560_n22142.n236 DGND 0.13fF $ **FLOATING
C5350 a_1560_n22142.n237 DGND 0.13fF $ **FLOATING
C5351 a_1560_n22142.n238 DGND 0.11fF $ **FLOATING
C5352 a_1560_n22142.n239 DGND 2.45fF $ **FLOATING
C5353 a_1560_n22142.t90 DGND 1.72fF
C5354 a_1560_n22142.t111 DGND 1.72fF
C5355 a_1560_n22142.n241 DGND 0.13fF $ **FLOATING
C5356 a_1560_n22142.n242 DGND 0.13fF $ **FLOATING
C5357 a_1560_n22142.n243 DGND 0.11fF $ **FLOATING
C5358 a_1560_n22142.t114 DGND 1.72fF
C5359 a_1560_n22142.t97 DGND 1.72fF
C5360 a_1560_n22142.n244 DGND 1.19fF $ **FLOATING
C5361 a_1560_n22142.t54 DGND 1.72fF
C5362 a_1560_n22142.t110 DGND 1.72fF
C5363 a_1560_n22142.t46 DGND 1.72fF
C5364 a_1560_n22142.t58 DGND 1.72fF
C5365 a_1560_n22142.n246 DGND 0.13fF $ **FLOATING
C5366 a_1560_n22142.n247 DGND 0.13fF $ **FLOATING
C5367 a_1560_n22142.n248 DGND 0.11fF $ **FLOATING
C5368 a_1560_n22142.n249 DGND 1.19fF $ **FLOATING
C5369 a_1560_n22142.t56 DGND 1.72fF
C5370 a_1560_n22142.t120 DGND 1.72fF
C5371 a_1560_n22142.n251 DGND 0.13fF $ **FLOATING
C5372 a_1560_n22142.n252 DGND 0.13fF $ **FLOATING
C5373 a_1560_n22142.n253 DGND 0.11fF $ **FLOATING
C5374 a_1560_n22142.n254 DGND 2.01fF $ **FLOATING
C5375 a_1560_n22142.n255 DGND 1.80fF $ **FLOATING
C5376 a_1560_n22142.n256 DGND 1.80fF $ **FLOATING
C5377 a_1560_n22142.t62 DGND 1.72fF
C5378 a_1560_n22142.t49 DGND 1.72fF
C5379 a_1560_n22142.t116 DGND 1.72fF
C5380 a_1560_n22142.t123 DGND 1.72fF
C5381 a_1560_n22142.n258 DGND 0.13fF $ **FLOATING
C5382 a_1560_n22142.n259 DGND 0.13fF $ **FLOATING
C5383 a_1560_n22142.n260 DGND 0.11fF $ **FLOATING
C5384 a_1560_n22142.n261 DGND 1.50fF $ **FLOATING
C5385 a_1560_n22142.n262 DGND 1.80fF $ **FLOATING
C5386 a_1560_n22142.n263 DGND 1.80fF $ **FLOATING
C5387 a_1560_n22142.t121 DGND 1.72fF
C5388 a_1560_n22142.t107 DGND 1.72fF
C5389 a_1560_n22142.n264 DGND 1.80fF $ **FLOATING
C5390 a_1560_n22142.t117 DGND 1.72fF
C5391 a_1560_n22142.t61 DGND 1.72fF
C5392 a_1560_n22142.n266 DGND 0.13fF $ **FLOATING
C5393 a_1560_n22142.n267 DGND 0.13fF $ **FLOATING
C5394 a_1560_n22142.n268 DGND 0.11fF $ **FLOATING
C5395 a_1560_n22142.n269 DGND 1.80fF $ **FLOATING
C5396 a_1560_n22142.t36 DGND 1.72fF
C5397 a_1560_n22142.t66 DGND 1.72fF
C5398 a_1560_n22142.n271 DGND 0.13fF $ **FLOATING
C5399 a_1560_n22142.n272 DGND 0.13fF $ **FLOATING
C5400 a_1560_n22142.n273 DGND 0.11fF $ **FLOATING
C5401 a_1560_n22142.t55 DGND 1.72fF
C5402 a_1560_n22142.t65 DGND 1.72fF
C5403 a_1560_n22142.n275 DGND 0.13fF $ **FLOATING
C5404 a_1560_n22142.n276 DGND 0.13fF $ **FLOATING
C5405 a_1560_n22142.n277 DGND 0.11fF $ **FLOATING
C5406 a_1560_n22142.n278 DGND 1.80fF $ **FLOATING
C5407 a_1560_n22142.t63 DGND 1.72fF
C5408 a_1560_n22142.t122 DGND 1.72fF
C5409 a_1560_n22142.n280 DGND 0.13fF $ **FLOATING
C5410 a_1560_n22142.n281 DGND 0.13fF $ **FLOATING
C5411 a_1560_n22142.n282 DGND 0.11fF $ **FLOATING
C5412 a_1560_n22142.n283 DGND 1.80fF $ **FLOATING
C5413 a_1560_n22142.t102 DGND 1.72fF
C5414 a_1560_n22142.t124 DGND 1.72fF
C5415 a_1560_n22142.n285 DGND 0.13fF $ **FLOATING
C5416 a_1560_n22142.n286 DGND 0.13fF $ **FLOATING
C5417 a_1560_n22142.n287 DGND 0.11fF $ **FLOATING
C5418 a_1560_n22142.n288 DGND 1.50fF $ **FLOATING
C5419 a_1560_n22142.n289 DGND 1.50fF $ **FLOATING
C5420 a_1560_n22142.t33 DGND 1.72fF
C5421 a_1560_n22142.t52 DGND 1.72fF
C5422 a_1560_n22142.n291 DGND 0.13fF $ **FLOATING
C5423 a_1560_n22142.n292 DGND 0.13fF $ **FLOATING
C5424 a_1560_n22142.n293 DGND 0.12fF $ **FLOATING
C5425 a_1560_n22142.t84 DGND 1.72fF
C5426 a_1560_n22142.t103 DGND 1.72fF
C5427 a_1560_n22142.n295 DGND 0.13fF $ **FLOATING
C5428 a_1560_n22142.n296 DGND 0.13fF $ **FLOATING
C5429 a_1560_n22142.n297 DGND 0.12fF $ **FLOATING
C5430 a_1560_n22142.t92 DGND 1.72fF
C5431 a_1560_n22142.t40 DGND 1.72fF
C5432 a_1560_n22142.n299 DGND 0.13fF $ **FLOATING
C5433 a_1560_n22142.n300 DGND 0.13fF $ **FLOATING
C5434 a_1560_n22142.n301 DGND 0.12fF $ **FLOATING
C5435 a_1560_n22142.t25 DGND 1.72fF
C5436 a_1560_n22142.t88 DGND 1.72fF
C5437 a_1560_n22142.n303 DGND 0.13fF $ **FLOATING
C5438 a_1560_n22142.n304 DGND 0.13fF $ **FLOATING
C5439 a_1560_n22142.n305 DGND 0.12fF $ **FLOATING
C5440 a_1560_n22142.n306 DGND 1.20fF $ **FLOATING
C5441 a_1560_n22142.t47 DGND 1.72fF
C5442 a_1560_n22142.t112 DGND 1.72fF
C5443 a_1560_n22142.n308 DGND 0.13fF $ **FLOATING
C5444 a_1560_n22142.n309 DGND 0.13fF $ **FLOATING
C5445 a_1560_n22142.n310 DGND 0.12fF $ **FLOATING
C5446 a_1560_n22142.t98 DGND 1.72fF
C5447 a_1560_n22142.t44 DGND 1.72fF
C5448 a_1560_n22142.n312 DGND 0.13fF $ **FLOATING
C5449 a_1560_n22142.n313 DGND 0.13fF $ **FLOATING
C5450 a_1560_n22142.n314 DGND 0.12fF $ **FLOATING
C5451 a_1560_n22142.n315 DGND 9.96fF $ **FLOATING
C5452 a_1560_n22142.n316 DGND 1.19fF $ **FLOATING
C5453 a_1560_n22142.n317 DGND 2.45fF $ **FLOATING
C5454 a_1560_n22142.n318 DGND 2.73fF $ **FLOATING
C5455 a_1560_n22142.n319 DGND 2.50fF $ **FLOATING
C5456 a_1560_n22142.n320 DGND 0.75fF $ **FLOATING
C5457 a_1560_n22142.n321 DGND 0.28fF $ **FLOATING
C5458 a_1560_n22142.t81 DGND 1.72fF
C5459 a_1560_n22142.t100 DGND 1.72fF
C5460 a_1560_n22142.n323 DGND 0.13fF $ **FLOATING
C5461 a_1560_n22142.n324 DGND 0.13fF $ **FLOATING
C5462 a_1560_n22142.n325 DGND 0.11fF $ **FLOATING
C5463 a_1560_n22142.t31 DGND 1.72fF
C5464 a_1560_n22142.t50 DGND 1.72fF
C5465 a_1560_n22142.n327 DGND 0.13fF $ **FLOATING
C5466 a_1560_n22142.n328 DGND 0.13fF $ **FLOATING
C5467 a_1560_n22142.n329 DGND 0.11fF $ **FLOATING
C5468 a_1560_n22142.n330 DGND 1.29fF $ **FLOATING
C5469 a_1560_n22142.n331 DGND 0.75fF $ **FLOATING
C5470 a_1560_n22142.n332 DGND 0.32fF $ **FLOATING
C5471 a_1560_n22142.n333 DGND 0.65fF $ **FLOATING
C5472 a_1560_n22142.n334 DGND 3.16fF $ **FLOATING
C5473 a_1560_n22142.n335 DGND 3.47fF $ **FLOATING
C5474 AVDD.n0 DGND 0.22fF $ **FLOATING
C5475 AVDD.n12 DGND 0.33fF $ **FLOATING
C5476 AVDD.n13 DGND 0.88fF $ **FLOATING
C5477 AVDD.n14 DGND 0.15fF $ **FLOATING
C5478 AVDD.n15 DGND 0.19fF $ **FLOATING
C5479 AVDD.n17 DGND 0.12fF $ **FLOATING
C5480 AVDD.n20 DGND 0.60fF $ **FLOATING
C5481 AVDD.n23 DGND 0.10fF $ **FLOATING
C5482 AVDD.n25 DGND 0.66fF $ **FLOATING
C5483 AVDD.n27 DGND 2.44fF $ **FLOATING
C5484 AVDD.n28 DGND 2.50fF $ **FLOATING
C5485 AVDD.n30 DGND 0.63fF $ **FLOATING
C5486 AVDD.t725 DGND 1.33fF
C5487 AVDD.n31 DGND 0.19fF $ **FLOATING
C5488 AVDD.n32 DGND 0.19fF $ **FLOATING
C5489 AVDD.n33 DGND 0.29fF $ **FLOATING
C5490 AVDD.n123 DGND 4.01fF $ **FLOATING
C5491 AVDD.n132 DGND 5.79fF $ **FLOATING
C5492 AVDD.t49 DGND 7.81fF
C5493 AVDD.n135 DGND 0.20fF $ **FLOATING
C5494 AVDD.n138 DGND 4.58fF $ **FLOATING
C5495 AVDD.t714 DGND 4.04fF
C5496 AVDD.n140 DGND 2.21fF $ **FLOATING
C5497 AVDD.n143 DGND 0.35fF $ **FLOATING
C5498 AVDD.n144 DGND 0.35fF $ **FLOATING
C5499 AVDD.n145 DGND 0.33fF $ **FLOATING
C5500 AVDD.n146 DGND 0.41fF $ **FLOATING
C5501 AVDD.n147 DGND 0.35fF $ **FLOATING
C5502 AVDD.n148 DGND 0.35fF $ **FLOATING
C5503 AVDD.n149 DGND 0.19fF $ **FLOATING
C5504 AVDD.n150 DGND 0.19fF $ **FLOATING
C5505 AVDD.n151 DGND 0.29fF $ **FLOATING
C5506 AVDD.n239 DGND 4.01fF $ **FLOATING
C5507 AVDD.n248 DGND 5.79fF $ **FLOATING
C5508 AVDD.t12 DGND 8.68fF
C5509 AVDD.n297 DGND 4.02fF $ **FLOATING
C5510 AVDD.n314 DGND 5.79fF $ **FLOATING
C5511 AVDD.t5 DGND 8.66fF
C5512 AVDD.n315 DGND 0.36fF $ **FLOATING
C5513 AVDD.n316 DGND 0.36fF $ **FLOATING
C5514 AVDD.n317 DGND 0.36fF $ **FLOATING
C5515 AVDD.n318 DGND 0.36fF $ **FLOATING
C5516 AVDD.n319 DGND 0.42fF $ **FLOATING
C5517 AVDD.n320 DGND 0.35fF $ **FLOATING
C5518 AVDD.n321 DGND 0.35fF $ **FLOATING
C5519 AVDD.n322 DGND 0.40fF $ **FLOATING
C5520 AVDD.n323 DGND 0.35fF $ **FLOATING
C5521 AVDD.n324 DGND 0.35fF $ **FLOATING
C5522 AVDD.n325 DGND 0.35fF $ **FLOATING
C5523 AVDD.n326 DGND 0.35fF $ **FLOATING
C5524 AVDD.n327 DGND 0.19fF $ **FLOATING
C5525 AVDD.n328 DGND 0.19fF $ **FLOATING
C5526 AVDD.n329 DGND 0.29fF $ **FLOATING
C5527 AVDD.n367 DGND 0.16fF $ **FLOATING
C5528 AVDD.n372 DGND 0.11fF $ **FLOATING
C5529 AVDD.t249 DGND 2.31fF
C5530 AVDD.n421 DGND 1.14fF $ **FLOATING
C5531 AVDD.n423 DGND 0.11fF $ **FLOATING
C5532 AVDD.n424 DGND 1.57fF $ **FLOATING
C5533 AVDD.t247 DGND 1.27fF
C5534 AVDD.n433 DGND 2.28fF $ **FLOATING
C5535 AVDD.t140 DGND 4.09fF
C5536 AVDD.t7 DGND 3.07fF
C5537 AVDD.n435 DGND 0.10fF $ **FLOATING
C5538 AVDD.n436 DGND 4.58fF $ **FLOATING
C5539 AVDD.n485 DGND 4.02fF $ **FLOATING
C5540 AVDD.n502 DGND 5.79fF $ **FLOATING
C5541 AVDD.t15 DGND 8.66fF
C5542 AVDD.n503 DGND 0.15fF $ **FLOATING
C5543 AVDD.n504 DGND 0.15fF $ **FLOATING
C5544 AVDD.n505 DGND 0.24fF $ **FLOATING
C5545 AVDD.n506 DGND 0.20fF $ **FLOATING
C5546 AVDD.n507 DGND 0.15fF $ **FLOATING
C5547 AVDD.n508 DGND 0.17fF $ **FLOATING
C5548 AVDD.n509 DGND 0.36fF $ **FLOATING
C5549 AVDD.n510 DGND 0.36fF $ **FLOATING
C5550 AVDD.n511 DGND 0.35fF $ **FLOATING
C5551 AVDD.n512 DGND 0.35fF $ **FLOATING
C5552 AVDD.n513 DGND 0.35fF $ **FLOATING
C5553 AVDD.n514 DGND 0.35fF $ **FLOATING
C5554 AVDD.n515 DGND 0.35fF $ **FLOATING
C5555 AVDD.n516 DGND 0.35fF $ **FLOATING
C5556 AVDD.n517 DGND 0.19fF $ **FLOATING
C5557 AVDD.n518 DGND 0.19fF $ **FLOATING
C5558 AVDD.n519 DGND 0.29fF $ **FLOATING
C5559 AVDD.t90 DGND 0.11fF
C5560 AVDD.n559 DGND 0.26fF $ **FLOATING
C5561 AVDD.n560 DGND 1.07fF $ **FLOATING
C5562 AVDD.n561 DGND 0.40fF $ **FLOATING
C5563 AVDD.n563 DGND 0.20fF $ **FLOATING
C5564 AVDD.n565 DGND 1.57fF $ **FLOATING
C5565 AVDD.t89 DGND 0.11fF
C5566 AVDD.n566 DGND 0.26fF $ **FLOATING
C5567 AVDD.n567 DGND 1.07fF $ **FLOATING
C5568 AVDD.n568 DGND 0.41fF $ **FLOATING
C5569 AVDD.n569 DGND 0.11fF $ **FLOATING
C5570 AVDD.n570 DGND 0.20fF $ **FLOATING
C5571 AVDD.n572 DGND 3.50fF $ **FLOATING
C5572 AVDD.n621 DGND 2.76fF $ **FLOATING
C5573 AVDD.n630 DGND 8.46fF $ **FLOATING
C5574 AVDD.t10 DGND 9.83fF
C5575 AVDD.n679 DGND 2.28fF $ **FLOATING
C5576 AVDD.t743 DGND 1.72fF
C5577 AVDD.n686 DGND 0.14fF $ **FLOATING
C5578 AVDD.n698 DGND 3.07fF $ **FLOATING
C5579 AVDD.n700 DGND 0.10fF $ **FLOATING
C5580 AVDD.n701 DGND 4.08fF $ **FLOATING
C5581 AVDD.t148 DGND 6.63fF
C5582 AVDD.n702 DGND 0.36fF $ **FLOATING
C5583 AVDD.n703 DGND 0.36fF $ **FLOATING
C5584 AVDD.n704 DGND 0.36fF $ **FLOATING
C5585 AVDD.n705 DGND 0.36fF $ **FLOATING
C5586 AVDD.n706 DGND 0.35fF $ **FLOATING
C5587 AVDD.n707 DGND 0.35fF $ **FLOATING
C5588 AVDD.n708 DGND 0.35fF $ **FLOATING
C5589 AVDD.n709 DGND 0.35fF $ **FLOATING
C5590 AVDD.n710 DGND 0.35fF $ **FLOATING
C5591 AVDD.n711 DGND 0.35fF $ **FLOATING
C5592 AVDD.n712 DGND 0.19fF $ **FLOATING
C5593 AVDD.n713 DGND 0.19fF $ **FLOATING
C5594 AVDD.n714 DGND 0.29fF $ **FLOATING
C5595 AVDD.n802 DGND 6.08fF $ **FLOATING
C5596 AVDD.n811 DGND 8.80fF $ **FLOATING
C5597 AVDD.t113 DGND 13.17fF
C5598 AVDD.n860 DGND 3.68fF $ **FLOATING
C5599 AVDD.n862 DGND 0.14fF $ **FLOATING
C5600 AVDD.n864 DGND 0.14fF $ **FLOATING
C5601 AVDD.n865 DGND 2.60fF $ **FLOATING
C5602 AVDD.n882 DGND 8.45fF $ **FLOATING
C5603 AVDD.t64 DGND 13.15fF
C5604 AVDD.n883 DGND 0.36fF $ **FLOATING
C5605 AVDD.n884 DGND 0.36fF $ **FLOATING
C5606 AVDD.n885 DGND 0.36fF $ **FLOATING
C5607 AVDD.n886 DGND 0.36fF $ **FLOATING
C5608 AVDD.n887 DGND 0.35fF $ **FLOATING
C5609 AVDD.n888 DGND 0.35fF $ **FLOATING
C5610 AVDD.n889 DGND 0.35fF $ **FLOATING
C5611 AVDD.n890 DGND 0.35fF $ **FLOATING
C5612 AVDD.n891 DGND 0.35fF $ **FLOATING
C5613 AVDD.n892 DGND 0.35fF $ **FLOATING
C5614 AVDD.n893 DGND 0.19fF $ **FLOATING
C5615 AVDD.n894 DGND 0.19fF $ **FLOATING
C5616 AVDD.n895 DGND 0.29fF $ **FLOATING
C5617 AVDD.n983 DGND 6.08fF $ **FLOATING
C5618 AVDD.n992 DGND 8.80fF $ **FLOATING
C5619 AVDD.t72 DGND 13.17fF
C5620 AVDD.n1041 DGND 6.11fF $ **FLOATING
C5621 AVDD.n1058 DGND 8.80fF $ **FLOATING
C5622 AVDD.t62 DGND 11.95fF
C5623 AVDD.n1059 DGND 8.36fF $ **FLOATING
C5624 AVDD.n1060 DGND 0.35fF $ **FLOATING
C5625 AVDD.n1061 DGND 0.35fF $ **FLOATING
C5626 AVDD.n1062 DGND 0.35fF $ **FLOATING
C5627 AVDD.n1063 DGND 0.35fF $ **FLOATING
C5628 AVDD.n1064 DGND 0.19fF $ **FLOATING
C5629 AVDD.n1065 DGND 0.19fF $ **FLOATING
C5630 AVDD.n1066 DGND 0.29fF $ **FLOATING
C5631 AVDD.t70 DGND 13.00fF
C5632 AVDD.n1146 DGND 6.11fF $ **FLOATING
C5633 AVDD.n1163 DGND 8.80fF $ **FLOATING
C5634 AVDD.t68 DGND 13.15fF
C5635 AVDD.n1164 DGND 0.36fF $ **FLOATING
C5636 AVDD.n1165 DGND 0.36fF $ **FLOATING
C5637 AVDD.t74 DGND 11.12fF
C5638 AVDD.n1166 DGND 0.13fF $ **FLOATING
C5639 AVDD.n1167 DGND 0.13fF $ **FLOATING
C5640 AVDD.n1168 DGND 0.13fF $ **FLOATING
C5641 AVDD.n1169 DGND 0.13fF $ **FLOATING
C5642 AVDD.n1170 DGND 0.13fF $ **FLOATING
C5643 AVDD.n1171 DGND 0.13fF $ **FLOATING
C5644 AVDD.n1172 DGND 0.13fF $ **FLOATING
C5645 AVDD.n1173 DGND 0.13fF $ **FLOATING
C5646 AVDD.n1174 DGND 0.50fF $ **FLOATING
C5647 AVDD.n1175 DGND 0.79fF $ **FLOATING
C5648 AVDD.n1176 DGND 0.13fF $ **FLOATING
C5649 AVDD.n1177 DGND 0.82fF $ **FLOATING
C5650 AVDD.n1178 DGND 0.13fF $ **FLOATING
C5651 AVDD.n1179 DGND 0.82fF $ **FLOATING
C5652 AVDD.n1180 DGND 0.13fF $ **FLOATING
C5653 AVDD.n1181 DGND 0.82fF $ **FLOATING
C5654 AVDD.n1182 DGND 0.13fF $ **FLOATING
C5655 AVDD.n1183 DGND 0.82fF $ **FLOATING
C5656 AVDD.n1184 DGND 0.13fF $ **FLOATING
C5657 AVDD.n1185 DGND 0.82fF $ **FLOATING
C5658 AVDD.n1186 DGND 0.13fF $ **FLOATING
C5659 AVDD.n1187 DGND 0.82fF $ **FLOATING
C5660 AVDD.n1188 DGND 0.13fF $ **FLOATING
C5661 AVDD.n1189 DGND 7.86fF $ **FLOATING
C5662 AVDD.n1190 DGND 0.82fF $ **FLOATING
C5663 AVDD.n1191 DGND 0.13fF $ **FLOATING
C5664 AVDD.n1192 DGND 0.82fF $ **FLOATING
C5665 AVDD.n1193 DGND 0.13fF $ **FLOATING
C5666 AVDD.n1194 DGND 0.13fF $ **FLOATING
C5667 AVDD.t394 DGND 6.22fF
C5668 AVDD.n1195 DGND 0.13fF $ **FLOATING
C5669 AVDD.n1196 DGND 0.64fF $ **FLOATING
C5670 AVDD.n1251 DGND 6.08fF $ **FLOATING
C5671 AVDD.n1260 DGND 4.64fF $ **FLOATING
C5672 AVDD.n1262 DGND 0.48fF $ **FLOATING
C5673 AVDD.n1263 DGND 0.13fF $ **FLOATING
C5674 AVDD.n1264 DGND 0.71fF $ **FLOATING
C5675 AVDD.n1265 DGND 1.17fF $ **FLOATING
C5676 AVDD.n1266 DGND 0.16fF $ **FLOATING
C5677 AVDD.n1267 DGND 0.32fF $ **FLOATING
C5678 AVDD.t138 DGND 0.11fF
C5679 AVDD.n1269 DGND 1.11fF $ **FLOATING
C5680 AVDD.n1270 DGND 0.26fF $ **FLOATING
C5681 AVDD.n1272 DGND 0.14fF $ **FLOATING
C5682 AVDD.t137 DGND 0.11fF
C5683 AVDD.n1273 DGND 1.12fF $ **FLOATING
C5684 AVDD.n1274 DGND 0.27fF $ **FLOATING
C5685 AVDD.n1277 DGND 0.14fF $ **FLOATING
C5686 AVDD.n1278 DGND 6.22fF $ **FLOATING
C5687 AVDD.n1295 DGND 2.76fF $ **FLOATING
C5688 AVDD.n1344 DGND 3.50fF $ **FLOATING
C5689 AVDD.n1347 DGND 0.20fF $ **FLOATING
C5690 AVDD.n1349 DGND 0.19fF $ **FLOATING
C5691 AVDD.n1351 DGND 0.94fF $ **FLOATING
C5692 AVDD.n1352 DGND 0.20fF $ **FLOATING
C5693 AVDD.n1354 DGND 0.20fF $ **FLOATING
C5694 AVDD.n1356 DGND 3.50fF $ **FLOATING
C5695 AVDD.n1406 DGND 5.19fF $ **FLOATING
C5696 AVDD.n1421 DGND 4.95fF $ **FLOATING
C5697 AVDD.n1423 DGND 0.51fF $ **FLOATING
C5698 AVDD.n1424 DGND 0.22fF $ **FLOATING
C5699 AVDD.n1425 DGND 0.77fF $ **FLOATING
C5700 AVDD.n1426 DGND 0.22fF $ **FLOATING
C5701 AVDD.n1427 DGND 0.14fF $ **FLOATING
C5702 AVDD.n1428 DGND 0.22fF $ **FLOATING
C5703 AVDD.n1429 DGND 0.22fF $ **FLOATING
C5704 AVDD.n1430 DGND 0.22fF $ **FLOATING
C5705 AVDD.n1431 DGND 0.77fF $ **FLOATING
C5706 AVDD.n1432 DGND 0.22fF $ **FLOATING
C5707 AVDD.n1433 DGND 0.14fF $ **FLOATING
C5708 AVDD.n1434 DGND 0.22fF $ **FLOATING
C5709 AVDD.n1435 DGND 0.77fF $ **FLOATING
C5710 AVDD.n1436 DGND 0.22fF $ **FLOATING
C5711 AVDD.n1437 DGND 0.14fF $ **FLOATING
C5712 AVDD.n1438 DGND 0.22fF $ **FLOATING
C5713 AVDD.n1439 DGND 0.22fF $ **FLOATING
C5714 AVDD.n1440 DGND 0.77fF $ **FLOATING
C5715 AVDD.n1441 DGND 0.22fF $ **FLOATING
C5716 AVDD.n1442 DGND 0.14fF $ **FLOATING
C5717 AVDD.n1443 DGND 0.22fF $ **FLOATING
C5718 AVDD.n1444 DGND 0.20fF $ **FLOATING
C5719 AVDD.n1445 DGND 0.77fF $ **FLOATING
C5720 AVDD.n1446 DGND 0.22fF $ **FLOATING
C5721 AVDD.n1447 DGND 0.14fF $ **FLOATING
C5722 AVDD.n1448 DGND 0.22fF $ **FLOATING
C5723 AVDD.n1449 DGND 0.22fF $ **FLOATING
C5724 AVDD.n1450 DGND 0.77fF $ **FLOATING
C5725 AVDD.n1451 DGND 0.22fF $ **FLOATING
C5726 AVDD.n1452 DGND 0.14fF $ **FLOATING
C5727 AVDD.n1453 DGND 0.22fF $ **FLOATING
C5728 AVDD.n1454 DGND 0.22fF $ **FLOATING
C5729 AVDD.n1455 DGND 0.77fF $ **FLOATING
C5730 AVDD.n1456 DGND 0.22fF $ **FLOATING
C5731 AVDD.n1457 DGND 0.14fF $ **FLOATING
C5732 AVDD.n1458 DGND 0.22fF $ **FLOATING
C5733 AVDD.n1459 DGND 0.77fF $ **FLOATING
C5734 AVDD.n1460 DGND 0.22fF $ **FLOATING
C5735 AVDD.n1461 DGND 0.14fF $ **FLOATING
C5736 AVDD.t125 DGND 10.81fF
C5737 AVDD.n1462 DGND 0.22fF $ **FLOATING
C5738 AVDD.n1463 DGND 0.19fF $ **FLOATING
C5739 AVDD.n1464 DGND 0.75fF $ **FLOATING
C5740 AVDD.n1465 DGND 0.21fF $ **FLOATING
C5741 AVDD.n1466 DGND 0.14fF $ **FLOATING
C5742 AVDD.n1467 DGND 6.19fF $ **FLOATING
C5743 AVDD.n1468 DGND 0.14fF $ **FLOATING
C5744 AVDD.n1469 DGND 0.55fF $ **FLOATING
C5745 AVDD.t452 DGND 0.46fF
C5746 AVDD.n1470 DGND 1.36fF $ **FLOATING
C5747 AVDD.t566 DGND 0.46fF
C5748 AVDD.n1471 DGND 0.64fF $ **FLOATING
C5749 AVDD.n1526 DGND 6.08fF $ **FLOATING
C5750 AVDD.n1535 DGND 8.80fF $ **FLOATING
C5751 AVDD.n1537 DGND 1.08fF $ **FLOATING
C5752 AVDD.n1538 DGND 1.37fF $ **FLOATING
C5753 AVDD.t76 DGND 10.85fF
C5754 AVDD.t680 DGND 0.46fF
C5755 AVDD.n1539 DGND 0.81fF $ **FLOATING
C5756 AVDD.n1540 DGND 0.19fF $ **FLOATING
C5757 AVDD.n1541 DGND 0.14fF $ **FLOATING
C5758 AVDD.n1543 DGND 0.14fF $ **FLOATING
C5759 AVDD.n1545 DGND 0.14fF $ **FLOATING
C5760 AVDD.n1547 DGND 0.14fF $ **FLOATING
C5761 AVDD.n1549 DGND 0.14fF $ **FLOATING
C5762 AVDD.n1551 DGND 0.14fF $ **FLOATING
C5763 AVDD.n1553 DGND 0.14fF $ **FLOATING
C5764 AVDD.n1555 DGND 0.14fF $ **FLOATING
C5765 AVDD.n1557 DGND 0.14fF $ **FLOATING
C5766 AVDD.n1558 DGND 6.96fF $ **FLOATING
C5767 AVDD.n1559 DGND 0.14fF $ **FLOATING
C5768 AVDD.n1560 DGND 0.55fF $ **FLOATING
C5769 AVDD.n1561 DGND 0.65fF $ **FLOATING
C5770 AVDD.n1610 DGND 6.11fF $ **FLOATING
C5771 AVDD.n1625 DGND 8.80fF $ **FLOATING
C5772 AVDD.n1627 DGND 1.11fF $ **FLOATING
C5773 AVDD.n1628 DGND 1.40fF $ **FLOATING
C5774 AVDD.t81 DGND 11.18fF
C5775 AVDD.t545 DGND 0.46fF
C5776 AVDD.n1629 DGND 0.81fF $ **FLOATING
C5777 AVDD.n1630 DGND 0.19fF $ **FLOATING
C5778 AVDD.n1631 DGND 0.14fF $ **FLOATING
C5779 AVDD.t404 DGND 0.46fF
C5780 AVDD.n1632 DGND 0.84fF $ **FLOATING
C5781 AVDD.n1633 DGND 0.24fF $ **FLOATING
C5782 AVDD.t599 DGND 0.46fF
C5783 AVDD.n1634 DGND 0.84fF $ **FLOATING
C5784 AVDD.n1635 DGND 0.24fF $ **FLOATING
C5785 AVDD.t638 DGND 0.46fF
C5786 AVDD.n1636 DGND 0.84fF $ **FLOATING
C5787 AVDD.n1637 DGND 0.24fF $ **FLOATING
C5788 AVDD.t497 DGND 0.46fF
C5789 AVDD.n1638 DGND 0.84fF $ **FLOATING
C5790 AVDD.n1639 DGND 0.24fF $ **FLOATING
C5791 AVDD.t683 DGND 0.46fF
C5792 AVDD.n1640 DGND 0.84fF $ **FLOATING
C5793 AVDD.n1641 DGND 0.24fF $ **FLOATING
C5794 AVDD.t527 DGND 0.46fF
C5795 AVDD.n1642 DGND 0.84fF $ **FLOATING
C5796 AVDD.n1643 DGND 0.24fF $ **FLOATING
C5797 AVDD.t393 DGND 0.46fF
C5798 AVDD.n1644 DGND 0.84fF $ **FLOATING
C5799 AVDD.n1645 DGND 0.24fF $ **FLOATING
C5800 AVDD.t590 DGND 0.46fF
C5801 AVDD.n1646 DGND 0.84fF $ **FLOATING
C5802 AVDD.n1647 DGND 0.24fF $ **FLOATING
C5803 AVDD.n1648 DGND 6.96fF $ **FLOATING
C5804 AVDD.n1649 DGND 0.14fF $ **FLOATING
C5805 AVDD.n1650 DGND 0.52fF $ **FLOATING
C5806 AVDD.n1651 DGND 0.36fF $ **FLOATING
C5807 AVDD.n1652 DGND 0.36fF $ **FLOATING
C5808 AVDD.n1653 DGND 0.35fF $ **FLOATING
C5809 AVDD.n1654 DGND 0.35fF $ **FLOATING
C5810 AVDD.n1655 DGND 0.36fF $ **FLOATING
C5811 AVDD.n1656 DGND 0.36fF $ **FLOATING
C5812 AVDD.t686 DGND 0.46fF
C5813 AVDD.n1657 DGND 0.61fF $ **FLOATING
C5814 AVDD.n1658 DGND 0.33fF $ **FLOATING
C5815 AVDD.n1707 DGND 3.81fF $ **FLOATING
C5816 AVDD.t485 DGND 0.46fF
C5817 AVDD.n1708 DGND 0.81fF $ **FLOATING
C5818 AVDD.n1709 DGND 0.19fF $ **FLOATING
C5819 AVDD.n1710 DGND 0.14fF $ **FLOATING
C5820 AVDD.n1712 DGND 0.14fF $ **FLOATING
C5821 AVDD.n1714 DGND 0.14fF $ **FLOATING
C5822 AVDD.n1716 DGND 0.14fF $ **FLOATING
C5823 AVDD.n1718 DGND 0.14fF $ **FLOATING
C5824 AVDD.n1720 DGND 0.14fF $ **FLOATING
C5825 AVDD.n1722 DGND 0.14fF $ **FLOATING
C5826 AVDD.n1724 DGND 0.14fF $ **FLOATING
C5827 AVDD.n1726 DGND 0.14fF $ **FLOATING
C5828 AVDD.n1727 DGND 2.58fF $ **FLOATING
C5829 AVDD.n1728 DGND 0.14fF $ **FLOATING
C5830 AVDD.n1729 DGND 0.27fF $ **FLOATING
C5831 AVDD.n1744 DGND 4.29fF $ **FLOATING
C5832 AVDD.n1746 DGND 0.44fF $ **FLOATING
C5833 AVDD.t85 DGND 11.16fF
C5834 AVDD.n1747 DGND 0.81fF $ **FLOATING
C5835 AVDD.n1748 DGND 0.19fF $ **FLOATING
C5836 AVDD.n1749 DGND 0.14fF $ **FLOATING
C5837 AVDD.n1751 DGND 0.14fF $ **FLOATING
C5838 AVDD.n1753 DGND 0.14fF $ **FLOATING
C5839 AVDD.n1755 DGND 0.14fF $ **FLOATING
C5840 AVDD.n1757 DGND 0.14fF $ **FLOATING
C5841 AVDD.n1759 DGND 0.14fF $ **FLOATING
C5842 AVDD.n1761 DGND 0.14fF $ **FLOATING
C5843 AVDD.n1763 DGND 0.14fF $ **FLOATING
C5844 AVDD.n1765 DGND 0.14fF $ **FLOATING
C5845 AVDD.n1766 DGND 6.22fF $ **FLOATING
C5846 AVDD.n1767 DGND 0.14fF $ **FLOATING
C5847 AVDD.n1768 DGND 0.52fF $ **FLOATING
C5848 AVDD.n1769 DGND 1.40fF $ **FLOATING
C5849 AVDD.n1770 DGND 0.65fF $ **FLOATING
C5850 AVDD.n1819 DGND 6.11fF $ **FLOATING
C5851 AVDD.n1834 DGND 4.99fF $ **FLOATING
C5852 AVDD.n1836 DGND 0.52fF $ **FLOATING
C5853 AVDD.n1838 DGND 0.13fF $ **FLOATING
C5854 AVDD.n1840 DGND 0.13fF $ **FLOATING
C5855 AVDD.n1842 DGND 0.13fF $ **FLOATING
C5856 AVDD.n1844 DGND 0.13fF $ **FLOATING
C5857 AVDD.n1846 DGND 0.13fF $ **FLOATING
C5858 AVDD.n1848 DGND 0.13fF $ **FLOATING
C5859 AVDD.n1850 DGND 0.13fF $ **FLOATING
C5860 AVDD.n1852 DGND 0.13fF $ **FLOATING
C5861 AVDD.n1853 DGND 1.19fF $ **FLOATING
C5862 AVDD.n1854 DGND 0.13fF $ **FLOATING
C5863 AVDD.t103 DGND 10.77fF
C5864 AVDD.n1856 DGND 0.13fF $ **FLOATING
C5865 AVDD.n1858 DGND 0.13fF $ **FLOATING
C5866 AVDD.n1860 DGND 0.13fF $ **FLOATING
C5867 AVDD.n1862 DGND 0.13fF $ **FLOATING
C5868 AVDD.n1864 DGND 0.13fF $ **FLOATING
C5869 AVDD.n1866 DGND 0.13fF $ **FLOATING
C5870 AVDD.n1868 DGND 0.13fF $ **FLOATING
C5871 AVDD.n1870 DGND 0.13fF $ **FLOATING
C5872 AVDD.n1872 DGND 0.13fF $ **FLOATING
C5873 AVDD.t34 DGND 6.19fF
C5874 AVDD.n1873 DGND 0.13fF $ **FLOATING
C5875 AVDD.n1874 DGND 0.13fF $ **FLOATING
C5876 AVDD.n1875 DGND 1.56fF $ **FLOATING
C5877 AVDD.n1877 DGND 0.13fF $ **FLOATING
C5878 AVDD.n1879 DGND 0.13fF $ **FLOATING
C5879 AVDD.n1881 DGND 0.13fF $ **FLOATING
C5880 AVDD.n1883 DGND 0.13fF $ **FLOATING
C5881 AVDD.n1885 DGND 0.13fF $ **FLOATING
C5882 AVDD.n1887 DGND 0.13fF $ **FLOATING
C5883 AVDD.n1889 DGND 0.13fF $ **FLOATING
C5884 AVDD.n1891 DGND 0.13fF $ **FLOATING
C5885 AVDD.t66 DGND 10.81fF
C5886 AVDD.n1893 DGND 0.13fF $ **FLOATING
C5887 AVDD.n1894 DGND 1.19fF $ **FLOATING
C5888 AVDD.n1895 DGND 0.13fF $ **FLOATING
C5889 AVDD.n1897 DGND 0.13fF $ **FLOATING
C5890 AVDD.n1899 DGND 0.13fF $ **FLOATING
C5891 AVDD.n1901 DGND 0.13fF $ **FLOATING
C5892 AVDD.n1903 DGND 0.13fF $ **FLOATING
C5893 AVDD.n1905 DGND 0.13fF $ **FLOATING
C5894 AVDD.n1907 DGND 0.13fF $ **FLOATING
C5895 AVDD.n1909 DGND 0.13fF $ **FLOATING
C5896 AVDD.n1911 DGND 0.13fF $ **FLOATING
C5897 AVDD.t24 DGND 6.96fF
C5898 AVDD.n1912 DGND 0.13fF $ **FLOATING
C5899 AVDD.n1913 DGND 0.64fF $ **FLOATING
C5900 AVDD.n1968 DGND 6.08fF $ **FLOATING
C5901 AVDD.n1977 DGND 8.80fF $ **FLOATING
C5902 AVDD.n1979 DGND 1.38fF $ **FLOATING
C5903 AVDD.n1980 DGND 0.13fF $ **FLOATING
C5904 AVDD.n1981 DGND 1.56fF $ **FLOATING
C5905 AVDD.n1982 DGND 0.37fF $ **FLOATING
C5906 AVDD.n2031 DGND 6.11fF $ **FLOATING
C5907 AVDD.n2046 DGND 8.80fF $ **FLOATING
C5908 AVDD.n2048 DGND 1.62fF $ **FLOATING
C5909 AVDD.t449 DGND 0.29fF
C5910 AVDD.n2049 DGND 0.32fF $ **FLOATING
C5911 AVDD.n2050 DGND 0.47fF $ **FLOATING
C5912 AVDD.t617 DGND 0.29fF
C5913 AVDD.t572 DGND 0.29fF
C5914 AVDD.n2051 DGND 0.34fF $ **FLOATING
C5915 AVDD.n2052 DGND 0.34fF $ **FLOATING
C5916 AVDD.n2053 DGND 0.52fF $ **FLOATING
C5917 AVDD.n2054 DGND 0.11fF $ **FLOATING
C5918 AVDD.n2055 DGND 0.28fF $ **FLOATING
C5919 AVDD.n2056 DGND 0.28fF $ **FLOATING
C5920 AVDD.t413 DGND 0.29fF
C5921 AVDD.n2057 DGND 0.33fF $ **FLOATING
C5922 AVDD.n2058 DGND 0.47fF $ **FLOATING
C5923 AVDD.n2060 DGND 0.59fF $ **FLOATING
C5924 AVDD.n2061 DGND 0.52fF $ **FLOATING
C5925 AVDD.n2110 DGND 6.11fF $ **FLOATING
C5926 AVDD.n2125 DGND 5.03fF $ **FLOATING
C5927 AVDD.n2127 DGND 0.31fF $ **FLOATING
C5928 AVDD.n2128 DGND 0.81fF $ **FLOATING
C5929 AVDD.n2129 DGND 0.19fF $ **FLOATING
C5930 AVDD.n2130 DGND 0.14fF $ **FLOATING
C5931 AVDD.n2132 DGND 0.14fF $ **FLOATING
C5932 AVDD.n2134 DGND 0.14fF $ **FLOATING
C5933 AVDD.n2136 DGND 0.14fF $ **FLOATING
C5934 AVDD.n2138 DGND 0.14fF $ **FLOATING
C5935 AVDD.n2140 DGND 0.14fF $ **FLOATING
C5936 AVDD.n2142 DGND 0.14fF $ **FLOATING
C5937 AVDD.n2144 DGND 0.14fF $ **FLOATING
C5938 AVDD.n2146 DGND 0.14fF $ **FLOATING
C5939 AVDD.n2147 DGND 6.19fF $ **FLOATING
C5940 AVDD.n2148 DGND 0.14fF $ **FLOATING
C5941 AVDD.n2149 DGND 0.69fF $ **FLOATING
C5942 AVDD.t130 DGND 4.29fF
C5943 AVDD.n2150 DGND 0.81fF $ **FLOATING
C5944 AVDD.n2151 DGND 0.19fF $ **FLOATING
C5945 AVDD.n2152 DGND 0.14fF $ **FLOATING
C5946 AVDD.n2154 DGND 0.14fF $ **FLOATING
C5947 AVDD.n2156 DGND 0.14fF $ **FLOATING
C5948 AVDD.n2158 DGND 0.14fF $ **FLOATING
C5949 AVDD.n2160 DGND 0.14fF $ **FLOATING
C5950 AVDD.n2162 DGND 0.14fF $ **FLOATING
C5951 AVDD.n2164 DGND 0.14fF $ **FLOATING
C5952 AVDD.n2166 DGND 0.14fF $ **FLOATING
C5953 AVDD.n2168 DGND 0.14fF $ **FLOATING
C5954 AVDD.n2169 DGND 6.96fF $ **FLOATING
C5955 AVDD.n2170 DGND 0.14fF $ **FLOATING
C5956 AVDD.n2171 DGND 0.75fF $ **FLOATING
C5957 AVDD.t491 DGND 0.46fF
C5958 AVDD.n2172 DGND 0.91fF $ **FLOATING
C5959 AVDD.n2174 DGND 0.13fF $ **FLOATING
C5960 AVDD.n2176 DGND 0.13fF $ **FLOATING
C5961 AVDD.n2178 DGND 0.13fF $ **FLOATING
C5962 AVDD.n2180 DGND 0.13fF $ **FLOATING
C5963 AVDD.n2182 DGND 0.13fF $ **FLOATING
C5964 AVDD.n2184 DGND 0.13fF $ **FLOATING
C5965 AVDD.n2186 DGND 0.13fF $ **FLOATING
C5966 AVDD.n2188 DGND 0.13fF $ **FLOATING
C5967 AVDD.n2189 DGND 1.19fF $ **FLOATING
C5968 AVDD.n2190 DGND 0.13fF $ **FLOATING
C5969 AVDD.n2239 DGND 3.76fF $ **FLOATING
C5970 AVDD.n2241 DGND 0.13fF $ **FLOATING
C5971 AVDD.n2243 DGND 0.13fF $ **FLOATING
C5972 AVDD.n2245 DGND 0.13fF $ **FLOATING
C5973 AVDD.n2247 DGND 0.13fF $ **FLOATING
C5974 AVDD.n2249 DGND 0.13fF $ **FLOATING
C5975 AVDD.n2251 DGND 0.13fF $ **FLOATING
C5976 AVDD.n2253 DGND 0.13fF $ **FLOATING
C5977 AVDD.n2255 DGND 0.13fF $ **FLOATING
C5978 AVDD.n2257 DGND 0.13fF $ **FLOATING
C5979 AVDD.t42 DGND 2.58fF
C5980 AVDD.n2258 DGND 0.13fF $ **FLOATING
C5981 AVDD.n2259 DGND 0.40fF $ **FLOATING
C5982 AVDD.n2260 DGND 0.13fF $ **FLOATING
C5983 AVDD.n2261 DGND 0.47fF $ **FLOATING
C5984 AVDD.n2276 DGND 8.53fF $ **FLOATING
C5985 AVDD.n2278 DGND 1.60fF $ **FLOATING
C5986 AVDD.n2279 DGND 0.36fF $ **FLOATING
C5987 AVDD.n2280 DGND 0.36fF $ **FLOATING
C5988 AVDD.n2281 DGND 0.36fF $ **FLOATING
C5989 AVDD.n2282 DGND 0.36fF $ **FLOATING
C5990 AVDD.n2283 DGND 0.35fF $ **FLOATING
C5991 AVDD.n2284 DGND 0.35fF $ **FLOATING
C5992 AVDD.t605 DGND 0.46fF
C5993 AVDD.n2285 DGND 0.64fF $ **FLOATING
C5994 AVDD.n2340 DGND 6.08fF $ **FLOATING
C5995 AVDD.n2349 DGND 8.80fF $ **FLOATING
C5996 AVDD.n2351 DGND 0.62fF $ **FLOATING
C5997 AVDD.n2352 DGND 0.92fF $ **FLOATING
C5998 AVDD.t377 DGND 0.46fF
C5999 AVDD.n2353 DGND 0.81fF $ **FLOATING
C6000 AVDD.n2354 DGND 0.19fF $ **FLOATING
C6001 AVDD.n2355 DGND 0.14fF $ **FLOATING
C6002 AVDD.t91 DGND 6.48fF
C6003 AVDD.n2357 DGND 0.14fF $ **FLOATING
C6004 AVDD.n2359 DGND 0.14fF $ **FLOATING
C6005 AVDD.n2361 DGND 0.14fF $ **FLOATING
C6006 AVDD.n2363 DGND 0.14fF $ **FLOATING
C6007 AVDD.n2365 DGND 0.14fF $ **FLOATING
C6008 AVDD.n2367 DGND 0.14fF $ **FLOATING
C6009 AVDD.n2369 DGND 0.14fF $ **FLOATING
C6010 AVDD.n2371 DGND 0.14fF $ **FLOATING
C6011 AVDD.n2372 DGND 4.55fF $ **FLOATING
C6012 AVDD.n2373 DGND 0.14fF $ **FLOATING
C6013 AVDD.n2374 DGND 0.75fF $ **FLOATING
C6014 AVDD.t596 DGND 0.46fF
C6015 AVDD.n2375 DGND 0.81fF $ **FLOATING
C6016 AVDD.n2376 DGND 0.19fF $ **FLOATING
C6017 AVDD.n2377 DGND 0.14fF $ **FLOATING
C6018 AVDD.n2379 DGND 0.14fF $ **FLOATING
C6019 AVDD.n2381 DGND 0.14fF $ **FLOATING
C6020 AVDD.n2383 DGND 0.14fF $ **FLOATING
C6021 AVDD.n2385 DGND 0.14fF $ **FLOATING
C6022 AVDD.n2387 DGND 0.14fF $ **FLOATING
C6023 AVDD.n2389 DGND 0.14fF $ **FLOATING
C6024 AVDD.n2391 DGND 0.14fF $ **FLOATING
C6025 AVDD.n2393 DGND 0.14fF $ **FLOATING
C6026 AVDD.n2394 DGND 6.70fF $ **FLOATING
C6027 AVDD.n2395 DGND 0.14fF $ **FLOATING
C6028 AVDD.n2396 DGND 0.69fF $ **FLOATING
C6029 AVDD.n2397 DGND 0.65fF $ **FLOATING
C6030 AVDD.n2446 DGND 6.11fF $ **FLOATING
C6031 AVDD.n2461 DGND 8.80fF $ **FLOATING
C6032 AVDD.n2463 DGND 1.56fF $ **FLOATING
C6033 AVDD.n2464 DGND 1.61fF $ **FLOATING
C6034 AVDD.n2465 DGND 0.52fF $ **FLOATING
C6035 AVDD.n2466 DGND 0.36fF $ **FLOATING
C6036 AVDD.n2467 DGND 0.28fF $ **FLOATING
C6037 AVDD.n2468 DGND 0.11fF $ **FLOATING
C6038 AVDD.t653 DGND 0.29fF
C6039 AVDD.n2469 DGND 0.33fF $ **FLOATING
C6040 AVDD.n2470 DGND 0.52fF $ **FLOATING
C6041 AVDD.n2471 DGND 0.40fF $ **FLOATING
C6042 AVDD.n2520 DGND 3.72fF $ **FLOATING
C6043 AVDD.n2521 DGND 0.64fF $ **FLOATING
C6044 AVDD.n2522 DGND 0.19fF $ **FLOATING
C6045 AVDD.n2523 DGND 0.14fF $ **FLOATING
C6046 AVDD.n2525 DGND 0.14fF $ **FLOATING
C6047 AVDD.n2527 DGND 0.14fF $ **FLOATING
C6048 AVDD.n2529 DGND 0.14fF $ **FLOATING
C6049 AVDD.n2531 DGND 0.14fF $ **FLOATING
C6050 AVDD.n2533 DGND 0.14fF $ **FLOATING
C6051 AVDD.n2535 DGND 0.14fF $ **FLOATING
C6052 AVDD.n2537 DGND 0.14fF $ **FLOATING
C6053 AVDD.n2539 DGND 0.14fF $ **FLOATING
C6054 AVDD.n2540 DGND 2.58fF $ **FLOATING
C6055 AVDD.n2541 DGND 0.14fF $ **FLOATING
C6056 AVDD.n2542 DGND 0.27fF $ **FLOATING
C6057 AVDD.n2557 DGND 8.58fF $ **FLOATING
C6058 AVDD.n2559 DGND 0.31fF $ **FLOATING
C6059 AVDD.n2560 DGND 1.61fF $ **FLOATING
C6060 AVDD.n2561 DGND 0.65fF $ **FLOATING
C6061 AVDD.n2610 DGND 6.11fF $ **FLOATING
C6062 AVDD.n2625 DGND 8.80fF $ **FLOATING
C6063 AVDD.n2627 DGND 0.97fF $ **FLOATING
C6064 AVDD.t14 DGND 6.76fF
C6065 AVDD.n2629 DGND 0.13fF $ **FLOATING
C6066 AVDD.n2631 DGND 0.13fF $ **FLOATING
C6067 AVDD.n2633 DGND 0.13fF $ **FLOATING
C6068 AVDD.n2635 DGND 0.13fF $ **FLOATING
C6069 AVDD.n2637 DGND 0.13fF $ **FLOATING
C6070 AVDD.n2639 DGND 0.13fF $ **FLOATING
C6071 AVDD.n2641 DGND 0.13fF $ **FLOATING
C6072 AVDD.n2643 DGND 0.13fF $ **FLOATING
C6073 AVDD.n2644 DGND 0.50fF $ **FLOATING
C6074 AVDD.n2645 DGND 0.88fF $ **FLOATING
C6075 AVDD.n2646 DGND 0.13fF $ **FLOATING
C6076 AVDD.n2648 DGND 0.13fF $ **FLOATING
C6077 AVDD.n2650 DGND 0.13fF $ **FLOATING
C6078 AVDD.n2652 DGND 0.13fF $ **FLOATING
C6079 AVDD.n2654 DGND 0.13fF $ **FLOATING
C6080 AVDD.n2656 DGND 0.13fF $ **FLOATING
C6081 AVDD.n2658 DGND 0.13fF $ **FLOATING
C6082 AVDD.n2660 DGND 0.13fF $ **FLOATING
C6083 AVDD.n2662 DGND 0.13fF $ **FLOATING
C6084 AVDD.n2664 DGND 0.13fF $ **FLOATING
C6085 AVDD.t23 DGND 6.96fF
C6086 AVDD.n2665 DGND 0.13fF $ **FLOATING
C6087 AVDD.n2666 DGND 0.13fF $ **FLOATING
C6088 AVDD.n2667 DGND 1.56fF $ **FLOATING
C6089 AVDD.n2668 DGND 0.36fF $ **FLOATING
C6090 AVDD.n2669 DGND 0.36fF $ **FLOATING
C6091 AVDD.n2670 DGND 0.35fF $ **FLOATING
C6092 AVDD.n2671 DGND 0.35fF $ **FLOATING
C6093 AVDD.n2672 DGND 0.36fF $ **FLOATING
C6094 AVDD.n2674 DGND 0.13fF $ **FLOATING
C6095 AVDD.n2676 DGND 0.13fF $ **FLOATING
C6096 AVDD.n2678 DGND 0.13fF $ **FLOATING
C6097 AVDD.n2680 DGND 0.13fF $ **FLOATING
C6098 AVDD.n2682 DGND 0.13fF $ **FLOATING
C6099 AVDD.n2684 DGND 0.13fF $ **FLOATING
C6100 AVDD.n2686 DGND 0.13fF $ **FLOATING
C6101 AVDD.n2688 DGND 0.13fF $ **FLOATING
C6102 AVDD.n2689 DGND 1.19fF $ **FLOATING
C6103 AVDD.n2690 DGND 0.13fF $ **FLOATING
C6104 AVDD.t208 DGND 6.43fF
C6105 AVDD.n2692 DGND 0.13fF $ **FLOATING
C6106 AVDD.n2694 DGND 0.13fF $ **FLOATING
C6107 AVDD.n2696 DGND 0.13fF $ **FLOATING
C6108 AVDD.n2698 DGND 0.13fF $ **FLOATING
C6109 AVDD.n2700 DGND 0.13fF $ **FLOATING
C6110 AVDD.n2702 DGND 0.13fF $ **FLOATING
C6111 AVDD.n2704 DGND 0.13fF $ **FLOATING
C6112 AVDD.n2706 DGND 0.13fF $ **FLOATING
C6113 AVDD.n2708 DGND 0.13fF $ **FLOATING
C6114 AVDD.t46 DGND 6.96fF
C6115 AVDD.n2709 DGND 0.13fF $ **FLOATING
C6116 AVDD.n2710 DGND 0.64fF $ **FLOATING
C6117 AVDD.n2765 DGND 6.08fF $ **FLOATING
C6118 AVDD.n2774 DGND 8.80fF $ **FLOATING
C6119 AVDD.n2776 DGND 0.93fF $ **FLOATING
C6120 AVDD.n2777 DGND 0.13fF $ **FLOATING
C6121 AVDD.n2778 DGND 1.56fF $ **FLOATING
C6122 AVDD.n2779 DGND 0.44fF $ **FLOATING
C6123 AVDD.n2828 DGND 4.07fF $ **FLOATING
C6124 AVDD.n2829 DGND 0.81fF $ **FLOATING
C6125 AVDD.n2830 DGND 0.19fF $ **FLOATING
C6126 AVDD.n2831 DGND 0.14fF $ **FLOATING
C6127 AVDD.n2833 DGND 0.14fF $ **FLOATING
C6128 AVDD.n2835 DGND 0.14fF $ **FLOATING
C6129 AVDD.n2837 DGND 0.14fF $ **FLOATING
C6130 AVDD.n2839 DGND 0.14fF $ **FLOATING
C6131 AVDD.n2841 DGND 0.14fF $ **FLOATING
C6132 AVDD.n2843 DGND 0.14fF $ **FLOATING
C6133 AVDD.n2845 DGND 0.14fF $ **FLOATING
C6134 AVDD.n2847 DGND 0.14fF $ **FLOATING
C6135 AVDD.n2848 DGND 2.60fF $ **FLOATING
C6136 AVDD.n2849 DGND 0.14fF $ **FLOATING
C6137 AVDD.n2850 DGND 0.27fF $ **FLOATING
C6138 AVDD.n2865 DGND 8.23fF $ **FLOATING
C6139 AVDD.n2867 DGND 0.31fF $ **FLOATING
C6140 AVDD.t671 DGND 0.46fF
C6141 AVDD.n2868 DGND 1.61fF $ **FLOATING
C6142 AVDD.n2869 DGND 0.36fF $ **FLOATING
C6143 AVDD.n2870 DGND 0.36fF $ **FLOATING
C6144 AVDD.n2871 DGND 0.35fF $ **FLOATING
C6145 AVDD.n2872 DGND 0.35fF $ **FLOATING
C6146 AVDD.t611 DGND 0.46fF
C6147 AVDD.n2873 DGND 0.64fF $ **FLOATING
C6148 AVDD.n2928 DGND 6.08fF $ **FLOATING
C6149 AVDD.n2937 DGND 8.80fF $ **FLOATING
C6150 AVDD.n2939 DGND 1.53fF $ **FLOATING
C6151 AVDD.n2940 DGND 1.61fF $ **FLOATING
C6152 AVDD.n2941 DGND 0.65fF $ **FLOATING
C6153 AVDD.n2990 DGND 6.11fF $ **FLOATING
C6154 AVDD.n3005 DGND 8.80fF $ **FLOATING
C6155 AVDD.n3007 DGND 0.66fF $ **FLOATING
C6156 AVDD.n3008 DGND 0.95fF $ **FLOATING
C6157 AVDD.t161 DGND 6.81fF
C6158 AVDD.t467 DGND 0.46fF
C6159 AVDD.n3009 DGND 0.81fF $ **FLOATING
C6160 AVDD.n3010 DGND 0.19fF $ **FLOATING
C6161 AVDD.n3011 DGND 0.14fF $ **FLOATING
C6162 AVDD.n3013 DGND 0.14fF $ **FLOATING
C6163 AVDD.n3015 DGND 0.14fF $ **FLOATING
C6164 AVDD.n3017 DGND 0.14fF $ **FLOATING
C6165 AVDD.n3019 DGND 0.14fF $ **FLOATING
C6166 AVDD.n3021 DGND 0.14fF $ **FLOATING
C6167 AVDD.n3023 DGND 0.14fF $ **FLOATING
C6168 AVDD.n3025 DGND 0.14fF $ **FLOATING
C6169 AVDD.n3027 DGND 0.14fF $ **FLOATING
C6170 AVDD.n3028 DGND 4.90fF $ **FLOATING
C6171 AVDD.n3029 DGND 0.14fF $ **FLOATING
C6172 AVDD.n3030 DGND 0.75fF $ **FLOATING
C6173 AVDD.t387 DGND 0.46fF
C6174 AVDD.n3031 DGND 0.81fF $ **FLOATING
C6175 AVDD.n3032 DGND 0.19fF $ **FLOATING
C6176 AVDD.n3033 DGND 0.14fF $ **FLOATING
C6177 AVDD.n3035 DGND 0.14fF $ **FLOATING
C6178 AVDD.n3037 DGND 0.14fF $ **FLOATING
C6179 AVDD.n3039 DGND 0.14fF $ **FLOATING
C6180 AVDD.n3041 DGND 0.14fF $ **FLOATING
C6181 AVDD.n3043 DGND 0.14fF $ **FLOATING
C6182 AVDD.n3045 DGND 0.14fF $ **FLOATING
C6183 AVDD.n3047 DGND 0.14fF $ **FLOATING
C6184 AVDD.n3049 DGND 0.14fF $ **FLOATING
C6185 AVDD.n3050 DGND 6.35fF $ **FLOATING
C6186 AVDD.n3051 DGND 0.14fF $ **FLOATING
C6187 AVDD.n3052 DGND 0.66fF $ **FLOATING
C6188 AVDD.t397 DGND 0.46fF
C6189 AVDD.n3053 DGND 0.55fF $ **FLOATING
C6190 AVDD.n3054 DGND 0.51fF $ **FLOATING
C6191 AVDD.n3109 DGND 6.08fF $ **FLOATING
C6192 AVDD.n3118 DGND 4.68fF $ **FLOATING
C6193 AVDD.n3120 DGND 0.31fF $ **FLOATING
C6194 AVDD.t509 DGND 0.46fF
C6195 AVDD.n3121 DGND 0.81fF $ **FLOATING
C6196 AVDD.n3122 DGND 0.19fF $ **FLOATING
C6197 AVDD.n3123 DGND 0.14fF $ **FLOATING
C6198 AVDD.n3125 DGND 0.14fF $ **FLOATING
C6199 AVDD.n3127 DGND 0.14fF $ **FLOATING
C6200 AVDD.n3129 DGND 0.14fF $ **FLOATING
C6201 AVDD.n3131 DGND 0.14fF $ **FLOATING
C6202 AVDD.n3133 DGND 0.14fF $ **FLOATING
C6203 AVDD.n3135 DGND 0.14fF $ **FLOATING
C6204 AVDD.n3137 DGND 0.14fF $ **FLOATING
C6205 AVDD.n3139 DGND 0.14fF $ **FLOATING
C6206 AVDD.n3140 DGND 6.22fF $ **FLOATING
C6207 AVDD.n3141 DGND 0.14fF $ **FLOATING
C6208 AVDD.n3142 DGND 0.66fF $ **FLOATING
C6209 AVDD.t172 DGND 4.29fF
C6210 AVDD.n3143 DGND 0.81fF $ **FLOATING
C6211 AVDD.n3144 DGND 0.19fF $ **FLOATING
C6212 AVDD.n3145 DGND 0.14fF $ **FLOATING
C6213 AVDD.n3147 DGND 0.14fF $ **FLOATING
C6214 AVDD.n3149 DGND 0.14fF $ **FLOATING
C6215 AVDD.n3151 DGND 0.14fF $ **FLOATING
C6216 AVDD.n3153 DGND 0.14fF $ **FLOATING
C6217 AVDD.n3155 DGND 0.14fF $ **FLOATING
C6218 AVDD.n3157 DGND 0.14fF $ **FLOATING
C6219 AVDD.n3159 DGND 0.14fF $ **FLOATING
C6220 AVDD.n3161 DGND 0.14fF $ **FLOATING
C6221 AVDD.n3162 DGND 6.96fF $ **FLOATING
C6222 AVDD.n3163 DGND 0.14fF $ **FLOATING
C6223 AVDD.n3164 DGND 0.75fF $ **FLOATING
C6224 AVDD.n3165 DGND 0.95fF $ **FLOATING
C6225 AVDD.n3166 DGND 0.44fF $ **FLOATING
C6226 AVDD.n3215 DGND 4.11fF $ **FLOATING
C6227 AVDD.n3217 DGND 0.13fF $ **FLOATING
C6228 AVDD.n3219 DGND 0.13fF $ **FLOATING
C6229 AVDD.n3221 DGND 0.13fF $ **FLOATING
C6230 AVDD.n3223 DGND 0.13fF $ **FLOATING
C6231 AVDD.n3225 DGND 0.13fF $ **FLOATING
C6232 AVDD.n3227 DGND 0.13fF $ **FLOATING
C6233 AVDD.n3229 DGND 0.13fF $ **FLOATING
C6234 AVDD.n3231 DGND 0.13fF $ **FLOATING
C6235 AVDD.n3232 DGND 1.19fF $ **FLOATING
C6236 AVDD.n3233 DGND 0.13fF $ **FLOATING
C6237 AVDD.n3235 DGND 0.13fF $ **FLOATING
C6238 AVDD.n3237 DGND 0.13fF $ **FLOATING
C6239 AVDD.n3239 DGND 0.13fF $ **FLOATING
C6240 AVDD.n3241 DGND 0.13fF $ **FLOATING
C6241 AVDD.n3243 DGND 0.13fF $ **FLOATING
C6242 AVDD.n3245 DGND 0.13fF $ **FLOATING
C6243 AVDD.n3247 DGND 0.13fF $ **FLOATING
C6244 AVDD.n3249 DGND 0.13fF $ **FLOATING
C6245 AVDD.n3251 DGND 0.13fF $ **FLOATING
C6246 AVDD.t25 DGND 2.60fF
C6247 AVDD.n3252 DGND 0.13fF $ **FLOATING
C6248 AVDD.n3253 DGND 0.13fF $ **FLOATING
C6249 AVDD.n3254 DGND 0.48fF $ **FLOATING
C6250 AVDD.n3269 DGND 8.18fF $ **FLOATING
C6251 AVDD.n3271 DGND 1.56fF $ **FLOATING
C6252 AVDD.n3272 DGND 0.61fF $ **FLOATING
C6253 AVDD.n3273 DGND 0.40fF $ **FLOATING
C6254 AVDD.n3328 DGND 6.08fF $ **FLOATING
C6255 AVDD.n3337 DGND 8.80fF $ **FLOATING
C6256 AVDD.n3339 DGND 1.62fF $ **FLOATING
C6257 AVDD.n3340 DGND 0.65fF $ **FLOATING
C6258 AVDD.n3389 DGND 6.11fF $ **FLOATING
C6259 AVDD.n3404 DGND 8.80fF $ **FLOATING
C6260 AVDD.n3406 DGND 1.42fF $ **FLOATING
C6261 AVDD.t159 DGND 11.14fF
C6262 AVDD.n3408 DGND 0.13fF $ **FLOATING
C6263 AVDD.n3410 DGND 0.13fF $ **FLOATING
C6264 AVDD.n3412 DGND 0.13fF $ **FLOATING
C6265 AVDD.n3414 DGND 0.13fF $ **FLOATING
C6266 AVDD.n3416 DGND 0.13fF $ **FLOATING
C6267 AVDD.n3418 DGND 0.13fF $ **FLOATING
C6268 AVDD.n3420 DGND 0.13fF $ **FLOATING
C6269 AVDD.n3422 DGND 0.13fF $ **FLOATING
C6270 AVDD.n3423 DGND 1.19fF $ **FLOATING
C6271 AVDD.n3424 DGND 0.13fF $ **FLOATING
C6272 AVDD.n3426 DGND 0.13fF $ **FLOATING
C6273 AVDD.n3428 DGND 0.13fF $ **FLOATING
C6274 AVDD.n3430 DGND 0.13fF $ **FLOATING
C6275 AVDD.n3432 DGND 0.13fF $ **FLOATING
C6276 AVDD.n3434 DGND 0.13fF $ **FLOATING
C6277 AVDD.n3436 DGND 0.13fF $ **FLOATING
C6278 AVDD.n3438 DGND 0.13fF $ **FLOATING
C6279 AVDD.n3440 DGND 0.13fF $ **FLOATING
C6280 AVDD.n3442 DGND 0.13fF $ **FLOATING
C6281 AVDD.t2 DGND 6.96fF
C6282 AVDD.n3443 DGND 0.13fF $ **FLOATING
C6283 AVDD.n3444 DGND 0.13fF $ **FLOATING
C6284 AVDD.n3445 DGND 1.56fF $ **FLOATING
C6285 AVDD.n3446 DGND 0.35fF $ **FLOATING
C6286 AVDD.n3447 DGND 0.35fF $ **FLOATING
C6287 AVDD.n3448 DGND 0.36fF $ **FLOATING
C6288 AVDD.n3449 DGND 0.36fF $ **FLOATING
C6289 AVDD.n3450 DGND 0.36fF $ **FLOATING
C6290 AVDD.n3451 DGND 0.36fF $ **FLOATING
C6291 AVDD.n3452 DGND 0.35fF $ **FLOATING
C6292 AVDD.n3453 DGND 0.35fF $ **FLOATING
C6293 AVDD.n3454 DGND 0.35fF $ **FLOATING
C6294 AVDD.n3455 DGND 0.35fF $ **FLOATING
C6295 AVDD.n3456 DGND 0.35fF $ **FLOATING
C6296 AVDD.n3457 DGND 0.65fF $ **FLOATING
C6297 AVDD.n3458 DGND 0.36fF $ **FLOATING
C6298 AVDD.n3460 DGND 0.23fF $ **FLOATING
C6299 AVDD.n3461 DGND 0.36fF $ **FLOATING
C6300 AVDD.n3462 DGND 0.35fF $ **FLOATING
C6301 AVDD.n3463 DGND 0.35fF $ **FLOATING
C6302 AVDD.n3464 DGND 0.65fF $ **FLOATING
C6303 AVDD.n3465 DGND 0.38fF $ **FLOATING
C6304 AVDD.n3468 DGND 0.17fF $ **FLOATING
C6305 AVDD.n3475 DGND 0.17fF $ **FLOATING
C6306 AVDD.n3478 DGND 0.19fF $ **FLOATING
C6307 AVDD.n3479 DGND 0.35fF $ **FLOATING
C6308 AVDD.n3480 DGND 0.14fF $ **FLOATING
C6309 AVDD.n3481 DGND 0.52fF $ **FLOATING
C6310 AVDD.n3482 DGND 0.32fF $ **FLOATING
C6311 AVDD.n3483 DGND 0.37fF $ **FLOATING
C6312 AVDD.n3484 DGND 0.25fF $ **FLOATING
C6313 AVDD.n3485 DGND 0.18fF $ **FLOATING
C6314 AVDD.n3486 DGND 0.15fF $ **FLOATING
C6315 AVDD.n3487 DGND 0.35fF $ **FLOATING
C6316 AVDD.n3488 DGND 0.16fF $ **FLOATING
C6317 AVDD.n3489 DGND 0.10fF $ **FLOATING
C6318 AVDD.n3490 DGND 0.24fF $ **FLOATING
C6319 AVDD.n3491 DGND 0.12fF $ **FLOATING
C6320 AVDD.n3493 DGND 0.91fF $ **FLOATING
C6321 AVDD.n3495 DGND 0.26fF $ **FLOATING
C6322 AVDD.n3496 DGND 0.22fF $ **FLOATING
C6323 AVDD.n3498 DGND 0.91fF $ **FLOATING
C6324 AVDD.n3499 DGND 0.23fF $ **FLOATING
C6325 AVDD.n3500 DGND 0.12fF $ **FLOATING
C6326 AVDD.n3503 DGND 0.83fF $ **FLOATING
C6327 AVDD.n3505 DGND 0.36fF $ **FLOATING
C6328 AVDD.n3507 DGND 0.21fF $ **FLOATING
C6329 AVDD.n3509 DGND 0.36fF $ **FLOATING
C6330 AVDD.n3511 DGND 0.21fF $ **FLOATING
C6331 AVDD.n3513 DGND 0.36fF $ **FLOATING
C6332 AVDD.n3515 DGND 0.21fF $ **FLOATING
C6333 AVDD.n3517 DGND 0.36fF $ **FLOATING
C6334 AVDD.n3519 DGND 0.21fF $ **FLOATING
C6335 AVDD.n3521 DGND 0.36fF $ **FLOATING
C6336 AVDD.n3523 DGND 0.36fF $ **FLOATING
C6337 AVDD.n3525 DGND 0.21fF $ **FLOATING
C6338 AVDD.n3527 DGND 0.36fF $ **FLOATING
C6339 AVDD.n3529 DGND 0.21fF $ **FLOATING
C6340 AVDD.n3531 DGND 0.36fF $ **FLOATING
C6341 AVDD.t374 DGND 11.16fF
C6342 AVDD.n3533 DGND 0.21fF $ **FLOATING
C6343 AVDD.n3535 DGND 0.23fF $ **FLOATING
C6344 AVDD.n3536 DGND 0.12fF $ **FLOATING
C6345 AVDD.n3539 DGND 0.35fF $ **FLOATING
C6346 AVDD.n3540 DGND 0.15fF $ **FLOATING
C6347 AVDD.n3541 DGND 0.62fF $ **FLOATING
C6348 AVDD.n3542 DGND 0.56fF $ **FLOATING
C6349 AVDD.n3543 DGND 0.25fF $ **FLOATING
C6350 AVDD.n3544 DGND 0.35fF $ **FLOATING
C6351 AVDD.n3545 DGND 0.18fF $ **FLOATING
C6352 AVDD.n3547 DGND 0.17fF $ **FLOATING
C6353 AVDD.n3554 DGND 0.17fF $ **FLOATING
C6354 AVDD.n3557 DGND 0.19fF $ **FLOATING
C6355 AVDD.n3558 DGND 0.15fF $ **FLOATING
C6356 AVDD.n3559 DGND 0.16fF $ **FLOATING
C6357 AVDD.n3560 DGND 0.10fF $ **FLOATING
C6358 AVDD.n3561 DGND 0.24fF $ **FLOATING
C6359 AVDD.n3562 DGND 0.12fF $ **FLOATING
C6360 AVDD.n3564 DGND 0.52fF $ **FLOATING
C6361 AVDD.n3565 DGND 0.97fF $ **FLOATING
C6362 AVDD.n3566 DGND 0.13fF $ **FLOATING
C6363 AVDD.n3567 DGND 0.15fF $ **FLOATING
C6364 AVDD.n3568 DGND 0.15fF $ **FLOATING
C6365 AVDD.n3570 DGND 0.15fF $ **FLOATING
C6366 AVDD.n3571 DGND 0.15fF $ **FLOATING
C6367 AVDD.n3573 DGND 0.15fF $ **FLOATING
C6368 AVDD.n3574 DGND 0.15fF $ **FLOATING
C6369 AVDD.n3576 DGND 0.20fF $ **FLOATING
C6370 AVDD.n3579 DGND 0.45fF $ **FLOATING
C6371 AVDD.n3585 DGND 0.10fF $ **FLOATING
C6372 AVDD.n3588 DGND 0.44fF $ **FLOATING
C6373 AVDD.n3591 DGND 0.12fF $ **FLOATING
C6374 AVDD.n3596 DGND 0.44fF $ **FLOATING
C6375 AVDD.n3599 DGND 0.12fF $ **FLOATING
C6376 AVDD.n3604 DGND 0.44fF $ **FLOATING
C6377 AVDD.n3607 DGND 0.12fF $ **FLOATING
C6378 AVDD.n3612 DGND 0.44fF $ **FLOATING
C6379 AVDD.n3615 DGND 0.12fF $ **FLOATING
C6380 AVDD.n3620 DGND 0.44fF $ **FLOATING
C6381 AVDD.n3623 DGND 0.12fF $ **FLOATING
C6382 AVDD.n3628 DGND 0.44fF $ **FLOATING
C6383 AVDD.n3631 DGND 0.12fF $ **FLOATING
C6384 AVDD.n3637 DGND 3.96fF $ **FLOATING
C6385 AVDD.n3638 DGND 0.13fF $ **FLOATING
C6386 AVDD.n3639 DGND 0.15fF $ **FLOATING
C6387 AVDD.n3641 DGND 0.15fF $ **FLOATING
C6388 AVDD.n3642 DGND 0.15fF $ **FLOATING
C6389 AVDD.n3644 DGND 0.15fF $ **FLOATING
C6390 AVDD.n3645 DGND 0.15fF $ **FLOATING
C6391 AVDD.n3647 DGND 0.15fF $ **FLOATING
C6392 AVDD.n3648 DGND 0.13fF $ **FLOATING
C6393 AVDD.n3650 DGND 4.60fF $ **FLOATING
C6394 AVDD.n3651 DGND 0.66fF $ **FLOATING
C6395 AVDD.n3652 DGND 0.24fF $ **FLOATING
C6396 AVDD.n3653 DGND 0.66fF $ **FLOATING
C6397 AVDD.n3654 DGND 0.24fF $ **FLOATING
C6398 AVDD.n3655 DGND 0.66fF $ **FLOATING
C6399 AVDD.n3656 DGND 0.24fF $ **FLOATING
C6400 AVDD.n3657 DGND 0.66fF $ **FLOATING
C6401 AVDD.n3658 DGND 0.24fF $ **FLOATING
C6402 AVDD.n3659 DGND 0.66fF $ **FLOATING
C6403 AVDD.n3660 DGND 0.24fF $ **FLOATING
C6404 AVDD.n3661 DGND 0.66fF $ **FLOATING
C6405 AVDD.n3662 DGND 0.24fF $ **FLOATING
C6406 AVDD.n3663 DGND 0.66fF $ **FLOATING
C6407 AVDD.n3664 DGND 0.24fF $ **FLOATING
C6408 AVDD.n3665 DGND 0.66fF $ **FLOATING
C6409 AVDD.n3666 DGND 0.24fF $ **FLOATING
C6410 AVDD.n3667 DGND 0.66fF $ **FLOATING
C6411 AVDD.n3668 DGND 0.24fF $ **FLOATING
C6412 AVDD.n3669 DGND 6.22fF $ **FLOATING
C6413 AVDD.n3670 DGND 0.14fF $ **FLOATING
C6414 AVDD.n3671 DGND 0.68fF $ **FLOATING
C6415 AVDD.n3672 DGND 0.52fF $ **FLOATING
C6416 AVDD.n3673 DGND 7.07fF $ **FLOATING
C6417 AVDD.n3674 DGND 0.22fF $ **FLOATING
C6418 AVDD.n3675 DGND 0.28fF $ **FLOATING
C6419 AVDD.n3676 DGND 0.13fF $ **FLOATING
C6420 AVDD.n3677 DGND 0.66fF $ **FLOATING
C6421 AVDD.n3678 DGND 0.13fF $ **FLOATING
C6422 AVDD.n3679 DGND 0.13fF $ **FLOATING
C6423 AVDD.n3680 DGND 0.66fF $ **FLOATING
C6424 AVDD.n3681 DGND 0.13fF $ **FLOATING
C6425 AVDD.n3682 DGND 0.13fF $ **FLOATING
C6426 AVDD.n3683 DGND 0.66fF $ **FLOATING
C6427 AVDD.n3684 DGND 0.13fF $ **FLOATING
C6428 AVDD.n3685 DGND 0.13fF $ **FLOATING
C6429 AVDD.n3686 DGND 0.44fF $ **FLOATING
C6430 AVDD.n3687 DGND 0.66fF $ **FLOATING
C6431 AVDD.n3688 DGND 0.13fF $ **FLOATING
C6432 AVDD.n3689 DGND 0.13fF $ **FLOATING
C6433 AVDD.t381 DGND 10.77fF
C6434 AVDD.n3690 DGND 0.66fF $ **FLOATING
C6435 AVDD.n3691 DGND 0.13fF $ **FLOATING
C6436 AVDD.n3692 DGND 0.13fF $ **FLOATING
C6437 AVDD.n3693 DGND 0.66fF $ **FLOATING
C6438 AVDD.n3694 DGND 0.13fF $ **FLOATING
C6439 AVDD.n3695 DGND 0.13fF $ **FLOATING
C6440 AVDD.n3696 DGND 0.66fF $ **FLOATING
C6441 AVDD.n3697 DGND 0.13fF $ **FLOATING
C6442 AVDD.n3698 DGND 0.13fF $ **FLOATING
C6443 AVDD.n3699 DGND 0.66fF $ **FLOATING
C6444 AVDD.n3700 DGND 0.13fF $ **FLOATING
C6445 AVDD.n3701 DGND 0.13fF $ **FLOATING
C6446 AVDD.n3702 DGND 0.66fF $ **FLOATING
C6447 AVDD.n3703 DGND 0.13fF $ **FLOATING
C6448 AVDD.n3704 DGND 0.13fF $ **FLOATING
C6449 AVDD.t366 DGND 6.19fF
C6450 AVDD.n3705 DGND 4.99fF $ **FLOATING
C6451 AVDD.n3707 DGND 0.26fF $ **FLOATING
C6452 AVDD.n3708 DGND 0.35fF $ **FLOATING
C6453 AVDD.n3709 DGND 0.14fF $ **FLOATING
C6454 AVDD.n3710 DGND 0.50fF $ **FLOATING
C6455 AVDD.n3711 DGND 0.32fF $ **FLOATING
C6456 AVDD.n3712 DGND 0.37fF $ **FLOATING
C6457 AVDD.n3713 DGND 0.25fF $ **FLOATING
C6458 AVDD.n3714 DGND 0.35fF $ **FLOATING
C6459 AVDD.n3715 DGND 0.18fF $ **FLOATING
C6460 AVDD.n3717 DGND 0.17fF $ **FLOATING
C6461 AVDD.n3724 DGND 0.17fF $ **FLOATING
C6462 AVDD.n3727 DGND 0.19fF $ **FLOATING
C6463 AVDD.n3728 DGND 0.15fF $ **FLOATING
C6464 AVDD.n3729 DGND 0.16fF $ **FLOATING
C6465 AVDD.n3730 DGND 0.10fF $ **FLOATING
C6466 AVDD.n3731 DGND 0.24fF $ **FLOATING
C6467 AVDD.n3732 DGND 0.12fF $ **FLOATING
C6468 AVDD.n3735 DGND 0.26fF $ **FLOATING
C6469 AVDD.n3737 DGND 0.16fF $ **FLOATING
C6470 AVDD.t838 DGND 3.08fF
C6471 AVDD.n3753 DGND 0.20fF $ **FLOATING
C6472 AVDD.n3756 DGND 2.11fF $ **FLOATING
C6473 AVDD.n3758 DGND 15.45fF $ **FLOATING
C6474 AVDD.t741 DGND 2.05fF
C6475 AVDD.t723 DGND 3.20fF
C6476 AVDD.n3778 DGND 0.15fF $ **FLOATING
C6477 AVDD.n3779 DGND 4.94fF $ **FLOATING
C6478 AVDD.n3783 DGND 0.32fF $ **FLOATING
C6479 AVDD.n3784 DGND 0.25fF $ **FLOATING
C6480 AVDD.n3791 DGND 0.19fF $ **FLOATING
C6481 AVDD.n3792 DGND 0.32fF $ **FLOATING
C6482 AVDD.t731 DGND 1.31fF
C6483 AVDD.n3796 DGND 0.20fF $ **FLOATING
C6484 AVDD.n3800 DGND 0.16fF $ **FLOATING
C6485 AVDD.t190 DGND 0.57fF
C6486 AVDD.n3812 DGND 0.16fF $ **FLOATING
C6487 AVDD.t763 DGND 0.59fF
C6488 level_shifter_up_2.VDD_HV DGND 0.16fF $ **FLOATING
C6489 AVDD.n3825 DGND 0.20fF $ **FLOATING
C6490 level_shifter_up_1.VDD_HV DGND 0.16fF $ **FLOATING
C6491 AVDD.n3829 DGND 0.32fF $ **FLOATING
C6492 AVDD.n3830 DGND 0.19fF $ **FLOATING
C6493 AVDD.n3831 DGND 0.42fF $ **FLOATING
C6494 AVDD.n3834 DGND 0.19fF $ **FLOATING
C6495 AVDD.t181 DGND 0.38fF
C6496 AVDD.n3843 DGND 0.39fF $ **FLOATING
C6497 AVDD.t767 DGND 0.59fF
C6498 AVDD.n3857 DGND 0.16fF $ **FLOATING
C6499 AVDD.t833 DGND 0.57fF
C6500 AVDD.n3872 DGND 0.16fF $ **FLOATING
C6501 AVDD.n3878 DGND 0.32fF $ **FLOATING
C6502 AVDD.n3879 DGND 0.25fF $ **FLOATING
C6503 AVDD.n3887 DGND 0.20fF $ **FLOATING
C6504 AVDD.t142 DGND 0.85fF
C6505 AVDD.n3896 DGND 0.23fF $ **FLOATING
C6506 AVDD.n3897 DGND 0.35fF $ **FLOATING
C6507 AVDD.n3901 DGND 0.10fF $ **FLOATING
C6508 AVDD.n3902 DGND 0.16fF $ **FLOATING
C6509 AVDD.t144 DGND 0.38fF
C6510 AVDD.n3910 DGND 0.39fF $ **FLOATING
C6511 AVDD.t707 DGND 0.59fF
C6512 AVDD.n3924 DGND 0.16fF $ **FLOATING
C6513 AVDD.t729 DGND 0.57fF
C6514 AVDD.n3939 DGND 0.16fF $ **FLOATING
C6515 AVDD.n3947 DGND 0.20fF $ **FLOATING
C6516 AVDD.n3948 DGND 0.37fF $ **FLOATING
C6517 AVDD.n3957 DGND 0.20fF $ **FLOATING
C6518 AVDD.n3958 DGND 0.19fF $ **FLOATING
C6519 AVDD.t262 DGND 0.85fF
C6520 AVDD.n3962 DGND 0.36fF $ **FLOATING
C6521 AVDD.n3963 DGND 0.35fF $ **FLOATING
C6522 AVDD.n3967 DGND 0.10fF $ **FLOATING
C6523 AVDD.n3968 DGND 0.16fF $ **FLOATING
C6524 AVDD.t0 DGND 0.38fF
C6525 AVDD.n3976 DGND 0.39fF $ **FLOATING
C6526 AVDD.n3984 DGND 0.16fF $ **FLOATING
C6527 AVDD.n3985 DGND 0.15fF $ **FLOATING
C6528 AVDD.n3989 DGND 0.44fF $ **FLOATING
C6529 AVDD.n3993 DGND 0.63fF $ **FLOATING
C6530 AVDD.n3994 DGND 0.21fF $ **FLOATING
C6531 AVDD.n3996 DGND 0.19fF $ **FLOATING
C6532 AVDD.n3997 DGND 0.14fF $ **FLOATING
C6533 AVDD.n3998 DGND 0.34fF $ **FLOATING
C6534 AVDD.n3999 DGND 0.15fF $ **FLOATING
C6535 AVDD.n4003 DGND 0.56fF $ **FLOATING
C6536 AVDD.n4007 DGND 0.11fF $ **FLOATING
C6537 AVDD.n4008 DGND 0.31fF $ **FLOATING
C6538 AVDD.n4009 DGND 0.12fF $ **FLOATING
C6539 AVDD.n4013 DGND 0.15fF $ **FLOATING
C6540 AVDD.n4017 DGND 0.54fF $ **FLOATING
C6541 AVDD.n4018 DGND 0.28fF $ **FLOATING
C6542 AVDD.n4021 DGND 0.34fF $ **FLOATING
C6543 AVDD.t718 DGND 0.47fF
C6544 AVDD.n4024 DGND 0.30fF $ **FLOATING
C6545 AVDD.n4026 DGND 0.33fF $ **FLOATING
C6546 AVDD.t717 DGND 0.33fF
C6547 AVDD.n4027 DGND 0.78fF $ **FLOATING
C6548 AVDD.n4028 DGND 0.34fF $ **FLOATING
C6549 AVDD.n4030 DGND 0.18fF $ **FLOATING
C6550 AVDD.n4031 DGND 0.58fF $ **FLOATING
C6551 AVDD.n4038 DGND 0.16fF $ **FLOATING
C6552 AVDD.n4040 DGND 0.20fF $ **FLOATING
C6553 AVDD.n4044 DGND 0.32fF $ **FLOATING
C6554 AVDD.n4045 DGND 0.19fF $ **FLOATING
C6555 AVDD.n4046 DGND 0.42fF $ **FLOATING
C6556 AVDD.n4049 DGND 0.19fF $ **FLOATING
C6557 AVDD.t29 DGND 0.38fF
C6558 AVDD.n4058 DGND 0.39fF $ **FLOATING
C6559 AVDD.t719 DGND 0.59fF
C6560 AVDD.n4072 DGND 0.16fF $ **FLOATING
C6561 AVDD.t40 DGND 0.57fF
C6562 AVDD.n4087 DGND 0.16fF $ **FLOATING
C6563 AVDD.n4093 DGND 0.32fF $ **FLOATING
C6564 AVDD.n4094 DGND 0.25fF $ **FLOATING
C6565 AVDD.n4102 DGND 0.20fF $ **FLOATING
C6566 AVDD.t745 DGND 0.85fF
C6567 AVDD.n4111 DGND 0.23fF $ **FLOATING
C6568 AVDD.n4112 DGND 0.35fF $ **FLOATING
C6569 AVDD.n4116 DGND 0.10fF $ **FLOATING
C6570 AVDD.n4117 DGND 0.16fF $ **FLOATING
C6571 AVDD.t215 DGND 0.38fF
C6572 AVDD.n4125 DGND 0.39fF $ **FLOATING
C6573 AVDD.t270 DGND 0.59fF
C6574 AVDD.n4139 DGND 0.16fF $ **FLOATING
C6575 AVDD.t54 DGND 0.57fF
C6576 AVDD.n4154 DGND 0.16fF $ **FLOATING
C6577 AVDD.n4162 DGND 0.20fF $ **FLOATING
C6578 AVDD.n4163 DGND 0.37fF $ **FLOATING
C6579 AVDD.n4172 DGND 0.20fF $ **FLOATING
C6580 AVDD.n4174 DGND 0.10fF $ **FLOATING
C6581 level_shifter_up_7.VDD_HV DGND 0.16fF $ **FLOATING
C6582 AVDD.n4175 DGND 0.19fF $ **FLOATING
C6583 AVDD.t765 DGND 0.85fF
C6584 AVDD.n4179 DGND 0.42fF $ **FLOATING
C6585 AVDD.n4181 DGND 0.18fF $ **FLOATING
C6586 AVDD.n4182 DGND 0.87fF $ **FLOATING
C6587 AVDD.n4185 DGND 1.09fF $ **FLOATING
C6588 AVDD.t749 DGND 1.74fF
C6589 AVDD.n4195 DGND 0.10fF $ **FLOATING
C6590 AVDD.n4198 DGND 0.17fF $ **FLOATING
C6591 AVDD.n4201 DGND 0.96fF $ **FLOATING
C6592 AVDD.n4202 DGND 0.22fF $ **FLOATING
C6593 AVDD.n4203 DGND 0.11fF $ **FLOATING
C6594 AVDD.t192 DGND 0.60fF
C6595 AVDD.n4207 DGND 0.91fF $ **FLOATING
C6596 AVDD.n4219 DGND 0.13fF $ **FLOATING
C6597 AVDD.n4220 DGND 0.17fF $ **FLOATING
C6598 AVDD.n4228 DGND 0.42fF $ **FLOATING
C6599 AVDD.t339 DGND 1.60fF
C6600 AVDD.n4239 DGND 0.19fF $ **FLOATING
C6601 AVDD.n4244 DGND 0.14fF $ **FLOATING
C6602 AVDD.n4245 DGND 1.60fF $ **FLOATING
C6603 AVDD.t760 DGND 0.45fF
C6604 AVDD.n4247 DGND 0.18fF $ **FLOATING
C6605 AVDD.n4248 DGND 0.80fF $ **FLOATING
C6606 AVDD.t806 DGND 0.58fF
C6607 AVDD.n4254 DGND 0.13fF $ **FLOATING
C6608 AVDD.n4255 DGND 0.19fF $ **FLOATING
C6609 AVDD.n4258 DGND 0.15fF $ **FLOATING
C6610 AVDD.n4262 DGND 0.47fF $ **FLOATING
C6611 AVDD.t56 DGND 0.41fF
C6612 AVDD.n4266 DGND 0.42fF $ **FLOATING
C6613 AVDD.n4269 DGND 0.15fF $ **FLOATING
C6614 AVDD.n4273 DGND 0.70fF $ **FLOATING
C6615 AVDD.t33 DGND 0.45fF
C6616 AVDD.n4279 DGND 0.15fF $ **FLOATING
C6617 AVDD.n4281 DGND 0.72fF $ **FLOATING
C6618 AVDD.n4284 DGND 0.15fF $ **FLOATING
C6619 AVDD.n4288 DGND 0.47fF $ **FLOATING
C6620 AVDD.t747 DGND 0.44fF
C6621 AVDD.t748 DGND 0.28fF
C6622 AVDD.t39 DGND 0.28fF
C6623 AVDD.n4294 DGND 0.19fF $ **FLOATING
C6624 AVDD.n4296 DGND 0.25fF $ **FLOATING
C6625 AVDD.n4297 DGND 0.13fF $ **FLOATING
C6626 AVDD.n4298 DGND 0.13fF $ **FLOATING
C6627 AVDD.t58 DGND 0.74fF
C6628 AVDD.t57 DGND 0.47fF
C6629 AVDD.t711 DGND 0.47fF
C6630 AVDD.n4301 DGND 0.31fF $ **FLOATING
C6631 AVDD.n4303 DGND 0.16fF $ **FLOATING
C6632 AVDD.n4304 DGND 0.17fF $ **FLOATING
C6633 AVDD.n4306 DGND 0.84fF $ **FLOATING
C6634 AVDD.n4308 DGND 0.19fF $ **FLOATING
C6635 AVDD.n4309 DGND 0.16fF $ **FLOATING
C6636 AVDD.t27 DGND 0.37fF
C6637 AVDD.n4310 DGND 0.16fF $ **FLOATING
C6638 AVDD.t28 DGND 0.34fF
C6639 AVDD.n4313 DGND 0.21fF $ **FLOATING
C6640 AVDD.n4315 DGND 0.20fF $ **FLOATING
C6641 AVDD.n4316 DGND 0.26fF $ **FLOATING
C6642 AVDD.n4319 DGND 0.26fF $ **FLOATING
C6643 AVDD.n4321 DGND 0.17fF $ **FLOATING
C6644 AVDD.t3 DGND 0.22fF
C6645 AVDD.n4322 DGND 0.31fF $ **FLOATING
C6646 AVDD.n4324 DGND 0.23fF $ **FLOATING
C6647 AVDD.t61 DGND 0.47fF
C6648 AVDD.n4326 DGND 0.64fF $ **FLOATING
C6649 AVDD.t721 DGND 0.61fF
C6650 AVDD.t716 DGND 0.34fF
C6651 AVDD.t153 DGND 0.74fF
C6652 AVDD.t154 DGND 0.47fF
C6653 AVDD.n4329 DGND 0.50fF $ **FLOATING
C6654 AVDD.n4331 DGND 0.15fF $ **FLOATING
C6655 AVDD.t36 DGND 0.44fF
C6656 AVDD.n4335 DGND 0.42fF $ **FLOATING
C6657 AVDD.n4341 DGND 0.15fF $ **FLOATING
C6658 AVDD.n4344 DGND 0.41fF $ **FLOATING
C6659 AVDD.n4347 DGND 0.11fF $ **FLOATING
C6660 AVDD.n4348 DGND 0.58fF $ **FLOATING
C6661 AVDD.t712 DGND 1.49fF
C6662 AVDD.n4350 DGND 0.36fF $ **FLOATING
C6663 AVDD.n4355 DGND 0.66fF $ **FLOATING
C6664 AVDD.n4359 DGND 0.62fF $ **FLOATING
C6665 AVDD.n4360 DGND 0.15fF $ **FLOATING
C6666 AVDD.n4363 DGND 0.34fF $ **FLOATING
C6667 AVDD.n4366 DGND 0.13fF $ **FLOATING
C6668 AVDD.n4368 DGND 0.12fF $ **FLOATING
C6669 AVDD.t37 DGND 0.28fF
C6670 AVDD.t722 DGND 0.44fF
C6671 AVDD.t38 DGND 0.28fF
C6672 AVDD.n4371 DGND 0.19fF $ **FLOATING
C6673 AVDD.n4373 DGND 0.19fF $ **FLOATING
C6674 AVDD.n4374 DGND 0.13fF $ **FLOATING
C6675 AVDD.n4375 DGND 0.13fF $ **FLOATING
C6676 AVDD.n4376 DGND 0.16fF $ **FLOATING
C6677 AVDD.n4378 DGND 0.25fF $ **FLOATING
C6678 AVDD.n4379 DGND 0.42fF $ **FLOATING
C6679 AVDD.t152 DGND 0.57fF
C6680 AVDD.t4 DGND 0.38fF
C6681 AVDD.n4381 DGND 0.19fF $ **FLOATING
C6682 AVDD.n4384 DGND 0.72fF $ **FLOATING
C6683 AVDD.n4386 DGND 0.53fF $ **FLOATING
C6684 AVDD.t185 DGND 0.44fF
C6685 AVDD.t709 DGND 2.22fF
C6686 AVDD.n4388 DGND 0.22fF $ **FLOATING
C6687 AVDD.n4389 DGND 0.27fF $ **FLOATING
C6688 AVDD.n4390 DGND 0.52fF $ **FLOATING
C6689 AVDD.n4391 DGND 0.16fF $ **FLOATING
C6690 level_shifter_up_6.VDD_HV DGND 0.35fF $ **FLOATING
C6691 AVDD.t739 DGND 2.02fF
C6692 AVDD.n4401 DGND 0.36fF $ **FLOATING
C6693 AVDD.n4404 DGND 0.60fF $ **FLOATING
C6694 AVDD.n4405 DGND 0.16fF $ **FLOATING
C6695 AVDD.n4407 DGND 0.21fF $ **FLOATING
C6696 AVDD.n4408 DGND 0.11fF $ **FLOATING
C6697 AVDD.n4409 DGND 2.51fF $ **FLOATING
C6698 AVDD.n4410 DGND 0.56fF $ **FLOATING
C6699 AVDD.n4411 DGND 9.86fF $ **FLOATING
C6700 AVDD.n4412 DGND 13.27fF $ **FLOATING
C6701 AVDD.n4413 DGND 1.60fF $ **FLOATING
C6702 AVDD.n4414 DGND 17.46fF $ **FLOATING
C6703 AVDD.n4415 DGND 0.35fF $ **FLOATING
C6704 AVDD.n4416 DGND 0.14fF $ **FLOATING
C6705 AVDD.n4417 DGND 0.50fF $ **FLOATING
C6706 AVDD.n4418 DGND 0.32fF $ **FLOATING
C6707 AVDD.n4419 DGND 0.37fF $ **FLOATING
C6708 AVDD.n4420 DGND 0.25fF $ **FLOATING
C6709 AVDD.n4421 DGND 0.35fF $ **FLOATING
C6710 AVDD.n4422 DGND 0.18fF $ **FLOATING
C6711 AVDD.n4424 DGND 0.17fF $ **FLOATING
C6712 AVDD.n4427 DGND 0.17fF $ **FLOATING
C6713 AVDD.n4430 DGND 0.19fF $ **FLOATING
C6714 AVDD.n4431 DGND 0.15fF $ **FLOATING
C6715 AVDD.n4433 DGND 0.10fF $ **FLOATING
C6716 AVDD.n4434 DGND 0.24fF $ **FLOATING
C6717 AVDD.n4435 DGND 0.12fF $ **FLOATING
C6718 AVDD.n4436 DGND 0.65fF $ **FLOATING
C6719 AVDD.n4438 DGND 0.36fF $ **FLOATING
C6720 AVDD.n4441 DGND 0.22fF $ **FLOATING
C6721 AVDD.n4442 DGND 0.26fF $ **FLOATING
C6722 AVDD.n4443 DGND 0.35fF $ **FLOATING
C6723 AVDD.n4444 DGND 0.14fF $ **FLOATING
C6724 AVDD.n4445 DGND 0.50fF $ **FLOATING
C6725 AVDD.n4446 DGND 0.32fF $ **FLOATING
C6726 AVDD.n4447 DGND 0.37fF $ **FLOATING
C6727 AVDD.n4448 DGND 0.25fF $ **FLOATING
C6728 AVDD.n4449 DGND 0.35fF $ **FLOATING
C6729 AVDD.n4450 DGND 0.18fF $ **FLOATING
C6730 AVDD.n4452 DGND 0.17fF $ **FLOATING
C6731 AVDD.t593 DGND 0.28fF
C6732 AVDD.n4460 DGND 0.21fF $ **FLOATING
C6733 AVDD.t390 DGND 0.28fF
C6734 AVDD.n4462 DGND 1.66fF $ **FLOATING
C6735 AVDD.t446 DGND 0.28fF
C6736 AVDD.n4464 DGND 0.21fF $ **FLOATING
C6737 AVDD.t563 DGND 0.28fF
C6738 AVDD.n4466 DGND 1.66fF $ **FLOATING
C6739 AVDD.t623 DGND 0.28fF
C6740 AVDD.n4470 DGND 0.21fF $ **FLOATING
C6741 AVDD.t425 DGND 0.28fF
C6742 AVDD.n4472 DGND 1.66fF $ **FLOATING
C6743 AVDD.t461 DGND 0.28fF
C6744 AVDD.t677 DGND 0.28fF
C6745 AVDD.n4476 DGND 0.33fF $ **FLOATING
C6746 AVDD.n4477 DGND 0.43fF $ **FLOATING
C6747 AVDD.n4479 DGND 0.48fF $ **FLOATING
C6748 AVDD.n4480 DGND 0.19fF $ **FLOATING
C6749 AVDD.n4481 DGND 0.38fF $ **FLOATING
C6750 AVDD.n4482 DGND 0.25fF $ **FLOATING
C6751 AVDD.n4483 DGND 2.09fF $ **FLOATING
C6752 AVDD.n4487 DGND 0.17fF $ **FLOATING
C6753 AVDD.n4490 DGND 0.17fF $ **FLOATING
C6754 AVDD.t569 DGND 0.20fF
C6755 AVDD.n4493 DGND 0.35fF $ **FLOATING
C6756 AVDD.n4494 DGND 2.79fF $ **FLOATING
C6757 AVDD.n4495 DGND 1.91fF $ **FLOATING
C6758 AVDD.n4496 DGND 0.35fF $ **FLOATING
C6759 AVDD.n4497 DGND 0.18fF $ **FLOATING
C6760 AVDD.n4498 DGND 0.14fF $ **FLOATING
C6761 AVDD.n4499 DGND 0.19fF $ **FLOATING
C6762 AVDD.n4501 DGND 6.11fF $ **FLOATING
C6763 AVDD.n4503 DGND 0.17fF $ **FLOATING
C6764 AVDD.n4506 DGND 0.19fF $ **FLOATING
C6765 AVDD.n4507 DGND 0.15fF $ **FLOATING
C6766 AVDD.n4508 DGND 0.16fF $ **FLOATING
C6767 AVDD.n4509 DGND 0.10fF $ **FLOATING
C6768 AVDD.n4510 DGND 0.24fF $ **FLOATING
C6769 AVDD.n4511 DGND 0.12fF $ **FLOATING
C6770 AVDD.n4512 DGND 0.65fF $ **FLOATING
C6771 AVDD.n4514 DGND 0.36fF $ **FLOATING
C6772 AVDD.n4517 DGND 0.22fF $ **FLOATING
C6773 AVDD.n4518 DGND 0.26fF $ **FLOATING
C6774 AVDD.n4519 DGND 0.35fF $ **FLOATING
C6775 AVDD.n4520 DGND 0.14fF $ **FLOATING
C6776 AVDD.n4521 DGND 0.50fF $ **FLOATING
C6777 AVDD.n4522 DGND 0.32fF $ **FLOATING
C6778 AVDD.n4523 DGND 0.37fF $ **FLOATING
C6779 AVDD.n4524 DGND 0.25fF $ **FLOATING
C6780 AVDD.n4525 DGND 0.35fF $ **FLOATING
C6781 AVDD.n4526 DGND 0.18fF $ **FLOATING
C6782 AVDD.n4528 DGND 0.17fF $ **FLOATING
C6783 AVDD.n4535 DGND 0.17fF $ **FLOATING
C6784 AVDD.n4538 DGND 0.19fF $ **FLOATING
C6785 AVDD.n4539 DGND 0.15fF $ **FLOATING
C6786 AVDD.n4540 DGND 0.16fF $ **FLOATING
C6787 AVDD.n4541 DGND 0.10fF $ **FLOATING
C6788 AVDD.n4542 DGND 0.24fF $ **FLOATING
C6789 AVDD.n4543 DGND 0.12fF $ **FLOATING
C6790 AVDD.n4546 DGND 0.26fF $ **FLOATING
C6791 AVDD.n4547 DGND 0.35fF $ **FLOATING
C6792 AVDD.n4548 DGND 0.14fF $ **FLOATING
C6793 AVDD.n4549 DGND 0.50fF $ **FLOATING
C6794 AVDD.n4550 DGND 0.32fF $ **FLOATING
C6795 AVDD.n4551 DGND 0.37fF $ **FLOATING
C6796 AVDD.n4552 DGND 0.25fF $ **FLOATING
C6797 AVDD.n4553 DGND 0.35fF $ **FLOATING
C6798 AVDD.n4554 DGND 0.18fF $ **FLOATING
C6799 AVDD.n4556 DGND 0.17fF $ **FLOATING
C6800 AVDD.t641 DGND 0.28fF
C6801 AVDD.n4560 DGND 0.21fF $ **FLOATING
C6802 AVDD.t440 DGND 0.28fF
C6803 AVDD.n4562 DGND 1.66fF $ **FLOATING
C6804 AVDD.t464 DGND 0.28fF
C6805 AVDD.n4564 DGND 0.21fF $ **FLOATING
C6806 AVDD.t584 DGND 0.28fF
C6807 AVDD.n4566 DGND 1.66fF $ **FLOATING
C6808 AVDD.t692 DGND 0.28fF
C6809 AVDD.t554 DGND 0.28fF
C6810 AVDD.n4570 DGND 1.96fF $ **FLOATING
C6811 AVDD.t518 DGND 0.28fF
C6812 AVDD.n4573 DGND 0.21fF $ **FLOATING
C6813 AVDD.n4574 DGND 0.10fF $ **FLOATING
C6814 AVDD.t380 DGND 0.28fF
C6815 AVDD.n4575 DGND 1.66fF $ **FLOATING
C6816 AVDD.n4583 DGND 6.08fF $ **FLOATING
C6817 AVDD.n4587 DGND 0.17fF $ **FLOATING
C6818 AVDD.n4590 DGND 0.19fF $ **FLOATING
C6819 AVDD.n4591 DGND 0.15fF $ **FLOATING
C6820 AVDD.n4592 DGND 0.16fF $ **FLOATING
C6821 AVDD.n4593 DGND 0.10fF $ **FLOATING
C6822 AVDD.n4595 DGND 0.22fF $ **FLOATING
C6823 AVDD.n4596 DGND 0.26fF $ **FLOATING
C6824 AVDD.n4597 DGND 18.37fF $ **FLOATING
C6825 AVDD.n4598 DGND 0.23fF $ **FLOATING
C6826 AVDD.n4599 DGND 0.36fF $ **FLOATING
C6827 AVDD.n4600 DGND 0.65fF $ **FLOATING
C6828 AVDD.n4601 DGND 0.36fF $ **FLOATING
C6829 AVDD.n4603 DGND 0.23fF $ **FLOATING
C6830 AVDD.n4604 DGND 0.36fF $ **FLOATING
C6831 AVDD.n4605 DGND 0.81fF $ **FLOATING
C6832 AVDD.n4606 DGND 0.19fF $ **FLOATING
C6833 AVDD.n4607 DGND 0.14fF $ **FLOATING
C6834 AVDD.n4609 DGND 0.14fF $ **FLOATING
C6835 AVDD.n4611 DGND 0.14fF $ **FLOATING
C6836 AVDD.n4613 DGND 0.14fF $ **FLOATING
C6837 AVDD.n4615 DGND 0.14fF $ **FLOATING
C6838 AVDD.n4617 DGND 0.14fF $ **FLOATING
C6839 AVDD.n4619 DGND 0.14fF $ **FLOATING
C6840 AVDD.n4621 DGND 0.14fF $ **FLOATING
C6841 AVDD.n4623 DGND 0.14fF $ **FLOATING
C6842 AVDD.n4624 DGND 0.29fF $ **FLOATING
C6843 AVDD.t701 DGND 0.46fF
C6844 AVDD.n4625 DGND 0.85fF $ **FLOATING
C6845 AVDD.n4626 DGND 0.14fF $ **FLOATING
C6846 AVDD.n4627 DGND 0.56fF $ **FLOATING
C6847 AVDD.t650 DGND 0.46fF
C6848 AVDD.n4628 DGND 0.85fF $ **FLOATING
C6849 AVDD.n4629 DGND 0.14fF $ **FLOATING
C6850 AVDD.n4630 DGND 0.24fF $ **FLOATING
C6851 AVDD.t668 DGND 0.46fF
C6852 AVDD.n4631 DGND 0.43fF $ **FLOATING
C6853 AVDD.n4632 DGND 0.19fF $ **FLOATING
C6854 AVDD.n4633 DGND 0.14fF $ **FLOATING
C6855 AVDD.n4634 DGND 0.56fF $ **FLOATING
C6856 AVDD.n4635 DGND 0.38fF $ **FLOATING
C6857 AVDD.t515 DGND 0.46fF
C6858 AVDD.n4636 DGND 0.85fF $ **FLOATING
C6859 AVDD.n4637 DGND 0.14fF $ **FLOATING
C6860 AVDD.t365 DGND 0.46fF
C6861 AVDD.n4638 DGND 0.85fF $ **FLOATING
C6862 AVDD.n4639 DGND 0.14fF $ **FLOATING
C6863 AVDD.n4640 DGND 0.56fF $ **FLOATING
C6864 AVDD.n4641 DGND 0.56fF $ **FLOATING
C6865 AVDD.t416 DGND 0.46fF
C6866 AVDD.n4642 DGND 0.85fF $ **FLOATING
C6867 AVDD.n4643 DGND 0.14fF $ **FLOATING
C6868 AVDD.t608 DGND 0.46fF
C6869 AVDD.n4644 DGND 0.85fF $ **FLOATING
C6870 AVDD.n4645 DGND 0.14fF $ **FLOATING
C6871 AVDD.t476 DGND 0.46fF
C6872 AVDD.n4646 DGND 0.56fF $ **FLOATING
C6873 AVDD.n4647 DGND 0.85fF $ **FLOATING
C6874 AVDD.n4648 DGND 0.14fF $ **FLOATING
C6875 AVDD.n4649 DGND 0.56fF $ **FLOATING
C6876 AVDD.n4650 DGND 0.56fF $ **FLOATING
C6877 AVDD.t503 DGND 0.46fF
C6878 AVDD.n4651 DGND 0.85fF $ **FLOATING
C6879 AVDD.n4652 DGND 0.14fF $ **FLOATING
C6880 AVDD.n4653 DGND 6.96fF $ **FLOATING
C6881 AVDD.n4654 DGND 0.14fF $ **FLOATING
C6882 AVDD.t548 DGND 0.46fF
C6883 AVDD.n4655 DGND 0.46fF $ **FLOATING
C6884 AVDD.n4656 DGND 2.11fF $ **FLOATING
C6885 AVDD.n4657 DGND 0.14fF $ **FLOATING
C6886 AVDD.n4658 DGND 6.96fF $ **FLOATING
C6887 AVDD.n4689 DGND 0.19fF $ **FLOATING
C6888 AVDD.n4690 DGND 0.30fF $ **FLOATING
C6889 AVDD.n4692 DGND 0.35fF $ **FLOATING
C6890 AVDD.n4699 DGND 0.32fF $ **FLOATING
C6891 AVDD.n4709 DGND 4.64fF $ **FLOATING
C6892 AVDD.n4758 DGND 6.08fF $ **FLOATING
C6893 AVDD.n4807 DGND 6.11fF $ **FLOATING
C6894 AVDD.t163 DGND 11.18fF
C6895 AVDD.n4822 DGND 8.80fF $ **FLOATING
C6896 AVDD.n4825 DGND 6.04fF $ **FLOATING
C6897 AVDD.n4826 DGND 0.36fF $ **FLOATING
C6898 AVDD.n4827 DGND 0.36fF $ **FLOATING
C6899 AVDD.n4828 DGND 0.24fF $ **FLOATING
C6900 AVDD.n4829 DGND 0.18fF $ **FLOATING
C6901 AVDD.n4830 DGND 0.13fF $ **FLOATING
C6902 AVDD.n4832 DGND 0.13fF $ **FLOATING
C6903 AVDD.n4834 DGND 0.13fF $ **FLOATING
C6904 AVDD.n4836 DGND 0.13fF $ **FLOATING
C6905 AVDD.n4838 DGND 0.13fF $ **FLOATING
C6906 AVDD.n4840 DGND 0.13fF $ **FLOATING
C6907 AVDD.n4842 DGND 0.13fF $ **FLOATING
C6908 AVDD.n4844 DGND 0.13fF $ **FLOATING
C6909 AVDD.n4846 DGND 0.13fF $ **FLOATING
C6910 AVDD.n4847 DGND 1.19fF $ **FLOATING
C6911 AVDD.n4848 DGND 0.13fF $ **FLOATING
C6912 AVDD.n4850 DGND 0.13fF $ **FLOATING
C6913 AVDD.n4852 DGND 0.13fF $ **FLOATING
C6914 AVDD.n4854 DGND 0.13fF $ **FLOATING
C6915 AVDD.n4856 DGND 0.13fF $ **FLOATING
C6916 AVDD.n4858 DGND 0.13fF $ **FLOATING
C6917 AVDD.n4860 DGND 0.13fF $ **FLOATING
C6918 AVDD.n4862 DGND 0.13fF $ **FLOATING
C6919 AVDD.n4864 DGND 0.13fF $ **FLOATING
C6920 AVDD.n4866 DGND 0.13fF $ **FLOATING
C6921 AVDD.n4867 DGND 0.24fF $ **FLOATING
C6922 AVDD.n4869 DGND 0.13fF $ **FLOATING
C6923 AVDD.t47 DGND 6.22fF
C6924 AVDD.t168 DGND 11.12fF
C6925 AVDD.n4900 DGND 0.19fF $ **FLOATING
C6926 AVDD.n4901 DGND 0.19fF $ **FLOATING
C6927 AVDD.n4902 DGND 0.29fF $ **FLOATING
C6928 AVDD.n4904 DGND 0.35fF $ **FLOATING
C6929 AVDD.n4905 DGND 0.35fF $ **FLOATING
C6930 AVDD.n4906 DGND 0.91fF $ **FLOATING
C6931 AVDD.n4908 DGND 0.23fF $ **FLOATING
C6932 AVDD.n4909 DGND 0.36fF $ **FLOATING
C6933 AVDD.t166 DGND 10.85fF
C6934 AVDD.n4924 DGND 8.80fF $ **FLOATING
C6935 AVDD.n4927 DGND 1.81fF $ **FLOATING
C6936 AVDD.n4928 DGND 0.36fF $ **FLOATING
C6937 AVDD.n4929 DGND 0.36fF $ **FLOATING
C6938 AVDD.n4930 DGND 0.33fF $ **FLOATING
C6939 AVDD.n4979 DGND 4.16fF $ **FLOATING
C6940 AVDD.n4980 DGND 0.81fF $ **FLOATING
C6941 AVDD.n4981 DGND 0.19fF $ **FLOATING
C6942 AVDD.n4982 DGND 0.14fF $ **FLOATING
C6943 AVDD.n4984 DGND 0.14fF $ **FLOATING
C6944 AVDD.n4986 DGND 0.14fF $ **FLOATING
C6945 AVDD.n4988 DGND 0.14fF $ **FLOATING
C6946 AVDD.n4990 DGND 0.14fF $ **FLOATING
C6947 AVDD.n4992 DGND 0.14fF $ **FLOATING
C6948 AVDD.n4994 DGND 0.14fF $ **FLOATING
C6949 AVDD.n4996 DGND 0.14fF $ **FLOATING
C6950 AVDD.n4998 DGND 0.14fF $ **FLOATING
C6951 AVDD.n4999 DGND 2.60fF $ **FLOATING
C6952 AVDD.n5000 DGND 0.14fF $ **FLOATING
C6953 AVDD.n5001 DGND 0.27fF $ **FLOATING
C6954 AVDD.n5016 DGND 4.29fF $ **FLOATING
C6955 AVDD.n5018 DGND 0.44fF $ **FLOATING
C6956 AVDD.t632 DGND 0.46fF
C6957 AVDD.n5019 DGND 0.81fF $ **FLOATING
C6958 AVDD.n5020 DGND 0.19fF $ **FLOATING
C6959 AVDD.n5021 DGND 0.14fF $ **FLOATING
C6960 AVDD.t157 DGND 10.81fF
C6961 AVDD.n5023 DGND 0.14fF $ **FLOATING
C6962 AVDD.n5025 DGND 0.14fF $ **FLOATING
C6963 AVDD.n5027 DGND 0.14fF $ **FLOATING
C6964 AVDD.n5029 DGND 0.14fF $ **FLOATING
C6965 AVDD.n5031 DGND 0.14fF $ **FLOATING
C6966 AVDD.n5033 DGND 0.14fF $ **FLOATING
C6967 AVDD.n5035 DGND 0.14fF $ **FLOATING
C6968 AVDD.n5037 DGND 0.14fF $ **FLOATING
C6969 AVDD.n5038 DGND 6.19fF $ **FLOATING
C6970 AVDD.n5039 DGND 0.14fF $ **FLOATING
C6971 AVDD.n5040 DGND 0.55fF $ **FLOATING
C6972 AVDD.t521 DGND 0.46fF
C6973 AVDD.n5041 DGND 1.32fF $ **FLOATING
C6974 AVDD.n5042 DGND 0.82fF $ **FLOATING
C6975 AVDD.n5043 DGND 3.97fF $ **FLOATING
C6976 AVDD.n5044 DGND 1.50fF $ **FLOATING
C6977 AVDD.n5045 DGND 0.40fF $ **FLOATING
C6978 AVDD.n5046 DGND 1.37fF $ **FLOATING
C6979 AVDD.n5047 DGND 16.93fF $ **FLOATING
C6980 AVDD.n5048 DGND 0.36fF $ **FLOATING
C6981 AVDD.n5049 DGND 0.36fF $ **FLOATING
C6982 AVDD.n5050 DGND 0.35fF $ **FLOATING
C6983 AVDD.n5051 DGND 0.35fF $ **FLOATING
C6984 AVDD.n5052 DGND 0.36fF $ **FLOATING
C6985 AVDD.n5053 DGND 0.36fF $ **FLOATING
C6986 AVDD.n5054 DGND 0.36fF $ **FLOATING
C6987 AVDD.n5055 DGND 0.36fF $ **FLOATING
C6988 AVDD.n5056 DGND 0.35fF $ **FLOATING
C6989 AVDD.n5057 DGND 0.35fF $ **FLOATING
C6990 AVDD.n5058 DGND 0.35fF $ **FLOATING
C6991 AVDD.n5059 DGND 0.35fF $ **FLOATING
C6992 AVDD.n5060 DGND 0.36fF $ **FLOATING
C6993 AVDD.n5061 DGND 0.36fF $ **FLOATING
C6994 AVDD.t196 DGND 13.17fF
C6995 AVDD.n5092 DGND 0.19fF $ **FLOATING
C6996 AVDD.n5093 DGND 0.19fF $ **FLOATING
C6997 AVDD.n5094 DGND 0.29fF $ **FLOATING
C6998 AVDD.n5096 DGND 0.35fF $ **FLOATING
C6999 AVDD.n5097 DGND 0.35fF $ **FLOATING
C7000 AVDD.n5098 DGND 12.44fF $ **FLOATING
C7001 AVDD.n5099 DGND 0.36fF $ **FLOATING
C7002 AVDD.n5100 DGND 0.36fF $ **FLOATING
C7003 AVDD.n5101 DGND 0.35fF $ **FLOATING
C7004 AVDD.n5102 DGND 0.35fF $ **FLOATING
C7005 AVDD.n5103 DGND 0.36fF $ **FLOATING
C7006 AVDD.n5104 DGND 0.36fF $ **FLOATING
C7007 AVDD.n5105 DGND 0.36fF $ **FLOATING
C7008 AVDD.n5106 DGND 0.36fF $ **FLOATING
C7009 AVDD.n5107 DGND 0.35fF $ **FLOATING
C7010 AVDD.n5108 DGND 0.35fF $ **FLOATING
C7011 AVDD.n5109 DGND 0.35fF $ **FLOATING
C7012 AVDD.n5110 DGND 0.35fF $ **FLOATING
C7013 AVDD.n5111 DGND 0.36fF $ **FLOATING
C7014 AVDD.n5112 DGND 0.36fF $ **FLOATING
C7015 AVDD.t155 DGND 13.15fF
C7016 AVDD.n5143 DGND 0.19fF $ **FLOATING
C7017 AVDD.n5144 DGND 0.19fF $ **FLOATING
C7018 AVDD.n5145 DGND 0.29fF $ **FLOATING
C7019 AVDD.n5147 DGND 0.35fF $ **FLOATING
C7020 AVDD.n5148 DGND 0.35fF $ **FLOATING
C7021 AVDD.n5149 DGND 17.39fF $ **FLOATING
C7022 AVDD.n5150 DGND 0.36fF $ **FLOATING
C7023 AVDD.n5151 DGND 0.36fF $ **FLOATING
C7024 AVDD.n5152 DGND 0.35fF $ **FLOATING
C7025 AVDD.n5153 DGND 0.35fF $ **FLOATING
C7026 AVDD.n5154 DGND 0.36fF $ **FLOATING
C7027 AVDD.n5155 DGND 0.36fF $ **FLOATING
C7028 AVDD.n5156 DGND 0.36fF $ **FLOATING
C7029 AVDD.n5157 DGND 0.36fF $ **FLOATING
C7030 AVDD.n5158 DGND 0.35fF $ **FLOATING
C7031 AVDD.n5159 DGND 0.35fF $ **FLOATING
C7032 AVDD.n5160 DGND 0.35fF $ **FLOATING
C7033 AVDD.n5161 DGND 0.35fF $ **FLOATING
C7034 AVDD.n5162 DGND 0.36fF $ **FLOATING
C7035 AVDD.n5163 DGND 0.36fF $ **FLOATING
C7036 AVDD.t194 DGND 13.17fF
C7037 AVDD.n5194 DGND 0.19fF $ **FLOATING
C7038 AVDD.n5195 DGND 0.19fF $ **FLOATING
C7039 AVDD.n5196 DGND 0.29fF $ **FLOATING
C7040 AVDD.n5198 DGND 0.35fF $ **FLOATING
C7041 AVDD.n5199 DGND 0.35fF $ **FLOATING
C7042 AVDD.n5200 DGND 11.23fF $ **FLOATING
C7043 AVDD.n5201 DGND 0.36fF $ **FLOATING
C7044 AVDD.n5202 DGND 0.36fF $ **FLOATING
C7045 AVDD.n5203 DGND 0.36fF $ **FLOATING
C7046 AVDD.n5204 DGND 0.36fF $ **FLOATING
C7047 AVDD.n5205 DGND 0.35fF $ **FLOATING
C7048 AVDD.n5206 DGND 0.35fF $ **FLOATING
C7049 AVDD.n5207 DGND 0.41fF $ **FLOATING
C7050 AVDD.n5208 DGND 0.35fF $ **FLOATING
C7051 AVDD.n5209 DGND 0.35fF $ **FLOATING
C7052 AVDD.n5210 DGND 0.36fF $ **FLOATING
C7053 AVDD.n5211 DGND 0.36fF $ **FLOATING
C7054 AVDD.t203 DGND 13.15fF
C7055 AVDD.n5242 DGND 0.19fF $ **FLOATING
C7056 AVDD.n5243 DGND 0.19fF $ **FLOATING
C7057 AVDD.n5244 DGND 0.29fF $ **FLOATING
C7058 AVDD.n5246 DGND 0.35fF $ **FLOATING
C7059 AVDD.n5247 DGND 0.35fF $ **FLOATING
C7060 AVDD.n5248 DGND 17.55fF $ **FLOATING
C7061 AVDD.n5249 DGND 0.36fF $ **FLOATING
C7062 AVDD.t488 DGND 0.29fF
C7063 AVDD.n5250 DGND 0.33fF $ **FLOATING
C7064 AVDD.n5251 DGND 0.52fF $ **FLOATING
C7065 AVDD.n5252 DGND 0.39fF $ **FLOATING
C7066 AVDD.t659 DGND 0.29fF
C7067 AVDD.n5253 DGND 0.31fF $ **FLOATING
C7068 AVDD.n5254 DGND 0.47fF $ **FLOATING
C7069 AVDD.n5255 DGND 0.36fF $ **FLOATING
C7070 AVDD.n5256 DGND 0.28fF $ **FLOATING
C7071 AVDD.n5257 DGND 0.10fF $ **FLOATING
C7072 AVDD.n5258 DGND 0.35fF $ **FLOATING
C7073 AVDD.n5259 DGND 0.35fF $ **FLOATING
C7074 AVDD.n5260 DGND 0.36fF $ **FLOATING
C7075 AVDD.n5261 DGND 0.36fF $ **FLOATING
C7076 AVDD.t43 DGND 13.17fF
C7077 AVDD.n5292 DGND 0.19fF $ **FLOATING
C7078 AVDD.n5293 DGND 0.19fF $ **FLOATING
C7079 AVDD.n5294 DGND 0.29fF $ **FLOATING
C7080 AVDD.t458 DGND 0.29fF
C7081 AVDD.n5296 DGND 0.34fF $ **FLOATING
C7082 AVDD.n5297 DGND 0.58fF $ **FLOATING
C7083 AVDD.n5298 DGND 0.35fF $ **FLOATING
C7084 AVDD.n5299 DGND 0.26fF $ **FLOATING
C7085 AVDD.n5300 DGND 0.14fF $ **FLOATING
C7086 AVDD.n5301 DGND 17.35fF $ **FLOATING
C7087 AVDD.n5302 DGND 0.39fF $ **FLOATING
C7088 AVDD.n5303 DGND 0.36fF $ **FLOATING
C7089 AVDD.t500 DGND 0.29fF
C7090 AVDD.n5304 DGND 0.32fF $ **FLOATING
C7091 AVDD.n5305 DGND 0.47fF $ **FLOATING
C7092 AVDD.n5306 DGND 0.10fF $ **FLOATING
C7093 AVDD.n5307 DGND 0.29fF $ **FLOATING
C7094 AVDD.n5308 DGND 0.36fF $ **FLOATING
C7095 AVDD.n5309 DGND 0.35fF $ **FLOATING
C7096 AVDD.n5310 DGND 0.35fF $ **FLOATING
C7097 AVDD.n5311 DGND 0.36fF $ **FLOATING
C7098 AVDD.n5312 DGND 0.36fF $ **FLOATING
C7099 AVDD.t93 DGND 13.15fF
C7100 AVDD.n5343 DGND 0.19fF $ **FLOATING
C7101 AVDD.n5344 DGND 0.19fF $ **FLOATING
C7102 AVDD.n5345 DGND 0.29fF $ **FLOATING
C7103 AVDD.n5347 DGND 0.36fF $ **FLOATING
C7104 AVDD.t629 DGND 0.29fF
C7105 AVDD.n5348 DGND 0.36fF $ **FLOATING
C7106 AVDD.n5349 DGND 0.55fF $ **FLOATING
C7107 AVDD.n5350 DGND 0.11fF $ **FLOATING
C7108 AVDD.n5351 DGND 0.27fF $ **FLOATING
C7109 AVDD.n5352 DGND 0.35fF $ **FLOATING
C7110 AVDD.n5353 DGND 11.77fF $ **FLOATING
C7111 AVDD.n5354 DGND 0.36fF $ **FLOATING
C7112 AVDD.n5355 DGND 0.29fF $ **FLOATING
C7113 AVDD.t662 DGND 0.29fF
C7114 AVDD.n5356 DGND 0.33fF $ **FLOATING
C7115 AVDD.n5357 DGND 0.55fF $ **FLOATING
C7116 AVDD.n5358 DGND 0.11fF $ **FLOATING
C7117 AVDD.t111 DGND 13.17fF
C7118 AVDD.n5389 DGND 0.19fF $ **FLOATING
C7119 AVDD.n5390 DGND 0.19fF $ **FLOATING
C7120 AVDD.n5391 DGND 0.29fF $ **FLOATING
C7121 AVDD.n5393 DGND 0.35fF $ **FLOATING
C7122 AVDD.n5394 DGND 0.35fF $ **FLOATING
C7123 AVDD.n5395 DGND 0.35fF $ **FLOATING
C7124 AVDD.n5396 DGND 0.35fF $ **FLOATING
C7125 AVDD.n5397 DGND 17.20fF $ **FLOATING
C7126 AVDD.n5398 DGND 0.38fF $ **FLOATING
C7127 AVDD.n5399 DGND 0.36fF $ **FLOATING
C7128 AVDD.n5400 DGND 0.41fF $ **FLOATING
C7129 AVDD.n5401 DGND 0.36fF $ **FLOATING
C7130 AVDD.n5402 DGND 0.36fF $ **FLOATING
C7131 AVDD.n5403 DGND 0.36fF $ **FLOATING
C7132 AVDD.n5404 DGND 0.36fF $ **FLOATING
C7133 AVDD.n5405 DGND 0.35fF $ **FLOATING
C7134 AVDD.n5406 DGND 0.35fF $ **FLOATING
C7135 AVDD.t695 DGND 0.29fF
C7136 AVDD.n5407 DGND 0.33fF $ **FLOATING
C7137 AVDD.n5408 DGND 0.55fF $ **FLOATING
C7138 AVDD.n5409 DGND 0.11fF $ **FLOATING
C7139 AVDD.n5410 DGND 0.28fF $ **FLOATING
C7140 AVDD.n5411 DGND 0.36fF $ **FLOATING
C7141 AVDD.t105 DGND 13.15fF
C7142 AVDD.n5442 DGND 0.19fF $ **FLOATING
C7143 AVDD.n5443 DGND 0.19fF $ **FLOATING
C7144 AVDD.n5444 DGND 0.29fF $ **FLOATING
C7145 AVDD.n5446 DGND 0.35fF $ **FLOATING
C7146 AVDD.n5447 DGND 0.35fF $ **FLOATING
C7147 AVDD.n5448 DGND 0.35fF $ **FLOATING
C7148 AVDD.n5449 DGND 0.35fF $ **FLOATING
C7149 AVDD.n5450 DGND 12.82fF $ **FLOATING
C7150 AVDD.n5451 DGND 0.36fF $ **FLOATING
C7151 AVDD.n5452 DGND 0.36fF $ **FLOATING
C7152 AVDD.n5453 DGND 0.35fF $ **FLOATING
C7153 AVDD.n5454 DGND 0.35fF $ **FLOATING
C7154 AVDD.n5455 DGND 0.36fF $ **FLOATING
C7155 AVDD.n5456 DGND 0.36fF $ **FLOATING
C7156 AVDD.n5457 DGND 0.36fF $ **FLOATING
C7157 AVDD.n5458 DGND 0.36fF $ **FLOATING
C7158 AVDD.n5459 DGND 0.35fF $ **FLOATING
C7159 AVDD.n5460 DGND 0.35fF $ **FLOATING
C7160 AVDD.n5461 DGND 0.36fF $ **FLOATING
C7161 AVDD.n5462 DGND 0.36fF $ **FLOATING
C7162 AVDD.n5493 DGND 0.19fF $ **FLOATING
C7163 AVDD.n5494 DGND 0.19fF $ **FLOATING
C7164 AVDD.n5495 DGND 0.29fF $ **FLOATING
C7165 AVDD.n5497 DGND 0.35fF $ **FLOATING
C7166 AVDD.n5498 DGND 0.35fF $ **FLOATING
C7167 AVDD.n5499 DGND 0.35fF $ **FLOATING
C7168 AVDD.n5500 DGND 0.35fF $ **FLOATING
C7169 AVDD.n5501 DGND 17.77fF $ **FLOATING
C7170 AVDD.n5502 DGND 0.36fF $ **FLOATING
C7171 AVDD.n5503 DGND 0.36fF $ **FLOATING
C7172 AVDD.n5504 DGND 0.35fF $ **FLOATING
C7173 AVDD.n5505 DGND 0.35fF $ **FLOATING
C7174 AVDD.n5506 DGND 0.36fF $ **FLOATING
C7175 AVDD.n5507 DGND 0.36fF $ **FLOATING
C7176 AVDD.n5538 DGND 0.19fF $ **FLOATING
C7177 AVDD.n5539 DGND 0.19fF $ **FLOATING
C7178 AVDD.n5540 DGND 0.29fF $ **FLOATING
C7179 AVDD.n5542 DGND 0.35fF $ **FLOATING
C7180 AVDD.n5543 DGND 0.35fF $ **FLOATING
C7181 AVDD.n5544 DGND 0.35fF $ **FLOATING
C7182 AVDD.n5545 DGND 0.35fF $ **FLOATING
C7183 AVDD.n5546 DGND 6.63fF $ **FLOATING
C7184 AVDD.n5547 DGND 0.36fF $ **FLOATING
C7185 AVDD.n5548 DGND 0.36fF $ **FLOATING
C7186 AVDD.n5549 DGND 0.35fF $ **FLOATING
C7187 AVDD.n5550 DGND 0.35fF $ **FLOATING
C7188 AVDD.n5551 DGND 0.36fF $ **FLOATING
C7189 AVDD.n5552 DGND 0.36fF $ **FLOATING
C7190 AVDD.n5553 DGND 0.36fF $ **FLOATING
C7191 AVDD.n5554 DGND 0.36fF $ **FLOATING
C7192 AVDD.n5555 DGND 0.35fF $ **FLOATING
C7193 AVDD.n5556 DGND 0.35fF $ **FLOATING
C7194 AVDD.n5557 DGND 0.36fF $ **FLOATING
C7195 AVDD.n5558 DGND 0.36fF $ **FLOATING
C7196 AVDD.n5589 DGND 0.19fF $ **FLOATING
C7197 AVDD.n5590 DGND 0.19fF $ **FLOATING
C7198 AVDD.n5591 DGND 0.29fF $ **FLOATING
C7199 AVDD.n5593 DGND 0.35fF $ **FLOATING
C7200 AVDD.n5594 DGND 0.35fF $ **FLOATING
C7201 AVDD.n5595 DGND 0.35fF $ **FLOATING
C7202 AVDD.n5596 DGND 0.35fF $ **FLOATING
C7203 AVDD.n5597 DGND 17.52fF $ **FLOATING
C7204 AVDD.n5598 DGND 0.36fF $ **FLOATING
C7205 AVDD.n5599 DGND 0.36fF $ **FLOATING
C7206 AVDD.n5600 DGND 0.35fF $ **FLOATING
C7207 AVDD.n5601 DGND 0.35fF $ **FLOATING
C7208 AVDD.n5602 DGND 0.36fF $ **FLOATING
C7209 AVDD.n5603 DGND 0.36fF $ **FLOATING
C7210 AVDD.n5604 DGND 0.36fF $ **FLOATING
C7211 AVDD.n5605 DGND 0.36fF $ **FLOATING
C7212 AVDD.n5606 DGND 0.35fF $ **FLOATING
C7213 AVDD.n5607 DGND 0.35fF $ **FLOATING
C7214 AVDD.n5608 DGND 15.85fF $ **FLOATING
C7215 AVDD.n5609 DGND 0.36fF $ **FLOATING
C7216 AVDD.n5610 DGND 0.36fF $ **FLOATING
C7217 AVDD.n5611 DGND 0.36fF $ **FLOATING
C7218 AVDD.n5612 DGND 0.36fF $ **FLOATING
C7219 AVDD.n5613 DGND 0.35fF $ **FLOATING
C7220 AVDD.n5614 DGND 0.35fF $ **FLOATING
C7221 AVDD.n5615 DGND 0.36fF $ **FLOATING
C7222 AVDD.n5616 DGND 0.36fF $ **FLOATING
C7223 AVDD.n5617 DGND 0.36fF $ **FLOATING
C7224 AVDD.n5618 DGND 0.36fF $ **FLOATING
C7225 AVDD.n5619 DGND 0.35fF $ **FLOATING
C7226 AVDD.n5620 DGND 0.35fF $ **FLOATING
C7227 AVDD.n5621 DGND 10.10fF $ **FLOATING
C7228 AVDD.n5622 DGND 0.36fF $ **FLOATING
C7229 AVDD.n5623 DGND 0.36fF $ **FLOATING
C7230 AVDD.n5624 DGND 0.36fF $ **FLOATING
C7231 AVDD.n5625 DGND 0.36fF $ **FLOATING
C7232 AVDD.n5626 DGND 0.35fF $ **FLOATING
C7233 AVDD.n5627 DGND 0.35fF $ **FLOATING
C7234 AVDD.n5628 DGND 15.85fF $ **FLOATING
C7235 AVDD.n5629 DGND 0.36fF $ **FLOATING
C7236 AVDD.n5630 DGND 0.36fF $ **FLOATING
C7237 AVDD.n5631 DGND 0.36fF $ **FLOATING
C7238 AVDD.n5632 DGND 0.36fF $ **FLOATING
C7239 AVDD.n5633 DGND 0.35fF $ **FLOATING
C7240 AVDD.n5634 DGND 0.35fF $ **FLOATING
C7241 AVDD.n5635 DGND 11.10fF $ **FLOATING
C7242 AVDD.n5636 DGND 0.36fF $ **FLOATING
C7243 AVDD.n5637 DGND 0.36fF $ **FLOATING
C7244 AVDD.n5638 DGND 0.36fF $ **FLOATING
C7245 AVDD.n5639 DGND 0.36fF $ **FLOATING
C7246 AVDD.n5640 DGND 0.35fF $ **FLOATING
C7247 AVDD.n5641 DGND 0.35fF $ **FLOATING
C7248 AVDD.n5642 DGND 9.97fF $ **FLOATING
C7249 AVDD.n5643 DGND 0.36fF $ **FLOATING
C7250 AVDD.n5644 DGND 0.36fF $ **FLOATING
C7251 AVDD.n5645 DGND 0.36fF $ **FLOATING
C7252 AVDD.n5646 DGND 0.36fF $ **FLOATING
C7253 AVDD.n5647 DGND 0.39fF $ **FLOATING
C7254 AVDD.n5648 DGND 0.35fF $ **FLOATING
C7255 AVDD.n5649 DGND 0.35fF $ **FLOATING
C7256 AVDD.n5650 DGND 11.10fF $ **FLOATING
C7257 AVDD.n5651 DGND 0.36fF $ **FLOATING
C7258 AVDD.n5652 DGND 0.36fF $ **FLOATING
C7259 AVDD.n5653 DGND 0.36fF $ **FLOATING
C7260 AVDD.n5654 DGND 0.36fF $ **FLOATING
C7261 AVDD.n5655 DGND 0.36fF $ **FLOATING
C7262 AVDD.n5656 DGND 0.36fF $ **FLOATING
C7263 AVDD.n5657 DGND 4.32fF $ **FLOATING
C7264 AVDD.n5658 DGND 0.36fF $ **FLOATING
C7265 AVDD.n5659 DGND 0.36fF $ **FLOATING
C7266 AVDD.n5660 DGND 0.36fF $ **FLOATING
C7267 AVDD.n5661 DGND 0.36fF $ **FLOATING
C7268 AVDD.n5663 DGND 0.19fF $ **FLOATING
C7269 AVDD.n5664 DGND 0.19fF $ **FLOATING
C7270 AVDD.n5665 DGND 0.29fF $ **FLOATING
C7271 AVDD.n5697 DGND 0.77fF $ **FLOATING
C7272 AVDD.n5698 DGND 0.53fF $ **FLOATING
C7273 AVDD.n5702 DGND 0.86fF $ **FLOATING
C7274 AVDD.t401 DGND 3.07fF
C7275 AVDD.t827 DGND 3.87fF
C7276 AVDD.t281 DGND 4.64fF
C7277 AVDD.n5704 DGND 2.28fF $ **FLOATING
C7278 AVDD.n5709 DGND 0.56fF $ **FLOATING
C7279 AVDD.n5710 DGND 0.30fF $ **FLOATING
C7280 AVDD.n5711 DGND 0.36fF $ **FLOATING
C7281 AVDD.n5712 DGND 0.36fF $ **FLOATING
C7282 AVDD.n5713 DGND 0.77fF $ **FLOATING
C7283 AVDD.n5714 DGND 0.53fF $ **FLOATING
C7284 AVDD.n5718 DGND 0.77fF $ **FLOATING
C7285 AVDD.n5719 DGND 0.42fF $ **FLOATING
C7286 AVDD.n5722 DGND 0.74fF $ **FLOATING
C7287 AVDD.n5726 DGND 0.77fF $ **FLOATING
C7288 AVDD.n5727 DGND 0.42fF $ **FLOATING
C7289 AVDD.n5730 DGND 0.74fF $ **FLOATING
C7290 AVDD.n5734 DGND 0.77fF $ **FLOATING
C7291 AVDD.n5735 DGND 0.42fF $ **FLOATING
C7292 AVDD.n5738 DGND 0.74fF $ **FLOATING
C7293 AVDD.t370 DGND 8.66fF
C7294 AVDD.n5740 DGND 5.79fF $ **FLOATING
C7295 AVDD.n5744 DGND 0.77fF $ **FLOATING
C7296 AVDD.n5745 DGND 0.41fF $ **FLOATING
C7297 AVDD.n5748 DGND 0.73fF $ **FLOATING
C7298 AVDD.n5753 DGND 0.20fF $ **FLOATING
C7299 AVDD.n5754 DGND 0.41fF $ **FLOATING
C7300 AVDD.n5755 DGND 0.43fF $ **FLOATING
C7301 AVDD.n5758 DGND 4.58fF $ **FLOATING
C7302 AVDD.n5767 DGND 0.25fF $ **FLOATING
C7303 AVDD.n5770 DGND 0.20fF $ **FLOATING
C7304 AVDD.n5771 DGND 0.41fF $ **FLOATING
C7305 AVDD.n5772 DGND 0.77fF $ **FLOATING
C7306 AVDD.n5773 DGND 0.42fF $ **FLOATING
C7307 AVDD.n5774 DGND 0.41fF $ **FLOATING
C7308 AVDD.n5784 DGND 0.25fF $ **FLOATING
C7309 AVDD.n5787 DGND 0.20fF $ **FLOATING
C7310 AVDD.n5788 DGND 0.41fF $ **FLOATING
C7311 AVDD.n5789 DGND 0.77fF $ **FLOATING
C7312 AVDD.n5790 DGND 0.42fF $ **FLOATING
C7313 AVDD.n5791 DGND 0.41fF $ **FLOATING
C7314 AVDD.n5795 DGND 0.20fF $ **FLOATING
C7315 AVDD.n5796 DGND 0.41fF $ **FLOATING
C7316 AVDD.n5797 DGND 0.43fF $ **FLOATING
C7317 AVDD.n5813 DGND 1.74fF $ **FLOATING
C7318 AVDD.n5814 DGND 0.11fF $ **FLOATING
C7319 AVDD.n5815 DGND 0.18fF $ **FLOATING
C7320 AVDD.n5816 DGND 0.81fF $ **FLOATING
C7321 AVDD.n5817 DGND 0.73fF $ **FLOATING
C7322 AVDD.n5827 DGND 0.99fF $ **FLOATING
C7323 level_shifter_up_5.VDD_HV DGND 0.29fF $ **FLOATING
C7324 AVDD.t52 DGND 7.15fF
C7325 AVDD.n5828 DGND 0.20fF $ **FLOATING
C7326 AVDD.n5832 DGND 0.16fF $ **FLOATING
C7327 AVDD.n5835 DGND 0.10fF $ **FLOATING
C7328 AVDD.n5837 DGND 0.63fF $ **FLOATING
C7329 AVDD.t341 DGND 0.89fF
C7330 AVDD.n5849 DGND 0.16fF $ **FLOATING
C7331 AVDD.n5858 DGND 0.51fF $ **FLOATING
C7332 AVDD.t287 DGND 4.07fF
C7333 AVDD.n5875 DGND 2.28fF $ **FLOATING
C7334 AVDD.t820 DGND 2.67fF
C7335 AVDD.n5876 DGND 0.76fF $ **FLOATING
C7336 AVDD.n5884 DGND 0.12fF $ **FLOATING
C7337 AVDD.n5885 DGND 0.16fF $ **FLOATING
C7338 AVDD.n5890 DGND 0.77fF $ **FLOATING
C7339 AVDD.t727 DGND 1.72fF
C7340 AVDD.n5893 DGND 0.76fF $ **FLOATING
C7341 AVDD.n5895 DGND 0.21fF $ **FLOATING
C7342 AVDD.n5898 DGND 0.13fF $ **FLOATING
C7343 AVDD.t20 DGND 2.09fF
C7344 AVDD.n5900 DGND 0.83fF $ **FLOATING
C7345 AVDD.t59 DGND 3.24fF
C7346 AVDD.t351 DGND 3.89fF
C7347 AVDD.t264 DGND 0.51fF
C7348 AVDD.n5915 DGND 1.12fF $ **FLOATING
C7349 AVDD.t147 DGND 2.44fF
C7350 AVDD.t279 DGND 4.87fF
C7351 AVDD.n5916 DGND 0.11fF $ **FLOATING
C7352 AVDD.n5917 DGND 0.46fF $ **FLOATING
C7353 AVDD.n5919 DGND 1.22fF $ **FLOATING
C7354 AVDD.t818 DGND 0.89fF
C7355 AVDD.n5927 DGND 0.16fF $ **FLOATING
C7356 AVDD.n5933 DGND 0.11fF $ **FLOATING
C7357 AVDD.n5934 DGND 0.18fF $ **FLOATING
C7358 AVDD.n5935 DGND 0.76fF $ **FLOATING
C7359 AVDD.n5952 DGND 2.28fF $ **FLOATING
C7360 AVDD.t814 DGND 2.51fF
C7361 AVDD.n6001 DGND 2.28fF $ **FLOATING
C7362 AVDD.n6051 DGND 2.28fF $ **FLOATING
C7363 AVDD.t829 DGND 3.08fF
C7364 AVDD.t95 DGND 0.76fF
C7365 AVDD.n6058 DGND 0.16fF $ **FLOATING
C7366 AVDD.n6062 DGND 0.20fF $ **FLOATING
C7367 AVDD.n6063 DGND 0.11fF $ **FLOATING
C7368 AVDD.n6064 DGND 0.18fF $ **FLOATING
C7369 AVDD.n6065 DGND 0.11fF $ **FLOATING
C7370 AVDD.n6066 DGND 0.18fF $ **FLOATING
C7371 AVDD.t344 DGND 0.75fF
C7372 AVDD.t361 DGND 3.54fF
C7373 AVDD.t21 DGND 2.28fF
C7374 AVDD.t357 DGND 5.06fF
C7375 AVDD.t275 DGND 1.12fF
C7376 level_shifter_up_0.VDD_HV DGND 0.13fF $ **FLOATING
C7377 AVDD.n6069 DGND 0.22fF $ **FLOATING
C7378 AVDD.n6071 DGND 0.12fF $ **FLOATING
C7379 AVDD.n6072 DGND 0.16fF $ **FLOATING
C7380 AVDD.t266 DGND 0.76fF
C7381 AVDD.t353 DGND 0.64fF
C7382 AVDD.n6086 DGND 0.11fF $ **FLOATING
C7383 AVDD.n6087 DGND 0.18fF $ **FLOATING
C7384 AVDD.n6088 DGND 0.11fF $ **FLOATING
C7385 AVDD.n6089 DGND 0.18fF $ **FLOATING
C7386 AVDD.t35 DGND 0.27fF
C7387 AVDD.t359 DGND 2.58fF
C7388 AVDD.t494 DGND 0.28fF
C7389 AVDD.t470 DGND 0.28fF
C7390 AVDD.n6095 DGND 0.21fF $ **FLOATING
C7391 AVDD.n6097 DGND 1.91fF $ **FLOATING
C7392 AVDD.t656 DGND 0.28fF
C7393 AVDD.t626 DGND 0.28fF
C7394 AVDD.n6099 DGND 0.21fF $ **FLOATING
C7395 AVDD.n6101 DGND 1.91fF $ **FLOATING
C7396 AVDD.n6105 DGND 2.28fF $ **FLOATING
C7397 AVDD.n6110 DGND 0.76fF $ **FLOATING
C7398 AVDD.t363 DGND 3.13fF
C7399 AVDD.t831 DGND 5.01fF
C7400 AVDD.t825 DGND 5.02fF
C7401 AVDD.t581 DGND 0.28fF
C7402 AVDD.t539 DGND 0.28fF
C7403 AVDD.n6123 DGND 0.21fF $ **FLOATING
C7404 AVDD.n6125 DGND 1.91fF $ **FLOATING
C7405 AVDD.n6128 DGND 0.21fF $ **FLOATING
C7406 AVDD.n6129 DGND 0.12fF $ **FLOATING
C7407 AVDD.t431 DGND 0.28fF
C7408 AVDD.t473 DGND 0.28fF
C7409 AVDD.n6131 DGND 1.91fF $ **FLOATING
C7410 AVDD.n6138 DGND 2.28fF $ **FLOATING
C7411 AVDD.n6142 DGND 0.25fF $ **FLOATING
C7412 AVDD.n6145 DGND 0.20fF $ **FLOATING
C7413 AVDD.n6146 DGND 0.41fF $ **FLOATING
C7414 AVDD.n6147 DGND 1.07fF $ **FLOATING
C7415 AVDD.n6148 DGND 0.41fF $ **FLOATING
C7416 AVDD.n6152 DGND 0.20fF $ **FLOATING
C7417 AVDD.n6153 DGND 0.41fF $ **FLOATING
C7418 AVDD.n6154 DGND 0.43fF $ **FLOATING
C7419 AVDD.t437 DGND 0.28fF
C7420 AVDD.t400 DGND 0.28fF
C7421 AVDD.n6163 DGND 0.21fF $ **FLOATING
C7422 AVDD.n6165 DGND 1.91fF $ **FLOATING
C7423 AVDD.n6169 DGND 0.21fF $ **FLOATING
C7424 AVDD.n6170 DGND 0.12fF $ **FLOATING
C7425 AVDD.t614 DGND 0.28fF
C7426 AVDD.t647 DGND 0.28fF
C7427 AVDD.n6172 DGND 1.91fF $ **FLOATING
C7428 AVDD.t506 DGND 0.28fF
C7429 AVDD.t479 DGND 0.28fF
C7430 AVDD.n6176 DGND 0.21fF $ **FLOATING
C7431 AVDD.n6178 DGND 1.91fF $ **FLOATING
C7432 AVDD.t560 DGND 0.28fF
C7433 AVDD.t428 DGND 0.28fF
C7434 AVDD.n6180 DGND 0.21fF $ **FLOATING
C7435 AVDD.n6182 DGND 1.90fF $ **FLOATING
C7436 AVDD.n6184 DGND 10.51fF $ **FLOATING
C7437 AVDD.n6186 DGND 0.25fF $ **FLOATING
C7438 AVDD.n6189 DGND 0.20fF $ **FLOATING
C7439 AVDD.n6190 DGND 0.41fF $ **FLOATING
C7440 AVDD.n6191 DGND 1.07fF $ **FLOATING
C7441 AVDD.n6192 DGND 0.41fF $ **FLOATING
C7442 AVDD.n6196 DGND 0.20fF $ **FLOATING
C7443 AVDD.n6197 DGND 0.41fF $ **FLOATING
C7444 AVDD.n6198 DGND 0.43fF $ **FLOATING
C7445 AVDD.n6208 DGND 0.25fF $ **FLOATING
C7446 AVDD.n6211 DGND 0.20fF $ **FLOATING
C7447 AVDD.n6212 DGND 0.41fF $ **FLOATING
C7448 AVDD.n6213 DGND 0.77fF $ **FLOATING
C7449 AVDD.n6214 DGND 0.42fF $ **FLOATING
C7450 AVDD.n6215 DGND 0.41fF $ **FLOATING
C7451 AVDD.n6219 DGND 0.20fF $ **FLOATING
C7452 AVDD.n6220 DGND 0.41fF $ **FLOATING
C7453 AVDD.n6221 DGND 0.43fF $ **FLOATING
C7454 AVDD.n6231 DGND 0.25fF $ **FLOATING
C7455 AVDD.n6234 DGND 0.20fF $ **FLOATING
C7456 AVDD.n6235 DGND 0.41fF $ **FLOATING
C7457 AVDD.n6236 DGND 0.77fF $ **FLOATING
C7458 AVDD.n6237 DGND 0.42fF $ **FLOATING
C7459 AVDD.n6238 DGND 0.41fF $ **FLOATING
C7460 AVDD.n6242 DGND 0.20fF $ **FLOATING
C7461 AVDD.n6243 DGND 0.41fF $ **FLOATING
C7462 AVDD.n6244 DGND 0.43fF $ **FLOATING
C7463 AVDD.n6254 DGND 0.25fF $ **FLOATING
C7464 AVDD.n6257 DGND 0.20fF $ **FLOATING
C7465 AVDD.n6258 DGND 0.41fF $ **FLOATING
C7466 AVDD.n6259 DGND 0.77fF $ **FLOATING
C7467 AVDD.n6260 DGND 0.42fF $ **FLOATING
C7468 AVDD.n6261 DGND 0.41fF $ **FLOATING
C7469 AVDD.n6265 DGND 0.20fF $ **FLOATING
C7470 AVDD.n6266 DGND 0.41fF $ **FLOATING
C7471 AVDD.n6267 DGND 0.43fF $ **FLOATING
C7472 AVDD.n6277 DGND 0.25fF $ **FLOATING
C7473 AVDD.n6280 DGND 0.19fF $ **FLOATING
C7474 AVDD.n6281 DGND 0.40fF $ **FLOATING
C7475 AVDD.n6282 DGND 0.74fF $ **FLOATING
C7476 AVDD.n6283 DGND 0.41fF $ **FLOATING
C7477 AVDD.n6284 DGND 0.41fF $ **FLOATING
C7478 AVDD.n6288 DGND 0.19fF $ **FLOATING
C7479 AVDD.n6289 DGND 0.40fF $ **FLOATING
C7480 AVDD.n6290 DGND 0.94fF $ **FLOATING
C7481 AVDD.n6292 DGND 0.77fF $ **FLOATING
C7482 AVDD.n6293 DGND 0.40fF $ **FLOATING
C7483 AVDD.n6294 DGND 0.19fF $ **FLOATING
C7484 AVDD.n6296 DGND 0.77fF $ **FLOATING
C7485 AVDD.n6297 DGND 0.42fF $ **FLOATING
C7486 AVDD.n6300 DGND 0.74fF $ **FLOATING
C7487 AVDD.n6303 DGND 7.67fF $ **FLOATING
C7488 AVDD.n6306 DGND 0.56fF $ **FLOATING
C7489 AVDD.n6307 DGND 0.30fF $ **FLOATING
C7490 AVDD.n6308 DGND 0.36fF $ **FLOATING
C7491 AVDD.n6309 DGND 0.36fF $ **FLOATING
C7492 AVDD.n6310 DGND 0.11fF $ **FLOATING
C7493 AVDD.n6311 DGND 0.18fF $ **FLOATING
C7494 AVDD.n6312 DGND 0.70fF $ **FLOATING
C7495 AVDD.n6315 DGND 0.37fF $ **FLOATING
C7496 AVDD.n6316 DGND 0.11fF $ **FLOATING
C7497 AVDD.n6317 DGND 0.18fF $ **FLOATING
C7498 AVDD.n6318 DGND 0.59fF $ **FLOATING
C7499 AVDD.n6321 DGND 0.26fF $ **FLOATING
C7500 AVDD.t48 DGND 2.28fF
C7501 AVDD.t285 DGND 3.31fF
C7502 AVDD.t816 DGND 3.81fF
C7503 AVDD.n6323 DGND 0.15fF $ **FLOATING
C7504 AVDD.n6324 DGND 1.83fF $ **FLOATING
C7505 AVDD.t283 DGND 3.86fF
C7506 AVDD.n6355 DGND 0.19fF $ **FLOATING
C7507 AVDD.n6356 DGND 0.30fF $ **FLOATING
C7508 AVDD.n6358 DGND 4.42fF $ **FLOATING
C7509 AVDD.n6359 DGND 4.39fF $ **FLOATING
C7510 AVDD.n6362 DGND 1.17fF $ **FLOATING
C7511 AVDD.n6366 DGND 0.14fF $ **FLOATING
C7512 AVDD.n6368 DGND 0.14fF $ **FLOATING
C7513 AVDD.n6369 DGND 0.30fF $ **FLOATING
C7514 AVDD.t97 DGND 2.38fF
C7515 AVDD.t9 DGND 1.14fF
C7516 AVDD.n6375 DGND 1.90fF $ **FLOATING
C7517 AVDD.t87 DGND 1.27fF
C7518 AVDD.n6376 DGND 2.26fF $ **FLOATING
C7519 AVDD.n6378 DGND 0.28fF $ **FLOATING
C7520 AVDD.n6389 DGND 0.18fF $ **FLOATING
C7521 AVDD.n6393 DGND 0.38fF $ **FLOATING
C7522 AVDD.n6394 DGND 0.64fF $ **FLOATING
C7523 AVDD.n6398 DGND 0.14fF $ **FLOATING
C7524 AVDD.t355 DGND 3.69fF
C7525 AVDD.n6403 DGND 0.38fF $ **FLOATING
C7526 AVDD.n6404 DGND 0.38fF $ **FLOATING
C7527 AVDD.n6405 DGND 0.50fF $ **FLOATING
C7528 AVDD.n6408 DGND 0.95fF $ **FLOATING
C7529 AVDD.n6409 DGND 0.51fF $ **FLOATING
C7530 AVDD.n6410 DGND 1.12fF $ **FLOATING
C7531 AVDD.n6411 DGND 1.27fF $ **FLOATING
C7532 AVDD.n6419 DGND 0.20fF $ **FLOATING
C7533 AVDD.n6422 DGND 2.28fF $ **FLOATING
C7534 AVDD.t808 DGND 2.27fF
C7535 AVDD.n6429 DGND 0.17fF $ **FLOATING
C7536 AVDD.n6430 DGND 0.12fF $ **FLOATING
C7537 AVDD.n6441 DGND 1.83fF $ **FLOATING
C7538 AVDD.n6490 DGND 2.15fF $ **FLOATING
C7539 AVDD.n6496 DGND 1.46fF $ **FLOATING
C7540 AVDD.t810 DGND 1.68fF
C7541 AVDD.n6500 DGND 1.73fF $ **FLOATING
C7542 AVDD.n6549 DGND 0.82fF $ **FLOATING
C7543 AVDD.n6567 DGND 2.15fF $ **FLOATING
C7544 AVDD.t99 DGND 1.30fF
C7545 AVDD.t812 DGND 2.26fF
C7546 AVDD.t31 DGND 1.12fF
C7547 level_shifter_up_4.VDD_HV DGND 0.13fF $ **FLOATING
C7548 a_1659_n4497.n0 DGND 1.61fF $ **FLOATING
C7549 a_1659_n4497.n1 DGND 1.64fF $ **FLOATING
C7550 a_1659_n4497.n2 DGND 1.34fF $ **FLOATING
C7551 a_1659_n4497.n3 DGND 1.61fF $ **FLOATING
C7552 a_1659_n4497.n4 DGND 1.64fF $ **FLOATING
C7553 a_1659_n4497.n5 DGND 1.61fF $ **FLOATING
C7554 a_1659_n4497.n6 DGND 1.64fF $ **FLOATING
C7555 a_1659_n4497.n7 DGND 1.34fF $ **FLOATING
C7556 a_1659_n4497.n8 DGND 2.03fF $ **FLOATING
C7557 a_1659_n4497.n9 DGND 1.61fF $ **FLOATING
C7558 a_1659_n4497.n10 DGND 1.64fF $ **FLOATING
C7559 a_1659_n4497.n11 DGND 2.03fF $ **FLOATING
C7560 a_1659_n4497.n12 DGND 1.77fF $ **FLOATING
C7561 a_1659_n4497.n13 DGND 1.77fF $ **FLOATING
C7562 a_1659_n4497.n14 DGND 1.64fF $ **FLOATING
C7563 a_1659_n4497.n15 DGND 1.64fF $ **FLOATING
C7564 a_1659_n4497.n16 DGND 1.77fF $ **FLOATING
C7565 a_1659_n4497.n17 DGND 1.34fF $ **FLOATING
C7566 a_1659_n4497.n18 DGND 1.64fF $ **FLOATING
C7567 a_1659_n4497.n19 DGND 1.77fF $ **FLOATING
C7568 a_1659_n4497.n20 DGND 1.34fF $ **FLOATING
C7569 a_1659_n4497.n21 DGND 1.77fF $ **FLOATING
C7570 a_1659_n4497.n22 DGND 1.64fF $ **FLOATING
C7571 a_1659_n4497.n23 DGND 1.64fF $ **FLOATING
C7572 a_1659_n4497.n24 DGND 1.77fF $ **FLOATING
C7573 a_1659_n4497.n25 DGND 1.34fF $ **FLOATING
C7574 a_1659_n4497.n26 DGND 1.64fF $ **FLOATING
C7575 a_1659_n4497.n27 DGND 1.77fF $ **FLOATING
C7576 a_1659_n4497.n28 DGND 1.34fF $ **FLOATING
C7577 a_1659_n4497.n29 DGND 1.77fF $ **FLOATING
C7578 a_1659_n4497.n30 DGND 1.64fF $ **FLOATING
C7579 a_1659_n4497.n31 DGND 1.64fF $ **FLOATING
C7580 a_1659_n4497.n32 DGND 1.77fF $ **FLOATING
C7581 a_1659_n4497.n33 DGND 2.03fF $ **FLOATING
C7582 a_1659_n4497.n34 DGND 1.64fF $ **FLOATING
C7583 a_1659_n4497.n35 DGND 1.77fF $ **FLOATING
C7584 a_1659_n4497.n36 DGND 2.03fF $ **FLOATING
C7585 a_1659_n4497.n37 DGND 2.63fF $ **FLOATING
C7586 a_1659_n4497.n38 DGND 1.77fF $ **FLOATING
C7587 a_1659_n4497.n39 DGND 1.34fF $ **FLOATING
C7588 a_1659_n4497.n40 DGND 1.64fF $ **FLOATING
C7589 a_1659_n4497.n41 DGND 1.77fF $ **FLOATING
C7590 a_1659_n4497.n42 DGND 1.34fF $ **FLOATING
C7591 a_1659_n4497.n43 DGND 1.64fF $ **FLOATING
C7592 a_1659_n4497.n44 DGND 1.77fF $ **FLOATING
C7593 a_1659_n4497.n45 DGND 1.34fF $ **FLOATING
C7594 a_1659_n4497.n46 DGND 2.63fF $ **FLOATING
C7595 a_1659_n4497.n47 DGND 1.77fF $ **FLOATING
C7596 a_1659_n4497.n48 DGND 1.34fF $ **FLOATING
C7597 a_1659_n4497.n49 DGND 1.64fF $ **FLOATING
C7598 a_1659_n4497.n50 DGND 1.77fF $ **FLOATING
C7599 a_1659_n4497.n51 DGND 2.03fF $ **FLOATING
C7600 a_1659_n4497.n52 DGND 1.64fF $ **FLOATING
C7601 a_1659_n4497.n53 DGND 1.77fF $ **FLOATING
C7602 a_1659_n4497.n54 DGND 2.03fF $ **FLOATING
C7603 a_1659_n4497.n55 DGND 1.92fF $ **FLOATING
C7604 a_1659_n4497.n56 DGND 1.92fF $ **FLOATING
C7605 a_1659_n4497.n57 DGND 1.64fF $ **FLOATING
C7606 a_1659_n4497.n58 DGND 1.77fF $ **FLOATING
C7607 a_1659_n4497.n59 DGND 2.03fF $ **FLOATING
C7608 a_1659_n4497.n60 DGND 1.64fF $ **FLOATING
C7609 a_1659_n4497.n61 DGND 1.77fF $ **FLOATING
C7610 a_1659_n4497.n62 DGND 2.03fF $ **FLOATING
C7611 a_1659_n4497.n63 DGND 1.64fF $ **FLOATING
C7612 a_1659_n4497.n64 DGND 1.77fF $ **FLOATING
C7613 a_1659_n4497.n65 DGND 2.03fF $ **FLOATING
C7614 a_1659_n4497.n66 DGND 1.64fF $ **FLOATING
C7615 a_1659_n4497.n67 DGND 1.77fF $ **FLOATING
C7616 a_1659_n4497.n68 DGND 2.03fF $ **FLOATING
C7617 a_1659_n4497.n69 DGND 1.64fF $ **FLOATING
C7618 Vxm.n0 DGND 0.79fF $ **FLOATING
C7619 Vxm.n1 DGND 1.63fF $ **FLOATING
C7620 Vxm.n2 DGND 1.32fF $ **FLOATING
C7621 Vxm.n3 DGND 1.63fF $ **FLOATING
C7622 Vxm.n4 DGND 0.79fF $ **FLOATING
C7623 Vxm.n5 DGND 2.02fF $ **FLOATING
C7624 Vxm.n6 DGND 1.63fF $ **FLOATING
C7625 Vxm.n7 DGND 0.79fF $ **FLOATING
C7626 Vxm.n8 DGND 2.02fF $ **FLOATING
C7627 Vxm.n9 DGND 1.63fF $ **FLOATING
C7628 Vxm.n10 DGND 0.79fF $ **FLOATING
C7629 Vxm.n11 DGND 2.35fF $ **FLOATING
C7630 Vxm.t22 DGND 0.19fF
C7631 Vxm.t20 DGND 0.19fF
C7632 Vxm.t10 DGND 0.19fF
C7633 Vxm.n12 DGND 4.63fF $ **FLOATING
C7634 Vxm.n13 DGND 4.63fF $ **FLOATING
C7635 Vxm.n14 DGND 4.45fF $ **FLOATING
C7636 Vxm.t15 DGND 0.19fF
C7637 Vxm.t29 DGND 0.19fF
C7638 Vxm.n15 DGND 4.63fF $ **FLOATING
C7639 Vxm.t0 DGND 0.19fF
C7640 Vxm.n16 DGND 4.63fF $ **FLOATING
C7641 Vxm.n17 DGND 4.85fF $ **FLOATING
C7642 Vxm.n18 DGND 3.77fF $ **FLOATING
C7643 Vxm.t43 DGND 0.19fF
C7644 Vxm.t32 DGND 0.19fF
C7645 Vxm.n19 DGND 4.63fF $ **FLOATING
C7646 Vxm.n20 DGND 5.04fF $ **FLOATING
C7647 Vxm.n21 DGND 2.29fF $ **FLOATING
C7648 Vxm.t39 DGND 0.19fF
C7649 Vxm.t7 DGND 0.19fF
C7650 Vxm.n22 DGND 4.63fF $ **FLOATING
C7651 Vxm.n23 DGND 5.04fF $ **FLOATING
C7652 Vxm.n24 DGND 2.29fF $ **FLOATING
C7653 Vxm.t12 DGND 0.19fF
C7654 Vxm.t101 DGND 0.19fF
C7655 Vxm.n25 DGND 4.63fF $ **FLOATING
C7656 Vxm.n26 DGND 5.04fF $ **FLOATING
C7657 Vxm.n27 DGND 2.29fF $ **FLOATING
C7658 Vxm.t102 DGND 0.19fF
C7659 Vxm.t24 DGND 0.19fF
C7660 Vxm.n28 DGND 4.63fF $ **FLOATING
C7661 Vxm.n29 DGND 5.04fF $ **FLOATING
C7662 Vxm.n30 DGND 2.29fF $ **FLOATING
C7663 Vxm.t40 DGND 0.19fF
C7664 Vxm.t33 DGND 0.19fF
C7665 Vxm.t16 DGND 0.19fF
C7666 Vxm.n31 DGND 4.63fF $ **FLOATING
C7667 Vxm.n32 DGND 4.63fF $ **FLOATING
C7668 Vxm.n33 DGND 4.45fF $ **FLOATING
C7669 Vxm.n34 DGND 1.80fF $ **FLOATING
C7670 Vxm.t13 DGND 0.19fF
C7671 Vxm.t2 DGND 0.19fF
C7672 Vxm.t11 DGND 0.19fF
C7673 Vxm.n35 DGND 4.63fF $ **FLOATING
C7674 Vxm.n36 DGND 4.63fF $ **FLOATING
C7675 Vxm.n37 DGND 4.45fF $ **FLOATING
C7676 Vxm.n38 DGND 11.77fF $ **FLOATING
C7677 Vxm.n39 DGND 12.97fF $ **FLOATING
C7678 Vxm.n40 DGND 0.79fF $ **FLOATING
C7679 Vxm.n41 DGND 0.91fF $ **FLOATING
C7680 Vxm.n42 DGND 0.91fF $ **FLOATING
C7681 Vxm.n43 DGND 0.79fF $ **FLOATING
C7682 Vxm.n44 DGND 1.32fF $ **FLOATING
C7683 Vxm.n45 DGND 2.02fF $ **FLOATING
C7684 Vxm.n46 DGND 0.91fF $ **FLOATING
C7685 Vxm.n47 DGND 0.79fF $ **FLOATING
C7686 Vxm.n48 DGND 2.02fF $ **FLOATING
C7687 Vxm.n49 DGND 0.91fF $ **FLOATING
C7688 Vxm.n50 DGND 0.79fF $ **FLOATING
C7689 Vxm.n51 DGND 2.35fF $ **FLOATING
C7690 Vxm.n52 DGND 3.90fF $ **FLOATING
C7691 Vxm.n53 DGND 0.91fF $ **FLOATING
C7692 Vxm.n54 DGND 0.79fF $ **FLOATING
C7693 Vxm.n55 DGND 1.32fF $ **FLOATING
C7694 Vxm.n56 DGND 0.91fF $ **FLOATING
C7695 Vxm.n57 DGND 0.79fF $ **FLOATING
C7696 Vxm.n58 DGND 2.02fF $ **FLOATING
C7697 Vxm.n59 DGND 0.91fF $ **FLOATING
C7698 Vxm.n60 DGND 0.79fF $ **FLOATING
C7699 Vxm.n61 DGND 2.02fF $ **FLOATING
C7700 Vxm.n62 DGND 0.91fF $ **FLOATING
C7701 Vxm.n63 DGND 0.79fF $ **FLOATING
C7702 Vxm.n64 DGND 2.35fF $ **FLOATING
C7703 Vxm.n65 DGND 3.23fF $ **FLOATING
C7704 Vxm.n66 DGND 2.16fF $ **FLOATING
C7705 Vxm.n67 DGND 1.90fF $ **FLOATING
C7706 Vxm.n68 DGND 2.29fF $ **FLOATING
C7707 Vxm.t44 DGND 0.19fF
C7708 Vxm.t14 DGND 0.19fF
C7709 Vxm.t45 DGND 0.19fF
C7710 Vxm.t103 DGND 0.19fF
C7711 Vxm.t6 DGND 0.19fF
C7712 Vxm.n69 DGND 4.63fF $ **FLOATING
C7713 Vxm.n70 DGND 4.63fF $ **FLOATING
C7714 Vxm.n71 DGND 4.63fF $ **FLOATING
C7715 Vxm.n72 DGND 4.63fF $ **FLOATING
C7716 Vxm.n73 DGND 4.45fF $ **FLOATING
C7717 Vxm.t21 DGND 0.19fF
C7718 Vxm.t23 DGND 0.19fF
C7719 Vxm.t9 DGND 0.19fF
C7720 Vxm.t99 DGND 0.19fF
C7721 Vxm.t95 DGND 0.19fF
C7722 Vxm.n74 DGND 4.63fF $ **FLOATING
C7723 Vxm.n75 DGND 4.63fF $ **FLOATING
C7724 Vxm.n76 DGND 4.63fF $ **FLOATING
C7725 Vxm.n77 DGND 4.63fF $ **FLOATING
C7726 Vxm.n78 DGND 4.45fF $ **FLOATING
C7727 Vxm.t27 DGND 0.19fF
C7728 Vxm.t28 DGND 0.19fF
C7729 Vxm.t5 DGND 0.19fF
C7730 Vxm.t4 DGND 0.19fF
C7731 Vxm.n79 DGND 4.63fF $ **FLOATING
C7732 Vxm.n80 DGND 4.63fF $ **FLOATING
C7733 Vxm.n81 DGND 4.63fF $ **FLOATING
C7734 Vxm.n82 DGND 5.04fF $ **FLOATING
C7735 Vxm.t42 DGND 0.19fF
C7736 Vxm.t17 DGND 0.19fF
C7737 Vxm.t96 DGND 0.19fF
C7738 Vxm.t3 DGND 0.19fF
C7739 Vxm.n83 DGND 4.63fF $ **FLOATING
C7740 Vxm.n84 DGND 4.63fF $ **FLOATING
C7741 Vxm.n85 DGND 4.63fF $ **FLOATING
C7742 Vxm.n86 DGND 5.04fF $ **FLOATING
C7743 Vxm.t18 DGND 0.19fF
C7744 Vxm.t31 DGND 0.19fF
C7745 Vxm.t1 DGND 0.19fF
C7746 Vxm.t26 DGND 0.19fF
C7747 Vxm.n87 DGND 4.63fF $ **FLOATING
C7748 Vxm.n88 DGND 4.63fF $ **FLOATING
C7749 Vxm.n89 DGND 4.63fF $ **FLOATING
C7750 Vxm.n90 DGND 5.04fF $ **FLOATING
C7751 Vxm.t8 DGND 0.19fF
C7752 Vxm.t19 DGND 0.19fF
C7753 Vxm.t36 DGND 0.19fF
C7754 Vxm.t35 DGND 0.19fF
C7755 Vxm.n91 DGND 4.63fF $ **FLOATING
C7756 Vxm.n92 DGND 4.63fF $ **FLOATING
C7757 Vxm.n93 DGND 4.63fF $ **FLOATING
C7758 Vxm.n94 DGND 5.04fF $ **FLOATING
C7759 Vxm.t98 DGND 0.19fF
C7760 Vxm.t94 DGND 0.19fF
C7761 Vxm.t37 DGND 0.19fF
C7762 Vxm.t30 DGND 0.19fF
C7763 Vxm.t41 DGND 0.19fF
C7764 Vxm.n95 DGND 4.63fF $ **FLOATING
C7765 Vxm.n96 DGND 4.63fF $ **FLOATING
C7766 Vxm.n97 DGND 4.63fF $ **FLOATING
C7767 Vxm.n98 DGND 4.63fF $ **FLOATING
C7768 Vxm.n99 DGND 4.85fF $ **FLOATING
C7769 Vxm.t38 DGND 0.19fF
C7770 Vxm.t34 DGND 0.19fF
C7771 Vxm.t97 DGND 0.19fF
C7772 Vxm.t25 DGND 0.19fF
C7773 Vxm.t100 DGND 0.19fF
C7774 Vxm.n100 DGND 4.63fF $ **FLOATING
C7775 Vxm.n101 DGND 4.63fF $ **FLOATING
C7776 Vxm.n102 DGND 4.63fF $ **FLOATING
C7777 Vxm.n103 DGND 4.63fF $ **FLOATING
C7778 Vxm.n104 DGND 4.45fF $ **FLOATING
C7779 Vxm.n105 DGND 3.77fF $ **FLOATING
C7780 Vxm.n106 DGND 2.29fF $ **FLOATING
C7781 Vxm.n107 DGND 2.29fF $ **FLOATING
C7782 Vxm.n108 DGND 2.29fF $ **FLOATING
C7783 Vxm.n109 DGND 2.29fF $ **FLOATING
C7784 Vxm.n110 DGND 1.80fF $ **FLOATING
C7785 Vxm.n111 DGND 2.54fF $ **FLOATING
C7786 Vxm.n112 DGND 4.63fF $ **FLOATING
C7787 Vxm.n113 DGND 0.91fF $ **FLOATING
C7788 Vxm.n114 DGND 0.79fF $ **FLOATING
C7789 Vxm.n115 DGND 1.87fF $ **FLOATING
C7790 Vxm.n116 DGND 0.79fF $ **FLOATING
C7791 Vxm.n117 DGND 1.32fF $ **FLOATING
C7792 Vxm.n118 DGND 0.91fF $ **FLOATING
C7793 Vxm.n119 DGND 0.79fF $ **FLOATING
C7794 Vxm.n120 DGND 2.02fF $ **FLOATING
C7795 Vxm.n121 DGND 2.02fF $ **FLOATING
C7796 Vxm.n122 DGND 0.91fF $ **FLOATING
C7797 Vxm.n123 DGND 0.79fF $ **FLOATING
C7798 Vxm.n124 DGND 2.35fF $ **FLOATING
C7799 Vxm.n125 DGND 3.52fF $ **FLOATING
C7800 Vxm.n126 DGND 0.91fF $ **FLOATING
C7801 Vxm.n127 DGND 0.91fF $ **FLOATING
C7802 Vxm.n128 DGND 0.79fF $ **FLOATING
C7803 Vxm.n129 DGND 1.32fF $ **FLOATING
C7804 Vxm.n130 DGND 0.91fF $ **FLOATING
C7805 Vxm.n131 DGND 0.91fF $ **FLOATING
C7806 Vxm.n132 DGND 0.79fF $ **FLOATING
C7807 Vxm.n133 DGND 2.02fF $ **FLOATING
C7808 Vxm.n134 DGND 0.91fF $ **FLOATING
C7809 Vxm.n135 DGND 0.91fF $ **FLOATING
C7810 Vxm.n136 DGND 0.79fF $ **FLOATING
C7811 Vxm.n137 DGND 2.02fF $ **FLOATING
C7812 Vxm.n138 DGND 0.91fF $ **FLOATING
C7813 Vxm.n139 DGND 0.91fF $ **FLOATING
C7814 Vxm.n140 DGND 0.79fF $ **FLOATING
C7815 Vxm.n141 DGND 2.35fF $ **FLOATING
C7816 Vxm.n142 DGND 3.27fF $ **FLOATING
C7817 casc_n.n0 DGND 1.29fF $ **FLOATING
C7818 casc_n.t88 DGND 0.30fF
C7819 casc_n.t165 DGND 0.27fF
C7820 casc_n.n1 DGND 2.40fF $ **FLOATING
C7821 casc_n.t184 DGND 0.27fF
C7822 casc_n.n2 DGND 1.29fF $ **FLOATING
C7823 casc_n.t113 DGND 0.27fF
C7824 casc_n.n3 DGND 1.29fF $ **FLOATING
C7825 casc_n.t141 DGND 0.27fF
C7826 casc_n.n4 DGND 1.29fF $ **FLOATING
C7827 casc_n.t42 DGND 0.27fF
C7828 casc_n.n5 DGND 1.29fF $ **FLOATING
C7829 casc_n.t65 DGND 0.27fF
C7830 casc_n.n6 DGND 1.29fF $ **FLOATING
C7831 casc_n.t160 DGND 0.27fF
C7832 casc_n.n7 DGND 1.29fF $ **FLOATING
C7833 casc_n.t100 DGND 0.27fF
C7834 casc_n.n8 DGND 1.29fF $ **FLOATING
C7835 casc_n.t196 DGND 0.27fF
C7836 casc_n.n9 DGND 1.29fF $ **FLOATING
C7837 casc_n.t52 DGND 0.27fF
C7838 casc_n.n10 DGND 1.29fF $ **FLOATING
C7839 casc_n.t128 DGND 0.27fF
C7840 casc_n.n11 DGND 1.29fF $ **FLOATING
C7841 casc_n.t153 DGND 0.27fF
C7842 casc_n.n12 DGND 1.29fF $ **FLOATING
C7843 casc_n.t72 DGND 0.27fF
C7844 casc_n.n13 DGND 1.29fF $ **FLOATING
C7845 casc_n.t89 DGND 0.27fF
C7846 casc_n.n14 DGND 1.29fF $ **FLOATING
C7847 casc_n.t166 DGND 0.27fF
C7848 casc_n.n15 DGND 1.29fF $ **FLOATING
C7849 casc_n.t185 DGND 0.27fF
C7850 casc_n.n16 DGND 1.29fF $ **FLOATING
C7851 casc_n.t114 DGND 0.27fF
C7852 casc_n.n17 DGND 1.29fF $ **FLOATING
C7853 casc_n.t142 DGND 0.27fF
C7854 casc_n.n18 DGND 1.29fF $ **FLOATING
C7855 casc_n.t60 DGND 0.27fF
C7856 casc_n.n19 DGND 1.29fF $ **FLOATING
C7857 casc_n.t175 DGND 0.27fF
C7858 casc_n.n20 DGND 1.29fF $ **FLOATING
C7859 casc_n.t82 DGND 0.27fF
C7860 casc_n.n21 DGND 1.29fF $ **FLOATING
C7861 casc_n.t101 DGND 0.27fF
C7862 casc_n.n22 DGND 1.29fF $ **FLOATING
C7863 casc_n.t197 DGND 0.27fF
C7864 casc_n.n23 DGND 1.29fF $ **FLOATING
C7865 casc_n.t53 DGND 0.27fF
C7866 casc_n.n24 DGND 1.29fF $ **FLOATING
C7867 casc_n.t129 DGND 0.27fF
C7868 casc_n.n25 DGND 1.03fF $ **FLOATING
C7869 casc_n.n26 DGND 0.87fF $ **FLOATING
C7870 casc_n.n27 DGND 0.54fF $ **FLOATING
C7871 casc_n.t13 DGND 0.27fF
C7872 casc_n.n28 DGND 0.44fF $ **FLOATING
C7873 casc_n.n29 DGND 0.45fF $ **FLOATING
C7874 casc_n.n30 DGND 0.54fF $ **FLOATING
C7875 casc_n.t22 DGND 0.27fF
C7876 casc_n.n31 DGND 0.86fF $ **FLOATING
C7877 casc_n.n32 DGND 1.65fF $ **FLOATING
C7878 casc_n.n33 DGND 1.02fF $ **FLOATING
C7879 casc_n.t87 DGND 0.30fF
C7880 casc_n.t103 DGND 0.27fF
C7881 casc_n.n34 DGND 2.39fF $ **FLOATING
C7882 casc_n.t44 DGND 0.27fF
C7883 casc_n.n35 DGND 1.29fF $ **FLOATING
C7884 casc_n.t96 DGND 0.27fF
C7885 casc_n.n36 DGND 1.29fF $ **FLOATING
C7886 casc_n.t39 DGND 0.27fF
C7887 casc_n.n37 DGND 1.29fF $ **FLOATING
C7888 casc_n.t54 DGND 0.27fF
C7889 casc_n.n38 DGND 1.29fF $ **FLOATING
C7890 casc_n.t161 DGND 0.27fF
C7891 casc_n.n39 DGND 1.29fF $ **FLOATING
C7892 casc_n.t168 DGND 0.27fF
C7893 casc_n.n40 DGND 1.29fF $ **FLOATING
C7894 casc_n.t104 DGND 0.27fF
C7895 casc_n.n41 DGND 1.29fF $ **FLOATING
C7896 casc_n.t163 DGND 0.27fF
C7897 casc_n.n42 DGND 1.29fF $ **FLOATING
C7898 casc_n.t97 DGND 0.27fF
C7899 casc_n.n43 DGND 1.29fF $ **FLOATING
C7900 casc_n.t110 DGND 0.27fF
C7901 casc_n.n44 DGND 1.03fF $ **FLOATING
C7902 casc_n.n45 DGND 0.86fF $ **FLOATING
C7903 casc_n.n46 DGND 0.54fF $ **FLOATING
C7904 casc_n.t28 DGND 0.27fF
C7905 casc_n.n47 DGND 0.45fF $ **FLOATING
C7906 casc_n.n48 DGND 0.45fF $ **FLOATING
C7907 casc_n.n49 DGND 0.54fF $ **FLOATING
C7908 casc_n.t19 DGND 0.27fF
C7909 casc_n.n50 DGND 0.46fF $ **FLOATING
C7910 casc_n.t198 DGND 0.30fF
C7911 casc_n.t180 DGND 0.27fF
C7912 casc_n.n51 DGND 2.36fF $ **FLOATING
C7913 casc_n.t79 DGND 0.27fF
C7914 casc_n.n52 DGND 1.29fF $ **FLOATING
C7915 casc_n.t187 DGND 0.27fF
C7916 casc_n.n53 DGND 1.29fF $ **FLOATING
C7917 casc_n.t83 DGND 0.27fF
C7918 casc_n.n54 DGND 1.29fF $ **FLOATING
C7919 casc_n.t73 DGND 0.27fF
C7920 casc_n.n55 DGND 1.29fF $ **FLOATING
C7921 casc_n.t140 DGND 0.27fF
C7922 casc_n.n56 DGND 1.29fF $ **FLOATING
C7923 casc_n.t78 DGND 0.27fF
C7924 casc_n.n57 DGND 1.29fF $ **FLOATING
C7925 casc_n.t146 DGND 0.27fF
C7926 casc_n.n58 DGND 1.29fF $ **FLOATING
C7927 casc_n.t131 DGND 0.27fF
C7928 casc_n.n59 DGND 1.29fF $ **FLOATING
C7929 casc_n.t137 DGND 0.27fF
C7930 casc_n.n60 DGND 1.29fF $ **FLOATING
C7931 casc_n.t118 DGND 0.27fF
C7932 casc_n.n61 DGND 1.29fF $ **FLOATING
C7933 casc_n.t177 DGND 0.27fF
C7934 casc_n.n62 DGND 1.29fF $ **FLOATING
C7935 casc_n.t130 DGND 0.27fF
C7936 casc_n.n63 DGND 1.29fF $ **FLOATING
C7937 casc_n.t181 DGND 0.27fF
C7938 casc_n.n64 DGND 1.29fF $ **FLOATING
C7939 casc_n.t171 DGND 0.27fF
C7940 casc_n.n65 DGND 1.29fF $ **FLOATING
C7941 casc_n.t69 DGND 0.27fF
C7942 casc_n.n66 DGND 1.29fF $ **FLOATING
C7943 casc_n.t176 DGND 0.27fF
C7944 casc_n.n67 DGND 1.29fF $ **FLOATING
C7945 casc_n.t74 DGND 0.27fF
C7946 casc_n.n68 DGND 1.29fF $ **FLOATING
C7947 casc_n.t62 DGND 0.27fF
C7948 casc_n.n69 DGND 1.29fF $ **FLOATING
C7949 casc_n.t127 DGND 0.27fF
C7950 casc_n.n70 DGND 1.29fF $ **FLOATING
C7951 casc_n.t105 DGND 0.27fF
C7952 casc_n.n71 DGND 1.29fF $ **FLOATING
C7953 casc_n.t116 DGND 0.27fF
C7954 casc_n.n72 DGND 1.29fF $ **FLOATING
C7955 casc_n.t59 DGND 0.27fF
C7956 casc_n.n73 DGND 1.29fF $ **FLOATING
C7957 casc_n.t124 DGND 0.27fF
C7958 casc_n.n74 DGND 1.29fF $ **FLOATING
C7959 casc_n.t102 DGND 0.27fF
C7960 casc_n.n75 DGND 1.29fF $ **FLOATING
C7961 casc_n.t167 DGND 0.27fF
C7962 casc_n.n76 DGND 1.29fF $ **FLOATING
C7963 casc_n.t115 DGND 0.27fF
C7964 casc_n.n77 DGND 1.03fF $ **FLOATING
C7965 casc_n.n78 DGND 0.86fF $ **FLOATING
C7966 casc_n.n79 DGND 0.54fF $ **FLOATING
C7967 casc_n.t4 DGND 0.27fF
C7968 casc_n.n80 DGND 0.45fF $ **FLOATING
C7969 casc_n.n81 DGND 0.45fF $ **FLOATING
C7970 casc_n.n82 DGND 0.54fF $ **FLOATING
C7971 casc_n.t10 DGND 0.27fF
C7972 casc_n.n83 DGND 0.61fF $ **FLOATING
C7973 casc_n.n84 DGND 0.61fF $ **FLOATING
C7974 casc_n.n85 DGND 0.54fF $ **FLOATING
C7975 casc_n.t25 DGND 0.27fF
C7976 casc_n.n86 DGND 0.45fF $ **FLOATING
C7977 casc_n.n87 DGND 0.45fF $ **FLOATING
C7978 casc_n.n88 DGND 0.54fF $ **FLOATING
C7979 casc_n.t31 DGND 0.27fF
C7980 casc_n.n89 DGND 0.56fF $ **FLOATING
C7981 casc_n.n90 DGND 0.82fF $ **FLOATING
C7982 casc_n.t34 DGND 0.27fF
C7983 casc_n.t145 DGND 0.30fF
C7984 casc_n.t47 DGND 0.27fF
C7985 casc_n.n91 DGND 2.39fF $ **FLOATING
C7986 casc_n.t189 DGND 0.27fF
C7987 casc_n.n92 DGND 1.29fF $ **FLOATING
C7988 casc_n.t122 DGND 0.27fF
C7989 casc_n.n93 DGND 1.29fF $ **FLOATING
C7990 casc_n.t91 DGND 0.27fF
C7991 casc_n.n94 DGND 1.29fF $ **FLOATING
C7992 casc_n.t172 DGND 0.27fF
C7993 casc_n.n95 DGND 1.29fF $ **FLOATING
C7994 casc_n.t155 DGND 0.27fF
C7995 casc_n.n96 DGND 1.29fF $ **FLOATING
C7996 casc_n.t61 DGND 0.27fF
C7997 casc_n.n97 DGND 1.29fF $ **FLOATING
C7998 casc_n.t37 DGND 0.27fF
C7999 casc_n.n98 DGND 1.29fF $ **FLOATING
C8000 casc_n.t135 DGND 0.27fF
C8001 casc_n.n99 DGND 1.29fF $ **FLOATING
C8002 casc_n.t106 DGND 0.27fF
C8003 casc_n.n100 DGND 1.29fF $ **FLOATING
C8004 casc_n.t51 DGND 0.27fF
C8005 casc_n.n101 DGND 1.29fF $ **FLOATING
C8006 casc_n.t195 DGND 0.27fF
C8007 casc_n.n102 DGND 1.28fF $ **FLOATING
C8008 casc_n.t126 DGND 0.27fF
C8009 casc_n.n103 DGND 0.74fF $ **FLOATING
C8010 casc_n.n104 DGND 1.02fF $ **FLOATING
C8011 casc_n.t7 DGND 0.27fF
C8012 casc_n.n105 DGND 0.63fF $ **FLOATING
C8013 casc_n.t80 DGND 0.27fF
C8014 casc_n.n106 DGND 1.11fF $ **FLOATING
C8015 casc_n.t98 DGND 0.27fF
C8016 casc_n.n107 DGND 1.29fF $ **FLOATING
C8017 casc_n.t192 DGND 0.27fF
C8018 casc_n.n108 DGND 1.29fF $ **FLOATING
C8019 casc_n.t49 DGND 0.27fF
C8020 casc_n.n109 DGND 1.29fF $ **FLOATING
C8021 casc_n.t125 DGND 0.27fF
C8022 casc_n.n110 DGND 1.29fF $ **FLOATING
C8023 casc_n.t152 DGND 0.27fF
C8024 casc_n.n111 DGND 1.29fF $ **FLOATING
C8025 casc_n.t71 DGND 0.27fF
C8026 casc_n.n112 DGND 1.29fF $ **FLOATING
C8027 casc_n.t182 DGND 0.27fF
C8028 casc_n.n113 DGND 1.29fF $ **FLOATING
C8029 casc_n.t109 DGND 0.27fF
C8030 casc_n.n114 DGND 1.29fF $ **FLOATING
C8031 casc_n.t138 DGND 0.27fF
C8032 casc_n.n115 DGND 1.29fF $ **FLOATING
C8033 casc_n.t40 DGND 0.27fF
C8034 casc_n.n116 DGND 1.29fF $ **FLOATING
C8035 casc_n.t63 DGND 0.27fF
C8036 casc_n.n117 DGND 1.29fF $ **FLOATING
C8037 casc_n.t157 DGND 0.27fF
C8038 casc_n.n118 DGND 1.29fF $ **FLOATING
C8039 casc_n.t173 DGND 0.27fF
C8040 casc_n.n119 DGND 1.29fF $ **FLOATING
C8041 casc_n.t81 DGND 0.27fF
C8042 casc_n.n120 DGND 1.29fF $ **FLOATING
C8043 casc_n.t99 DGND 0.27fF
C8044 casc_n.n121 DGND 1.29fF $ **FLOATING
C8045 casc_n.t194 DGND 0.27fF
C8046 casc_n.n122 DGND 1.29fF $ **FLOATING
C8047 casc_n.t50 DGND 0.27fF
C8048 casc_n.n123 DGND 1.29fF $ **FLOATING
C8049 casc_n.t149 DGND 0.27fF
C8050 casc_n.n124 DGND 1.29fF $ **FLOATING
C8051 casc_n.t86 DGND 0.27fF
C8052 casc_n.n125 DGND 1.29fF $ **FLOATING
C8053 casc_n.t164 DGND 0.27fF
C8054 casc_n.n126 DGND 1.29fF $ **FLOATING
C8055 casc_n.t183 DGND 0.27fF
C8056 casc_n.n127 DGND 1.29fF $ **FLOATING
C8057 casc_n.t112 DGND 0.27fF
C8058 casc_n.n128 DGND 1.29fF $ **FLOATING
C8059 casc_n.t139 DGND 0.27fF
C8060 casc_n.n129 DGND 1.29fF $ **FLOATING
C8061 casc_n.t41 DGND 0.27fF
C8062 casc_n.n130 DGND 1.29fF $ **FLOATING
C8063 casc_n.t64 DGND 0.27fF
C8064 casc_n.n131 DGND 1.29fF $ **FLOATING
C8065 casc_n.t159 DGND 0.27fF
C8066 casc_n.n132 DGND 1.29fF $ **FLOATING
C8067 casc_n.t174 DGND 0.27fF
C8068 casc_n.n133 DGND 1.29fF $ **FLOATING
C8069 casc_n.t95 DGND 0.27fF
C8070 casc_n.n134 DGND 0.95fF $ **FLOATING
C8071 casc_n.t66 DGND 0.30fF
C8072 casc_n.t144 DGND 0.27fF
C8073 casc_n.n135 DGND 2.39fF $ **FLOATING
C8074 casc_n.t117 DGND 0.27fF
C8075 casc_n.n136 DGND 1.29fF $ **FLOATING
C8076 casc_n.t43 DGND 0.27fF
C8077 casc_n.n137 DGND 1.29fF $ **FLOATING
C8078 casc_n.t186 DGND 0.27fF
C8079 casc_n.n138 DGND 1.29fF $ **FLOATING
C8080 casc_n.t90 DGND 0.27fF
C8081 casc_n.n139 DGND 1.29fF $ **FLOATING
C8082 casc_n.t75 DGND 0.27fF
C8083 casc_n.n140 DGND 1.29fF $ **FLOATING
C8084 casc_n.t154 DGND 0.27fF
C8085 casc_n.n141 DGND 1.29fF $ **FLOATING
C8086 casc_n.t132 DGND 0.27fF
C8087 casc_n.n142 DGND 1.29fF $ **FLOATING
C8088 casc_n.t55 DGND 0.27fF
C8089 casc_n.n143 DGND 1.29fF $ **FLOATING
C8090 casc_n.t199 DGND 0.27fF
C8091 casc_n.n144 DGND 1.29fF $ **FLOATING
C8092 casc_n.t150 DGND 0.27fF
C8093 casc_n.n145 DGND 1.29fF $ **FLOATING
C8094 casc_n.t121 DGND 0.27fF
C8095 casc_n.n146 DGND 1.28fF $ **FLOATING
C8096 casc_n.t46 DGND 0.27fF
C8097 casc_n.n147 DGND 0.74fF $ **FLOATING
C8098 casc_n.t92 DGND 0.30fF
C8099 casc_n.t169 DGND 0.27fF
C8100 casc_n.n148 DGND 2.40fF $ **FLOATING
C8101 casc_n.t191 DGND 0.27fF
C8102 casc_n.n149 DGND 1.29fF $ **FLOATING
C8103 casc_n.t119 DGND 0.27fF
C8104 casc_n.n150 DGND 1.29fF $ **FLOATING
C8105 casc_n.t147 DGND 0.27fF
C8106 casc_n.n151 DGND 1.29fF $ **FLOATING
C8107 casc_n.t45 DGND 0.27fF
C8108 casc_n.n152 DGND 1.29fF $ **FLOATING
C8109 casc_n.t70 DGND 0.27fF
C8110 casc_n.n153 DGND 1.29fF $ **FLOATING
C8111 casc_n.t162 DGND 0.27fF
C8112 casc_n.n154 DGND 1.29fF $ **FLOATING
C8113 casc_n.t108 DGND 0.27fF
C8114 casc_n.n155 DGND 1.29fF $ **FLOATING
C8115 casc_n.t200 DGND 0.27fF
C8116 casc_n.n156 DGND 1.29fF $ **FLOATING
C8117 casc_n.t57 DGND 0.27fF
C8118 casc_n.n157 DGND 1.29fF $ **FLOATING
C8119 casc_n.t133 DGND 0.27fF
C8120 casc_n.n158 DGND 1.29fF $ **FLOATING
C8121 casc_n.t156 DGND 0.27fF
C8122 casc_n.n159 DGND 1.29fF $ **FLOATING
C8123 casc_n.t76 DGND 0.27fF
C8124 casc_n.n160 DGND 1.29fF $ **FLOATING
C8125 casc_n.t93 DGND 0.27fF
C8126 casc_n.n161 DGND 1.29fF $ **FLOATING
C8127 casc_n.t170 DGND 0.27fF
C8128 casc_n.n162 DGND 1.29fF $ **FLOATING
C8129 casc_n.t193 DGND 0.27fF
C8130 casc_n.n163 DGND 1.29fF $ **FLOATING
C8131 casc_n.t120 DGND 0.27fF
C8132 casc_n.n164 DGND 1.29fF $ **FLOATING
C8133 casc_n.t148 DGND 0.27fF
C8134 casc_n.n165 DGND 1.29fF $ **FLOATING
C8135 casc_n.t67 DGND 0.27fF
C8136 casc_n.n166 DGND 1.29fF $ **FLOATING
C8137 casc_n.t179 DGND 0.27fF
C8138 casc_n.n167 DGND 1.29fF $ **FLOATING
C8139 casc_n.t84 DGND 0.27fF
C8140 casc_n.n168 DGND 1.29fF $ **FLOATING
C8141 casc_n.t111 DGND 0.27fF
C8142 casc_n.n169 DGND 1.29fF $ **FLOATING
C8143 casc_n.t201 DGND 0.27fF
C8144 casc_n.n170 DGND 1.29fF $ **FLOATING
C8145 casc_n.t58 DGND 0.27fF
C8146 casc_n.n171 DGND 1.29fF $ **FLOATING
C8147 casc_n.t134 DGND 0.27fF
C8148 casc_n.n172 DGND 1.29fF $ **FLOATING
C8149 casc_n.t158 DGND 0.27fF
C8150 casc_n.n173 DGND 1.29fF $ **FLOATING
C8151 casc_n.t77 DGND 0.27fF
C8152 casc_n.n174 DGND 1.29fF $ **FLOATING
C8153 casc_n.t94 DGND 0.27fF
C8154 casc_n.n175 DGND 1.29fF $ **FLOATING
C8155 casc_n.t188 DGND 0.27fF
C8156 casc_n.n176 DGND 0.95fF $ **FLOATING
C8157 casc_n.n177 DGND 1.60fF $ **FLOATING
C8158 casc_n.n178 DGND 2.15fF $ **FLOATING
C8159 casc_n.t16 DGND 0.27fF
C8160 casc_n.t56 DGND 0.30fF
C8161 casc_n.t136 DGND 0.27fF
C8162 casc_n.n179 DGND 2.39fF $ **FLOATING
C8163 casc_n.t107 DGND 0.27fF
C8164 casc_n.n180 DGND 1.29fF $ **FLOATING
C8165 casc_n.t38 DGND 0.27fF
C8166 casc_n.n181 DGND 1.29fF $ **FLOATING
C8167 casc_n.t178 DGND 0.27fF
C8168 casc_n.n182 DGND 1.29fF $ **FLOATING
C8169 casc_n.t85 DGND 0.27fF
C8170 casc_n.n183 DGND 1.29fF $ **FLOATING
C8171 casc_n.t68 DGND 0.27fF
C8172 casc_n.n184 DGND 1.29fF $ **FLOATING
C8173 casc_n.t151 DGND 0.27fF
C8174 casc_n.n185 DGND 1.29fF $ **FLOATING
C8175 casc_n.t123 DGND 0.27fF
C8176 casc_n.n186 DGND 1.29fF $ **FLOATING
C8177 casc_n.t48 DGND 0.27fF
C8178 casc_n.n187 DGND 1.29fF $ **FLOATING
C8179 casc_n.t190 DGND 0.27fF
C8180 casc_n.n188 DGND 1.29fF $ **FLOATING
C8181 casc_n.t143 DGND 0.27fF
C8182 casc_n.n189 DGND 1.03fF $ **FLOATING
C8183 casc_n.n190 DGND 0.86fF $ **FLOATING
C8184 casc_n.n191 DGND 0.54fF $ **FLOATING
C8185 casc_n.n192 DGND 0.46fF $ **FLOATING
C8186 casc_n.n193 DGND 0.44fF $ **FLOATING
C8187 casc_n.n194 DGND 0.53fF $ **FLOATING
C8188 casc_n.n195 DGND 0.11fF $ **FLOATING
C8189 casc_n.n196 DGND 1.07fF $ **FLOATING
.ends

