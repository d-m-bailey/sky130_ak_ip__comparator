magic
tech sky130A
magscale 1 2
timestamp 1713228438
<< nwell >>
rect -1516 -815 1516 815
<< mvpmos >>
rect -1258 118 -458 518
rect -400 118 400 518
rect 458 118 1258 518
rect -1258 -518 -458 -118
rect -400 -518 400 -118
rect 458 -518 1258 -118
<< mvpdiff >>
rect -1316 506 -1258 518
rect -1316 130 -1304 506
rect -1270 130 -1258 506
rect -1316 118 -1258 130
rect -458 506 -400 518
rect -458 130 -446 506
rect -412 130 -400 506
rect -458 118 -400 130
rect 400 506 458 518
rect 400 130 412 506
rect 446 130 458 506
rect 400 118 458 130
rect 1258 506 1316 518
rect 1258 130 1270 506
rect 1304 130 1316 506
rect 1258 118 1316 130
rect -1316 -130 -1258 -118
rect -1316 -506 -1304 -130
rect -1270 -506 -1258 -130
rect -1316 -518 -1258 -506
rect -458 -130 -400 -118
rect -458 -506 -446 -130
rect -412 -506 -400 -130
rect -458 -518 -400 -506
rect 400 -130 458 -118
rect 400 -506 412 -130
rect 446 -506 458 -130
rect 400 -518 458 -506
rect 1258 -130 1316 -118
rect 1258 -506 1270 -130
rect 1304 -506 1316 -130
rect 1258 -518 1316 -506
<< mvpdiffc >>
rect -1304 130 -1270 506
rect -446 130 -412 506
rect 412 130 446 506
rect 1270 130 1304 506
rect -1304 -506 -1270 -130
rect -446 -506 -412 -130
rect 412 -506 446 -130
rect 1270 -506 1304 -130
<< mvnsubdiff >>
rect -1450 737 1450 749
rect -1450 703 -1342 737
rect 1342 703 1450 737
rect -1450 691 1450 703
rect -1450 641 -1392 691
rect -1450 -641 -1438 641
rect -1404 -641 -1392 641
rect 1392 641 1450 691
rect -1450 -691 -1392 -641
rect 1392 -641 1404 641
rect 1438 -641 1450 641
rect 1392 -691 1450 -641
rect -1450 -703 1450 -691
rect -1450 -737 -1342 -703
rect 1342 -737 1450 -703
rect -1450 -749 1450 -737
<< mvnsubdiffcont >>
rect -1342 703 1342 737
rect -1438 -641 -1404 641
rect 1404 -641 1438 641
rect -1342 -737 1342 -703
<< poly >>
rect -1258 599 -458 615
rect -1258 565 -1242 599
rect -474 565 -458 599
rect -1258 518 -458 565
rect -400 599 400 615
rect -400 565 -384 599
rect 384 565 400 599
rect -400 518 400 565
rect 458 599 1258 615
rect 458 565 474 599
rect 1242 565 1258 599
rect 458 518 1258 565
rect -1258 71 -458 118
rect -1258 37 -1242 71
rect -474 37 -458 71
rect -1258 21 -458 37
rect -400 71 400 118
rect -400 37 -384 71
rect 384 37 400 71
rect -400 21 400 37
rect 458 71 1258 118
rect 458 37 474 71
rect 1242 37 1258 71
rect 458 21 1258 37
rect -1258 -37 -458 -21
rect -1258 -71 -1242 -37
rect -474 -71 -458 -37
rect -1258 -118 -458 -71
rect -400 -37 400 -21
rect -400 -71 -384 -37
rect 384 -71 400 -37
rect -400 -118 400 -71
rect 458 -37 1258 -21
rect 458 -71 474 -37
rect 1242 -71 1258 -37
rect 458 -118 1258 -71
rect -1258 -565 -458 -518
rect -1258 -599 -1242 -565
rect -474 -599 -458 -565
rect -1258 -615 -458 -599
rect -400 -565 400 -518
rect -400 -599 -384 -565
rect 384 -599 400 -565
rect -400 -615 400 -599
rect 458 -565 1258 -518
rect 458 -599 474 -565
rect 1242 -599 1258 -565
rect 458 -615 1258 -599
<< polycont >>
rect -1242 565 -474 599
rect -384 565 384 599
rect 474 565 1242 599
rect -1242 37 -474 71
rect -384 37 384 71
rect 474 37 1242 71
rect -1242 -71 -474 -37
rect -384 -71 384 -37
rect 474 -71 1242 -37
rect -1242 -599 -474 -565
rect -384 -599 384 -565
rect 474 -599 1242 -565
<< locali >>
rect -1438 703 -1342 737
rect 1342 703 1438 737
rect -1438 641 -1404 703
rect 1404 641 1438 703
rect -1258 565 -1242 599
rect -474 565 -458 599
rect -400 565 -384 599
rect 384 565 400 599
rect 458 565 474 599
rect 1242 565 1258 599
rect -1304 506 -1270 522
rect -1304 114 -1270 130
rect -446 506 -412 522
rect -446 114 -412 130
rect 412 506 446 522
rect 412 114 446 130
rect 1270 506 1304 522
rect 1270 114 1304 130
rect -1258 37 -1242 71
rect -474 37 -458 71
rect -400 37 -384 71
rect 384 37 400 71
rect 458 37 474 71
rect 1242 37 1258 71
rect -1258 -71 -1242 -37
rect -474 -71 -458 -37
rect -400 -71 -384 -37
rect 384 -71 400 -37
rect 458 -71 474 -37
rect 1242 -71 1258 -37
rect -1304 -130 -1270 -114
rect -1304 -522 -1270 -506
rect -446 -130 -412 -114
rect -446 -522 -412 -506
rect 412 -130 446 -114
rect 412 -522 446 -506
rect 1270 -130 1304 -114
rect 1270 -522 1304 -506
rect -1258 -599 -1242 -565
rect -474 -599 -458 -565
rect -400 -599 -384 -565
rect 384 -599 400 -565
rect 458 -599 474 -565
rect 1242 -599 1258 -565
rect -1438 -703 -1404 -641
rect 1404 -703 1438 -641
rect -1438 -737 -1342 -703
rect 1342 -737 1438 -703
<< viali >>
rect -1123 703 1123 737
rect -1242 565 -474 599
rect -384 565 384 599
rect 474 565 1242 599
rect -1438 -562 -1404 562
rect -1304 130 -1270 506
rect -446 130 -412 506
rect 412 130 446 506
rect 1270 130 1304 506
rect -1242 37 -474 71
rect -384 37 384 71
rect 474 37 1242 71
rect -1242 -71 -474 -37
rect -384 -71 384 -37
rect 474 -71 1242 -37
rect -1304 -506 -1270 -130
rect -446 -506 -412 -130
rect 412 -506 446 -130
rect 1270 -506 1304 -130
rect 1404 -562 1438 562
rect -1242 -599 -474 -565
rect -384 -599 384 -565
rect 474 -599 1242 -565
rect -1123 -737 1123 -703
<< metal1 >>
rect -1135 737 1135 743
rect -1135 703 -1123 737
rect 1123 703 1135 737
rect -1135 697 1135 703
rect -1254 599 -462 605
rect -1444 562 -1398 574
rect -1444 -562 -1438 562
rect -1404 -562 -1398 562
rect -1254 565 -1242 599
rect -474 565 -462 599
rect -1254 559 -462 565
rect -396 599 396 605
rect -396 565 -384 599
rect 384 565 396 599
rect -396 559 396 565
rect 462 599 1254 605
rect 462 565 474 599
rect 1242 565 1254 599
rect 462 559 1254 565
rect 1398 562 1444 574
rect -1310 506 -1264 518
rect -1310 130 -1304 506
rect -1270 130 -1264 506
rect -1310 118 -1264 130
rect -452 506 -406 518
rect -452 130 -446 506
rect -412 130 -406 506
rect -452 118 -406 130
rect 406 506 452 518
rect 406 130 412 506
rect 446 130 452 506
rect 406 118 452 130
rect 1264 506 1310 518
rect 1264 130 1270 506
rect 1304 130 1310 506
rect 1264 118 1310 130
rect -1254 71 -462 77
rect -1254 37 -1242 71
rect -474 37 -462 71
rect -1254 31 -462 37
rect -396 71 396 77
rect -396 37 -384 71
rect 384 37 396 71
rect -396 31 396 37
rect 462 71 1254 77
rect 462 37 474 71
rect 1242 37 1254 71
rect 462 31 1254 37
rect -1254 -37 -462 -31
rect -1254 -71 -1242 -37
rect -474 -71 -462 -37
rect -1254 -77 -462 -71
rect -396 -37 396 -31
rect -396 -71 -384 -37
rect 384 -71 396 -37
rect -396 -77 396 -71
rect 462 -37 1254 -31
rect 462 -71 474 -37
rect 1242 -71 1254 -37
rect 462 -77 1254 -71
rect -1310 -130 -1264 -118
rect -1310 -506 -1304 -130
rect -1270 -506 -1264 -130
rect -1310 -518 -1264 -506
rect -452 -130 -406 -118
rect -452 -506 -446 -130
rect -412 -506 -406 -130
rect -452 -518 -406 -506
rect 406 -130 452 -118
rect 406 -506 412 -130
rect 446 -506 452 -130
rect 406 -518 452 -506
rect 1264 -130 1310 -118
rect 1264 -506 1270 -130
rect 1304 -506 1310 -130
rect 1264 -518 1310 -506
rect -1444 -574 -1398 -562
rect -1254 -565 -462 -559
rect -1254 -599 -1242 -565
rect -474 -599 -462 -565
rect -1254 -605 -462 -599
rect -396 -565 396 -559
rect -396 -599 -384 -565
rect 384 -599 396 -565
rect -396 -605 396 -599
rect 462 -565 1254 -559
rect 462 -599 474 -565
rect 1242 -599 1254 -565
rect 1398 -562 1404 562
rect 1438 -562 1444 562
rect 1398 -574 1444 -562
rect 462 -605 1254 -599
rect -1135 -703 1135 -697
rect -1135 -737 -1123 -703
rect 1123 -737 1135 -703
rect -1135 -743 1135 -737
<< properties >>
string FIXED_BBOX -1421 -720 1421 720
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 2 l 4 m 2 nf 3 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 80 viagr 80 viagl 80 viagt 80
<< end >>
