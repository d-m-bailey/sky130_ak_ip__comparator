magic
tech sky130A
magscale 1 2
timestamp 1713585847
<< error_p >>
rect -111 145 -47 151
rect 47 145 111 151
rect -111 111 -99 145
rect 47 111 59 145
rect -111 105 -47 111
rect 47 105 111 111
<< nwell >>
rect -387 -362 387 362
<< mvpmos >>
rect -129 -136 -29 64
rect 29 -136 129 64
<< mvpdiff >>
rect -187 52 -129 64
rect -187 -124 -175 52
rect -141 -124 -129 52
rect -187 -136 -129 -124
rect -29 52 29 64
rect -29 -124 -17 52
rect 17 -124 29 52
rect -29 -136 29 -124
rect 129 52 187 64
rect 129 -124 141 52
rect 175 -124 187 52
rect 129 -136 187 -124
<< mvpdiffc >>
rect -175 -124 -141 52
rect -17 -124 17 52
rect 141 -124 175 52
<< mvnsubdiff >>
rect -321 284 321 296
rect -321 250 -213 284
rect 213 250 321 284
rect -321 238 321 250
rect -321 188 -263 238
rect -321 -188 -309 188
rect -275 -188 -263 188
rect 263 188 321 238
rect -321 -238 -263 -188
rect 263 -188 275 188
rect 309 -188 321 188
rect 263 -238 321 -188
rect -321 -250 321 -238
rect -321 -284 -213 -250
rect 213 -284 321 -250
rect -321 -296 321 -284
<< mvnsubdiffcont >>
rect -213 250 213 284
rect -309 -188 -275 188
rect 275 -188 309 188
rect -213 -284 213 -250
<< poly >>
rect -129 145 -29 161
rect -129 111 -113 145
rect -45 111 -29 145
rect -129 64 -29 111
rect 29 145 129 161
rect 29 111 45 145
rect 113 111 129 145
rect 29 64 129 111
rect -129 -162 -29 -136
rect 29 -162 129 -136
<< polycont >>
rect -113 111 -45 145
rect 45 111 113 145
<< locali >>
rect -309 250 -213 284
rect 213 250 309 284
rect -309 200 -275 250
rect 275 200 309 250
rect -129 111 -113 145
rect -45 111 -29 145
rect 29 111 45 145
rect 113 111 129 145
rect -175 52 -141 68
rect -175 -140 -141 -124
rect -17 52 17 68
rect -17 -140 17 -124
rect 141 52 175 68
rect 141 -140 175 -124
rect -309 -250 -275 -200
rect 275 -250 309 -200
rect -309 -284 -220 -250
rect 220 -284 309 -250
<< viali >>
rect -309 188 -275 200
rect -309 -188 -275 188
rect 275 188 309 200
rect -99 111 -59 145
rect 59 111 99 145
rect -175 -124 -141 52
rect -17 -124 17 52
rect 141 -124 175 52
rect -309 -200 -275 -188
rect 275 -188 309 188
rect 275 -200 309 -188
rect -220 -284 -213 -250
rect -213 -284 213 -250
rect 213 -284 220 -250
<< metal1 >>
rect -315 200 -269 212
rect -315 -200 -309 200
rect -275 -200 -269 200
rect 269 200 315 212
rect -111 145 -47 151
rect -111 111 -99 145
rect -59 111 -47 145
rect -111 105 -47 111
rect 47 145 111 151
rect 47 111 59 145
rect 99 111 111 145
rect 47 105 111 111
rect -181 52 -135 64
rect -181 -124 -175 52
rect -141 -124 -135 52
rect -181 -136 -135 -124
rect -23 52 23 64
rect -23 -124 -17 52
rect 17 -124 23 52
rect -23 -136 23 -124
rect 135 52 181 64
rect 135 -124 141 52
rect 175 -124 181 52
rect 135 -136 181 -124
rect -315 -212 -269 -200
rect 269 -200 275 200
rect 309 -200 315 200
rect 269 -212 315 -200
rect -232 -250 232 -244
rect -232 -284 -220 -250
rect 220 -284 232 -250
rect -232 -290 232 -284
<< properties >>
string FIXED_BBOX -292 -267 292 267
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 1 l 0.50 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 60 viagb 80 viagr 80 viagl 80 viagt 0
<< end >>
