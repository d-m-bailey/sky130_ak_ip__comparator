magic
tech sky130A
magscale 1 2
timestamp 1713548572
<< error_p >>
rect -266 281 -208 287
rect -108 281 -50 287
rect 50 281 108 287
rect 208 281 266 287
rect -266 247 -254 281
rect -108 247 -96 281
rect 50 247 62 281
rect 208 247 220 281
rect -266 241 -208 247
rect -108 241 -50 247
rect 50 241 108 247
rect 208 241 266 247
rect -266 -247 -208 -241
rect -108 -247 -50 -241
rect 50 -247 108 -241
rect 208 -247 266 -241
rect -266 -281 -254 -247
rect -108 -281 -96 -247
rect 50 -281 62 -247
rect 208 -281 220 -247
rect -266 -287 -208 -281
rect -108 -287 -50 -281
rect 50 -287 108 -281
rect 208 -287 266 -281
<< nwell >>
rect -545 -497 545 497
<< mvpmos >>
rect -287 -200 -187 200
rect -129 -200 -29 200
rect 29 -200 129 200
rect 187 -200 287 200
<< mvpdiff >>
rect -345 188 -287 200
rect -345 -188 -333 188
rect -299 -188 -287 188
rect -345 -200 -287 -188
rect -187 188 -129 200
rect -187 -188 -175 188
rect -141 -188 -129 188
rect -187 -200 -129 -188
rect -29 188 29 200
rect -29 -188 -17 188
rect 17 -188 29 188
rect -29 -200 29 -188
rect 129 188 187 200
rect 129 -188 141 188
rect 175 -188 187 188
rect 129 -200 187 -188
rect 287 188 345 200
rect 287 -188 299 188
rect 333 -188 345 188
rect 287 -200 345 -188
<< mvpdiffc >>
rect -333 -188 -299 188
rect -175 -188 -141 188
rect -17 -188 17 188
rect 141 -188 175 188
rect 299 -188 333 188
<< mvnsubdiff >>
rect -479 419 479 431
rect -479 385 -371 419
rect 371 385 479 419
rect -479 373 479 385
rect -479 323 -421 373
rect -479 -323 -467 323
rect -433 -323 -421 323
rect 421 323 479 373
rect -479 -373 -421 -323
rect 421 -323 433 323
rect 467 -323 479 323
rect 421 -373 479 -323
rect -479 -385 479 -373
rect -479 -419 -371 -385
rect 371 -419 479 -385
rect -479 -431 479 -419
<< mvnsubdiffcont >>
rect -371 385 371 419
rect -467 -323 -433 323
rect 433 -323 467 323
rect -371 -419 371 -385
<< poly >>
rect -287 281 -187 297
rect -287 247 -271 281
rect -203 247 -187 281
rect -287 200 -187 247
rect -129 281 -29 297
rect -129 247 -113 281
rect -45 247 -29 281
rect -129 200 -29 247
rect 29 281 129 297
rect 29 247 45 281
rect 113 247 129 281
rect 29 200 129 247
rect 187 281 287 297
rect 187 247 203 281
rect 271 247 287 281
rect 187 200 287 247
rect -287 -247 -187 -200
rect -287 -281 -271 -247
rect -203 -281 -187 -247
rect -287 -297 -187 -281
rect -129 -247 -29 -200
rect -129 -281 -113 -247
rect -45 -281 -29 -247
rect -129 -297 -29 -281
rect 29 -247 129 -200
rect 29 -281 45 -247
rect 113 -281 129 -247
rect 29 -297 129 -281
rect 187 -247 287 -200
rect 187 -281 203 -247
rect 271 -281 287 -247
rect 187 -297 287 -281
<< polycont >>
rect -271 247 -203 281
rect -113 247 -45 281
rect 45 247 113 281
rect 203 247 271 281
rect -271 -281 -203 -247
rect -113 -281 -45 -247
rect 45 -281 113 -247
rect 203 -281 271 -247
<< locali >>
rect -467 385 -371 419
rect 371 385 467 419
rect -467 323 -433 385
rect 433 323 467 385
rect -287 247 -271 281
rect -203 247 -187 281
rect -129 247 -113 281
rect -45 247 -29 281
rect 29 247 45 281
rect 113 247 129 281
rect 187 247 203 281
rect 271 247 287 281
rect -333 188 -299 204
rect -333 -204 -299 -188
rect -175 188 -141 204
rect -175 -204 -141 -188
rect -17 188 17 204
rect -17 -204 17 -188
rect 141 188 175 204
rect 141 -204 175 -188
rect 299 188 333 204
rect 299 -204 333 -188
rect -287 -281 -271 -247
rect -203 -281 -187 -247
rect -129 -281 -113 -247
rect -45 -281 -29 -247
rect 29 -281 45 -247
rect 113 -281 129 -247
rect 187 -281 203 -247
rect 271 -281 287 -247
rect -467 -385 -433 -323
rect 433 -385 467 -323
rect -467 -419 -371 -385
rect 371 -419 467 -385
<< viali >>
rect -467 -308 -433 308
rect -254 247 -220 281
rect -96 247 -62 281
rect 62 247 96 281
rect 220 247 254 281
rect -333 -188 -299 188
rect -175 -188 -141 188
rect -17 -188 17 188
rect 141 -188 175 188
rect 299 -188 333 188
rect -254 -281 -220 -247
rect -96 -281 -62 -247
rect 62 -281 96 -247
rect 220 -281 254 -247
rect 433 -308 467 308
rect -346 -419 346 -385
<< metal1 >>
rect -473 308 -427 320
rect -473 -308 -467 308
rect -433 -308 -427 308
rect 427 308 473 320
rect -266 281 -208 287
rect -266 247 -254 281
rect -220 247 -208 281
rect -266 241 -208 247
rect -108 281 -50 287
rect -108 247 -96 281
rect -62 247 -50 281
rect -108 241 -50 247
rect 50 281 108 287
rect 50 247 62 281
rect 96 247 108 281
rect 50 241 108 247
rect 208 281 266 287
rect 208 247 220 281
rect 254 247 266 281
rect 208 241 266 247
rect -339 188 -293 200
rect -339 -188 -333 188
rect -299 -188 -293 188
rect -339 -200 -293 -188
rect -181 188 -135 200
rect -181 -188 -175 188
rect -141 -188 -135 188
rect -181 -200 -135 -188
rect -23 188 23 200
rect -23 -188 -17 188
rect 17 -188 23 188
rect -23 -200 23 -188
rect 135 188 181 200
rect 135 -188 141 188
rect 175 -188 181 188
rect 135 -200 181 -188
rect 293 188 339 200
rect 293 -188 299 188
rect 333 -188 339 188
rect 293 -200 339 -188
rect -266 -247 -208 -241
rect -266 -281 -254 -247
rect -220 -281 -208 -247
rect -266 -287 -208 -281
rect -108 -247 -50 -241
rect -108 -281 -96 -247
rect -62 -281 -50 -247
rect -108 -287 -50 -281
rect 50 -247 108 -241
rect 50 -281 62 -247
rect 96 -281 108 -247
rect 50 -287 108 -281
rect 208 -247 266 -241
rect 208 -281 220 -247
rect 254 -281 266 -247
rect 208 -287 266 -281
rect -473 -320 -427 -308
rect 427 -308 433 308
rect 467 -308 473 308
rect 427 -320 473 -308
rect -358 -385 358 -379
rect -358 -419 -346 -385
rect 346 -419 358 -385
rect -358 -425 358 -419
<< properties >>
string FIXED_BBOX -450 -402 450 402
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 2 l 0.5 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 80 viagr 80 viagl 80 viagt 0
<< end >>
