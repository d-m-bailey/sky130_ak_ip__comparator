magic
tech sky130A
magscale 1 2
timestamp 1713548572
<< nwell >>
rect -1261 -697 1261 697
<< mvpmos >>
rect -1003 -400 -803 400
rect -745 -400 -545 400
rect -487 -400 -287 400
rect -229 -400 -29 400
rect 29 -400 229 400
rect 287 -400 487 400
rect 545 -400 745 400
rect 803 -400 1003 400
<< mvpdiff >>
rect -1061 388 -1003 400
rect -1061 -388 -1049 388
rect -1015 -388 -1003 388
rect -1061 -400 -1003 -388
rect -803 388 -745 400
rect -803 -388 -791 388
rect -757 -388 -745 388
rect -803 -400 -745 -388
rect -545 388 -487 400
rect -545 -388 -533 388
rect -499 -388 -487 388
rect -545 -400 -487 -388
rect -287 388 -229 400
rect -287 -388 -275 388
rect -241 -388 -229 388
rect -287 -400 -229 -388
rect -29 388 29 400
rect -29 -388 -17 388
rect 17 -388 29 388
rect -29 -400 29 -388
rect 229 388 287 400
rect 229 -388 241 388
rect 275 -388 287 388
rect 229 -400 287 -388
rect 487 388 545 400
rect 487 -388 499 388
rect 533 -388 545 388
rect 487 -400 545 -388
rect 745 388 803 400
rect 745 -388 757 388
rect 791 -388 803 388
rect 745 -400 803 -388
rect 1003 388 1061 400
rect 1003 -388 1015 388
rect 1049 -388 1061 388
rect 1003 -400 1061 -388
<< mvpdiffc >>
rect -1049 -388 -1015 388
rect -791 -388 -757 388
rect -533 -388 -499 388
rect -275 -388 -241 388
rect -17 -388 17 388
rect 241 -388 275 388
rect 499 -388 533 388
rect 757 -388 791 388
rect 1015 -388 1049 388
<< mvnsubdiff >>
rect -1195 619 1195 631
rect -1195 585 -1087 619
rect 1087 585 1195 619
rect -1195 573 1195 585
rect -1195 523 -1137 573
rect -1195 -523 -1183 523
rect -1149 -523 -1137 523
rect 1137 523 1195 573
rect -1195 -573 -1137 -523
rect 1137 -523 1149 523
rect 1183 -523 1195 523
rect 1137 -573 1195 -523
rect -1195 -585 1195 -573
rect -1195 -619 -1087 -585
rect 1087 -619 1195 -585
rect -1195 -631 1195 -619
<< mvnsubdiffcont >>
rect -1087 585 1087 619
rect -1183 -523 -1149 523
rect 1149 -523 1183 523
rect -1087 -619 1087 -585
<< poly >>
rect -1003 481 -803 497
rect -1003 447 -987 481
rect -819 447 -803 481
rect -1003 400 -803 447
rect -745 481 -545 497
rect -745 447 -729 481
rect -561 447 -545 481
rect -745 400 -545 447
rect -487 481 -287 497
rect -487 447 -471 481
rect -303 447 -287 481
rect -487 400 -287 447
rect -229 481 -29 497
rect -229 447 -213 481
rect -45 447 -29 481
rect -229 400 -29 447
rect 29 481 229 497
rect 29 447 45 481
rect 213 447 229 481
rect 29 400 229 447
rect 287 481 487 497
rect 287 447 303 481
rect 471 447 487 481
rect 287 400 487 447
rect 545 481 745 497
rect 545 447 561 481
rect 729 447 745 481
rect 545 400 745 447
rect 803 481 1003 497
rect 803 447 819 481
rect 987 447 1003 481
rect 803 400 1003 447
rect -1003 -447 -803 -400
rect -1003 -481 -987 -447
rect -819 -481 -803 -447
rect -1003 -497 -803 -481
rect -745 -447 -545 -400
rect -745 -481 -729 -447
rect -561 -481 -545 -447
rect -745 -497 -545 -481
rect -487 -447 -287 -400
rect -487 -481 -471 -447
rect -303 -481 -287 -447
rect -487 -497 -287 -481
rect -229 -447 -29 -400
rect -229 -481 -213 -447
rect -45 -481 -29 -447
rect -229 -497 -29 -481
rect 29 -447 229 -400
rect 29 -481 45 -447
rect 213 -481 229 -447
rect 29 -497 229 -481
rect 287 -447 487 -400
rect 287 -481 303 -447
rect 471 -481 487 -447
rect 287 -497 487 -481
rect 545 -447 745 -400
rect 545 -481 561 -447
rect 729 -481 745 -447
rect 545 -497 745 -481
rect 803 -447 1003 -400
rect 803 -481 819 -447
rect 987 -481 1003 -447
rect 803 -497 1003 -481
<< polycont >>
rect -987 447 -819 481
rect -729 447 -561 481
rect -471 447 -303 481
rect -213 447 -45 481
rect 45 447 213 481
rect 303 447 471 481
rect 561 447 729 481
rect 819 447 987 481
rect -987 -481 -819 -447
rect -729 -481 -561 -447
rect -471 -481 -303 -447
rect -213 -481 -45 -447
rect 45 -481 213 -447
rect 303 -481 471 -447
rect 561 -481 729 -447
rect 819 -481 987 -447
<< locali >>
rect -1183 585 -1087 619
rect 1087 585 1183 619
rect -1183 523 -1149 585
rect 1149 523 1183 585
rect -1003 447 -987 481
rect -819 447 -803 481
rect -745 447 -729 481
rect -561 447 -545 481
rect -487 447 -471 481
rect -303 447 -287 481
rect -229 447 -213 481
rect -45 447 -29 481
rect 29 447 45 481
rect 213 447 229 481
rect 287 447 303 481
rect 471 447 487 481
rect 545 447 561 481
rect 729 447 745 481
rect 803 447 819 481
rect 987 447 1003 481
rect -1049 388 -1015 404
rect -1049 -404 -1015 -388
rect -791 388 -757 404
rect -791 -404 -757 -388
rect -533 388 -499 404
rect -533 -404 -499 -388
rect -275 388 -241 404
rect -275 -404 -241 -388
rect -17 388 17 404
rect -17 -404 17 -388
rect 241 388 275 404
rect 241 -404 275 -388
rect 499 388 533 404
rect 499 -404 533 -388
rect 757 388 791 404
rect 757 -404 791 -388
rect 1015 388 1049 404
rect 1015 -404 1049 -388
rect -1003 -481 -987 -447
rect -819 -481 -803 -447
rect -745 -481 -729 -447
rect -561 -481 -545 -447
rect -487 -481 -471 -447
rect -303 -481 -287 -447
rect -229 -481 -213 -447
rect -45 -481 -29 -447
rect 29 -481 45 -447
rect 213 -481 229 -447
rect 287 -481 303 -447
rect 471 -481 487 -447
rect 545 -481 561 -447
rect 729 -481 745 -447
rect 803 -481 819 -447
rect 987 -481 1003 -447
rect -1183 -585 -1149 -523
rect 1149 -585 1183 -523
rect -1183 -619 -1087 -585
rect 1087 -619 1183 -585
<< viali >>
rect -970 447 -836 481
rect -712 447 -578 481
rect -454 447 -320 481
rect -196 447 -62 481
rect 62 447 196 481
rect 320 447 454 481
rect 578 447 712 481
rect 836 447 970 481
rect -1049 -388 -1015 388
rect -791 -388 -757 388
rect -533 -388 -499 388
rect -275 -388 -241 388
rect -17 -388 17 388
rect 241 -388 275 388
rect 499 -388 533 388
rect 757 -388 791 388
rect 1015 -388 1049 388
rect -970 -481 -836 -447
rect -712 -481 -578 -447
rect -454 -481 -320 -447
rect -196 -481 -62 -447
rect 62 -481 196 -447
rect 320 -481 454 -447
rect 578 -481 712 -447
rect 836 -481 970 -447
<< metal1 >>
rect -982 481 -824 487
rect -982 447 -970 481
rect -836 447 -824 481
rect -982 441 -824 447
rect -724 481 -566 487
rect -724 447 -712 481
rect -578 447 -566 481
rect -724 441 -566 447
rect -466 481 -308 487
rect -466 447 -454 481
rect -320 447 -308 481
rect -466 441 -308 447
rect -208 481 -50 487
rect -208 447 -196 481
rect -62 447 -50 481
rect -208 441 -50 447
rect 50 481 208 487
rect 50 447 62 481
rect 196 447 208 481
rect 50 441 208 447
rect 308 481 466 487
rect 308 447 320 481
rect 454 447 466 481
rect 308 441 466 447
rect 566 481 724 487
rect 566 447 578 481
rect 712 447 724 481
rect 566 441 724 447
rect 824 481 982 487
rect 824 447 836 481
rect 970 447 982 481
rect 824 441 982 447
rect -1055 388 -1009 400
rect -1055 -388 -1049 388
rect -1015 -388 -1009 388
rect -1055 -400 -1009 -388
rect -797 388 -751 400
rect -797 -388 -791 388
rect -757 -388 -751 388
rect -797 -400 -751 -388
rect -539 388 -493 400
rect -539 -388 -533 388
rect -499 -388 -493 388
rect -539 -400 -493 -388
rect -281 388 -235 400
rect -281 -388 -275 388
rect -241 -388 -235 388
rect -281 -400 -235 -388
rect -23 388 23 400
rect -23 -388 -17 388
rect 17 -388 23 388
rect -23 -400 23 -388
rect 235 388 281 400
rect 235 -388 241 388
rect 275 -388 281 388
rect 235 -400 281 -388
rect 493 388 539 400
rect 493 -388 499 388
rect 533 -388 539 388
rect 493 -400 539 -388
rect 751 388 797 400
rect 751 -388 757 388
rect 791 -388 797 388
rect 751 -400 797 -388
rect 1009 388 1055 400
rect 1009 -388 1015 388
rect 1049 -388 1055 388
rect 1009 -400 1055 -388
rect -982 -447 -824 -441
rect -982 -481 -970 -447
rect -836 -481 -824 -447
rect -982 -487 -824 -481
rect -724 -447 -566 -441
rect -724 -481 -712 -447
rect -578 -481 -566 -447
rect -724 -487 -566 -481
rect -466 -447 -308 -441
rect -466 -481 -454 -447
rect -320 -481 -308 -447
rect -466 -487 -308 -481
rect -208 -447 -50 -441
rect -208 -481 -196 -447
rect -62 -481 -50 -447
rect -208 -487 -50 -481
rect 50 -447 208 -441
rect 50 -481 62 -447
rect 196 -481 208 -447
rect 50 -487 208 -481
rect 308 -447 466 -441
rect 308 -481 320 -447
rect 454 -481 466 -447
rect 308 -487 466 -481
rect 566 -447 724 -441
rect 566 -481 578 -447
rect 712 -481 724 -447
rect 566 -487 724 -481
rect 824 -447 982 -441
rect 824 -481 836 -447
rect 970 -481 982 -447
rect 824 -487 982 -481
<< properties >>
string FIXED_BBOX -1166 -602 1166 602
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 4 l 1 m 1 nf 8 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 80 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
