magic
tech sky130A
magscale 1 2
timestamp 1713548572
<< error_p >>
rect -190 172 -126 178
rect -32 172 32 178
rect 126 172 190 178
rect -190 138 -178 172
rect -32 138 -20 172
rect 126 138 138 172
rect -190 132 -126 138
rect -32 132 32 138
rect 126 132 190 138
rect -190 -138 -126 -132
rect -32 -138 32 -132
rect 126 -138 190 -132
rect -190 -172 -178 -138
rect -32 -172 -20 -138
rect 126 -172 138 -138
rect -190 -178 -126 -172
rect -32 -178 32 -172
rect 126 -178 190 -172
<< pwell >>
rect -436 -358 436 358
<< mvnmos >>
rect -208 -100 -108 100
rect -50 -100 50 100
rect 108 -100 208 100
<< mvndiff >>
rect -266 88 -208 100
rect -266 -88 -254 88
rect -220 -88 -208 88
rect -266 -100 -208 -88
rect -108 88 -50 100
rect -108 -88 -96 88
rect -62 -88 -50 88
rect -108 -100 -50 -88
rect 50 88 108 100
rect 50 -88 62 88
rect 96 -88 108 88
rect 50 -100 108 -88
rect 208 88 266 100
rect 208 -88 220 88
rect 254 -88 266 88
rect 208 -100 266 -88
<< mvndiffc >>
rect -254 -88 -220 88
rect -96 -88 -62 88
rect 62 -88 96 88
rect 220 -88 254 88
<< mvpsubdiff >>
rect -400 310 400 322
rect -400 276 -292 310
rect 292 276 400 310
rect -400 264 400 276
rect -400 214 -342 264
rect -400 -214 -388 214
rect -354 -214 -342 214
rect 342 214 400 264
rect -400 -264 -342 -214
rect 342 -214 354 214
rect 388 -214 400 214
rect 342 -264 400 -214
rect -400 -276 400 -264
rect -400 -310 -292 -276
rect 292 -310 400 -276
rect -400 -322 400 -310
<< mvpsubdiffcont >>
rect -292 276 292 310
rect -388 -214 -354 214
rect 354 -214 388 214
rect -292 -310 292 -276
<< poly >>
rect -208 172 -108 188
rect -208 138 -192 172
rect -124 138 -108 172
rect -208 100 -108 138
rect -50 172 50 188
rect -50 138 -34 172
rect 34 138 50 172
rect -50 100 50 138
rect 108 172 208 188
rect 108 138 124 172
rect 192 138 208 172
rect 108 100 208 138
rect -208 -138 -108 -100
rect -208 -172 -192 -138
rect -124 -172 -108 -138
rect -208 -188 -108 -172
rect -50 -138 50 -100
rect -50 -172 -34 -138
rect 34 -172 50 -138
rect -50 -188 50 -172
rect 108 -138 208 -100
rect 108 -172 124 -138
rect 192 -172 208 -138
rect 108 -188 208 -172
<< polycont >>
rect -192 138 -124 172
rect -34 138 34 172
rect 124 138 192 172
rect -192 -172 -124 -138
rect -34 -172 34 -138
rect 124 -172 192 -138
<< locali >>
rect -388 276 -292 310
rect 292 276 388 310
rect -388 221 -354 276
rect 354 214 388 276
rect -208 138 -192 172
rect -124 138 -108 172
rect -50 138 -34 172
rect 34 138 50 172
rect 108 138 124 172
rect 192 138 208 172
rect -254 88 -220 104
rect -254 -104 -220 -88
rect -96 88 -62 104
rect -96 -104 -62 -88
rect 62 88 96 104
rect 62 -104 96 -88
rect 220 88 254 104
rect 220 -104 254 -88
rect -208 -172 -192 -138
rect -124 -172 -108 -138
rect -50 -172 -34 -138
rect 34 -172 50 -138
rect 108 -172 124 -138
rect 192 -172 208 -138
rect -388 -276 -354 -221
rect 354 -276 388 -214
rect -388 -310 -292 -276
rect 292 -310 388 -276
<< viali >>
rect -388 214 -354 221
rect -388 -214 -354 214
rect -178 138 -138 172
rect -20 138 20 172
rect 138 138 178 172
rect -254 -88 -220 88
rect -96 -88 -62 88
rect 62 -88 96 88
rect 220 -88 254 88
rect -178 -172 -138 -138
rect -20 -172 20 -138
rect 138 -172 178 -138
rect -388 -221 -354 -214
rect -283 -310 283 -276
<< metal1 >>
rect -394 221 -348 233
rect -394 -221 -388 221
rect -354 -221 -348 221
rect -190 172 -126 178
rect -190 138 -178 172
rect -138 138 -126 172
rect -190 132 -126 138
rect -32 172 32 178
rect -32 138 -20 172
rect 20 138 32 172
rect -32 132 32 138
rect 126 172 190 178
rect 126 138 138 172
rect 178 138 190 172
rect 126 132 190 138
rect -260 88 -214 100
rect -260 -88 -254 88
rect -220 -88 -214 88
rect -260 -100 -214 -88
rect -102 88 -56 100
rect -102 -88 -96 88
rect -62 -88 -56 88
rect -102 -100 -56 -88
rect 56 88 102 100
rect 56 -88 62 88
rect 96 -88 102 88
rect 56 -100 102 -88
rect 214 88 260 100
rect 214 -88 220 88
rect 254 -88 260 88
rect 214 -100 260 -88
rect -190 -138 -126 -132
rect -190 -172 -178 -138
rect -138 -172 -126 -138
rect -190 -178 -126 -172
rect -32 -138 32 -132
rect -32 -172 -20 -138
rect 20 -172 32 -138
rect -32 -178 32 -172
rect 126 -138 190 -132
rect 126 -172 138 -138
rect 178 -172 190 -138
rect 126 -178 190 -172
rect -394 -233 -348 -221
rect -295 -276 295 -270
rect -295 -310 -283 -276
rect 283 -310 295 -276
rect -295 -316 295 -310
<< properties >>
string FIXED_BBOX -371 -293 371 293
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 1 l 0.5 m 1 nf 3 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 60 viagb 80 viagr 0 viagl 80 viagt 0
<< end >>
