magic
tech sky130A
magscale 1 2
timestamp 1713585847
<< pwell >>
rect -278 -358 278 358
<< mvnmos >>
rect -50 -100 50 100
<< mvndiff >>
rect -108 88 -50 100
rect -108 -88 -96 88
rect -62 -88 -50 88
rect -108 -100 -50 -88
rect 50 88 108 100
rect 50 -88 62 88
rect 96 -88 108 88
rect 50 -100 108 -88
<< mvndiffc >>
rect -96 -88 -62 88
rect 62 -88 96 88
<< mvpsubdiff >>
rect -242 310 242 322
rect -242 276 -134 310
rect 134 276 242 310
rect -242 264 242 276
rect -242 -264 -184 264
rect 184 -264 242 264
rect -242 -276 242 -264
rect -242 -310 -134 -276
rect 134 -310 242 -276
rect -242 -322 242 -310
<< mvpsubdiffcont >>
rect -134 276 134 310
rect -134 -310 134 -276
<< poly >>
rect -50 172 50 188
rect -50 138 -34 172
rect 34 138 50 172
rect -50 100 50 138
rect -50 -138 50 -100
rect -50 -172 -34 -138
rect 34 -172 50 -138
rect -50 -188 50 -172
<< polycont >>
rect -34 138 34 172
rect -34 -172 34 -138
<< locali >>
rect -230 276 -157 310
rect 157 276 230 310
rect -230 -276 -196 276
rect -50 138 -34 172
rect 34 138 50 172
rect -96 88 -62 104
rect -96 -104 -62 -88
rect 62 88 96 104
rect 62 -104 96 -88
rect -50 -172 -34 -138
rect 34 -172 50 -138
rect 196 -276 230 276
rect -230 -310 -157 -276
rect 157 -310 230 -276
<< viali >>
rect -157 276 -134 310
rect -134 276 134 310
rect 134 276 157 310
rect -34 138 34 172
rect -96 -88 -62 88
rect 62 -88 96 88
rect -34 -172 34 -138
rect -157 -310 -134 -276
rect -134 -310 134 -276
rect 134 -310 157 -276
<< metal1 >>
rect -169 310 169 316
rect -169 276 -157 310
rect 157 276 169 310
rect -169 270 169 276
rect -46 172 46 178
rect -46 138 -34 172
rect 34 138 46 172
rect -46 132 46 138
rect -102 88 -56 100
rect -102 -88 -96 88
rect -62 -88 -56 88
rect -102 -100 -56 -88
rect 56 88 102 100
rect 56 -88 62 88
rect 96 -88 102 88
rect 56 -100 102 -88
rect -46 -138 46 -132
rect -46 -172 -34 -138
rect 34 -172 46 -138
rect -46 -178 46 -172
rect -169 -276 169 -270
rect -169 -310 -157 -276
rect 157 -310 169 -276
rect -169 -316 169 -310
<< properties >>
string FIXED_BBOX -213 -293 213 293
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 1 l 0.50 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 0 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 80 viagr 0 viagl 0 viagt 80
<< end >>
