magic
tech sky130A
magscale 1 2
timestamp 1713074216
<< nwell >>
rect -545 -697 545 697
<< mvpmos >>
rect -287 -400 -187 400
rect -129 -400 -29 400
rect 29 -400 129 400
rect 187 -400 287 400
<< mvpdiff >>
rect -345 388 -287 400
rect -345 -388 -333 388
rect -299 -388 -287 388
rect -345 -400 -287 -388
rect -187 388 -129 400
rect -187 -388 -175 388
rect -141 -388 -129 388
rect -187 -400 -129 -388
rect -29 388 29 400
rect -29 -388 -17 388
rect 17 -388 29 388
rect -29 -400 29 -388
rect 129 388 187 400
rect 129 -388 141 388
rect 175 -388 187 388
rect 129 -400 187 -388
rect 287 388 345 400
rect 287 -388 299 388
rect 333 -388 345 388
rect 287 -400 345 -388
<< mvpdiffc >>
rect -333 -388 -299 388
rect -175 -388 -141 388
rect -17 -388 17 388
rect 141 -388 175 388
rect 299 -388 333 388
<< mvnsubdiff >>
rect -479 619 479 631
rect -479 585 -371 619
rect 371 585 479 619
rect -479 573 479 585
rect -479 523 -421 573
rect -479 -523 -467 523
rect -433 -523 -421 523
rect 421 523 479 573
rect -479 -573 -421 -523
rect 421 -523 433 523
rect 467 -523 479 523
rect 421 -573 479 -523
rect -479 -585 479 -573
rect -479 -619 -371 -585
rect 371 -619 479 -585
rect -479 -631 479 -619
<< mvnsubdiffcont >>
rect -371 585 371 619
rect -467 -523 -433 523
rect 433 -523 467 523
rect -371 -619 371 -585
<< poly >>
rect -287 481 -187 497
rect -287 447 -271 481
rect -203 447 -187 481
rect -287 400 -187 447
rect -129 481 -29 497
rect -129 447 -113 481
rect -45 447 -29 481
rect -129 400 -29 447
rect 29 481 129 497
rect 29 447 45 481
rect 113 447 129 481
rect 29 400 129 447
rect 187 481 287 497
rect 187 447 203 481
rect 271 447 287 481
rect 187 400 287 447
rect -287 -447 -187 -400
rect -287 -481 -271 -447
rect -203 -481 -187 -447
rect -287 -497 -187 -481
rect -129 -447 -29 -400
rect -129 -481 -113 -447
rect -45 -481 -29 -447
rect -129 -497 -29 -481
rect 29 -447 129 -400
rect 29 -481 45 -447
rect 113 -481 129 -447
rect 29 -497 129 -481
rect 187 -447 287 -400
rect 187 -481 203 -447
rect 271 -481 287 -447
rect 187 -497 287 -481
<< polycont >>
rect -271 447 -203 481
rect -113 447 -45 481
rect 45 447 113 481
rect 203 447 271 481
rect -271 -481 -203 -447
rect -113 -481 -45 -447
rect 45 -481 113 -447
rect 203 -481 271 -447
<< locali >>
rect -467 585 -371 619
rect 371 585 467 619
rect -467 523 -433 585
rect 433 523 467 585
rect -287 447 -271 481
rect -203 447 -187 481
rect -129 447 -113 481
rect -45 447 -29 481
rect 29 447 45 481
rect 113 447 129 481
rect 187 447 203 481
rect 271 447 287 481
rect -333 388 -299 404
rect -333 -404 -299 -388
rect -175 388 -141 404
rect -175 -404 -141 -388
rect -17 388 17 404
rect -17 -404 17 -388
rect 141 388 175 404
rect 141 -404 175 -388
rect 299 388 333 404
rect 299 -404 333 -388
rect -287 -481 -271 -447
rect -203 -481 -187 -447
rect -129 -481 -113 -447
rect -45 -481 -29 -447
rect 29 -481 45 -447
rect 113 -481 129 -447
rect 187 -481 203 -447
rect 271 -481 287 -447
rect -467 -585 -433 -523
rect 433 -585 467 -523
rect -467 -619 -371 -585
rect 371 -619 467 -585
<< viali >>
rect -264 447 -210 481
rect -106 447 -52 481
rect 52 447 106 481
rect 210 447 264 481
rect -333 -388 -299 388
rect -175 -388 -141 388
rect -17 -388 17 388
rect 141 -388 175 388
rect 299 -388 333 388
rect -264 -481 -210 -447
rect -106 -481 -52 -447
rect 52 -481 106 -447
rect 210 -481 264 -447
<< metal1 >>
rect -276 481 -198 487
rect -276 447 -264 481
rect -210 447 -198 481
rect -276 441 -198 447
rect -118 481 -40 487
rect -118 447 -106 481
rect -52 447 -40 481
rect -118 441 -40 447
rect 40 481 118 487
rect 40 447 52 481
rect 106 447 118 481
rect 40 441 118 447
rect 198 481 276 487
rect 198 447 210 481
rect 264 447 276 481
rect 198 441 276 447
rect -339 388 -293 400
rect -339 -388 -333 388
rect -299 -388 -293 388
rect -339 -400 -293 -388
rect -181 388 -135 400
rect -181 -388 -175 388
rect -141 -388 -135 388
rect -181 -400 -135 -388
rect -23 388 23 400
rect -23 -388 -17 388
rect 17 -388 23 388
rect -23 -400 23 -388
rect 135 388 181 400
rect 135 -388 141 388
rect 175 -388 181 388
rect 135 -400 181 -388
rect 293 388 339 400
rect 293 -388 299 388
rect 333 -388 339 388
rect 293 -400 339 -388
rect -276 -447 -198 -441
rect -276 -481 -264 -447
rect -210 -481 -198 -447
rect -276 -487 -198 -481
rect -118 -447 -40 -441
rect -118 -481 -106 -447
rect -52 -481 -40 -447
rect -118 -487 -40 -481
rect 40 -447 118 -441
rect 40 -481 52 -447
rect 106 -481 118 -447
rect 40 -487 118 -481
rect 198 -447 276 -441
rect 198 -481 210 -447
rect 264 -481 276 -447
rect 198 -487 276 -481
<< properties >>
string FIXED_BBOX -450 -602 450 602
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 4 l 0.5 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 80 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
